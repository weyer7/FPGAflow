magic
tech sky130A
magscale 1 2
timestamp 1737231330
<< viali >>
rect 7021 37281 7055 37315
rect 8125 37281 8159 37315
rect 10241 37281 10275 37315
rect 11253 37281 11287 37315
rect 12817 37281 12851 37315
rect 17233 37281 17267 37315
rect 17509 37281 17543 37315
rect 6837 37213 6871 37247
rect 7941 37213 7975 37247
rect 10057 37213 10091 37247
rect 11069 37213 11103 37247
rect 12633 37213 12667 37247
rect 17141 37213 17175 37247
rect 6745 37145 6779 37179
rect 6377 37077 6411 37111
rect 7481 37077 7515 37111
rect 7849 37077 7883 37111
rect 9597 37077 9631 37111
rect 9965 37077 9999 37111
rect 10609 37077 10643 37111
rect 10977 37077 11011 37111
rect 12173 37077 12207 37111
rect 12541 37077 12575 37111
rect 4445 36805 4479 36839
rect 8677 36805 8711 36839
rect 10793 36805 10827 36839
rect 11897 36805 11931 36839
rect 6193 36737 6227 36771
rect 17417 36737 17451 36771
rect 18153 36737 18187 36771
rect 18705 36737 18739 36771
rect 19165 36737 19199 36771
rect 4169 36669 4203 36703
rect 6653 36669 6687 36703
rect 6929 36669 6963 36703
rect 8769 36669 8803 36703
rect 9045 36669 9079 36703
rect 11621 36669 11655 36703
rect 13645 36669 13679 36703
rect 14013 36669 14047 36703
rect 14289 36669 14323 36703
rect 15761 36669 15795 36703
rect 17509 36669 17543 36703
rect 18245 36669 18279 36703
rect 19441 36669 19475 36703
rect 19625 36669 19659 36703
rect 19901 36669 19935 36703
rect 21649 36669 21683 36703
rect 22845 36669 22879 36703
rect 23121 36669 23155 36703
rect 24869 36669 24903 36703
rect 24961 36669 24995 36703
rect 25237 36669 25271 36703
rect 17785 36601 17819 36635
rect 17049 36533 17083 36567
rect 26709 36533 26743 36567
rect 8953 36329 8987 36363
rect 18153 36329 18187 36363
rect 19993 36329 20027 36363
rect 25145 36329 25179 36363
rect 19441 36261 19475 36295
rect 19717 36261 19751 36295
rect 6469 36193 6503 36227
rect 6745 36193 6779 36227
rect 8493 36193 8527 36227
rect 9597 36193 9631 36227
rect 10609 36193 10643 36227
rect 12357 36193 12391 36227
rect 13185 36193 13219 36227
rect 14933 36193 14967 36227
rect 15117 36193 15151 36227
rect 17969 36193 18003 36227
rect 19533 36193 19567 36227
rect 19625 36193 19659 36227
rect 20637 36193 20671 36227
rect 23397 36193 23431 36227
rect 25697 36193 25731 36227
rect 9413 36125 9447 36159
rect 10333 36125 10367 36159
rect 13277 36125 13311 36159
rect 14657 36125 14691 36159
rect 14749 36125 14783 36159
rect 15025 36125 15059 36159
rect 17141 36125 17175 36159
rect 17325 36125 17359 36159
rect 17877 36125 17911 36159
rect 19257 36125 19291 36159
rect 19349 36125 19383 36159
rect 19809 36125 19843 36159
rect 19901 36125 19935 36159
rect 24041 36125 24075 36159
rect 24225 36125 24259 36159
rect 24593 36125 24627 36159
rect 25605 36125 25639 36159
rect 26065 36125 26099 36159
rect 26249 36125 26283 36159
rect 26341 36125 26375 36159
rect 26525 36125 26559 36159
rect 9321 36057 9355 36091
rect 15393 36057 15427 36091
rect 23121 36057 23155 36091
rect 24409 36057 24443 36091
rect 26433 36057 26467 36091
rect 13645 35989 13679 36023
rect 14473 35989 14507 36023
rect 16865 35989 16899 36023
rect 17233 35989 17267 36023
rect 17509 35989 17543 36023
rect 20361 35989 20395 36023
rect 20453 35989 20487 36023
rect 21649 35989 21683 36023
rect 24225 35989 24259 36023
rect 24777 35989 24811 36023
rect 25513 35989 25547 36023
rect 26157 35989 26191 36023
rect 9597 35785 9631 35819
rect 13001 35785 13035 35819
rect 13737 35785 13771 35819
rect 15025 35785 15059 35819
rect 17969 35785 18003 35819
rect 19441 35785 19475 35819
rect 20177 35785 20211 35819
rect 22477 35785 22511 35819
rect 23213 35785 23247 35819
rect 23581 35785 23615 35819
rect 24317 35785 24351 35819
rect 24685 35785 24719 35819
rect 25897 35785 25931 35819
rect 26525 35785 26559 35819
rect 13645 35717 13679 35751
rect 16221 35717 16255 35751
rect 17417 35717 17451 35751
rect 18153 35717 18187 35751
rect 22845 35717 22879 35751
rect 25697 35717 25731 35751
rect 9229 35649 9263 35683
rect 9873 35649 9907 35683
rect 12449 35649 12483 35683
rect 12633 35649 12667 35683
rect 12723 35649 12757 35683
rect 12909 35649 12943 35683
rect 13185 35649 13219 35683
rect 14289 35649 14323 35683
rect 14381 35649 14415 35683
rect 14473 35649 14507 35683
rect 15209 35649 15243 35683
rect 15577 35649 15611 35683
rect 15761 35649 15795 35683
rect 15853 35649 15887 35683
rect 16037 35649 16071 35683
rect 16681 35649 16715 35683
rect 17049 35649 17083 35683
rect 17141 35649 17175 35683
rect 17877 35649 17911 35683
rect 19165 35649 19199 35683
rect 19901 35649 19935 35683
rect 20545 35649 20579 35683
rect 21281 35649 21315 35683
rect 21833 35649 21867 35683
rect 21926 35649 21960 35683
rect 22063 35649 22097 35683
rect 22201 35649 22235 35683
rect 22339 35649 22373 35683
rect 22569 35649 22603 35683
rect 22662 35649 22696 35683
rect 22937 35649 22971 35683
rect 23034 35649 23068 35683
rect 23305 35649 23339 35683
rect 23489 35649 23523 35683
rect 23949 35649 23983 35683
rect 24225 35649 24259 35683
rect 24501 35649 24535 35683
rect 24777 35649 24811 35683
rect 24961 35649 24995 35683
rect 25053 35649 25087 35683
rect 25329 35649 25363 35683
rect 26157 35649 26191 35683
rect 26341 35649 26375 35683
rect 6377 35581 6411 35615
rect 6653 35581 6687 35615
rect 8401 35581 8435 35615
rect 9321 35581 9355 35615
rect 9965 35581 9999 35615
rect 13829 35581 13863 35615
rect 14197 35581 14231 35615
rect 15393 35581 15427 35615
rect 15485 35581 15519 35615
rect 19809 35581 19843 35615
rect 20637 35581 20671 35615
rect 20821 35581 20855 35615
rect 21189 35581 21223 35615
rect 21649 35581 21683 35615
rect 24041 35581 24075 35615
rect 24869 35581 24903 35615
rect 10241 35513 10275 35547
rect 13185 35513 13219 35547
rect 13277 35513 13311 35547
rect 18153 35513 18187 35547
rect 26065 35513 26099 35547
rect 12725 35445 12759 35479
rect 14657 35445 14691 35479
rect 16865 35445 16899 35479
rect 16957 35445 16991 35479
rect 19073 35445 19107 35479
rect 20085 35445 20119 35479
rect 23397 35445 23431 35479
rect 25421 35445 25455 35479
rect 25605 35445 25639 35479
rect 25881 35445 25915 35479
rect 7021 35241 7055 35275
rect 9321 35241 9355 35275
rect 9873 35241 9907 35275
rect 12633 35241 12667 35275
rect 12817 35241 12851 35275
rect 13461 35241 13495 35275
rect 14197 35241 14231 35275
rect 14565 35241 14599 35275
rect 20085 35241 20119 35275
rect 21741 35241 21775 35275
rect 22661 35241 22695 35275
rect 22753 35241 22787 35275
rect 25237 35241 25271 35275
rect 25513 35241 25547 35275
rect 26065 35241 26099 35275
rect 26341 35241 26375 35275
rect 26525 35241 26559 35275
rect 26985 35241 27019 35275
rect 13277 35173 13311 35207
rect 23029 35173 23063 35207
rect 4905 35105 4939 35139
rect 6929 35105 6963 35139
rect 7481 35105 7515 35139
rect 7573 35105 7607 35139
rect 11437 35105 11471 35139
rect 12541 35105 12575 35139
rect 14105 35105 14139 35139
rect 16773 35105 16807 35139
rect 17049 35105 17083 35139
rect 19901 35105 19935 35139
rect 22845 35105 22879 35139
rect 25605 35105 25639 35139
rect 26801 35105 26835 35139
rect 9229 35037 9263 35071
rect 9413 35037 9447 35071
rect 9689 35037 9723 35071
rect 9873 35037 9907 35071
rect 10149 35037 10183 35071
rect 11345 35037 11379 35071
rect 12633 35037 12667 35071
rect 12725 35037 12759 35071
rect 13001 35037 13035 35071
rect 13369 35037 13403 35071
rect 13645 35037 13679 35071
rect 14381 35037 14415 35071
rect 16681 35037 16715 35071
rect 17877 35037 17911 35071
rect 18153 35037 18187 35071
rect 18245 35037 18279 35071
rect 18337 35037 18371 35071
rect 18521 35037 18555 35071
rect 18613 35037 18647 35071
rect 19809 35037 19843 35071
rect 21747 35037 21781 35071
rect 21925 35037 21959 35071
rect 22293 35037 22327 35071
rect 22569 35037 22603 35071
rect 22937 35037 22971 35071
rect 23121 35037 23155 35071
rect 24777 35037 24811 35071
rect 24869 35037 24903 35071
rect 25053 35037 25087 35071
rect 25329 35037 25363 35071
rect 25421 35037 25455 35071
rect 26525 35037 26559 35071
rect 26709 35037 26743 35071
rect 27077 35037 27111 35071
rect 5181 34969 5215 35003
rect 13093 34969 13127 35003
rect 13277 34969 13311 35003
rect 13829 34969 13863 35003
rect 22109 34969 22143 35003
rect 22477 34969 22511 35003
rect 25881 34969 25915 35003
rect 26097 34969 26131 35003
rect 26801 34969 26835 35003
rect 7389 34901 7423 34935
rect 11713 34901 11747 34935
rect 12265 34901 12299 34935
rect 26249 34901 26283 34935
rect 6377 34697 6411 34731
rect 6837 34697 6871 34731
rect 9137 34697 9171 34731
rect 9597 34697 9631 34731
rect 11529 34697 11563 34731
rect 13001 34697 13035 34731
rect 19257 34697 19291 34731
rect 10149 34629 10183 34663
rect 22661 34629 22695 34663
rect 6745 34561 6779 34595
rect 8309 34561 8343 34595
rect 9229 34561 9263 34595
rect 9965 34561 9999 34595
rect 10057 34561 10091 34595
rect 10241 34561 10275 34595
rect 11897 34561 11931 34595
rect 12357 34561 12391 34595
rect 12817 34561 12851 34595
rect 13001 34561 13035 34595
rect 15025 34561 15059 34595
rect 15209 34561 15243 34595
rect 15853 34561 15887 34595
rect 16773 34561 16807 34595
rect 16957 34561 16991 34595
rect 17693 34561 17727 34595
rect 18429 34561 18463 34595
rect 18521 34561 18555 34595
rect 18705 34561 18739 34595
rect 18889 34561 18923 34595
rect 18981 34561 19015 34595
rect 22201 34561 22235 34595
rect 22293 34561 22327 34595
rect 22477 34561 22511 34595
rect 23213 34561 23247 34595
rect 23305 34561 23339 34595
rect 23489 34561 23523 34595
rect 25605 34561 25639 34595
rect 25881 34561 25915 34595
rect 25973 34561 26007 34595
rect 26426 34561 26460 34595
rect 7021 34493 7055 34527
rect 8401 34493 8435 34527
rect 9413 34493 9447 34527
rect 9873 34493 9907 34527
rect 11989 34493 12023 34527
rect 12081 34493 12115 34527
rect 12449 34493 12483 34527
rect 14933 34493 14967 34527
rect 15761 34493 15795 34527
rect 16865 34493 16899 34527
rect 17601 34493 17635 34527
rect 18061 34493 18095 34527
rect 19257 34493 19291 34527
rect 26525 34493 26559 34527
rect 26801 34493 26835 34527
rect 8677 34425 8711 34459
rect 8769 34425 8803 34459
rect 12725 34425 12759 34459
rect 18613 34425 18647 34459
rect 19073 34425 19107 34459
rect 25697 34425 25731 34459
rect 9965 34357 9999 34391
rect 12357 34357 12391 34391
rect 15393 34357 15427 34391
rect 15485 34357 15519 34391
rect 15669 34357 15703 34391
rect 18245 34357 18279 34391
rect 23673 34357 23707 34391
rect 26157 34357 26191 34391
rect 10057 34153 10091 34187
rect 11529 34153 11563 34187
rect 17969 34153 18003 34187
rect 23121 34153 23155 34187
rect 27537 34153 27571 34187
rect 21649 34085 21683 34119
rect 6745 34017 6779 34051
rect 8769 34017 8803 34051
rect 10241 34017 10275 34051
rect 11161 34017 11195 34051
rect 11989 34017 12023 34051
rect 15393 34017 15427 34051
rect 17233 34017 17267 34051
rect 17509 34017 17543 34051
rect 19257 34017 19291 34051
rect 22661 34017 22695 34051
rect 25789 34017 25823 34051
rect 26065 34017 26099 34051
rect 8953 33949 8987 33983
rect 9413 33949 9447 33983
rect 9898 33949 9932 33983
rect 10149 33949 10183 33983
rect 10885 33949 10919 33983
rect 11897 33949 11931 33983
rect 12081 33949 12115 33983
rect 14197 33949 14231 33983
rect 14657 33949 14691 33983
rect 14841 33949 14875 33983
rect 14933 33949 14967 33983
rect 15025 33949 15059 33983
rect 15209 33949 15243 33983
rect 17601 33949 17635 33983
rect 17785 33949 17819 33983
rect 18429 33949 18463 33983
rect 18522 33949 18556 33983
rect 18797 33949 18831 33983
rect 18894 33949 18928 33983
rect 21281 33949 21315 33983
rect 21833 33949 21867 33983
rect 21925 33949 21959 33983
rect 22753 33949 22787 33983
rect 23489 33949 23523 33983
rect 7021 33881 7055 33915
rect 11370 33881 11404 33915
rect 14381 33881 14415 33915
rect 14565 33881 14599 33915
rect 15485 33881 15519 33915
rect 18705 33881 18739 33915
rect 19540 33881 19574 33915
rect 24133 33881 24167 33915
rect 9137 33813 9171 33847
rect 9689 33813 9723 33847
rect 9781 33813 9815 33847
rect 11253 33813 11287 33847
rect 19073 33813 19107 33847
rect 24041 33813 24075 33847
rect 8861 33609 8895 33643
rect 9597 33609 9631 33643
rect 11729 33609 11763 33643
rect 11897 33609 11931 33643
rect 14841 33609 14875 33643
rect 15117 33609 15151 33643
rect 16957 33609 16991 33643
rect 23029 33609 23063 33643
rect 9965 33541 9999 33575
rect 10149 33541 10183 33575
rect 11529 33541 11563 33575
rect 12265 33541 12299 33575
rect 15577 33541 15611 33575
rect 22753 33541 22787 33575
rect 23397 33541 23431 33575
rect 25237 33541 25271 33575
rect 25421 33541 25455 33575
rect 6377 33473 6411 33507
rect 8493 33473 8527 33507
rect 8677 33473 8711 33507
rect 8769 33473 8803 33507
rect 8953 33473 8987 33507
rect 9781 33473 9815 33507
rect 9873 33473 9907 33507
rect 11069 33473 11103 33507
rect 11161 33473 11195 33507
rect 11345 33473 11379 33507
rect 11989 33473 12023 33507
rect 14289 33473 14323 33507
rect 14657 33473 14691 33507
rect 16865 33473 16899 33507
rect 17049 33473 17083 33507
rect 21189 33473 21223 33507
rect 21373 33473 21407 33507
rect 21649 33473 21683 33507
rect 21833 33473 21867 33507
rect 22109 33473 22143 33507
rect 22477 33473 22511 33507
rect 22661 33473 22695 33507
rect 22845 33473 22879 33507
rect 23121 33473 23155 33507
rect 25053 33473 25087 33507
rect 6653 33405 6687 33439
rect 8401 33405 8435 33439
rect 8585 33405 8619 33439
rect 12081 33405 12115 33439
rect 14013 33405 14047 33439
rect 14473 33405 14507 33439
rect 24869 33405 24903 33439
rect 11345 33337 11379 33371
rect 15301 33337 15335 33371
rect 22109 33337 22143 33371
rect 11713 33269 11747 33303
rect 21005 33269 21039 33303
rect 21557 33269 21591 33303
rect 7021 33065 7055 33099
rect 10885 33065 10919 33099
rect 11161 33065 11195 33099
rect 11253 33065 11287 33099
rect 13461 33065 13495 33099
rect 22477 33065 22511 33099
rect 18889 32997 18923 33031
rect 7665 32929 7699 32963
rect 13185 32929 13219 32963
rect 13277 32929 13311 32963
rect 15301 32929 15335 32963
rect 18705 32929 18739 32963
rect 20177 32929 20211 32963
rect 23029 32929 23063 32963
rect 25237 32929 25271 32963
rect 27629 32929 27663 32963
rect 29561 32929 29595 32963
rect 7481 32861 7515 32895
rect 10793 32861 10827 32895
rect 10885 32861 10919 32895
rect 11253 32861 11287 32895
rect 11437 32861 11471 32895
rect 14381 32861 14415 32895
rect 14565 32861 14599 32895
rect 14657 32861 14691 32895
rect 14841 32861 14875 32895
rect 14933 32861 14967 32895
rect 15117 32861 15151 32895
rect 15393 32861 15427 32895
rect 15485 32861 15519 32895
rect 15669 32861 15703 32895
rect 17877 32861 17911 32895
rect 18061 32861 18095 32895
rect 18153 32861 18187 32895
rect 18245 32861 18279 32895
rect 18429 32861 18463 32895
rect 18981 32861 19015 32895
rect 23489 32861 23523 32895
rect 24409 32861 24443 32895
rect 29193 32861 29227 32895
rect 29929 32861 29963 32895
rect 12817 32793 12851 32827
rect 14473 32793 14507 32827
rect 14749 32793 14783 32827
rect 18705 32793 18739 32827
rect 20453 32793 20487 32827
rect 24225 32793 24259 32827
rect 25053 32793 25087 32827
rect 25605 32793 25639 32827
rect 27353 32793 27387 32827
rect 7389 32725 7423 32759
rect 15577 32725 15611 32759
rect 18613 32725 18647 32759
rect 21925 32725 21959 32759
rect 22845 32725 22879 32759
rect 22937 32725 22971 32759
rect 24501 32725 24535 32759
rect 24685 32725 24719 32759
rect 25145 32725 25179 32759
rect 28641 32725 28675 32759
rect 31355 32725 31389 32759
rect 11069 32521 11103 32555
rect 11897 32521 11931 32555
rect 12541 32521 12575 32555
rect 15209 32521 15243 32555
rect 17509 32521 17543 32555
rect 19993 32521 20027 32555
rect 20545 32521 20579 32555
rect 22569 32521 22603 32555
rect 25329 32521 25363 32555
rect 5089 32453 5123 32487
rect 8401 32453 8435 32487
rect 14841 32453 14875 32487
rect 14933 32453 14967 32487
rect 23489 32453 23523 32487
rect 24685 32453 24719 32487
rect 4905 32385 4939 32419
rect 5181 32385 5215 32419
rect 8953 32385 8987 32419
rect 9413 32385 9447 32419
rect 9597 32385 9631 32419
rect 10609 32385 10643 32419
rect 10885 32385 10919 32419
rect 11161 32385 11195 32419
rect 11529 32385 11563 32419
rect 11713 32385 11747 32419
rect 12173 32385 12207 32419
rect 13001 32385 13035 32419
rect 14749 32385 14783 32419
rect 15117 32385 15151 32419
rect 15485 32385 15519 32419
rect 15577 32385 15611 32419
rect 15669 32385 15703 32419
rect 15853 32385 15887 32419
rect 15945 32385 15979 32419
rect 16129 32385 16163 32419
rect 16681 32385 16715 32419
rect 17141 32385 17175 32419
rect 17325 32385 17359 32419
rect 17693 32385 17727 32419
rect 17785 32385 17819 32419
rect 17969 32385 18003 32419
rect 18245 32385 18279 32419
rect 20729 32385 20763 32419
rect 20913 32385 20947 32419
rect 22017 32385 22051 32419
rect 22109 32385 22143 32419
rect 22201 32385 22235 32419
rect 22753 32385 22787 32419
rect 23029 32385 23063 32419
rect 24225 32385 24259 32419
rect 24409 32385 24443 32419
rect 24501 32385 24535 32419
rect 24961 32385 24995 32419
rect 25421 32385 25455 32419
rect 25605 32385 25639 32419
rect 25697 32385 25731 32419
rect 25973 32385 26007 32419
rect 30573 32385 30607 32419
rect 30665 32385 30699 32419
rect 31125 32385 31159 32419
rect 31309 32385 31343 32419
rect 31493 32385 31527 32419
rect 32137 32385 32171 32419
rect 6377 32317 6411 32351
rect 6653 32317 6687 32351
rect 9045 32317 9079 32351
rect 9505 32317 9539 32351
rect 10701 32317 10735 32351
rect 12081 32317 12115 32351
rect 12817 32317 12851 32351
rect 12909 32317 12943 32351
rect 13093 32317 13127 32351
rect 16957 32317 16991 32351
rect 17877 32317 17911 32351
rect 21005 32317 21039 32351
rect 21833 32317 21867 32351
rect 24869 32317 24903 32351
rect 26985 32317 27019 32351
rect 27261 32317 27295 32351
rect 30297 32317 30331 32351
rect 30941 32317 30975 32351
rect 32505 32317 32539 32351
rect 33931 32317 33965 32351
rect 34621 32317 34655 32351
rect 9321 32249 9355 32283
rect 11253 32249 11287 32283
rect 14565 32249 14599 32283
rect 16865 32249 16899 32283
rect 22385 32249 22419 32283
rect 26065 32249 26099 32283
rect 28825 32249 28859 32283
rect 4721 32181 4755 32215
rect 10885 32181 10919 32215
rect 11529 32181 11563 32215
rect 12633 32181 12667 32215
rect 15393 32181 15427 32215
rect 15853 32181 15887 32215
rect 16129 32181 16163 32215
rect 16773 32181 16807 32215
rect 17325 32181 17359 32215
rect 18508 32181 18542 32215
rect 21925 32181 21959 32215
rect 22937 32181 22971 32215
rect 25421 32181 25455 32215
rect 25789 32181 25823 32215
rect 28733 32181 28767 32215
rect 34069 32181 34103 32215
rect 7113 31977 7147 32011
rect 9505 31977 9539 32011
rect 9597 31977 9631 32011
rect 10425 31977 10459 32011
rect 11161 31977 11195 32011
rect 11989 31977 12023 32011
rect 12344 31977 12378 32011
rect 13829 31977 13863 32011
rect 15393 31977 15427 32011
rect 17969 31977 18003 32011
rect 18061 31977 18095 32011
rect 18797 31977 18831 32011
rect 20821 31977 20855 32011
rect 22753 31977 22787 32011
rect 24409 31977 24443 32011
rect 25145 31977 25179 32011
rect 27445 31977 27479 32011
rect 28457 31977 28491 32011
rect 29009 31977 29043 32011
rect 30573 31977 30607 32011
rect 6377 31909 6411 31943
rect 8953 31909 8987 31943
rect 10609 31909 10643 31943
rect 15945 31909 15979 31943
rect 16313 31909 16347 31943
rect 16865 31909 16899 31943
rect 17601 31909 17635 31943
rect 18429 31909 18463 31943
rect 22109 31909 22143 31943
rect 23121 31909 23155 31943
rect 24041 31909 24075 31943
rect 24133 31909 24167 31943
rect 24961 31909 24995 31943
rect 29377 31909 29411 31943
rect 5549 31841 5583 31875
rect 5825 31841 5859 31875
rect 7573 31841 7607 31875
rect 7757 31841 7791 31875
rect 8401 31841 8435 31875
rect 11345 31841 11379 31875
rect 11529 31841 11563 31875
rect 16681 31841 16715 31875
rect 16773 31841 16807 31875
rect 18889 31841 18923 31875
rect 20361 31841 20395 31875
rect 23949 31841 23983 31875
rect 28089 31841 28123 31875
rect 29101 31841 29135 31875
rect 30297 31841 30331 31875
rect 32045 31841 32079 31875
rect 32321 31841 32355 31875
rect 32781 31841 32815 31875
rect 33057 31841 33091 31875
rect 34529 31841 34563 31875
rect 35265 31841 35299 31875
rect 3801 31773 3835 31807
rect 6561 31773 6595 31807
rect 6745 31773 6779 31807
rect 6837 31773 6871 31807
rect 8125 31773 8159 31807
rect 8585 31773 8619 31807
rect 8677 31773 8711 31807
rect 9965 31773 9999 31807
rect 10333 31773 10367 31807
rect 10425 31773 10459 31807
rect 10701 31773 10735 31807
rect 10793 31773 10827 31807
rect 10977 31773 11011 31807
rect 11621 31773 11655 31807
rect 12081 31773 12115 31807
rect 15025 31773 15059 31807
rect 15209 31773 15243 31807
rect 15853 31773 15887 31807
rect 16037 31773 16071 31807
rect 16129 31773 16163 31807
rect 16543 31773 16577 31807
rect 17049 31773 17083 31807
rect 17141 31773 17175 31807
rect 17417 31773 17451 31807
rect 17877 31773 17911 31807
rect 18199 31773 18233 31807
rect 18337 31773 18371 31807
rect 18613 31773 18647 31807
rect 19257 31773 19291 31807
rect 19441 31773 19475 31807
rect 19625 31773 19659 31807
rect 19717 31773 19751 31807
rect 19993 31773 20027 31807
rect 20085 31773 20119 31807
rect 20269 31773 20303 31807
rect 20453 31773 20487 31807
rect 21005 31773 21039 31807
rect 21189 31773 21223 31807
rect 21373 31773 21407 31807
rect 21465 31773 21499 31807
rect 21649 31773 21683 31807
rect 22293 31773 22327 31807
rect 22477 31773 22511 31807
rect 23029 31773 23063 31807
rect 23213 31773 23247 31807
rect 23581 31773 23615 31807
rect 24225 31773 24259 31807
rect 24593 31773 24627 31807
rect 24869 31773 24903 31807
rect 27629 31773 27663 31807
rect 28733 31773 28767 31807
rect 29193 31773 29227 31807
rect 29561 31773 29595 31807
rect 32689 31773 32723 31807
rect 28411 31739 28445 31773
rect 9321 31705 9355 31739
rect 9781 31705 9815 31739
rect 10149 31705 10183 31739
rect 21097 31705 21131 31739
rect 22937 31705 22971 31739
rect 25329 31705 25363 31739
rect 27721 31705 27755 31739
rect 27813 31705 27847 31739
rect 27951 31705 27985 31739
rect 28641 31705 28675 31739
rect 7481 31637 7515 31671
rect 8033 31637 8067 31671
rect 8677 31637 8711 31671
rect 9137 31637 9171 31671
rect 9229 31637 9263 31671
rect 15669 31637 15703 31671
rect 19809 31637 19843 31671
rect 21833 31637 21867 31671
rect 22569 31637 22603 31671
rect 22737 31637 22771 31671
rect 24777 31637 24811 31671
rect 25119 31637 25153 31671
rect 28273 31637 28307 31671
rect 32505 31637 32539 31671
rect 34713 31637 34747 31671
rect 5273 31433 5307 31467
rect 7573 31433 7607 31467
rect 9873 31433 9907 31467
rect 11161 31433 11195 31467
rect 11897 31433 11931 31467
rect 15669 31433 15703 31467
rect 18889 31433 18923 31467
rect 19441 31433 19475 31467
rect 19625 31433 19659 31467
rect 24685 31433 24719 31467
rect 28365 31433 28399 31467
rect 32321 31433 32355 31467
rect 33517 31433 33551 31467
rect 33885 31433 33919 31467
rect 6469 31365 6503 31399
rect 8033 31365 8067 31399
rect 9689 31365 9723 31399
rect 10793 31365 10827 31399
rect 11529 31365 11563 31399
rect 11713 31365 11747 31399
rect 13277 31365 13311 31399
rect 18153 31365 18187 31399
rect 22569 31365 22603 31399
rect 23857 31365 23891 31399
rect 24593 31365 24627 31399
rect 27353 31365 27387 31399
rect 27629 31365 27663 31399
rect 27997 31365 28031 31399
rect 28089 31365 28123 31399
rect 32597 31365 32631 31399
rect 34437 31365 34471 31399
rect 6101 31297 6135 31331
rect 7297 31297 7331 31331
rect 7757 31297 7791 31331
rect 7941 31297 7975 31331
rect 9229 31297 9263 31331
rect 9505 31297 9539 31331
rect 9965 31297 9999 31331
rect 10333 31297 10367 31331
rect 10977 31297 11011 31331
rect 11805 31297 11839 31331
rect 11897 31297 11931 31331
rect 12081 31297 12115 31331
rect 13093 31297 13127 31331
rect 13369 31297 13403 31331
rect 13461 31297 13495 31331
rect 13737 31297 13771 31331
rect 15577 31297 15611 31331
rect 15761 31297 15795 31331
rect 18429 31297 18463 31331
rect 18705 31297 18739 31331
rect 19349 31297 19383 31331
rect 19441 31297 19475 31331
rect 19533 31297 19567 31331
rect 19717 31297 19751 31331
rect 20085 31297 20119 31331
rect 20269 31297 20303 31331
rect 20361 31297 20395 31331
rect 20545 31297 20579 31331
rect 20821 31297 20855 31331
rect 21281 31297 21315 31331
rect 21465 31297 21499 31331
rect 22017 31297 22051 31331
rect 22477 31297 22511 31331
rect 22661 31297 22695 31331
rect 23673 31297 23707 31331
rect 24225 31297 24259 31331
rect 24409 31297 24443 31331
rect 24685 31297 24719 31331
rect 24869 31297 24903 31331
rect 25881 31297 25915 31331
rect 27537 31297 27571 31331
rect 27721 31297 27755 31331
rect 27813 31297 27847 31331
rect 28181 31297 28215 31331
rect 29009 31297 29043 31331
rect 29193 31297 29227 31331
rect 31953 31297 31987 31331
rect 32505 31297 32539 31331
rect 32689 31297 32723 31331
rect 32873 31297 32907 31331
rect 33701 31297 33735 31331
rect 33977 31297 34011 31331
rect 34253 31297 34287 31331
rect 5089 31229 5123 31263
rect 5181 31229 5215 31263
rect 9413 31229 9447 31263
rect 10241 31229 10275 31263
rect 14013 31229 14047 31263
rect 15485 31229 15519 31263
rect 18521 31229 18555 31263
rect 19165 31229 19199 31263
rect 21097 31229 21131 31263
rect 21925 31229 21959 31263
rect 22385 31229 22419 31263
rect 23489 31229 23523 31263
rect 25697 31229 25731 31263
rect 28457 31229 28491 31263
rect 29561 31229 29595 31263
rect 29837 31229 29871 31263
rect 9321 31161 9355 31195
rect 9689 31161 9723 31195
rect 10701 31161 10735 31195
rect 11805 31161 11839 31195
rect 34069 31161 34103 31195
rect 5641 31093 5675 31127
rect 9045 31093 9079 31127
rect 13645 31093 13679 31127
rect 16681 31093 16715 31127
rect 19901 31093 19935 31127
rect 21005 31093 21039 31127
rect 26065 31093 26099 31127
rect 27077 31093 27111 31127
rect 29377 31093 29411 31127
rect 31309 31093 31343 31127
rect 9413 30889 9447 30923
rect 14565 30889 14599 30923
rect 16865 30889 16899 30923
rect 17417 30889 17451 30923
rect 17785 30889 17819 30923
rect 21005 30889 21039 30923
rect 21189 30889 21223 30923
rect 22845 30889 22879 30923
rect 25145 30889 25179 30923
rect 29653 30889 29687 30923
rect 9597 30821 9631 30855
rect 9965 30821 9999 30855
rect 23489 30821 23523 30855
rect 27997 30821 28031 30855
rect 29377 30821 29411 30855
rect 29745 30821 29779 30855
rect 6929 30753 6963 30787
rect 16773 30753 16807 30787
rect 25053 30753 25087 30787
rect 25605 30753 25639 30787
rect 25973 30753 26007 30787
rect 28825 30753 28859 30787
rect 29561 30753 29595 30787
rect 30757 30753 30791 30787
rect 32597 30753 32631 30787
rect 5181 30685 5215 30719
rect 7205 30685 7239 30719
rect 8585 30685 8619 30719
rect 8953 30685 8987 30719
rect 9045 30685 9079 30719
rect 9229 30685 9263 30719
rect 9597 30685 9631 30719
rect 9781 30685 9815 30719
rect 9873 30685 9907 30719
rect 10057 30675 10091 30709
rect 11161 30685 11195 30719
rect 14197 30685 14231 30719
rect 14381 30685 14415 30719
rect 17236 30685 17270 30719
rect 17693 30685 17727 30719
rect 20637 30685 20671 30719
rect 21097 30685 21131 30719
rect 21281 30685 21315 30719
rect 23121 30685 23155 30719
rect 23305 30685 23339 30719
rect 23581 30685 23615 30719
rect 24685 30685 24719 30719
rect 24869 30685 24903 30719
rect 25237 30685 25271 30719
rect 25329 30685 25363 30719
rect 27721 30685 27755 30719
rect 28733 30685 28767 30719
rect 29252 30685 29286 30719
rect 29837 30685 29871 30719
rect 30941 30685 30975 30719
rect 7665 30617 7699 30651
rect 7849 30617 7883 30651
rect 20821 30617 20855 30651
rect 24593 30617 24627 30651
rect 28181 30617 28215 30651
rect 29929 30617 29963 30651
rect 32873 30617 32907 30651
rect 7389 30549 7423 30583
rect 11253 30549 11287 30583
rect 17233 30549 17267 30583
rect 23213 30549 23247 30583
rect 27399 30549 27433 30583
rect 29193 30549 29227 30583
rect 31125 30549 31159 30583
rect 34345 30549 34379 30583
rect 9137 30345 9171 30379
rect 31033 30345 31067 30379
rect 32689 30345 32723 30379
rect 3709 30277 3743 30311
rect 5457 30277 5491 30311
rect 17969 30277 18003 30311
rect 18889 30277 18923 30311
rect 26525 30277 26559 30311
rect 26709 30277 26743 30311
rect 27997 30277 28031 30311
rect 28181 30277 28215 30311
rect 30757 30277 30791 30311
rect 31125 30277 31159 30311
rect 33149 30277 33183 30311
rect 33793 30277 33827 30311
rect 36185 30277 36219 30311
rect 5733 30209 5767 30243
rect 6377 30209 6411 30243
rect 8217 30209 8251 30243
rect 8401 30209 8435 30243
rect 8585 30209 8619 30243
rect 8769 30209 8803 30243
rect 9045 30209 9079 30243
rect 9229 30209 9263 30243
rect 9781 30209 9815 30243
rect 9965 30209 9999 30243
rect 17877 30209 17911 30243
rect 18245 30209 18279 30243
rect 18613 30209 18647 30243
rect 22937 30209 22971 30243
rect 23029 30209 23063 30243
rect 23305 30209 23339 30243
rect 23673 30209 23707 30243
rect 23857 30209 23891 30243
rect 27353 30209 27387 30243
rect 27537 30209 27571 30243
rect 27813 30209 27847 30243
rect 30297 30209 30331 30243
rect 30389 30209 30423 30243
rect 30482 30209 30516 30243
rect 30665 30209 30699 30243
rect 30895 30209 30929 30243
rect 31309 30209 31343 30243
rect 31493 30209 31527 30243
rect 31585 30209 31619 30243
rect 31769 30209 31803 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 32413 30209 32447 30243
rect 32505 30209 32539 30243
rect 32781 30209 32815 30243
rect 32965 30209 32999 30243
rect 33241 30209 33275 30243
rect 33425 30209 33459 30243
rect 33517 30209 33551 30243
rect 33701 30209 33735 30243
rect 33885 30209 33919 30243
rect 6653 30141 6687 30175
rect 18429 30141 18463 30175
rect 20637 30141 20671 30175
rect 23765 30141 23799 30175
rect 25697 30141 25731 30175
rect 25973 30141 26007 30175
rect 28273 30141 28307 30175
rect 30021 30141 30055 30175
rect 34161 30141 34195 30175
rect 34437 30141 34471 30175
rect 8217 30073 8251 30107
rect 9965 30073 9999 30107
rect 27629 30073 27663 30107
rect 33333 30073 33367 30107
rect 34069 30073 34103 30107
rect 8125 30005 8159 30039
rect 8953 30005 8987 30039
rect 24225 30005 24259 30039
rect 26341 30005 26375 30039
rect 31861 30005 31895 30039
rect 6285 29801 6319 29835
rect 9965 29801 9999 29835
rect 16681 29801 16715 29835
rect 17509 29801 17543 29835
rect 18797 29801 18831 29835
rect 22109 29801 22143 29835
rect 24961 29801 24995 29835
rect 25881 29801 25915 29835
rect 29377 29801 29411 29835
rect 30297 29801 30331 29835
rect 32873 29801 32907 29835
rect 35081 29801 35115 29835
rect 9321 29733 9355 29767
rect 10517 29733 10551 29767
rect 14933 29733 14967 29767
rect 28733 29733 28767 29767
rect 34529 29733 34563 29767
rect 3065 29665 3099 29699
rect 4905 29665 4939 29699
rect 6837 29665 6871 29699
rect 8217 29665 8251 29699
rect 11069 29665 11103 29699
rect 22477 29665 22511 29699
rect 22753 29665 22787 29699
rect 26985 29665 27019 29699
rect 30113 29665 30147 29699
rect 30481 29665 30515 29699
rect 30941 29665 30975 29699
rect 31677 29665 31711 29699
rect 2881 29597 2915 29631
rect 5181 29597 5215 29631
rect 6653 29597 6687 29631
rect 7665 29597 7699 29631
rect 7849 29597 7883 29631
rect 8401 29597 8435 29631
rect 8585 29597 8619 29631
rect 9137 29597 9171 29631
rect 9321 29597 9355 29631
rect 10149 29597 10183 29631
rect 10333 29597 10367 29631
rect 10425 29597 10459 29631
rect 10701 29597 10735 29631
rect 10793 29597 10827 29631
rect 12720 29597 12754 29631
rect 13092 29597 13126 29631
rect 13185 29597 13219 29631
rect 15112 29597 15146 29631
rect 15484 29597 15518 29631
rect 15577 29597 15611 29631
rect 17693 29597 17727 29631
rect 17785 29597 17819 29631
rect 17969 29597 18003 29631
rect 18061 29597 18095 29631
rect 18153 29597 18187 29631
rect 18246 29597 18280 29631
rect 18618 29597 18652 29631
rect 20453 29597 20487 29631
rect 20913 29597 20947 29631
rect 21649 29597 21683 29631
rect 21925 29597 21959 29631
rect 22201 29597 22235 29631
rect 22293 29597 22327 29631
rect 22845 29597 22879 29631
rect 24409 29597 24443 29631
rect 24681 29597 24715 29631
rect 24777 29597 24811 29631
rect 26249 29597 26283 29631
rect 26709 29597 26743 29631
rect 28825 29597 28859 29631
rect 29193 29597 29227 29631
rect 30573 29597 30607 29631
rect 31217 29597 31251 29631
rect 31401 29597 31435 29631
rect 32137 29597 32171 29631
rect 32505 29597 32539 29631
rect 32781 29597 32815 29631
rect 34345 29597 34379 29631
rect 34529 29597 34563 29631
rect 34897 29597 34931 29631
rect 34989 29597 35023 29631
rect 35633 29597 35667 29631
rect 4721 29529 4755 29563
rect 6745 29529 6779 29563
rect 11161 29529 11195 29563
rect 12817 29529 12851 29563
rect 12909 29529 12943 29563
rect 15209 29529 15243 29563
rect 15301 29529 15335 29563
rect 16649 29529 16683 29563
rect 16865 29529 16899 29563
rect 18429 29529 18463 29563
rect 18521 29529 18555 29563
rect 21189 29529 21223 29563
rect 24593 29529 24627 29563
rect 26065 29529 26099 29563
rect 26341 29529 26375 29563
rect 26893 29529 26927 29563
rect 27261 29529 27295 29563
rect 29009 29529 29043 29563
rect 29101 29529 29135 29563
rect 31033 29529 31067 29563
rect 31309 29529 31343 29563
rect 31539 29529 31573 29563
rect 34805 29529 34839 29563
rect 35817 29529 35851 29563
rect 2421 29461 2455 29495
rect 2789 29461 2823 29495
rect 4261 29461 4295 29495
rect 4629 29461 4663 29495
rect 5733 29461 5767 29495
rect 7113 29461 7147 29495
rect 12541 29461 12575 29495
rect 16497 29461 16531 29495
rect 21741 29461 21775 29495
rect 29561 29461 29595 29495
rect 30665 29461 30699 29495
rect 30849 29461 30883 29495
rect 32229 29461 32263 29495
rect 35449 29461 35483 29495
rect 36093 29461 36127 29495
rect 5825 29257 5859 29291
rect 6745 29257 6779 29291
rect 7757 29257 7791 29291
rect 7849 29257 7883 29291
rect 9229 29257 9263 29291
rect 9321 29257 9355 29291
rect 10057 29257 10091 29291
rect 16681 29257 16715 29291
rect 18337 29257 18371 29291
rect 23765 29257 23799 29291
rect 25421 29257 25455 29291
rect 26985 29257 27019 29291
rect 27997 29257 28031 29291
rect 30573 29257 30607 29291
rect 31861 29257 31895 29291
rect 32781 29257 32815 29291
rect 34069 29257 34103 29291
rect 1777 29189 1811 29223
rect 3893 29189 3927 29223
rect 5917 29189 5951 29223
rect 6837 29189 6871 29223
rect 7481 29189 7515 29223
rect 8861 29189 8895 29223
rect 9689 29189 9723 29223
rect 11897 29189 11931 29223
rect 12653 29189 12687 29223
rect 13277 29189 13311 29223
rect 13369 29189 13403 29223
rect 14381 29189 14415 29223
rect 16221 29189 16255 29223
rect 17417 29189 17451 29223
rect 20821 29189 20855 29223
rect 22201 29189 22235 29223
rect 26801 29189 26835 29223
rect 27813 29189 27847 29223
rect 30849 29189 30883 29223
rect 32505 29189 32539 29223
rect 32873 29189 32907 29223
rect 33425 29189 33459 29223
rect 7205 29121 7239 29155
rect 7389 29121 7423 29155
rect 7573 29121 7607 29155
rect 7987 29121 8021 29155
rect 8125 29121 8159 29155
rect 8217 29121 8251 29155
rect 8345 29121 8379 29155
rect 8468 29121 8502 29155
rect 8574 29121 8608 29155
rect 8733 29121 8767 29155
rect 8953 29121 8987 29155
rect 9091 29121 9125 29155
rect 9505 29121 9539 29155
rect 9597 29121 9631 29155
rect 9873 29121 9907 29155
rect 10241 29121 10275 29155
rect 10425 29121 10459 29155
rect 10517 29121 10551 29155
rect 10885 29121 10919 29155
rect 11161 29121 11195 29155
rect 11621 29121 11655 29155
rect 11805 29121 11839 29155
rect 11989 29121 12023 29155
rect 12265 29121 12299 29155
rect 12358 29121 12392 29155
rect 12541 29121 12575 29155
rect 12769 29121 12803 29155
rect 13180 29121 13214 29155
rect 13552 29121 13586 29155
rect 13645 29121 13679 29155
rect 14105 29121 14139 29155
rect 14289 29121 14323 29155
rect 14473 29121 14507 29155
rect 14749 29121 14783 29155
rect 15025 29121 15059 29155
rect 15301 29121 15335 29155
rect 15485 29121 15519 29155
rect 16129 29121 16163 29155
rect 16313 29121 16347 29155
rect 16477 29121 16511 29155
rect 18337 29121 18371 29155
rect 19809 29121 19843 29155
rect 19901 29121 19935 29155
rect 19993 29121 20027 29155
rect 20085 29121 20119 29155
rect 20545 29121 20579 29155
rect 20637 29121 20671 29155
rect 20913 29121 20947 29155
rect 21097 29121 21131 29155
rect 21189 29121 21223 29155
rect 21373 29121 21407 29155
rect 21465 29121 21499 29155
rect 22063 29121 22097 29155
rect 22293 29121 22327 29155
rect 22448 29121 22482 29155
rect 22569 29121 22603 29155
rect 22845 29121 22879 29155
rect 23029 29121 23063 29155
rect 23397 29121 23431 29155
rect 23949 29121 23983 29155
rect 24041 29121 24075 29155
rect 24501 29121 24535 29155
rect 24593 29121 24627 29155
rect 24777 29121 24811 29155
rect 24869 29121 24903 29155
rect 25329 29121 25363 29155
rect 26157 29121 26191 29155
rect 26341 29121 26375 29155
rect 26433 29121 26467 29155
rect 26525 29121 26559 29155
rect 27164 29121 27198 29155
rect 27261 29121 27295 29155
rect 27353 29121 27387 29155
rect 27536 29121 27570 29155
rect 27629 29121 27663 29155
rect 27721 29121 27755 29155
rect 28181 29121 28215 29155
rect 28273 29121 28307 29155
rect 28365 29121 28399 29155
rect 28483 29121 28517 29155
rect 28641 29121 28675 29155
rect 28917 29121 28951 29155
rect 29469 29121 29503 29155
rect 29653 29121 29687 29155
rect 30021 29121 30055 29155
rect 30113 29121 30147 29155
rect 30297 29121 30331 29155
rect 30389 29121 30423 29155
rect 30481 29121 30515 29155
rect 30757 29121 30791 29155
rect 30941 29121 30975 29155
rect 31855 29121 31889 29155
rect 32295 29121 32329 29155
rect 32413 29121 32447 29155
rect 32597 29121 32631 29155
rect 32965 29121 32999 29155
rect 33149 29121 33183 29155
rect 33793 29121 33827 29155
rect 33885 29121 33919 29155
rect 1501 29053 1535 29087
rect 3617 29053 3651 29087
rect 6101 29053 6135 29087
rect 6929 29053 6963 29087
rect 10793 29053 10827 29087
rect 11253 29053 11287 29087
rect 15117 29053 15151 29087
rect 16865 29053 16899 29087
rect 16957 29053 16991 29087
rect 18613 29053 18647 29087
rect 22661 29053 22695 29087
rect 23489 29053 23523 29087
rect 24225 29053 24259 29087
rect 24317 29053 24351 29087
rect 29377 29053 29411 29087
rect 31585 29053 31619 29087
rect 32137 29053 32171 29087
rect 34161 29053 34195 29087
rect 34437 29053 34471 29087
rect 36185 29053 36219 29087
rect 3249 28985 3283 29019
rect 5457 28985 5491 29019
rect 10609 28985 10643 29019
rect 12909 28985 12943 29019
rect 14657 28985 14691 29019
rect 15209 28985 15243 29019
rect 17417 28985 17451 29019
rect 18153 28985 18187 29019
rect 18429 28985 18463 29019
rect 20269 28985 20303 29019
rect 20361 28985 20395 29019
rect 21925 28985 21959 29019
rect 24133 28985 24167 29019
rect 31769 28985 31803 29019
rect 5365 28917 5399 28951
rect 6377 28917 6411 28951
rect 12173 28917 12207 28951
rect 13001 28917 13035 28951
rect 15945 28917 15979 28951
rect 20821 28917 20855 28951
rect 23489 28917 23523 28951
rect 29193 28917 29227 28951
rect 29837 28917 29871 28951
rect 33517 28917 33551 28951
rect 3801 28713 3835 28747
rect 7573 28713 7607 28747
rect 8309 28713 8343 28747
rect 16773 28713 16807 28747
rect 17233 28713 17267 28747
rect 18245 28713 18279 28747
rect 20453 28713 20487 28747
rect 24961 28713 24995 28747
rect 27353 28713 27387 28747
rect 28181 28713 28215 28747
rect 28825 28713 28859 28747
rect 34805 28713 34839 28747
rect 9413 28645 9447 28679
rect 10241 28645 10275 28679
rect 10977 28645 11011 28679
rect 12541 28645 12575 28679
rect 20913 28645 20947 28679
rect 25329 28645 25363 28679
rect 26893 28645 26927 28679
rect 32781 28645 32815 28679
rect 33609 28645 33643 28679
rect 5273 28577 5307 28611
rect 5549 28577 5583 28611
rect 5825 28577 5859 28611
rect 6101 28577 6135 28611
rect 10701 28577 10735 28611
rect 11161 28577 11195 28611
rect 11621 28577 11655 28611
rect 12173 28577 12207 28611
rect 25237 28577 25271 28611
rect 25421 28577 25455 28611
rect 26433 28577 26467 28611
rect 34069 28577 34103 28611
rect 35173 28577 35207 28611
rect 35817 28577 35851 28611
rect 1409 28509 1443 28543
rect 7665 28509 7699 28543
rect 7758 28509 7792 28543
rect 8033 28509 8067 28543
rect 8130 28509 8164 28543
rect 11253 28509 11287 28543
rect 12081 28509 12115 28543
rect 12265 28509 12299 28543
rect 12357 28509 12391 28543
rect 12720 28509 12754 28543
rect 13092 28509 13126 28543
rect 13185 28509 13219 28543
rect 17693 28509 17727 28543
rect 17969 28509 18003 28543
rect 18061 28509 18095 28543
rect 19533 28509 19567 28543
rect 19717 28509 19751 28543
rect 20637 28509 20671 28543
rect 20821 28509 20855 28543
rect 21092 28509 21126 28543
rect 21464 28509 21498 28543
rect 21557 28509 21591 28543
rect 22196 28509 22230 28543
rect 22385 28509 22419 28543
rect 22568 28509 22602 28543
rect 22661 28509 22695 28543
rect 23305 28509 23339 28543
rect 23581 28509 23615 28543
rect 25697 28509 25731 28543
rect 26157 28509 26191 28543
rect 26249 28509 26283 28543
rect 26709 28509 26743 28543
rect 26801 28509 26835 28543
rect 26985 28509 27019 28543
rect 27721 28509 27755 28543
rect 27997 28509 28031 28543
rect 29101 28509 29135 28543
rect 31953 28509 31987 28543
rect 32137 28509 32171 28543
rect 32229 28509 32263 28543
rect 32505 28509 32539 28543
rect 32689 28509 32723 28543
rect 32873 28509 32907 28543
rect 33241 28509 33275 28543
rect 33425 28509 33459 28543
rect 33517 28509 33551 28543
rect 33793 28509 33827 28543
rect 34253 28509 34287 28543
rect 34989 28509 35023 28543
rect 35081 28509 35115 28543
rect 35265 28509 35299 28543
rect 1685 28441 1719 28475
rect 7941 28441 7975 28475
rect 9689 28441 9723 28475
rect 9965 28441 9999 28475
rect 10793 28441 10827 28475
rect 11529 28441 11563 28475
rect 12817 28441 12851 28475
rect 12909 28441 12943 28475
rect 16741 28441 16775 28475
rect 16957 28441 16991 28475
rect 17049 28441 17083 28475
rect 17877 28441 17911 28475
rect 21189 28441 21223 28475
rect 21281 28441 21315 28475
rect 22293 28441 22327 28475
rect 27261 28441 27295 28475
rect 28457 28441 28491 28475
rect 35541 28441 35575 28475
rect 3157 28373 3191 28407
rect 9873 28373 9907 28407
rect 10701 28373 10735 28407
rect 11897 28373 11931 28407
rect 16589 28373 16623 28407
rect 17249 28373 17283 28407
rect 17417 28373 17451 28407
rect 19349 28373 19383 28407
rect 22017 28373 22051 28407
rect 23121 28373 23155 28407
rect 23489 28373 23523 28407
rect 25605 28373 25639 28407
rect 25789 28373 25823 28407
rect 26525 28373 26559 28407
rect 27813 28373 27847 28407
rect 28834 28373 28868 28407
rect 32045 28373 32079 28407
rect 32505 28373 32539 28407
rect 33333 28373 33367 28407
rect 34437 28373 34471 28407
rect 2421 28169 2455 28203
rect 5089 28169 5123 28203
rect 8493 28169 8527 28203
rect 10241 28169 10275 28203
rect 16681 28169 16715 28203
rect 17785 28169 17819 28203
rect 19073 28169 19107 28203
rect 29101 28169 29135 28203
rect 29729 28169 29763 28203
rect 30757 28169 30791 28203
rect 32505 28169 32539 28203
rect 33523 28169 33557 28203
rect 3985 28101 4019 28135
rect 4077 28101 4111 28135
rect 4721 28101 4755 28135
rect 10793 28101 10827 28135
rect 10885 28101 10919 28135
rect 16957 28101 16991 28135
rect 29929 28101 29963 28135
rect 30665 28101 30699 28135
rect 33307 28101 33341 28135
rect 33422 28101 33456 28135
rect 33103 28067 33137 28101
rect 2789 28033 2823 28067
rect 2881 28033 2915 28067
rect 3801 28033 3835 28067
rect 4169 28033 4203 28067
rect 4445 28033 4479 28067
rect 4629 28033 4663 28067
rect 4813 28033 4847 28067
rect 5641 28033 5675 28067
rect 6745 28033 6779 28067
rect 7113 28033 7147 28067
rect 7297 28033 7331 28067
rect 7573 28033 7607 28067
rect 8401 28033 8435 28067
rect 8585 28033 8619 28067
rect 10517 28033 10551 28067
rect 12633 28033 12667 28067
rect 16819 28033 16853 28067
rect 17049 28033 17083 28067
rect 17232 28033 17266 28067
rect 17325 28033 17359 28067
rect 17693 28033 17727 28067
rect 17877 28033 17911 28067
rect 18153 28033 18187 28067
rect 18337 28033 18371 28067
rect 18429 28033 18463 28067
rect 18613 28033 18647 28067
rect 18889 28033 18923 28067
rect 19533 28033 19567 28067
rect 21005 28033 21039 28067
rect 21097 28033 21131 28067
rect 23673 28033 23707 28067
rect 24225 28033 24259 28067
rect 24409 28033 24443 28067
rect 26065 28033 26099 28067
rect 28089 28033 28123 28067
rect 28457 28033 28491 28067
rect 28917 28033 28951 28067
rect 29101 28033 29135 28067
rect 30205 28033 30239 28067
rect 30297 28033 30331 28067
rect 31493 28033 31527 28067
rect 31769 28033 31803 28067
rect 31953 28033 31987 28067
rect 32413 28033 32447 28067
rect 32597 28033 32631 28067
rect 33609 28033 33643 28067
rect 33701 28033 33735 28067
rect 34621 28033 34655 28067
rect 34989 28033 35023 28067
rect 35081 28033 35115 28067
rect 35265 28033 35299 28067
rect 36185 28033 36219 28067
rect 3065 27965 3099 27999
rect 10425 27965 10459 27999
rect 12909 27965 12943 27999
rect 17969 27965 18003 27999
rect 18705 27965 18739 27999
rect 19625 27965 19659 27999
rect 20821 27965 20855 27999
rect 23489 27965 23523 27999
rect 24685 27965 24719 27999
rect 26341 27965 26375 27999
rect 27445 27965 27479 27999
rect 28365 27965 28399 27999
rect 28825 27965 28859 27999
rect 30573 27965 30607 27999
rect 30941 27965 30975 27999
rect 31033 27965 31067 27999
rect 32873 27965 32907 27999
rect 7389 27897 7423 27931
rect 19901 27897 19935 27931
rect 24501 27897 24535 27931
rect 31953 27897 31987 27931
rect 36001 27897 36035 27931
rect 4353 27829 4387 27863
rect 4997 27829 5031 27863
rect 12449 27829 12483 27863
rect 12817 27829 12851 27863
rect 19533 27829 19567 27863
rect 24041 27829 24075 27863
rect 24593 27829 24627 27863
rect 25881 27829 25915 27863
rect 26249 27829 26283 27863
rect 28181 27829 28215 27863
rect 29561 27829 29595 27863
rect 29745 27829 29779 27863
rect 30021 27829 30055 27863
rect 31217 27829 31251 27863
rect 31401 27829 31435 27863
rect 32137 27829 32171 27863
rect 32781 27829 32815 27863
rect 32965 27829 32999 27863
rect 33149 27829 33183 27863
rect 34437 27829 34471 27863
rect 34897 27829 34931 27863
rect 35173 27829 35207 27863
rect 8953 27625 8987 27659
rect 13185 27625 13219 27659
rect 16221 27625 16255 27659
rect 24869 27625 24903 27659
rect 25237 27625 25271 27659
rect 26893 27625 26927 27659
rect 28377 27625 28411 27659
rect 29193 27625 29227 27659
rect 30205 27625 30239 27659
rect 34989 27625 35023 27659
rect 36001 27625 36035 27659
rect 9965 27557 9999 27591
rect 10517 27557 10551 27591
rect 15393 27557 15427 27591
rect 16497 27557 16531 27591
rect 24133 27557 24167 27591
rect 3157 27489 3191 27523
rect 7021 27489 7055 27523
rect 8677 27489 8711 27523
rect 11161 27489 11195 27523
rect 23305 27489 23339 27523
rect 24501 27489 24535 27523
rect 28641 27489 28675 27523
rect 30113 27489 30147 27523
rect 34253 27489 34287 27523
rect 34345 27489 34379 27523
rect 34529 27489 34563 27523
rect 1409 27421 1443 27455
rect 4629 27421 4663 27455
rect 4997 27421 5031 27455
rect 7757 27421 7791 27455
rect 8033 27421 8067 27455
rect 8217 27421 8251 27455
rect 8493 27421 8527 27455
rect 9091 27421 9125 27455
rect 9504 27421 9538 27455
rect 9597 27421 9631 27455
rect 10149 27421 10183 27455
rect 10425 27421 10459 27455
rect 10701 27421 10735 27455
rect 10793 27421 10827 27455
rect 11069 27421 11103 27455
rect 12357 27421 12391 27455
rect 12541 27421 12575 27455
rect 12725 27421 12759 27455
rect 12817 27421 12851 27455
rect 12909 27421 12943 27455
rect 13093 27421 13127 27455
rect 13323 27421 13357 27455
rect 13681 27421 13715 27455
rect 13829 27421 13863 27455
rect 14841 27421 14875 27455
rect 15209 27421 15243 27455
rect 16676 27421 16710 27455
rect 16773 27421 16807 27455
rect 16865 27421 16899 27455
rect 16993 27421 17027 27455
rect 17141 27421 17175 27455
rect 17417 27421 17451 27455
rect 17509 27421 17543 27455
rect 17693 27421 17727 27455
rect 17785 27421 17819 27455
rect 17877 27421 17911 27455
rect 18153 27421 18187 27455
rect 19349 27421 19383 27455
rect 19441 27421 19475 27455
rect 19533 27421 19567 27455
rect 19809 27421 19843 27455
rect 19901 27421 19935 27455
rect 20085 27421 20119 27455
rect 21097 27421 21131 27455
rect 21373 27421 21407 27455
rect 21833 27421 21867 27455
rect 23029 27421 23063 27455
rect 23121 27421 23155 27455
rect 24409 27421 24443 27455
rect 24593 27421 24627 27455
rect 24685 27421 24719 27455
rect 25053 27421 25087 27455
rect 25329 27421 25363 27455
rect 25513 27421 25547 27455
rect 29837 27421 29871 27455
rect 30389 27421 30423 27455
rect 30481 27421 30515 27455
rect 30665 27421 30699 27455
rect 30757 27421 30791 27455
rect 31033 27421 31067 27455
rect 31217 27421 31251 27455
rect 31861 27421 31895 27455
rect 31973 27421 32007 27455
rect 34069 27421 34103 27455
rect 34161 27421 34195 27455
rect 34713 27421 34747 27455
rect 35173 27421 35207 27455
rect 35265 27421 35299 27455
rect 35449 27421 35483 27455
rect 35541 27421 35575 27455
rect 36185 27421 36219 27455
rect 29239 27387 29273 27421
rect 1685 27353 1719 27387
rect 3801 27353 3835 27387
rect 4813 27353 4847 27387
rect 4905 27353 4939 27387
rect 6745 27353 6779 27387
rect 9229 27353 9263 27387
rect 9321 27353 9355 27387
rect 13461 27353 13495 27387
rect 13553 27353 13587 27387
rect 15025 27353 15059 27387
rect 15117 27353 15151 27387
rect 16037 27353 16071 27387
rect 18245 27353 18279 27387
rect 18521 27353 18555 27387
rect 18705 27353 18739 27387
rect 19717 27353 19751 27387
rect 21649 27353 21683 27387
rect 24133 27353 24167 27387
rect 25881 27353 25915 27387
rect 26065 27353 26099 27387
rect 29009 27353 29043 27387
rect 29745 27353 29779 27387
rect 29929 27353 29963 27387
rect 31677 27353 31711 27387
rect 32229 27353 32263 27387
rect 5181 27285 5215 27319
rect 5273 27285 5307 27319
rect 7113 27285 7147 27319
rect 10333 27285 10367 27319
rect 16237 27285 16271 27319
rect 16405 27285 16439 27319
rect 17233 27285 17267 27319
rect 18889 27285 18923 27319
rect 20269 27285 20303 27319
rect 20913 27285 20947 27319
rect 21281 27285 21315 27319
rect 21465 27285 21499 27319
rect 23305 27285 23339 27319
rect 23397 27285 23431 27319
rect 23581 27285 23615 27319
rect 23673 27285 23707 27319
rect 25697 27285 25731 27319
rect 26249 27285 26283 27319
rect 29377 27285 29411 27319
rect 29561 27285 29595 27319
rect 30941 27285 30975 27319
rect 32045 27285 32079 27319
rect 34805 27285 34839 27319
rect 2237 27081 2271 27115
rect 2697 27081 2731 27115
rect 6377 27081 6411 27115
rect 6745 27081 6779 27115
rect 7573 27081 7607 27115
rect 12449 27081 12483 27115
rect 21991 27081 22025 27115
rect 24041 27081 24075 27115
rect 24225 27081 24259 27115
rect 25973 27081 26007 27115
rect 28457 27081 28491 27115
rect 31493 27081 31527 27115
rect 2605 27013 2639 27047
rect 8401 27013 8435 27047
rect 8493 27013 8527 27047
rect 10425 27013 10459 27047
rect 11253 27013 11287 27047
rect 11345 27013 11379 27047
rect 13829 27013 13863 27047
rect 17969 27013 18003 27047
rect 22201 27013 22235 27047
rect 23673 27013 23707 27047
rect 24593 27013 24627 27047
rect 26433 27013 26467 27047
rect 30389 27013 30423 27047
rect 30573 27013 30607 27047
rect 31125 27013 31159 27047
rect 31341 27013 31375 27047
rect 32933 27013 32967 27047
rect 33149 27013 33183 27047
rect 33425 27013 33459 27047
rect 34621 27013 34655 27047
rect 35265 27013 35299 27047
rect 36001 27013 36035 27047
rect 3249 26945 3283 26979
rect 5825 26945 5859 26979
rect 7481 26945 7515 26979
rect 7849 26945 7883 26979
rect 8263 26945 8297 26979
rect 8676 26945 8710 26979
rect 8769 26945 8803 26979
rect 10517 26945 10551 26979
rect 10885 26945 10919 26979
rect 10977 26945 11011 26979
rect 12265 26945 12299 26979
rect 12541 26945 12575 26979
rect 12817 26945 12851 26979
rect 13001 26945 13035 26979
rect 13185 26945 13219 26979
rect 13369 26945 13403 26979
rect 13461 26945 13495 26979
rect 13554 26945 13588 26979
rect 13737 26945 13771 26979
rect 13926 26945 13960 26979
rect 18245 26945 18279 26979
rect 19717 26945 19751 26979
rect 20269 26945 20303 26979
rect 20453 26945 20487 26979
rect 20913 26945 20947 26979
rect 21373 26945 21407 26979
rect 22293 26945 22327 26979
rect 23857 26945 23891 26979
rect 24409 26945 24443 26979
rect 24685 26945 24719 26979
rect 25053 26945 25087 26979
rect 26801 26945 26835 26979
rect 28365 26945 28399 26979
rect 28549 26945 28583 26979
rect 29929 26945 29963 26979
rect 30803 26945 30837 26979
rect 31033 26945 31067 26979
rect 33241 26945 33275 26979
rect 33701 26945 33735 26979
rect 33885 26945 33919 26979
rect 34345 26945 34379 26979
rect 34437 26945 34471 26979
rect 34805 26945 34839 26979
rect 34897 26945 34931 26979
rect 35541 26945 35575 26979
rect 35725 26945 35759 26979
rect 35909 26945 35943 26979
rect 2881 26877 2915 26911
rect 3525 26877 3559 26911
rect 4997 26877 5031 26911
rect 6837 26877 6871 26911
rect 7021 26877 7055 26911
rect 8033 26877 8067 26911
rect 10425 26877 10459 26911
rect 13093 26877 13127 26911
rect 22385 26877 22419 26911
rect 22569 26877 22603 26911
rect 24777 26877 24811 26911
rect 26985 26877 27019 26911
rect 27261 26877 27295 26911
rect 29745 26877 29779 26911
rect 10701 26809 10735 26843
rect 12173 26809 12207 26843
rect 18153 26809 18187 26843
rect 20085 26809 20119 26843
rect 26065 26809 26099 26843
rect 26617 26809 26651 26843
rect 30205 26809 30239 26843
rect 30757 26809 30791 26843
rect 33609 26809 33643 26843
rect 34161 26809 34195 26843
rect 35817 26809 35851 26843
rect 5181 26741 5215 26775
rect 8125 26741 8159 26775
rect 9965 26741 9999 26775
rect 12633 26741 12667 26775
rect 14105 26741 14139 26775
rect 18061 26741 18095 26775
rect 21833 26741 21867 26775
rect 22017 26741 22051 26775
rect 22293 26741 22327 26775
rect 30113 26741 30147 26775
rect 31309 26741 31343 26775
rect 32781 26741 32815 26775
rect 32965 26741 32999 26775
rect 33701 26741 33735 26775
rect 35265 26741 35299 26775
rect 35449 26741 35483 26775
rect 4813 26537 4847 26571
rect 8033 26537 8067 26571
rect 8953 26537 8987 26571
rect 9689 26537 9723 26571
rect 17785 26537 17819 26571
rect 21097 26537 21131 26571
rect 21925 26537 21959 26571
rect 26249 26537 26283 26571
rect 26709 26537 26743 26571
rect 26985 26537 27019 26571
rect 30205 26537 30239 26571
rect 32597 26537 32631 26571
rect 33701 26537 33735 26571
rect 35081 26537 35115 26571
rect 5641 26469 5675 26503
rect 13369 26469 13403 26503
rect 14841 26469 14875 26503
rect 15301 26469 15335 26503
rect 21281 26469 21315 26503
rect 33793 26469 33827 26503
rect 36001 26469 36035 26503
rect 3893 26401 3927 26435
rect 5365 26401 5399 26435
rect 14933 26401 14967 26435
rect 21373 26401 21407 26435
rect 21741 26401 21775 26435
rect 26341 26401 26375 26435
rect 35541 26401 35575 26435
rect 4721 26333 4755 26367
rect 5825 26333 5859 26367
rect 5917 26333 5951 26367
rect 6193 26333 6227 26367
rect 6929 26333 6963 26367
rect 7941 26333 7975 26367
rect 8171 26333 8205 26367
rect 8401 26333 8435 26367
rect 8584 26333 8618 26367
rect 8677 26333 8711 26367
rect 9137 26333 9171 26367
rect 9505 26333 9539 26367
rect 9873 26333 9907 26367
rect 10149 26333 10183 26367
rect 12541 26333 12575 26367
rect 12725 26333 12759 26367
rect 12817 26333 12851 26367
rect 12909 26333 12943 26367
rect 13093 26333 13127 26367
rect 13553 26333 13587 26367
rect 13645 26333 13679 26367
rect 13921 26333 13955 26367
rect 14197 26333 14231 26367
rect 14345 26333 14379 26367
rect 14473 26333 14507 26367
rect 14662 26333 14696 26367
rect 15117 26333 15151 26367
rect 15393 26333 15427 26367
rect 16773 26333 16807 26367
rect 17049 26333 17083 26367
rect 17233 26333 17267 26367
rect 17412 26333 17446 26367
rect 17509 26333 17543 26367
rect 22385 26333 22419 26367
rect 22477 26333 22511 26367
rect 22661 26333 22695 26367
rect 22753 26333 22787 26367
rect 25881 26333 25915 26367
rect 26525 26333 26559 26367
rect 27445 26333 27479 26367
rect 27813 26333 27847 26367
rect 27905 26333 27939 26367
rect 28181 26333 28215 26367
rect 28365 26333 28399 26367
rect 30573 26333 30607 26367
rect 30849 26333 30883 26367
rect 32781 26333 32815 26367
rect 32873 26333 32907 26367
rect 32965 26333 32999 26367
rect 33241 26333 33275 26367
rect 33333 26333 33367 26367
rect 33609 26333 33643 26367
rect 33885 26333 33919 26367
rect 34069 26333 34103 26367
rect 34713 26333 34747 26367
rect 34897 26333 34931 26367
rect 35265 26333 35299 26367
rect 35449 26333 35483 26367
rect 36185 26333 36219 26367
rect 5181 26265 5215 26299
rect 6009 26265 6043 26299
rect 6745 26265 6779 26299
rect 8309 26265 8343 26299
rect 9229 26265 9263 26299
rect 9321 26265 9355 26299
rect 12357 26265 12391 26299
rect 13737 26265 13771 26299
rect 14565 26265 14599 26299
rect 17601 26265 17635 26299
rect 17785 26265 17819 26299
rect 20913 26265 20947 26299
rect 21113 26265 21147 26299
rect 22201 26265 22235 26299
rect 26065 26265 26099 26299
rect 26893 26265 26927 26299
rect 28273 26265 28307 26299
rect 30389 26265 30423 26299
rect 33083 26265 33117 26299
rect 34805 26265 34839 26299
rect 5273 26197 5307 26231
rect 7297 26197 7331 26231
rect 10057 26197 10091 26231
rect 16589 26197 16623 26231
rect 21557 26197 21591 26231
rect 27261 26197 27295 26231
rect 27997 26197 28031 26231
rect 30757 26197 30791 26231
rect 3157 25993 3191 26027
rect 4997 25993 5031 26027
rect 8217 25993 8251 26027
rect 9781 25993 9815 26027
rect 18889 25993 18923 26027
rect 19625 25993 19659 26027
rect 23413 25993 23447 26027
rect 23581 25993 23615 26027
rect 24961 25993 24995 26027
rect 32689 25993 32723 26027
rect 33517 25993 33551 26027
rect 6009 25925 6043 25959
rect 9873 25925 9907 25959
rect 10701 25925 10735 25959
rect 10793 25925 10827 25959
rect 12817 25925 12851 25959
rect 18236 25925 18270 25959
rect 23213 25925 23247 25959
rect 24133 25925 24167 25959
rect 24225 25925 24259 25959
rect 29009 25925 29043 25959
rect 30113 25925 30147 25959
rect 30297 25925 30331 25959
rect 31585 25925 31619 25959
rect 32229 25925 32263 25959
rect 33977 25925 34011 25959
rect 8401 25857 8435 25891
rect 8493 25857 8527 25891
rect 8585 25857 8619 25891
rect 8769 25857 8803 25891
rect 10333 25857 10367 25891
rect 10609 25857 10643 25891
rect 10977 25857 11011 25891
rect 11529 25857 11563 25891
rect 11713 25857 11747 25891
rect 12081 25857 12115 25891
rect 12265 25857 12299 25891
rect 12449 25857 12483 25891
rect 12542 25857 12576 25891
rect 12725 25857 12759 25891
rect 12955 25857 12989 25891
rect 15761 25857 15795 25891
rect 15945 25857 15979 25891
rect 16221 25857 16255 25891
rect 16313 25857 16347 25891
rect 17141 25857 17175 25891
rect 17509 25857 17543 25891
rect 17693 25857 17727 25891
rect 17969 25857 18003 25891
rect 18613 25857 18647 25891
rect 18705 25857 18739 25891
rect 18981 25857 19015 25891
rect 19625 25857 19659 25891
rect 23857 25857 23891 25891
rect 24005 25857 24039 25891
rect 24322 25857 24356 25891
rect 24777 25857 24811 25891
rect 25053 25857 25087 25891
rect 25605 25857 25639 25891
rect 25789 25857 25823 25891
rect 26157 25857 26191 25891
rect 26249 25857 26283 25891
rect 26341 25857 26375 25891
rect 26525 25857 26559 25891
rect 27169 25857 27203 25891
rect 27261 25857 27295 25891
rect 27445 25857 27479 25891
rect 27537 25857 27571 25891
rect 28779 25857 28813 25891
rect 28917 25857 28951 25891
rect 29101 25857 29135 25891
rect 29561 25857 29595 25891
rect 29745 25857 29779 25891
rect 31769 25857 31803 25891
rect 31953 25857 31987 25891
rect 32413 25857 32447 25891
rect 32873 25857 32907 25891
rect 33149 25857 33183 25891
rect 33333 25857 33367 25891
rect 33701 25857 33735 25891
rect 34437 25857 34471 25891
rect 34529 25857 34563 25891
rect 34713 25857 34747 25891
rect 35173 25857 35207 25891
rect 35449 25857 35483 25891
rect 1409 25789 1443 25823
rect 1685 25789 1719 25823
rect 3249 25789 3283 25823
rect 3525 25789 3559 25823
rect 5181 25789 5215 25823
rect 6377 25789 6411 25823
rect 6653 25789 6687 25823
rect 9781 25789 9815 25823
rect 10241 25789 10275 25823
rect 11161 25789 11195 25823
rect 11805 25789 11839 25823
rect 11897 25789 11931 25823
rect 16037 25789 16071 25823
rect 16681 25789 16715 25823
rect 17049 25789 17083 25823
rect 19441 25789 19475 25823
rect 19993 25789 20027 25823
rect 28641 25789 28675 25823
rect 31861 25789 31895 25823
rect 33057 25789 33091 25823
rect 33793 25789 33827 25823
rect 34345 25789 34379 25823
rect 10057 25721 10091 25755
rect 16313 25721 16347 25755
rect 16773 25721 16807 25755
rect 24501 25721 24535 25755
rect 25881 25721 25915 25755
rect 29469 25721 29503 25755
rect 8125 25653 8159 25687
rect 9321 25653 9355 25687
rect 13093 25653 13127 25687
rect 15577 25653 15611 25687
rect 18245 25653 18279 25687
rect 18705 25653 18739 25687
rect 23397 25653 23431 25687
rect 24593 25653 24627 25687
rect 26985 25653 27019 25687
rect 29285 25653 29319 25687
rect 29929 25653 29963 25687
rect 30113 25653 30147 25687
rect 31493 25653 31527 25687
rect 33333 25653 33367 25687
rect 33977 25653 34011 25687
rect 34069 25653 34103 25687
rect 34253 25653 34287 25687
rect 34529 25653 34563 25687
rect 35357 25653 35391 25687
rect 2237 25449 2271 25483
rect 3893 25449 3927 25483
rect 6837 25449 6871 25483
rect 9781 25449 9815 25483
rect 11253 25449 11287 25483
rect 17233 25449 17267 25483
rect 19625 25449 19659 25483
rect 23489 25449 23523 25483
rect 24225 25449 24259 25483
rect 29745 25449 29779 25483
rect 30941 25449 30975 25483
rect 35081 25449 35115 25483
rect 35541 25449 35575 25483
rect 8493 25381 8527 25415
rect 8953 25381 8987 25415
rect 14105 25381 14139 25415
rect 17417 25381 17451 25415
rect 20821 25381 20855 25415
rect 25789 25381 25823 25415
rect 32321 25381 32355 25415
rect 33885 25381 33919 25415
rect 35909 25381 35943 25415
rect 2881 25313 2915 25347
rect 4445 25313 4479 25347
rect 5365 25313 5399 25347
rect 6285 25313 6319 25347
rect 6377 25313 6411 25347
rect 7849 25313 7883 25347
rect 9321 25313 9355 25347
rect 10333 25313 10367 25347
rect 10425 25313 10459 25347
rect 21005 25313 21039 25347
rect 21189 25313 21223 25347
rect 23673 25313 23707 25347
rect 25053 25313 25087 25347
rect 27353 25313 27387 25347
rect 27721 25313 27755 25347
rect 31677 25313 31711 25347
rect 32045 25313 32079 25347
rect 32137 25313 32171 25347
rect 2697 25245 2731 25279
rect 5641 25245 5675 25279
rect 5733 25245 5767 25279
rect 6009 25245 6043 25279
rect 6469 25245 6503 25279
rect 7113 25245 7147 25279
rect 7271 25245 7305 25279
rect 7573 25245 7607 25279
rect 8309 25245 8343 25279
rect 9137 25245 9171 25279
rect 9965 25245 9999 25279
rect 10057 25245 10091 25279
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 10793 25245 10827 25279
rect 10977 25245 11011 25279
rect 11069 25245 11103 25279
rect 11897 25245 11931 25279
rect 12081 25245 12115 25279
rect 12633 25245 12667 25279
rect 13093 25245 13127 25279
rect 13185 25245 13219 25279
rect 13369 25245 13403 25279
rect 13461 25245 13495 25279
rect 14289 25245 14323 25279
rect 14473 25245 14507 25279
rect 14657 25245 14691 25279
rect 15117 25245 15151 25279
rect 15301 25245 15335 25279
rect 15393 25245 15427 25279
rect 15485 25245 15519 25279
rect 17601 25245 17635 25279
rect 17877 25245 17911 25279
rect 18245 25245 18279 25279
rect 18521 25245 18555 25279
rect 18889 25245 18923 25279
rect 19257 25245 19291 25279
rect 19441 25245 19475 25279
rect 19809 25245 19843 25279
rect 20085 25245 20119 25279
rect 20269 25245 20303 25279
rect 21281 25245 21315 25279
rect 21649 25245 21683 25279
rect 22017 25245 22051 25279
rect 22477 25245 22511 25279
rect 23121 25245 23155 25279
rect 23949 25245 23983 25279
rect 24041 25245 24075 25279
rect 24961 25245 24995 25279
rect 25605 25245 25639 25279
rect 30849 25245 30883 25279
rect 31125 25245 31159 25279
rect 31217 25245 31251 25279
rect 31309 25245 31343 25279
rect 31493 25245 31527 25279
rect 31585 25245 31619 25279
rect 31861 25245 31895 25279
rect 31953 25245 31987 25279
rect 32505 25245 32539 25279
rect 32781 25245 32815 25279
rect 32873 25245 32907 25279
rect 32965 25245 32999 25279
rect 33057 25245 33091 25279
rect 33149 25245 33183 25279
rect 33517 25245 33551 25279
rect 33701 25245 33735 25279
rect 33793 25245 33827 25279
rect 33977 25245 34011 25279
rect 35081 25245 35115 25279
rect 35265 25245 35299 25279
rect 35725 25245 35759 25279
rect 36093 25245 36127 25279
rect 5825 25177 5859 25211
rect 7389 25177 7423 25211
rect 7481 25177 7515 25211
rect 8007 25177 8041 25211
rect 8125 25177 8159 25211
rect 8217 25177 8251 25211
rect 14381 25177 14415 25211
rect 16865 25177 16899 25211
rect 19349 25177 19383 25211
rect 22937 25177 22971 25211
rect 23581 25177 23615 25211
rect 27997 25177 28031 25211
rect 29929 25177 29963 25211
rect 2605 25109 2639 25143
rect 4261 25109 4295 25143
rect 4353 25109 4387 25143
rect 4721 25109 4755 25143
rect 5457 25109 5491 25143
rect 7757 25109 7791 25143
rect 10885 25109 10919 25143
rect 12541 25109 12575 25143
rect 12909 25109 12943 25143
rect 15669 25109 15703 25143
rect 17242 25109 17276 25143
rect 21373 25109 21407 25143
rect 23213 25109 23247 25143
rect 23305 25109 23339 25143
rect 25927 25109 25961 25143
rect 27905 25109 27939 25143
rect 29561 25109 29595 25143
rect 29729 25109 29763 25143
rect 30757 25109 30791 25143
rect 32689 25109 32723 25143
rect 33241 25109 33275 25143
rect 3249 24905 3283 24939
rect 5917 24905 5951 24939
rect 9689 24905 9723 24939
rect 12173 24905 12207 24939
rect 15853 24905 15887 24939
rect 17417 24905 17451 24939
rect 18153 24905 18187 24939
rect 27353 24905 27387 24939
rect 28825 24905 28859 24939
rect 31509 24905 31543 24939
rect 32137 24905 32171 24939
rect 33057 24905 33091 24939
rect 3617 24837 3651 24871
rect 19073 24837 19107 24871
rect 19993 24837 20027 24871
rect 21649 24837 21683 24871
rect 22661 24837 22695 24871
rect 30731 24837 30765 24871
rect 31309 24837 31343 24871
rect 21419 24803 21453 24837
rect 9686 24769 9720 24803
rect 12357 24769 12391 24803
rect 12449 24769 12483 24803
rect 12725 24769 12759 24803
rect 13277 24769 13311 24803
rect 13369 24769 13403 24803
rect 13553 24769 13587 24803
rect 13645 24769 13679 24803
rect 15577 24769 15611 24803
rect 15945 24769 15979 24803
rect 17601 24769 17635 24803
rect 17877 24769 17911 24803
rect 18521 24769 18555 24803
rect 18797 24769 18831 24803
rect 18981 24769 19015 24803
rect 19257 24769 19291 24803
rect 19901 24769 19935 24803
rect 20085 24769 20119 24803
rect 20269 24769 20303 24803
rect 22109 24769 22143 24803
rect 23305 24769 23339 24803
rect 23397 24769 23431 24803
rect 23765 24769 23799 24803
rect 24869 24769 24903 24803
rect 26157 24769 26191 24803
rect 26433 24769 26467 24803
rect 28089 24769 28123 24803
rect 28273 24769 28307 24803
rect 28549 24769 28583 24803
rect 29101 24769 29135 24803
rect 29193 24769 29227 24803
rect 29377 24769 29411 24803
rect 29469 24769 29503 24803
rect 30849 24769 30883 24803
rect 30941 24769 30975 24803
rect 31033 24769 31067 24803
rect 32321 24769 32355 24803
rect 32413 24769 32447 24803
rect 32505 24769 32539 24803
rect 32689 24769 32723 24803
rect 32873 24769 32907 24803
rect 33057 24769 33091 24803
rect 33701 24769 33735 24803
rect 33793 24769 33827 24803
rect 34161 24769 34195 24803
rect 1409 24701 1443 24735
rect 1685 24701 1719 24735
rect 3709 24701 3743 24735
rect 3801 24701 3835 24735
rect 4169 24701 4203 24735
rect 4445 24701 4479 24735
rect 6469 24701 6503 24735
rect 6745 24701 6779 24735
rect 8217 24701 8251 24735
rect 8953 24701 8987 24735
rect 10149 24701 10183 24735
rect 11621 24701 11655 24735
rect 11713 24701 11747 24735
rect 11805 24701 11839 24735
rect 11897 24701 11931 24735
rect 12081 24701 12115 24735
rect 15209 24701 15243 24735
rect 17785 24701 17819 24735
rect 19441 24701 19475 24735
rect 22017 24701 22051 24735
rect 22201 24701 22235 24735
rect 22293 24701 22327 24735
rect 22937 24701 22971 24735
rect 24685 24701 24719 24735
rect 24961 24701 24995 24735
rect 25053 24701 25087 24735
rect 25145 24701 25179 24735
rect 26341 24701 26375 24735
rect 27169 24701 27203 24735
rect 27261 24701 27295 24735
rect 28181 24701 28215 24735
rect 30573 24701 30607 24735
rect 33609 24701 33643 24735
rect 33885 24701 33919 24735
rect 34437 24701 34471 24735
rect 36185 24701 36219 24735
rect 18613 24633 18647 24667
rect 21281 24633 21315 24667
rect 27721 24633 27755 24667
rect 31677 24633 31711 24667
rect 3157 24565 3191 24599
rect 8309 24565 8343 24599
rect 9505 24565 9539 24599
rect 10057 24565 10091 24599
rect 12633 24565 12667 24599
rect 13093 24565 13127 24599
rect 15485 24565 15519 24599
rect 15669 24565 15703 24599
rect 17877 24565 17911 24599
rect 17969 24565 18003 24599
rect 18153 24565 18187 24599
rect 19717 24565 19751 24599
rect 21465 24565 21499 24599
rect 21833 24565 21867 24599
rect 25973 24565 26007 24599
rect 29653 24565 29687 24599
rect 31217 24565 31251 24599
rect 31493 24565 31527 24599
rect 34069 24565 34103 24599
rect 4721 24361 4755 24395
rect 7297 24361 7331 24395
rect 11437 24361 11471 24395
rect 12173 24361 12207 24395
rect 12357 24361 12391 24395
rect 14105 24361 14139 24395
rect 15761 24361 15795 24395
rect 15945 24361 15979 24395
rect 22385 24361 22419 24395
rect 23397 24361 23431 24395
rect 26019 24361 26053 24395
rect 26157 24361 26191 24395
rect 27629 24361 27663 24395
rect 28733 24361 28767 24395
rect 29009 24361 29043 24395
rect 29193 24361 29227 24395
rect 33333 24361 33367 24395
rect 33793 24361 33827 24395
rect 34713 24361 34747 24395
rect 35817 24361 35851 24395
rect 8401 24293 8435 24327
rect 10241 24293 10275 24327
rect 16221 24293 16255 24327
rect 20085 24293 20119 24327
rect 32689 24293 32723 24327
rect 33609 24293 33643 24327
rect 35357 24293 35391 24327
rect 5365 24225 5399 24259
rect 6101 24225 6135 24259
rect 7849 24225 7883 24259
rect 8769 24225 8803 24259
rect 10701 24225 10735 24259
rect 11621 24225 11655 24259
rect 11989 24225 12023 24259
rect 22569 24225 22603 24259
rect 22937 24225 22971 24259
rect 33885 24225 33919 24259
rect 3433 24157 3467 24191
rect 4537 24157 4571 24191
rect 5181 24157 5215 24191
rect 6469 24157 6503 24191
rect 6561 24157 6595 24191
rect 6837 24157 6871 24191
rect 7665 24157 7699 24191
rect 8585 24157 8619 24191
rect 9597 24157 9631 24191
rect 9965 24157 9999 24191
rect 10333 24157 10367 24191
rect 10793 24157 10827 24191
rect 11164 24157 11198 24191
rect 11713 24157 11747 24191
rect 12725 24157 12759 24191
rect 12818 24157 12852 24191
rect 13001 24157 13035 24191
rect 13231 24157 13265 24191
rect 14289 24157 14323 24191
rect 14473 24157 14507 24191
rect 14657 24157 14691 24191
rect 16405 24157 16439 24191
rect 16589 24157 16623 24191
rect 16773 24157 16807 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20361 24157 20395 24191
rect 22293 24157 22327 24191
rect 22753 24157 22787 24191
rect 22845 24157 22879 24191
rect 23029 24157 23063 24191
rect 24501 24157 24535 24191
rect 24685 24157 24719 24191
rect 24777 24157 24811 24191
rect 24961 24157 24995 24191
rect 25053 24157 25087 24191
rect 25145 24157 25179 24191
rect 25329 24157 25363 24191
rect 25881 24157 25915 24191
rect 26341 24157 26375 24191
rect 27261 24157 27295 24191
rect 28181 24157 28215 24191
rect 28365 24157 28399 24191
rect 28549 24157 28583 24191
rect 31033 24157 31067 24191
rect 32505 24157 32539 24191
rect 32689 24157 32723 24191
rect 33057 24157 33091 24191
rect 33977 24157 34011 24191
rect 34897 24157 34931 24191
rect 34989 24157 35023 24191
rect 35265 24157 35299 24191
rect 36093 24157 36127 24191
rect 5089 24089 5123 24123
rect 5549 24089 5583 24123
rect 6653 24089 6687 24123
rect 8217 24089 8251 24123
rect 12081 24089 12115 24123
rect 12541 24089 12575 24123
rect 13093 24089 13127 24123
rect 14381 24089 14415 24123
rect 16129 24089 16163 24123
rect 16497 24089 16531 24123
rect 20085 24089 20119 24123
rect 23581 24089 23615 24123
rect 25513 24089 25547 24123
rect 27629 24089 27663 24123
rect 28457 24089 28491 24123
rect 28871 24089 28905 24123
rect 29041 24089 29075 24123
rect 33175 24089 33209 24123
rect 33365 24089 33399 24123
rect 35081 24089 35115 24123
rect 35541 24089 35575 24123
rect 2789 24021 2823 24055
rect 3985 24021 4019 24055
rect 6285 24021 6319 24055
rect 7757 24021 7791 24055
rect 11161 24021 11195 24055
rect 11345 24021 11379 24055
rect 12341 24021 12375 24055
rect 13369 24021 13403 24055
rect 15945 24021 15979 24055
rect 19533 24021 19567 24055
rect 19901 24021 19935 24055
rect 20269 24021 20303 24055
rect 23213 24021 23247 24055
rect 23381 24021 23415 24055
rect 26249 24021 26283 24055
rect 27813 24021 27847 24055
rect 31217 24021 31251 24055
rect 32873 24021 32907 24055
rect 33517 24021 33551 24055
rect 2329 23817 2363 23851
rect 4537 23817 4571 23851
rect 10057 23817 10091 23851
rect 10241 23817 10275 23851
rect 15945 23817 15979 23851
rect 16405 23817 16439 23851
rect 17417 23817 17451 23851
rect 18061 23817 18095 23851
rect 19718 23817 19752 23851
rect 21833 23817 21867 23851
rect 28273 23817 28307 23851
rect 30465 23817 30499 23851
rect 31049 23817 31083 23851
rect 33977 23817 34011 23851
rect 5549 23749 5583 23783
rect 9229 23749 9263 23783
rect 12357 23749 12391 23783
rect 13829 23749 13863 23783
rect 13921 23749 13955 23783
rect 16681 23749 16715 23783
rect 17058 23749 17092 23783
rect 24501 23749 24535 23783
rect 25881 23749 25915 23783
rect 30665 23749 30699 23783
rect 30849 23749 30883 23783
rect 31585 23749 31619 23783
rect 2789 23681 2823 23715
rect 5181 23681 5215 23715
rect 5274 23681 5308 23715
rect 5457 23681 5491 23715
rect 5687 23681 5721 23715
rect 8953 23681 8987 23715
rect 9137 23681 9171 23715
rect 9326 23681 9360 23715
rect 10116 23681 10150 23715
rect 11345 23681 11379 23715
rect 11897 23681 11931 23715
rect 12541 23681 12575 23715
rect 12725 23681 12759 23715
rect 13093 23681 13127 23715
rect 13185 23681 13219 23715
rect 13369 23681 13403 23715
rect 13737 23681 13771 23715
rect 14105 23681 14139 23715
rect 15393 23681 15427 23715
rect 15945 23681 15979 23715
rect 16313 23681 16347 23715
rect 16497 23681 16531 23715
rect 17325 23681 17359 23715
rect 17601 23681 17635 23715
rect 18245 23681 18279 23715
rect 18521 23681 18555 23715
rect 18705 23681 18739 23715
rect 19658 23681 19692 23715
rect 22109 23681 22143 23715
rect 22569 23681 22603 23715
rect 23029 23681 23063 23715
rect 23397 23681 23431 23715
rect 24685 23681 24719 23715
rect 24777 23681 24811 23715
rect 24961 23681 24995 23715
rect 25053 23681 25087 23715
rect 25329 23681 25363 23715
rect 25421 23681 25455 23715
rect 25605 23681 25639 23715
rect 25697 23681 25731 23715
rect 25789 23681 25823 23715
rect 26065 23681 26099 23715
rect 28089 23681 28123 23715
rect 28641 23681 28675 23715
rect 28733 23681 28767 23715
rect 31309 23681 31343 23715
rect 31402 23681 31436 23715
rect 31677 23681 31711 23715
rect 31815 23681 31849 23715
rect 33057 23681 33091 23715
rect 33793 23681 33827 23715
rect 35173 23681 35207 23715
rect 36185 23681 36219 23715
rect 2421 23613 2455 23647
rect 2605 23613 2639 23647
rect 3065 23613 3099 23647
rect 6377 23613 6411 23647
rect 6653 23613 6687 23647
rect 8125 23613 8159 23647
rect 8769 23613 8803 23647
rect 9597 23613 9631 23647
rect 11785 23613 11819 23647
rect 12173 23613 12207 23647
rect 12265 23613 12299 23647
rect 15485 23613 15519 23647
rect 17693 23613 17727 23647
rect 17785 23613 17819 23647
rect 17877 23613 17911 23647
rect 18981 23613 19015 23647
rect 19073 23613 19107 23647
rect 19441 23613 19475 23647
rect 20177 23613 20211 23647
rect 22017 23613 22051 23647
rect 22201 23613 22235 23647
rect 22293 23613 22327 23647
rect 27905 23613 27939 23647
rect 33609 23613 33643 23647
rect 35265 23613 35299 23647
rect 8953 23545 8987 23579
rect 9689 23545 9723 23579
rect 11253 23545 11287 23579
rect 13277 23545 13311 23579
rect 13553 23545 13587 23579
rect 25145 23545 25179 23579
rect 26065 23545 26099 23579
rect 31217 23545 31251 23579
rect 33425 23545 33459 23579
rect 36001 23545 36035 23579
rect 1961 23477 1995 23511
rect 5825 23477 5859 23511
rect 8217 23477 8251 23511
rect 11621 23477 11655 23511
rect 12909 23477 12943 23511
rect 17049 23477 17083 23511
rect 18797 23477 18831 23511
rect 19533 23477 19567 23511
rect 20085 23477 20119 23511
rect 22845 23477 22879 23511
rect 28457 23477 28491 23511
rect 28917 23477 28951 23511
rect 30297 23477 30331 23511
rect 30481 23477 30515 23511
rect 31033 23477 31067 23511
rect 31953 23477 31987 23511
rect 33517 23477 33551 23511
rect 35173 23477 35207 23511
rect 35541 23477 35575 23511
rect 3801 23273 3835 23307
rect 9137 23273 9171 23307
rect 9689 23273 9723 23307
rect 13737 23273 13771 23307
rect 14749 23273 14783 23307
rect 17325 23273 17359 23307
rect 22845 23273 22879 23307
rect 24869 23273 24903 23307
rect 26617 23273 26651 23307
rect 27077 23273 27111 23307
rect 27169 23273 27203 23307
rect 27353 23273 27387 23307
rect 28181 23273 28215 23307
rect 28641 23273 28675 23307
rect 3157 23205 3191 23239
rect 7113 23205 7147 23239
rect 8033 23205 8067 23239
rect 12909 23205 12943 23239
rect 21235 23205 21269 23239
rect 23121 23205 23155 23239
rect 28365 23205 28399 23239
rect 29653 23205 29687 23239
rect 1409 23137 1443 23171
rect 1685 23137 1719 23171
rect 4353 23137 4387 23171
rect 7665 23137 7699 23171
rect 10057 23137 10091 23171
rect 10609 23137 10643 23171
rect 14657 23137 14691 23171
rect 17141 23137 17175 23171
rect 19257 23137 19291 23171
rect 20545 23137 20579 23171
rect 21649 23137 21683 23171
rect 22201 23137 22235 23171
rect 22569 23137 22603 23171
rect 22686 23137 22720 23171
rect 25973 23137 26007 23171
rect 31677 23137 31711 23171
rect 4169 23069 4203 23103
rect 4629 23069 4663 23103
rect 4722 23069 4756 23103
rect 4905 23069 4939 23103
rect 5133 23069 5167 23103
rect 7481 23069 7515 23103
rect 9045 23069 9079 23103
rect 9413 23069 9447 23103
rect 9597 23069 9631 23103
rect 9873 23069 9907 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 10425 23069 10459 23103
rect 10517 23069 10551 23103
rect 10701 23069 10735 23103
rect 11345 23069 11379 23103
rect 11529 23069 11563 23103
rect 12265 23069 12299 23103
rect 12449 23069 12483 23103
rect 12633 23069 12667 23103
rect 12725 23069 12759 23103
rect 13001 23069 13035 23103
rect 13185 23069 13219 23103
rect 13921 23069 13955 23103
rect 14105 23069 14139 23103
rect 14289 23069 14323 23103
rect 14749 23069 14783 23103
rect 15761 23069 15795 23103
rect 16037 23069 16071 23103
rect 16405 23069 16439 23103
rect 16497 23069 16531 23103
rect 16681 23069 16715 23103
rect 16773 23069 16807 23103
rect 16866 23069 16900 23103
rect 17509 23069 17543 23103
rect 17601 23069 17635 23103
rect 17693 23069 17727 23103
rect 18889 23069 18923 23103
rect 19073 23069 19107 23103
rect 19441 23069 19475 23103
rect 19533 23069 19567 23103
rect 19625 23069 19659 23103
rect 19809 23069 19843 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 20913 23069 20947 23103
rect 21097 23069 21131 23103
rect 21373 23069 21407 23103
rect 21741 23069 21775 23103
rect 21833 23069 21867 23103
rect 22109 23069 22143 23103
rect 23280 23069 23314 23103
rect 23765 23069 23799 23103
rect 25053 23069 25087 23103
rect 25329 23069 25363 23103
rect 26157 23069 26191 23103
rect 26249 23069 26283 23103
rect 26801 23069 26835 23103
rect 26893 23069 26927 23103
rect 28457 23069 28491 23103
rect 29837 23069 29871 23103
rect 30021 23069 30055 23103
rect 30297 23069 30331 23103
rect 30389 23069 30423 23103
rect 30573 23069 30607 23103
rect 30665 23069 30699 23103
rect 31217 23069 31251 23103
rect 31401 23069 31435 23103
rect 31519 23069 31553 23103
rect 31769 23069 31803 23103
rect 32321 23069 32355 23103
rect 35265 23069 35299 23103
rect 4261 23001 4295 23035
rect 4997 23001 5031 23035
rect 7573 23001 7607 23035
rect 8309 23001 8343 23035
rect 11713 23001 11747 23035
rect 14473 23001 14507 23035
rect 15117 23001 15151 23035
rect 22477 23001 22511 23035
rect 25237 23001 25271 23035
rect 25973 23001 26007 23035
rect 27077 23001 27111 23035
rect 27537 23001 27571 23035
rect 27997 23001 28031 23035
rect 31033 23001 31067 23035
rect 31309 23001 31343 23035
rect 35081 23001 35115 23035
rect 5273 22933 5307 22967
rect 12265 22933 12299 22967
rect 13001 22933 13035 22967
rect 14197 22933 14231 22967
rect 14933 22933 14967 22967
rect 18889 22933 18923 22967
rect 19257 22933 19291 22967
rect 19717 22933 19751 22967
rect 20913 22933 20947 22967
rect 22017 22933 22051 22967
rect 23397 22933 23431 22967
rect 23489 22933 23523 22967
rect 27337 22933 27371 22967
rect 28207 22933 28241 22967
rect 29929 22933 29963 22967
rect 30205 22933 30239 22967
rect 30849 22933 30883 22967
rect 31953 22933 31987 22967
rect 32137 22933 32171 22967
rect 35449 22933 35483 22967
rect 2973 22729 3007 22763
rect 9965 22729 9999 22763
rect 10057 22729 10091 22763
rect 13001 22729 13035 22763
rect 15301 22729 15335 22763
rect 19441 22729 19475 22763
rect 22201 22729 22235 22763
rect 23121 22729 23155 22763
rect 25237 22729 25271 22763
rect 26985 22729 27019 22763
rect 27997 22729 28031 22763
rect 30941 22729 30975 22763
rect 7665 22661 7699 22695
rect 7941 22661 7975 22695
rect 11345 22661 11379 22695
rect 13636 22661 13670 22695
rect 22017 22661 22051 22695
rect 22569 22661 22603 22695
rect 28273 22661 28307 22695
rect 28365 22661 28399 22695
rect 32137 22661 32171 22695
rect 32781 22661 32815 22695
rect 33149 22661 33183 22695
rect 34253 22661 34287 22695
rect 34345 22661 34379 22695
rect 2881 22593 2915 22627
rect 3341 22593 3375 22627
rect 4353 22593 4387 22627
rect 4445 22593 4479 22627
rect 4629 22593 4663 22627
rect 4721 22593 4755 22627
rect 4813 22593 4847 22627
rect 4997 22593 5031 22627
rect 5181 22593 5215 22627
rect 5457 22593 5491 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 6193 22593 6227 22627
rect 7849 22593 7883 22627
rect 8038 22593 8072 22627
rect 9781 22593 9815 22627
rect 10977 22593 11011 22627
rect 11989 22593 12023 22627
rect 12449 22593 12483 22627
rect 12541 22593 12575 22627
rect 12633 22593 12667 22627
rect 13060 22593 13094 22627
rect 14013 22593 14047 22627
rect 14381 22593 14415 22627
rect 14565 22593 14599 22627
rect 14657 22593 14691 22627
rect 15577 22593 15611 22627
rect 15761 22593 15795 22627
rect 16129 22593 16163 22627
rect 16865 22593 16899 22627
rect 17141 22593 17175 22627
rect 17600 22593 17634 22627
rect 17693 22593 17727 22627
rect 17785 22593 17819 22627
rect 17969 22593 18003 22627
rect 19165 22593 19199 22627
rect 19349 22593 19383 22627
rect 19625 22593 19659 22627
rect 19901 22593 19935 22627
rect 20085 22593 20119 22627
rect 20177 22593 20211 22627
rect 20361 22593 20395 22627
rect 21005 22593 21039 22627
rect 21189 22593 21223 22627
rect 21373 22593 21407 22627
rect 21833 22593 21867 22627
rect 22109 22593 22143 22627
rect 22385 22593 22419 22627
rect 22661 22593 22695 22627
rect 23121 22593 23155 22627
rect 24133 22593 24167 22627
rect 24317 22593 24351 22627
rect 24409 22593 24443 22627
rect 24501 22593 24535 22627
rect 25329 22593 25363 22627
rect 27261 22593 27295 22627
rect 27353 22593 27387 22627
rect 27445 22593 27479 22627
rect 27629 22593 27663 22627
rect 28176 22593 28210 22627
rect 28548 22593 28582 22627
rect 28641 22593 28675 22627
rect 29377 22593 29411 22627
rect 29469 22593 29503 22627
rect 29929 22593 29963 22627
rect 30021 22593 30055 22627
rect 30205 22593 30239 22627
rect 30389 22593 30423 22627
rect 30481 22593 30515 22627
rect 30665 22593 30699 22627
rect 30757 22593 30791 22627
rect 31217 22593 31251 22627
rect 32413 22593 32447 22627
rect 32873 22593 32907 22627
rect 33057 22593 33091 22627
rect 33241 22593 33275 22627
rect 34161 22593 34195 22627
rect 34529 22593 34563 22627
rect 34897 22593 34931 22627
rect 35173 22593 35207 22627
rect 3157 22525 3191 22559
rect 3985 22525 4019 22559
rect 4169 22525 4203 22559
rect 9597 22525 9631 22559
rect 10149 22525 10183 22559
rect 11161 22525 11195 22559
rect 11897 22525 11931 22559
rect 17325 22525 17359 22559
rect 19257 22525 19291 22559
rect 22753 22525 22787 22559
rect 23305 22525 23339 22559
rect 29193 22525 29227 22559
rect 29285 22525 29319 22559
rect 30113 22525 30147 22559
rect 31125 22525 31159 22559
rect 31309 22525 31343 22559
rect 31401 22525 31435 22559
rect 32229 22525 32263 22559
rect 35909 22525 35943 22559
rect 36185 22525 36219 22559
rect 6101 22457 6135 22491
rect 13461 22457 13495 22491
rect 21833 22457 21867 22491
rect 29745 22457 29779 22491
rect 33425 22457 33459 22491
rect 35173 22457 35207 22491
rect 2513 22389 2547 22423
rect 4905 22389 4939 22423
rect 7665 22389 7699 22423
rect 11253 22389 11287 22423
rect 13185 22389 13219 22423
rect 13645 22389 13679 22423
rect 14197 22389 14231 22423
rect 20269 22389 20303 22423
rect 24777 22389 24811 22423
rect 29653 22389 29687 22423
rect 31585 22389 31619 22423
rect 32137 22389 32171 22423
rect 32597 22389 32631 22423
rect 33977 22389 34011 22423
rect 1672 22185 1706 22219
rect 4629 22185 4663 22219
rect 8125 22185 8159 22219
rect 8309 22185 8343 22219
rect 14289 22185 14323 22219
rect 15485 22185 15519 22219
rect 29929 22185 29963 22219
rect 30113 22185 30147 22219
rect 30849 22185 30883 22219
rect 31033 22185 31067 22219
rect 8953 22117 8987 22151
rect 11713 22117 11747 22151
rect 18245 22117 18279 22151
rect 18429 22117 18463 22151
rect 19349 22117 19383 22151
rect 23673 22117 23707 22151
rect 1409 22049 1443 22083
rect 3157 22049 3191 22083
rect 4261 22049 4295 22083
rect 4353 22049 4387 22083
rect 6745 22049 6779 22083
rect 7665 22049 7699 22083
rect 7757 22049 7791 22083
rect 15853 22049 15887 22083
rect 16037 22049 16071 22083
rect 23765 22049 23799 22083
rect 24409 22049 24443 22083
rect 26157 22049 26191 22083
rect 26893 22049 26927 22083
rect 4808 21981 4842 22015
rect 5180 21981 5214 22015
rect 5273 21981 5307 22015
rect 5365 21981 5399 22015
rect 5549 21981 5583 22015
rect 5733 21981 5767 22015
rect 6009 21981 6043 22015
rect 6101 21981 6135 22015
rect 6285 21981 6319 22015
rect 6377 21981 6411 22015
rect 6561 21981 6595 22015
rect 6653 21981 6687 22015
rect 6837 21981 6871 22015
rect 7481 21981 7515 22015
rect 7573 21981 7607 22015
rect 8677 21981 8711 22015
rect 9228 21959 9262 21993
rect 9321 21981 9355 22015
rect 9413 21981 9447 22015
rect 9597 21981 9631 22015
rect 9873 21981 9907 22015
rect 10149 21981 10183 22015
rect 10885 21981 10919 22015
rect 11069 21981 11103 22015
rect 11161 21981 11195 22015
rect 11345 21981 11379 22015
rect 11897 21981 11931 22015
rect 12081 21981 12115 22015
rect 12173 21981 12207 22015
rect 13093 21981 13127 22015
rect 13277 21981 13311 22015
rect 13553 21981 13587 22015
rect 13829 21981 13863 22015
rect 14381 21981 14415 22015
rect 14473 21981 14507 22015
rect 15669 21981 15703 22015
rect 15945 21981 15979 22015
rect 16129 21981 16163 22015
rect 17969 21981 18003 22015
rect 18061 21981 18095 22015
rect 18561 21981 18595 22015
rect 18797 21981 18831 22015
rect 18981 21981 19015 22015
rect 19533 21981 19567 22015
rect 23397 21981 23431 22015
rect 23673 21981 23707 22015
rect 24225 21981 24259 22015
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 25053 21981 25087 22015
rect 25329 21981 25363 22015
rect 25697 21981 25731 22015
rect 26433 21981 26467 22015
rect 26525 21981 26559 22015
rect 26617 21981 26651 22015
rect 26801 21981 26835 22015
rect 27077 21981 27111 22015
rect 27169 21981 27203 22015
rect 27537 21981 27571 22015
rect 27629 21981 27663 22015
rect 4905 21913 4939 21947
rect 4997 21913 5031 21947
rect 5641 21913 5675 21947
rect 8300 21913 8334 21947
rect 12909 21913 12943 21947
rect 13737 21913 13771 21947
rect 17509 21913 17543 21947
rect 18705 21913 18739 21947
rect 29745 21913 29779 21947
rect 30665 21913 30699 21947
rect 3801 21845 3835 21879
rect 4169 21845 4203 21879
rect 5917 21845 5951 21879
rect 7941 21845 7975 21879
rect 9689 21845 9723 21879
rect 10057 21845 10091 21879
rect 10977 21845 11011 21879
rect 11253 21845 11287 21879
rect 13369 21845 13403 21879
rect 14105 21845 14139 21879
rect 23489 21845 23523 21879
rect 24041 21845 24075 21879
rect 24133 21845 24167 21879
rect 27353 21845 27387 21879
rect 29945 21845 29979 21879
rect 30865 21845 30899 21879
rect 4445 21641 4479 21675
rect 12265 21641 12299 21675
rect 15577 21641 15611 21675
rect 17325 21641 17359 21675
rect 19533 21641 19567 21675
rect 20545 21641 20579 21675
rect 21833 21641 21867 21675
rect 22585 21641 22619 21675
rect 22753 21641 22787 21675
rect 24225 21641 24259 21675
rect 25037 21641 25071 21675
rect 1777 21573 1811 21607
rect 13737 21573 13771 21607
rect 16957 21573 16991 21607
rect 17049 21573 17083 21607
rect 18429 21573 18463 21607
rect 19349 21573 19383 21607
rect 20085 21573 20119 21607
rect 20637 21573 20671 21607
rect 21985 21573 22019 21607
rect 22201 21573 22235 21607
rect 22385 21573 22419 21607
rect 25237 21573 25271 21607
rect 28319 21573 28353 21607
rect 28549 21573 28583 21607
rect 1501 21505 1535 21539
rect 3893 21505 3927 21539
rect 4537 21505 4571 21539
rect 4629 21505 4663 21539
rect 4813 21505 4847 21539
rect 4905 21505 4939 21539
rect 5089 21505 5123 21539
rect 5181 21505 5215 21539
rect 5365 21505 5399 21539
rect 7941 21505 7975 21539
rect 8493 21505 8527 21539
rect 8769 21505 8803 21539
rect 9229 21505 9263 21539
rect 9551 21505 9585 21539
rect 9873 21505 9907 21539
rect 10425 21505 10459 21539
rect 10701 21505 10735 21539
rect 11069 21505 11103 21539
rect 11161 21505 11195 21539
rect 11339 21505 11373 21539
rect 11897 21505 11931 21539
rect 12173 21505 12207 21539
rect 14013 21505 14047 21539
rect 14473 21505 14507 21539
rect 14841 21505 14875 21539
rect 15577 21505 15611 21539
rect 16865 21505 16899 21539
rect 17233 21505 17267 21539
rect 17509 21505 17543 21539
rect 17601 21505 17635 21539
rect 17693 21505 17727 21539
rect 17969 21505 18003 21539
rect 18061 21505 18095 21539
rect 18245 21505 18279 21539
rect 19073 21505 19107 21539
rect 20361 21505 20395 21539
rect 20913 21505 20947 21539
rect 24133 21505 24167 21539
rect 24317 21505 24351 21539
rect 24593 21505 24627 21539
rect 27169 21505 27203 21539
rect 28181 21505 28215 21539
rect 28457 21505 28491 21539
rect 28641 21505 28675 21539
rect 3249 21437 3283 21471
rect 5273 21437 5307 21471
rect 10517 21437 10551 21471
rect 11529 21437 11563 21471
rect 12081 21437 12115 21471
rect 15301 21437 15335 21471
rect 15485 21437 15519 21471
rect 17785 21437 17819 21471
rect 19257 21437 19291 21471
rect 20177 21437 20211 21471
rect 20729 21437 20763 21471
rect 23857 21437 23891 21471
rect 27353 21437 27387 21471
rect 9321 21369 9355 21403
rect 10977 21369 11011 21403
rect 11345 21369 11379 21403
rect 11621 21369 11655 21403
rect 18889 21369 18923 21403
rect 19717 21369 19751 21403
rect 21097 21369 21131 21403
rect 16681 21301 16715 21335
rect 18797 21301 18831 21335
rect 19533 21301 19567 21335
rect 20085 21301 20119 21335
rect 20729 21301 20763 21335
rect 22017 21301 22051 21335
rect 22569 21301 22603 21335
rect 24501 21301 24535 21335
rect 24869 21301 24903 21335
rect 25053 21301 25087 21335
rect 26985 21301 27019 21335
rect 28825 21301 28859 21335
rect 5733 21097 5767 21131
rect 13185 21097 13219 21131
rect 15669 21097 15703 21131
rect 17877 21097 17911 21131
rect 18705 21097 18739 21131
rect 20545 21097 20579 21131
rect 22753 21097 22787 21131
rect 23397 21097 23431 21131
rect 30205 21097 30239 21131
rect 33333 21097 33367 21131
rect 34897 21097 34931 21131
rect 7941 21029 7975 21063
rect 11897 21029 11931 21063
rect 16405 21029 16439 21063
rect 30941 21029 30975 21063
rect 35541 21029 35575 21063
rect 3157 20961 3191 20995
rect 7113 20961 7147 20995
rect 7297 20961 7331 20995
rect 7757 20961 7791 20995
rect 8493 20961 8527 20995
rect 8677 20961 8711 20995
rect 10241 20961 10275 20995
rect 10609 20961 10643 20995
rect 11161 20961 11195 20995
rect 11437 20961 11471 20995
rect 12173 20961 12207 20995
rect 13093 20961 13127 20995
rect 14657 20961 14691 20995
rect 16221 20961 16255 20995
rect 19257 20961 19291 20995
rect 22017 20961 22051 20995
rect 28641 20961 28675 20995
rect 30297 20961 30331 20995
rect 32597 20961 32631 20995
rect 32781 20961 32815 20995
rect 4353 20893 4387 20927
rect 4537 20893 4571 20927
rect 4721 20893 4755 20927
rect 4813 20893 4847 20927
rect 4905 20893 4939 20927
rect 5365 20893 5399 20927
rect 5549 20893 5583 20927
rect 5641 20893 5675 20927
rect 5825 20893 5859 20927
rect 7021 20893 7055 20927
rect 7205 20893 7239 20927
rect 7573 20893 7607 20927
rect 7941 20893 7975 20927
rect 8953 20893 8987 20927
rect 9689 20893 9723 20927
rect 10057 20893 10091 20927
rect 10793 20893 10827 20927
rect 11345 20893 11379 20927
rect 12265 20893 12299 20927
rect 12633 20893 12667 20927
rect 13185 20893 13219 20927
rect 14473 20893 14507 20927
rect 15485 20893 15519 20927
rect 15761 20893 15795 20927
rect 15853 20893 15887 20927
rect 16129 20893 16163 20927
rect 16313 20893 16347 20927
rect 17233 20893 17267 20927
rect 17326 20893 17360 20927
rect 17739 20893 17773 20927
rect 17969 20893 18003 20927
rect 18153 20893 18187 20927
rect 18245 20893 18279 20927
rect 18337 20893 18371 20927
rect 18429 20893 18463 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 19625 20893 19659 20927
rect 19717 20893 19751 20927
rect 19901 20893 19935 20927
rect 20049 20893 20083 20927
rect 20407 20893 20441 20927
rect 21557 20893 21591 20927
rect 22109 20893 22143 20927
rect 22477 20893 22511 20927
rect 22594 20893 22628 20927
rect 23213 20893 23247 20927
rect 28181 20887 28215 20921
rect 28273 20893 28307 20927
rect 28365 20893 28399 20927
rect 29561 20893 29595 20927
rect 29719 20893 29753 20927
rect 29929 20893 29963 20927
rect 30021 20893 30055 20927
rect 30757 20893 30791 20927
rect 31125 20893 31159 20927
rect 31309 20893 31343 20927
rect 31861 20893 31895 20927
rect 33517 20893 33551 20927
rect 33609 20893 33643 20927
rect 34897 20893 34931 20927
rect 34989 20893 35023 20927
rect 35449 20893 35483 20927
rect 35725 20893 35759 20927
rect 35817 20893 35851 20927
rect 7665 20825 7699 20859
rect 8401 20825 8435 20859
rect 12541 20825 12575 20859
rect 14289 20825 14323 20859
rect 15577 20825 15611 20859
rect 17509 20825 17543 20859
rect 17601 20825 17635 20859
rect 20177 20825 20211 20859
rect 20269 20825 20303 20859
rect 22845 20825 22879 20859
rect 28483 20825 28517 20859
rect 29837 20825 29871 20859
rect 30435 20825 30469 20859
rect 30573 20825 30607 20859
rect 30665 20825 30699 20859
rect 33333 20825 33367 20859
rect 35357 20825 35391 20859
rect 2513 20757 2547 20791
rect 2881 20757 2915 20791
rect 2973 20757 3007 20791
rect 3801 20757 3835 20791
rect 5089 20757 5123 20791
rect 5549 20757 5583 20791
rect 7481 20757 7515 20791
rect 8033 20757 8067 20791
rect 9137 20757 9171 20791
rect 9505 20757 9539 20791
rect 9597 20757 9631 20791
rect 9873 20757 9907 20791
rect 11069 20757 11103 20791
rect 11437 20757 11471 20791
rect 12817 20757 12851 20791
rect 14105 20757 14139 20791
rect 14381 20757 14415 20791
rect 15301 20757 15335 20791
rect 16037 20757 16071 20791
rect 16405 20757 16439 20791
rect 21649 20757 21683 20791
rect 21741 20757 21775 20791
rect 22385 20757 22419 20791
rect 23029 20757 23063 20791
rect 23121 20757 23155 20791
rect 27997 20757 28031 20791
rect 31493 20757 31527 20791
rect 31677 20757 31711 20791
rect 32873 20757 32907 20791
rect 33241 20757 33275 20791
rect 33793 20757 33827 20791
rect 34713 20757 34747 20791
rect 36001 20757 36035 20791
rect 3801 20553 3835 20587
rect 5273 20553 5307 20587
rect 6469 20553 6503 20587
rect 7757 20553 7791 20587
rect 8217 20553 8251 20587
rect 16221 20553 16255 20587
rect 17049 20553 17083 20587
rect 18705 20553 18739 20587
rect 20821 20553 20855 20587
rect 22109 20553 22143 20587
rect 23029 20553 23063 20587
rect 26341 20553 26375 20587
rect 26509 20553 26543 20587
rect 5733 20485 5767 20519
rect 7113 20485 7147 20519
rect 7205 20485 7239 20519
rect 13277 20485 13311 20519
rect 16865 20485 16899 20519
rect 17693 20485 17727 20519
rect 18337 20485 18371 20519
rect 18537 20485 18571 20519
rect 18797 20485 18831 20519
rect 21465 20485 21499 20519
rect 23581 20485 23615 20519
rect 26709 20485 26743 20519
rect 29745 20485 29779 20519
rect 31401 20485 31435 20519
rect 1593 20417 1627 20451
rect 4537 20417 4571 20451
rect 4721 20417 4755 20451
rect 4905 20417 4939 20451
rect 4997 20417 5031 20451
rect 5365 20417 5399 20451
rect 5458 20417 5492 20451
rect 5641 20417 5675 20451
rect 5871 20417 5905 20451
rect 6653 20417 6687 20451
rect 6837 20417 6871 20451
rect 6929 20417 6963 20451
rect 7317 20417 7351 20451
rect 8125 20417 8159 20451
rect 8769 20417 8803 20451
rect 8953 20417 8987 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 13185 20417 13219 20451
rect 13369 20417 13403 20451
rect 13645 20417 13679 20451
rect 16037 20417 16071 20451
rect 16681 20417 16715 20451
rect 17601 20417 17635 20451
rect 17785 20417 17819 20451
rect 17969 20417 18003 20451
rect 20637 20417 20671 20451
rect 20729 20417 20763 20451
rect 20913 20417 20947 20451
rect 21005 20417 21039 20451
rect 21097 20417 21131 20451
rect 21281 20417 21315 20451
rect 21557 20417 21591 20451
rect 22293 20417 22327 20451
rect 22937 20417 22971 20451
rect 23133 20417 23167 20451
rect 23949 20417 23983 20451
rect 24777 20417 24811 20451
rect 25053 20417 25087 20451
rect 25881 20417 25915 20451
rect 27261 20417 27295 20451
rect 27537 20417 27571 20451
rect 27721 20417 27755 20451
rect 27997 20417 28031 20451
rect 28181 20417 28215 20451
rect 29561 20417 29595 20451
rect 29837 20417 29871 20451
rect 29929 20417 29963 20451
rect 30665 20417 30699 20451
rect 30849 20417 30883 20451
rect 31283 20417 31317 20451
rect 31493 20417 31527 20451
rect 31585 20417 31619 20451
rect 32597 20417 32631 20451
rect 32873 20417 32907 20451
rect 33517 20417 33551 20451
rect 33609 20417 33643 20451
rect 33793 20417 33827 20451
rect 33885 20417 33919 20451
rect 34621 20417 34655 20451
rect 34805 20417 34839 20451
rect 1869 20349 1903 20383
rect 3893 20349 3927 20383
rect 4077 20349 4111 20383
rect 8401 20349 8435 20383
rect 12541 20349 12575 20383
rect 13737 20349 13771 20383
rect 14013 20349 14047 20383
rect 14289 20349 14323 20383
rect 15853 20349 15887 20383
rect 22477 20349 22511 20383
rect 23765 20349 23799 20383
rect 23857 20349 23891 20383
rect 24961 20349 24995 20383
rect 25605 20349 25639 20383
rect 27445 20349 27479 20383
rect 28089 20349 28123 20383
rect 31125 20349 31159 20383
rect 32781 20349 32815 20383
rect 33333 20349 33367 20383
rect 3433 20281 3467 20315
rect 6929 20281 6963 20315
rect 8585 20281 8619 20315
rect 17417 20281 17451 20315
rect 21281 20281 21315 20315
rect 25145 20281 25179 20315
rect 27077 20281 27111 20315
rect 3341 20213 3375 20247
rect 4813 20213 4847 20247
rect 6009 20213 6043 20247
rect 6837 20213 6871 20247
rect 8953 20213 8987 20247
rect 11529 20213 11563 20247
rect 13921 20213 13955 20247
rect 15761 20213 15795 20247
rect 18521 20213 18555 20247
rect 20085 20213 20119 20247
rect 23765 20213 23799 20247
rect 24593 20213 24627 20247
rect 26525 20213 26559 20247
rect 27629 20213 27663 20247
rect 30113 20213 30147 20247
rect 30665 20213 30699 20247
rect 31033 20213 31067 20247
rect 31769 20213 31803 20247
rect 32413 20213 32447 20247
rect 32597 20213 32631 20247
rect 34713 20213 34747 20247
rect 3801 20009 3835 20043
rect 5089 20009 5123 20043
rect 5549 20009 5583 20043
rect 7113 20009 7147 20043
rect 7481 20009 7515 20043
rect 12173 20009 12207 20043
rect 14657 20009 14691 20043
rect 15485 20009 15519 20043
rect 17233 20009 17267 20043
rect 19625 20009 19659 20043
rect 20453 20009 20487 20043
rect 24225 20009 24259 20043
rect 31493 20009 31527 20043
rect 3157 19941 3191 19975
rect 6193 19941 6227 19975
rect 14841 19941 14875 19975
rect 19441 19941 19475 19975
rect 27905 19941 27939 19975
rect 1409 19873 1443 19907
rect 1685 19873 1719 19907
rect 4445 19873 4479 19907
rect 5181 19873 5215 19907
rect 7205 19873 7239 19907
rect 7941 19873 7975 19907
rect 8125 19873 8159 19907
rect 11253 19873 11287 19907
rect 13645 19873 13679 19907
rect 16405 19873 16439 19907
rect 25421 19873 25455 19907
rect 27997 19873 28031 19907
rect 28089 19873 28123 19907
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 4813 19805 4847 19839
rect 4905 19805 4939 19839
rect 5365 19805 5399 19839
rect 6285 19805 6319 19839
rect 6469 19805 6503 19839
rect 7297 19805 7331 19839
rect 11437 19805 11471 19839
rect 11529 19805 11563 19839
rect 13921 19805 13955 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 14473 19805 14507 19839
rect 14749 19805 14783 19839
rect 14933 19805 14967 19839
rect 15209 19805 15243 19839
rect 15301 19805 15335 19839
rect 16301 19805 16335 19839
rect 16497 19805 16531 19839
rect 17049 19805 17083 19839
rect 17233 19805 17267 19839
rect 23765 19805 23799 19839
rect 23857 19805 23891 19839
rect 24041 19805 24075 19839
rect 24409 19805 24443 19839
rect 24593 19805 24627 19839
rect 24869 19805 24903 19839
rect 26709 19805 26743 19839
rect 26893 19805 26927 19839
rect 27813 19805 27847 19839
rect 28273 19805 28307 19839
rect 31309 19805 31343 19839
rect 7021 19737 7055 19771
rect 7849 19737 7883 19771
rect 9781 19737 9815 19771
rect 14381 19737 14415 19771
rect 19809 19737 19843 19771
rect 20085 19737 20119 19771
rect 20269 19737 20303 19771
rect 10057 19669 10091 19703
rect 11253 19669 11287 19703
rect 19609 19669 19643 19703
rect 26525 19669 26559 19703
rect 27629 19669 27663 19703
rect 10333 19465 10367 19499
rect 13737 19465 13771 19499
rect 17325 19465 17359 19499
rect 18797 19465 18831 19499
rect 23765 19465 23799 19499
rect 24501 19465 24535 19499
rect 25053 19465 25087 19499
rect 28917 19465 28951 19499
rect 30113 19465 30147 19499
rect 30849 19465 30883 19499
rect 3249 19397 3283 19431
rect 12173 19397 12207 19431
rect 12357 19397 12391 19431
rect 27629 19397 27663 19431
rect 29745 19397 29779 19431
rect 30481 19397 30515 19431
rect 3157 19329 3191 19363
rect 3617 19329 3651 19363
rect 4261 19329 4295 19363
rect 5365 19329 5399 19363
rect 8493 19329 8527 19363
rect 11713 19329 11747 19363
rect 11805 19329 11839 19363
rect 11897 19329 11931 19363
rect 12081 19329 12115 19363
rect 13921 19329 13955 19363
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17877 19329 17911 19363
rect 18061 19329 18095 19363
rect 18153 19329 18187 19363
rect 18301 19329 18335 19363
rect 18429 19329 18463 19363
rect 18521 19329 18555 19363
rect 18659 19329 18693 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 19165 19329 19199 19363
rect 20545 19329 20579 19363
rect 20821 19329 20855 19363
rect 21005 19329 21039 19363
rect 21264 19329 21298 19363
rect 21373 19329 21407 19363
rect 21649 19329 21683 19363
rect 24041 19329 24075 19363
rect 24146 19329 24180 19363
rect 24246 19332 24280 19366
rect 24409 19329 24443 19363
rect 24685 19329 24719 19363
rect 24869 19329 24903 19363
rect 24961 19329 24995 19363
rect 25237 19329 25271 19363
rect 25421 19329 25455 19363
rect 25513 19329 25547 19363
rect 26065 19329 26099 19363
rect 27169 19329 27203 19363
rect 28273 19329 28307 19363
rect 28366 19329 28400 19363
rect 28549 19329 28583 19363
rect 28641 19329 28675 19363
rect 28738 19329 28772 19363
rect 29469 19329 29503 19363
rect 29562 19329 29596 19363
rect 29837 19329 29871 19363
rect 29934 19329 29968 19363
rect 30205 19329 30239 19363
rect 30298 19329 30332 19363
rect 30573 19329 30607 19363
rect 30711 19329 30745 19363
rect 3341 19261 3375 19295
rect 8769 19261 8803 19295
rect 10241 19261 10275 19295
rect 10885 19261 10919 19295
rect 14105 19261 14139 19295
rect 17785 19261 17819 19295
rect 20269 19261 20303 19295
rect 26157 19261 26191 19295
rect 27261 19261 27295 19295
rect 11529 19193 11563 19227
rect 19349 19193 19383 19227
rect 26985 19193 27019 19227
rect 2789 19125 2823 19159
rect 4813 19125 4847 19159
rect 12541 19125 12575 19159
rect 17601 19125 17635 19159
rect 17693 19125 17727 19159
rect 18889 19125 18923 19159
rect 20637 19125 20671 19159
rect 20729 19125 20763 19159
rect 21097 19125 21131 19159
rect 21557 19125 21591 19159
rect 26157 19125 26191 19159
rect 26433 19125 26467 19159
rect 27537 19125 27571 19159
rect 3617 18921 3651 18955
rect 6561 18921 6595 18955
rect 8309 18921 8343 18955
rect 8585 18921 8619 18955
rect 8953 18921 8987 18955
rect 9965 18921 9999 18955
rect 17141 18921 17175 18955
rect 19441 18921 19475 18955
rect 19993 18921 20027 18955
rect 22109 18921 22143 18955
rect 22293 18921 22327 18955
rect 22661 18921 22695 18955
rect 25053 18921 25087 18955
rect 25237 18921 25271 18955
rect 26525 18921 26559 18955
rect 31953 18921 31987 18955
rect 32413 18921 32447 18955
rect 32505 18921 32539 18955
rect 32873 18921 32907 18955
rect 33333 18921 33367 18955
rect 35909 18921 35943 18955
rect 6653 18853 6687 18887
rect 19257 18853 19291 18887
rect 22753 18853 22787 18887
rect 26893 18853 26927 18887
rect 1869 18785 1903 18819
rect 4537 18785 4571 18819
rect 5089 18785 5123 18819
rect 7297 18785 7331 18819
rect 8033 18785 8067 18819
rect 9413 18785 9447 18819
rect 9505 18785 9539 18819
rect 10977 18785 11011 18819
rect 11713 18785 11747 18819
rect 12449 18785 12483 18819
rect 12633 18785 12667 18819
rect 18061 18785 18095 18819
rect 18613 18785 18647 18819
rect 19073 18785 19107 18819
rect 22569 18785 22603 18819
rect 26709 18785 26743 18819
rect 32137 18785 32171 18819
rect 32597 18785 32631 18819
rect 33517 18785 33551 18819
rect 4813 18717 4847 18751
rect 8217 18717 8251 18751
rect 8677 18717 8711 18751
rect 10241 18717 10275 18751
rect 10793 18717 10827 18751
rect 11621 18717 11655 18751
rect 14105 18717 14139 18751
rect 16589 18717 16623 18751
rect 16865 18717 16899 18751
rect 17049 18717 17083 18751
rect 17325 18717 17359 18751
rect 17417 18717 17451 18751
rect 18889 18717 18923 18751
rect 19441 18717 19475 18751
rect 19533 18717 19567 18751
rect 20821 18717 20855 18751
rect 21005 18717 21039 18751
rect 21097 18717 21131 18751
rect 21189 18717 21223 18751
rect 21281 18717 21315 18751
rect 21465 18717 21499 18751
rect 21649 18717 21683 18751
rect 22845 18717 22879 18751
rect 26157 18717 26191 18751
rect 26341 18717 26375 18751
rect 26617 18717 26651 18751
rect 32229 18717 32263 18751
rect 32505 18717 32539 18751
rect 33241 18717 33275 18751
rect 33701 18717 33735 18751
rect 34805 18717 34839 18751
rect 34898 18717 34932 18751
rect 35270 18717 35304 18751
rect 35725 18717 35759 18751
rect 19947 18683 19981 18717
rect 2145 18649 2179 18683
rect 4353 18649 4387 18683
rect 7021 18649 7055 18683
rect 7481 18649 7515 18683
rect 9965 18649 9999 18683
rect 10701 18649 10735 18683
rect 11529 18649 11563 18683
rect 14381 18649 14415 18683
rect 19717 18649 19751 18683
rect 20177 18649 20211 18683
rect 21557 18649 21591 18683
rect 22261 18649 22295 18683
rect 22477 18649 22511 18683
rect 25221 18649 25255 18683
rect 25421 18649 25455 18683
rect 27169 18649 27203 18683
rect 31953 18649 31987 18683
rect 35081 18649 35115 18683
rect 35173 18649 35207 18683
rect 35541 18649 35575 18683
rect 3985 18581 4019 18615
rect 4445 18581 4479 18615
rect 7113 18581 7147 18615
rect 9321 18581 9355 18615
rect 10149 18581 10183 18615
rect 10333 18581 10367 18615
rect 11161 18581 11195 18615
rect 11989 18581 12023 18615
rect 12357 18581 12391 18615
rect 15853 18581 15887 18615
rect 15945 18581 15979 18615
rect 16681 18581 16715 18615
rect 19809 18581 19843 18615
rect 20637 18581 20671 18615
rect 21373 18581 21407 18615
rect 25881 18581 25915 18615
rect 26249 18581 26283 18615
rect 33885 18581 33919 18615
rect 35449 18581 35483 18615
rect 3157 18377 3191 18411
rect 5181 18377 5215 18411
rect 5917 18377 5951 18411
rect 9321 18377 9355 18411
rect 9689 18377 9723 18411
rect 10885 18377 10919 18411
rect 10977 18377 11011 18411
rect 11897 18377 11931 18411
rect 12081 18377 12115 18411
rect 12541 18377 12575 18411
rect 14749 18377 14783 18411
rect 15117 18377 15151 18411
rect 18889 18377 18923 18411
rect 19717 18377 19751 18411
rect 21097 18377 21131 18411
rect 23213 18377 23247 18411
rect 23381 18377 23415 18411
rect 26249 18377 26283 18411
rect 31217 18377 31251 18411
rect 3709 18309 3743 18343
rect 9781 18309 9815 18343
rect 11713 18309 11747 18343
rect 13369 18309 13403 18343
rect 13553 18309 13587 18343
rect 18521 18309 18555 18343
rect 22661 18309 22695 18343
rect 23581 18309 23615 18343
rect 25329 18309 25363 18343
rect 25545 18309 25579 18343
rect 28181 18309 28215 18343
rect 28273 18309 28307 18343
rect 28549 18309 28583 18343
rect 30757 18309 30791 18343
rect 1409 18241 1443 18275
rect 5825 18241 5859 18275
rect 7021 18241 7055 18275
rect 11529 18241 11563 18275
rect 12173 18241 12207 18275
rect 12909 18241 12943 18275
rect 13737 18241 13771 18275
rect 18245 18241 18279 18275
rect 18393 18241 18427 18275
rect 18613 18241 18647 18275
rect 18751 18241 18785 18275
rect 20085 18241 20119 18275
rect 20269 18241 20303 18275
rect 20453 18241 20487 18275
rect 20729 18241 20763 18275
rect 21281 18241 21315 18275
rect 21465 18241 21499 18275
rect 23029 18241 23063 18275
rect 23121 18241 23155 18275
rect 23949 18241 23983 18275
rect 24133 18241 24167 18275
rect 24961 18241 24995 18275
rect 25145 18241 25179 18275
rect 25881 18241 25915 18275
rect 28043 18241 28077 18275
rect 28365 18241 28399 18275
rect 28917 18241 28951 18275
rect 31033 18241 31067 18275
rect 1685 18173 1719 18207
rect 3433 18173 3467 18207
rect 6101 18173 6135 18207
rect 7297 18173 7331 18207
rect 9965 18173 9999 18207
rect 11161 18173 11195 18207
rect 13001 18173 13035 18207
rect 13093 18173 13127 18207
rect 15209 18173 15243 18207
rect 15393 18173 15427 18207
rect 21005 18173 21039 18207
rect 22753 18173 22787 18207
rect 24593 18173 24627 18207
rect 25973 18173 26007 18207
rect 27905 18173 27939 18207
rect 30849 18173 30883 18207
rect 24685 18105 24719 18139
rect 5457 18037 5491 18071
rect 8769 18037 8803 18071
rect 10517 18037 10551 18071
rect 19993 18037 20027 18071
rect 20177 18037 20211 18071
rect 20545 18037 20579 18071
rect 20913 18037 20947 18071
rect 22845 18037 22879 18071
rect 23397 18037 23431 18071
rect 23765 18037 23799 18071
rect 24317 18037 24351 18071
rect 25513 18037 25547 18071
rect 25697 18037 25731 18071
rect 26065 18037 26099 18071
rect 28733 18037 28767 18071
rect 30757 18037 30791 18071
rect 2145 17833 2179 17867
rect 7665 17833 7699 17867
rect 13093 17833 13127 17867
rect 15301 17833 15335 17867
rect 15945 17833 15979 17867
rect 22385 17833 22419 17867
rect 22569 17833 22603 17867
rect 24225 17833 24259 17867
rect 25237 17833 25271 17867
rect 18429 17765 18463 17799
rect 20913 17765 20947 17799
rect 23673 17765 23707 17799
rect 25421 17765 25455 17799
rect 2605 17697 2639 17731
rect 2697 17697 2731 17731
rect 3525 17697 3559 17731
rect 5549 17697 5583 17731
rect 5825 17697 5859 17731
rect 7297 17697 7331 17731
rect 8217 17697 8251 17731
rect 9505 17697 9539 17731
rect 17785 17697 17819 17731
rect 25513 17697 25547 17731
rect 26249 17697 26283 17731
rect 2973 17629 3007 17663
rect 4445 17629 4479 17663
rect 10977 17629 11011 17663
rect 11161 17629 11195 17663
rect 12265 17629 12299 17663
rect 12449 17629 12483 17663
rect 12817 17629 12851 17663
rect 13001 17629 13035 17663
rect 13093 17629 13127 17663
rect 13277 17629 13311 17663
rect 13737 17629 13771 17663
rect 14473 17629 14507 17663
rect 15117 17629 15151 17663
rect 15209 17629 15243 17663
rect 15945 17629 15979 17663
rect 16037 17629 16071 17663
rect 16313 17629 16347 17663
rect 17233 17629 17267 17663
rect 17325 17629 17359 17663
rect 17601 17629 17635 17663
rect 18705 17629 18739 17663
rect 18797 17629 18831 17663
rect 18889 17629 18923 17663
rect 19073 17629 19107 17663
rect 19993 17629 20027 17663
rect 21373 17629 21407 17663
rect 23489 17629 23523 17663
rect 24041 17629 24075 17663
rect 25697 17629 25731 17663
rect 25973 17629 26007 17663
rect 26341 17629 26375 17663
rect 2513 17561 2547 17595
rect 3801 17561 3835 17595
rect 8033 17561 8067 17595
rect 8953 17561 8987 17595
rect 14657 17561 14691 17595
rect 14841 17561 14875 17595
rect 15393 17561 15427 17595
rect 16129 17561 16163 17595
rect 16497 17561 16531 17595
rect 17417 17561 17451 17595
rect 18061 17561 18095 17595
rect 21097 17561 21131 17595
rect 21281 17561 21315 17595
rect 21557 17561 21591 17595
rect 21741 17561 21775 17595
rect 22753 17561 22787 17595
rect 23857 17561 23891 17595
rect 25053 17561 25087 17595
rect 8125 17493 8159 17527
rect 11069 17493 11103 17527
rect 12357 17493 12391 17527
rect 12817 17493 12851 17527
rect 13553 17493 13587 17527
rect 14933 17493 14967 17527
rect 15669 17493 15703 17527
rect 17049 17493 17083 17527
rect 17969 17493 18003 17527
rect 18521 17493 18555 17527
rect 19809 17493 19843 17527
rect 22553 17493 22587 17527
rect 25253 17493 25287 17527
rect 25513 17493 25547 17527
rect 2697 17289 2731 17323
rect 6653 17289 6687 17323
rect 8769 17289 8803 17323
rect 9597 17289 9631 17323
rect 10149 17289 10183 17323
rect 12725 17289 12759 17323
rect 14089 17289 14123 17323
rect 14381 17289 14415 17323
rect 19809 17289 19843 17323
rect 20821 17289 20855 17323
rect 22569 17289 22603 17323
rect 22753 17289 22787 17323
rect 23305 17289 23339 17323
rect 25697 17289 25731 17323
rect 25881 17289 25915 17323
rect 27077 17289 27111 17323
rect 29485 17289 29519 17323
rect 29653 17289 29687 17323
rect 2789 17221 2823 17255
rect 10885 17221 10919 17255
rect 14289 17221 14323 17255
rect 16037 17221 16071 17255
rect 20453 17221 20487 17255
rect 23489 17221 23523 17255
rect 29285 17221 29319 17255
rect 34253 17221 34287 17255
rect 34345 17221 34379 17255
rect 34483 17221 34517 17255
rect 6101 17153 6135 17187
rect 7297 17153 7331 17187
rect 8033 17153 8067 17187
rect 8125 17153 8159 17187
rect 10057 17153 10091 17187
rect 10793 17153 10827 17187
rect 11805 17153 11839 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 12817 17153 12851 17187
rect 13645 17153 13679 17187
rect 14565 17153 14599 17187
rect 14841 17153 14875 17187
rect 15209 17153 15243 17187
rect 15301 17153 15335 17187
rect 15485 17153 15519 17187
rect 16313 17153 16347 17187
rect 16957 17153 16991 17187
rect 17049 17153 17083 17187
rect 17141 17153 17175 17187
rect 17233 17153 17267 17187
rect 17601 17153 17635 17187
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 19993 17153 20027 17187
rect 20637 17153 20671 17187
rect 20913 17153 20947 17187
rect 21061 17153 21095 17187
rect 21189 17153 21223 17187
rect 21281 17153 21315 17187
rect 21419 17153 21453 17187
rect 22293 17153 22327 17187
rect 22661 17153 22695 17187
rect 22845 17153 22879 17187
rect 23673 17153 23707 17187
rect 23949 17153 23983 17187
rect 24225 17153 24259 17187
rect 24409 17153 24443 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 32137 17153 32171 17187
rect 32229 17153 32263 17187
rect 32413 17153 32447 17187
rect 32873 17153 32907 17187
rect 32965 17153 32999 17187
rect 33149 17153 33183 17187
rect 33977 17153 34011 17187
rect 34161 17153 34195 17187
rect 2973 17085 3007 17119
rect 3617 17085 3651 17119
rect 3893 17085 3927 17119
rect 5365 17085 5399 17119
rect 8861 17085 8895 17119
rect 9045 17085 9079 17119
rect 9689 17085 9723 17119
rect 9873 17085 9907 17119
rect 11069 17085 11103 17119
rect 12633 17085 12667 17119
rect 13829 17085 13863 17119
rect 15025 17085 15059 17119
rect 16129 17085 16163 17119
rect 16773 17085 16807 17119
rect 17693 17085 17727 17119
rect 20177 17085 20211 17119
rect 22569 17085 22603 17119
rect 34621 17085 34655 17119
rect 8309 17017 8343 17051
rect 10425 17017 10459 17051
rect 15393 17017 15427 17051
rect 17969 17017 18003 17051
rect 24041 17017 24075 17051
rect 24133 17017 24167 17051
rect 24593 17017 24627 17051
rect 25329 17017 25363 17051
rect 2329 16949 2363 16983
rect 5457 16949 5491 16983
rect 8401 16949 8435 16983
rect 9229 16949 9263 16983
rect 11529 16949 11563 16983
rect 13185 16949 13219 16983
rect 13461 16949 13495 16983
rect 13921 16949 13955 16983
rect 14105 16949 14139 16983
rect 14749 16949 14783 16983
rect 16037 16949 16071 16983
rect 16497 16949 16531 16983
rect 17601 16949 17635 16983
rect 19165 16949 19199 16983
rect 19625 16949 19659 16983
rect 21557 16949 21591 16983
rect 22385 16949 22419 16983
rect 23765 16949 23799 16983
rect 25697 16949 25731 16983
rect 29469 16949 29503 16983
rect 32597 16949 32631 16983
rect 32689 16949 32723 16983
rect 32873 16949 32907 16983
rect 2132 16745 2166 16779
rect 4353 16745 4387 16779
rect 7941 16745 7975 16779
rect 10425 16745 10459 16779
rect 15393 16745 15427 16779
rect 15669 16745 15703 16779
rect 16129 16745 16163 16779
rect 17141 16745 17175 16779
rect 17417 16745 17451 16779
rect 19257 16745 19291 16779
rect 21097 16745 21131 16779
rect 21281 16745 21315 16779
rect 29745 16745 29779 16779
rect 32505 16745 32539 16779
rect 33425 16745 33459 16779
rect 25881 16677 25915 16711
rect 26065 16677 26099 16711
rect 28273 16677 28307 16711
rect 1869 16609 1903 16643
rect 4905 16609 4939 16643
rect 5641 16609 5675 16643
rect 5917 16609 5951 16643
rect 10885 16609 10919 16643
rect 10977 16609 11011 16643
rect 12817 16609 12851 16643
rect 16037 16609 16071 16643
rect 25513 16609 25547 16643
rect 29837 16609 29871 16643
rect 32413 16609 32447 16643
rect 4721 16541 4755 16575
rect 8492 16541 8526 16575
rect 8585 16541 8619 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9229 16541 9263 16575
rect 9413 16541 9447 16575
rect 9689 16541 9723 16575
rect 9873 16541 9907 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 10793 16541 10827 16575
rect 11253 16541 11287 16575
rect 11437 16541 11471 16575
rect 11713 16541 11747 16575
rect 12265 16541 12299 16575
rect 12633 16541 12667 16575
rect 13001 16541 13035 16575
rect 13277 16541 13311 16575
rect 13553 16541 13587 16575
rect 14105 16541 14139 16575
rect 14657 16541 14691 16575
rect 15485 16541 15519 16575
rect 15577 16541 15611 16575
rect 15853 16541 15887 16575
rect 17049 16541 17083 16575
rect 17141 16541 17175 16575
rect 17325 16541 17359 16575
rect 17601 16541 17635 16575
rect 17693 16541 17727 16575
rect 18153 16541 18187 16575
rect 19441 16541 19475 16575
rect 19533 16541 19567 16575
rect 19809 16541 19843 16575
rect 19901 16541 19935 16575
rect 20085 16541 20119 16575
rect 20177 16541 20211 16575
rect 20361 16541 20395 16575
rect 23305 16541 23339 16575
rect 23489 16541 23523 16575
rect 23581 16541 23615 16575
rect 23673 16541 23707 16575
rect 24961 16541 24995 16575
rect 25237 16541 25271 16575
rect 25421 16541 25455 16575
rect 25697 16541 25731 16575
rect 25973 16541 26007 16575
rect 26525 16541 26559 16575
rect 27629 16541 27663 16575
rect 27777 16541 27811 16575
rect 27905 16541 27939 16575
rect 28135 16541 28169 16575
rect 30021 16541 30055 16575
rect 32505 16541 32539 16575
rect 33609 16541 33643 16575
rect 33793 16541 33827 16575
rect 34989 16541 35023 16575
rect 35357 16541 35391 16575
rect 7925 16473 7959 16507
rect 8125 16473 8159 16507
rect 10241 16473 10275 16507
rect 16129 16473 16163 16507
rect 17417 16473 17451 16507
rect 17969 16473 18003 16507
rect 18337 16473 18371 16507
rect 19625 16473 19659 16507
rect 20913 16473 20947 16507
rect 24409 16473 24443 16507
rect 27997 16473 28031 16507
rect 29745 16473 29779 16507
rect 32229 16473 32263 16507
rect 35173 16473 35207 16507
rect 35265 16473 35299 16507
rect 3617 16405 3651 16439
rect 4813 16405 4847 16439
rect 7389 16405 7423 16439
rect 7757 16405 7791 16439
rect 8217 16405 8251 16439
rect 9137 16405 9171 16439
rect 9229 16405 9263 16439
rect 9781 16405 9815 16439
rect 11897 16405 11931 16439
rect 14197 16405 14231 16439
rect 15209 16405 15243 16439
rect 16865 16405 16899 16439
rect 17877 16405 17911 16439
rect 20545 16405 20579 16439
rect 21123 16405 21157 16439
rect 23949 16405 23983 16439
rect 26341 16405 26375 16439
rect 30205 16405 30239 16439
rect 32689 16405 32723 16439
rect 35541 16405 35575 16439
rect 6377 16201 6411 16235
rect 6745 16201 6779 16235
rect 12725 16201 12759 16235
rect 14289 16201 14323 16235
rect 15577 16201 15611 16235
rect 17233 16201 17267 16235
rect 19165 16201 19199 16235
rect 24133 16201 24167 16235
rect 25789 16201 25823 16235
rect 27629 16201 27663 16235
rect 29469 16201 29503 16235
rect 1685 16133 1719 16167
rect 17601 16133 17635 16167
rect 18705 16133 18739 16167
rect 19625 16133 19659 16167
rect 25037 16133 25071 16167
rect 25237 16133 25271 16167
rect 26249 16133 26283 16167
rect 29101 16133 29135 16167
rect 31309 16133 31343 16167
rect 1409 16065 1443 16099
rect 3801 16065 3835 16099
rect 3893 16065 3927 16099
rect 6193 16065 6227 16099
rect 6837 16065 6871 16099
rect 8217 16065 8251 16099
rect 8401 16065 8435 16099
rect 10793 16065 10827 16099
rect 10885 16065 10919 16099
rect 11069 16065 11103 16099
rect 11161 16065 11195 16099
rect 12173 16065 12207 16099
rect 12541 16065 12575 16099
rect 12633 16065 12667 16099
rect 12909 16065 12943 16099
rect 13461 16065 13495 16099
rect 13829 16065 13863 16099
rect 14105 16065 14139 16099
rect 15117 16065 15151 16099
rect 15393 16065 15427 16099
rect 17417 16065 17451 16099
rect 17509 16065 17543 16099
rect 17785 16065 17819 16099
rect 18981 16065 19015 16099
rect 19257 16065 19291 16099
rect 19405 16065 19439 16099
rect 19533 16065 19567 16099
rect 19722 16065 19756 16099
rect 22017 16065 22051 16099
rect 22201 16065 22235 16099
rect 22293 16065 22327 16099
rect 23489 16087 23523 16121
rect 23673 16065 23707 16099
rect 24317 16065 24351 16099
rect 24409 16065 24443 16099
rect 24501 16065 24535 16099
rect 24619 16065 24653 16099
rect 25605 16065 25639 16099
rect 25789 16065 25823 16099
rect 26433 16065 26467 16099
rect 26525 16065 26559 16099
rect 26709 16065 26743 16099
rect 26801 16065 26835 16099
rect 27813 16065 27847 16099
rect 27905 16065 27939 16099
rect 27997 16065 28031 16099
rect 28181 16065 28215 16099
rect 28917 16065 28951 16099
rect 29193 16065 29227 16099
rect 29285 16065 29319 16099
rect 30665 16065 30699 16099
rect 30849 16065 30883 16099
rect 31125 16065 31159 16099
rect 31401 16065 31435 16099
rect 31493 16065 31527 16099
rect 3157 15997 3191 16031
rect 4077 15997 4111 16031
rect 5917 15997 5951 16031
rect 6929 15997 6963 16031
rect 7757 15997 7791 16031
rect 13001 15997 13035 16031
rect 15301 15997 15335 16031
rect 18797 15997 18831 16031
rect 19993 15997 20027 16031
rect 20269 15997 20303 16031
rect 21833 15997 21867 16031
rect 24777 15997 24811 16031
rect 26157 15997 26191 16031
rect 3433 15929 3467 15963
rect 12081 15929 12115 15963
rect 13369 15929 13403 15963
rect 19901 15929 19935 15963
rect 23857 15929 23891 15963
rect 4445 15861 4479 15895
rect 7205 15861 7239 15895
rect 8309 15861 8343 15895
rect 10609 15861 10643 15895
rect 12265 15861 12299 15895
rect 15393 15861 15427 15895
rect 18981 15861 19015 15895
rect 23489 15861 23523 15895
rect 24869 15861 24903 15895
rect 25053 15861 25087 15895
rect 30665 15861 30699 15895
rect 31033 15861 31067 15895
rect 31677 15861 31711 15895
rect 3801 15657 3835 15691
rect 6101 15657 6135 15691
rect 12909 15657 12943 15691
rect 15025 15657 15059 15691
rect 15485 15657 15519 15691
rect 16313 15657 16347 15691
rect 17509 15657 17543 15691
rect 20453 15657 20487 15691
rect 21741 15657 21775 15691
rect 22661 15657 22695 15691
rect 25973 15657 26007 15691
rect 26525 15657 26559 15691
rect 27261 15657 27295 15691
rect 31493 15657 31527 15691
rect 8125 15589 8159 15623
rect 15853 15589 15887 15623
rect 26341 15589 26375 15623
rect 4445 15521 4479 15555
rect 6745 15521 6779 15555
rect 7757 15521 7791 15555
rect 8585 15521 8619 15555
rect 9413 15521 9447 15555
rect 12357 15521 12391 15555
rect 12725 15521 12759 15555
rect 15301 15521 15335 15555
rect 17877 15521 17911 15555
rect 17969 15521 18003 15555
rect 6469 15453 6503 15487
rect 6561 15453 6595 15487
rect 8493 15453 8527 15487
rect 8677 15453 8711 15487
rect 9137 15453 9171 15487
rect 9229 15453 9263 15487
rect 9321 15453 9355 15487
rect 9689 15453 9723 15487
rect 9873 15453 9907 15487
rect 9965 15453 9999 15487
rect 10149 15453 10183 15487
rect 10333 15453 10367 15487
rect 10517 15453 10551 15487
rect 10671 15453 10705 15487
rect 12265 15453 12299 15487
rect 12449 15453 12483 15487
rect 12541 15453 12575 15487
rect 13001 15453 13035 15487
rect 15393 15453 15427 15487
rect 15761 15453 15795 15487
rect 16037 15453 16071 15487
rect 16129 15453 16163 15487
rect 17693 15453 17727 15487
rect 19809 15453 19843 15487
rect 19993 15453 20027 15487
rect 20085 15453 20119 15487
rect 20177 15453 20211 15487
rect 22017 15453 22051 15487
rect 22109 15453 22143 15487
rect 22201 15453 22235 15487
rect 22477 15453 22511 15487
rect 26157 15453 26191 15487
rect 26433 15453 26467 15487
rect 26709 15453 26743 15487
rect 26893 15453 26927 15487
rect 26985 15453 27019 15487
rect 27077 15453 27111 15487
rect 27261 15453 27295 15487
rect 28549 15453 28583 15487
rect 28641 15453 28675 15487
rect 28917 15453 28951 15487
rect 31493 15453 31527 15487
rect 31585 15453 31619 15487
rect 33236 15453 33270 15487
rect 33425 15453 33459 15487
rect 33608 15453 33642 15487
rect 33701 15453 33735 15487
rect 12725 15385 12759 15419
rect 16313 15385 16347 15419
rect 22753 15385 22787 15419
rect 28733 15385 28767 15419
rect 31769 15385 31803 15419
rect 33333 15385 33367 15419
rect 8217 15317 8251 15351
rect 8953 15317 8987 15351
rect 10241 15317 10275 15351
rect 10885 15317 10919 15351
rect 12081 15317 12115 15351
rect 15669 15317 15703 15351
rect 22385 15317 22419 15351
rect 28365 15317 28399 15351
rect 31309 15317 31343 15351
rect 33057 15317 33091 15351
rect 4721 15113 4755 15147
rect 7389 15113 7423 15147
rect 7757 15113 7791 15147
rect 10793 15113 10827 15147
rect 12633 15113 12667 15147
rect 12817 15113 12851 15147
rect 13553 15113 13587 15147
rect 15945 15113 15979 15147
rect 17325 15113 17359 15147
rect 17877 15113 17911 15147
rect 18797 15113 18831 15147
rect 18889 15113 18923 15147
rect 19057 15113 19091 15147
rect 19349 15113 19383 15147
rect 20253 15113 20287 15147
rect 22477 15113 22511 15147
rect 26341 15113 26375 15147
rect 27721 15113 27755 15147
rect 29193 15113 29227 15147
rect 14565 15045 14599 15079
rect 15209 15045 15243 15079
rect 19257 15045 19291 15079
rect 20453 15045 20487 15079
rect 22661 15045 22695 15079
rect 23765 15045 23799 15079
rect 23857 15045 23891 15079
rect 28825 15045 28859 15079
rect 29285 15045 29319 15079
rect 31217 15045 31251 15079
rect 35173 15045 35207 15079
rect 2973 14977 3007 15011
rect 5089 14977 5123 15011
rect 5273 14977 5307 15011
rect 6837 14977 6871 15011
rect 7021 14977 7055 15011
rect 7113 14977 7147 15011
rect 8861 14977 8895 15011
rect 8953 14977 8987 15011
rect 9229 14977 9263 15011
rect 10425 14977 10459 15011
rect 10796 14977 10830 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12081 14977 12115 15011
rect 12357 14977 12391 15011
rect 12541 14977 12575 15011
rect 12758 14977 12792 15011
rect 13277 14977 13311 15011
rect 14289 14977 14323 15011
rect 14933 14977 14967 15011
rect 15025 14977 15059 15011
rect 15761 14977 15795 15011
rect 16037 14977 16071 15011
rect 17509 14977 17543 15011
rect 18061 14977 18095 15011
rect 18153 14977 18187 15011
rect 18337 14977 18371 15011
rect 18521 14977 18555 15011
rect 18613 14977 18647 15011
rect 19625 14977 19659 15011
rect 19717 14977 19751 15011
rect 19809 14977 19843 15011
rect 19993 14977 20027 15011
rect 21465 14977 21499 15011
rect 22109 14977 22143 15011
rect 22201 14977 22235 15011
rect 22569 14977 22603 15011
rect 22845 14977 22879 15011
rect 23029 14977 23063 15011
rect 23121 14977 23155 15011
rect 23305 14977 23339 15011
rect 23647 14977 23681 15011
rect 23949 14977 23983 15011
rect 24133 14977 24167 15011
rect 24501 14977 24535 15011
rect 24777 14977 24811 15011
rect 26433 14977 26467 15011
rect 26617 14977 26651 15011
rect 27077 14977 27111 15011
rect 27353 14977 27387 15011
rect 27629 14977 27663 15011
rect 27721 14977 27755 15011
rect 28549 14977 28583 15011
rect 28642 14977 28676 15011
rect 28917 14977 28951 15011
rect 29014 14977 29048 15011
rect 29561 14977 29595 15011
rect 29837 14977 29871 15011
rect 30021 14977 30055 15011
rect 31677 14977 31711 15011
rect 32413 14977 32447 15011
rect 32505 14977 32539 15011
rect 32597 14977 32631 15011
rect 32781 14977 32815 15011
rect 34943 14977 34977 15011
rect 35081 14977 35115 15011
rect 35301 14977 35335 15011
rect 35449 14977 35483 15011
rect 3249 14909 3283 14943
rect 7849 14909 7883 14943
rect 8033 14909 8067 14943
rect 10333 14909 10367 14943
rect 12173 14909 12207 14943
rect 13369 14909 13403 14943
rect 13737 14909 13771 14943
rect 14381 14909 14415 14943
rect 15301 14909 15335 14943
rect 17785 14909 17819 14943
rect 21189 14909 21223 14943
rect 23489 14909 23523 14943
rect 24409 14909 24443 14943
rect 24869 14909 24903 14943
rect 29469 14909 29503 14943
rect 31033 14909 31067 14943
rect 13185 14841 13219 14875
rect 14105 14841 14139 14875
rect 17693 14841 17727 14875
rect 20085 14841 20119 14875
rect 22937 14841 22971 14875
rect 27077 14841 27111 14875
rect 29745 14841 29779 14875
rect 5181 14773 5215 14807
rect 6653 14773 6687 14807
rect 8677 14773 8711 14807
rect 9137 14773 9171 14807
rect 10977 14773 11011 14807
rect 13921 14773 13955 14807
rect 14565 14773 14599 14807
rect 14749 14773 14783 14807
rect 14933 14773 14967 14807
rect 15577 14773 15611 14807
rect 15669 14773 15703 14807
rect 18061 14773 18095 14807
rect 19073 14773 19107 14807
rect 20269 14773 20303 14807
rect 21281 14773 21315 14807
rect 21649 14773 21683 14807
rect 21833 14773 21867 14807
rect 22293 14773 22327 14807
rect 24225 14773 24259 14807
rect 29285 14773 29319 14807
rect 30021 14773 30055 14807
rect 31493 14773 31527 14807
rect 32229 14773 32263 14807
rect 34805 14773 34839 14807
rect 4169 14569 4203 14603
rect 7113 14569 7147 14603
rect 7849 14569 7883 14603
rect 10333 14569 10367 14603
rect 12725 14569 12759 14603
rect 12909 14569 12943 14603
rect 16313 14569 16347 14603
rect 19533 14569 19567 14603
rect 19993 14569 20027 14603
rect 21373 14569 21407 14603
rect 21465 14569 21499 14603
rect 21557 14569 21591 14603
rect 22477 14569 22511 14603
rect 28365 14569 28399 14603
rect 13369 14501 13403 14535
rect 13737 14501 13771 14535
rect 16129 14501 16163 14535
rect 17141 14501 17175 14535
rect 17601 14501 17635 14535
rect 17693 14501 17727 14535
rect 18521 14501 18555 14535
rect 19901 14501 19935 14535
rect 5089 14433 5123 14467
rect 5733 14433 5767 14467
rect 6561 14433 6595 14467
rect 7205 14433 7239 14467
rect 7665 14433 7699 14467
rect 8677 14433 8711 14467
rect 9505 14433 9539 14467
rect 11345 14433 11379 14467
rect 12081 14433 12115 14467
rect 17233 14433 17267 14467
rect 19809 14433 19843 14467
rect 22753 14433 22787 14467
rect 26893 14433 26927 14467
rect 4353 14365 4387 14399
rect 4721 14365 4755 14399
rect 4997 14365 5031 14399
rect 5181 14365 5215 14399
rect 5273 14365 5307 14399
rect 5641 14365 5675 14399
rect 7573 14365 7607 14399
rect 8033 14365 8067 14399
rect 8217 14365 8251 14399
rect 8309 14365 8343 14399
rect 8585 14365 8619 14399
rect 8769 14365 8803 14399
rect 9781 14365 9815 14399
rect 10241 14365 10275 14399
rect 11897 14365 11931 14399
rect 12449 14365 12483 14399
rect 12541 14365 12575 14399
rect 13001 14365 13035 14399
rect 13093 14365 13127 14399
rect 13553 14365 13587 14399
rect 13645 14365 13679 14399
rect 13829 14365 13863 14399
rect 14657 14365 14691 14399
rect 15209 14365 15243 14399
rect 15577 14365 15611 14399
rect 15669 14365 15703 14399
rect 16313 14365 16347 14399
rect 16405 14365 16439 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 17509 14365 17543 14399
rect 17785 14365 17819 14399
rect 17972 14343 18006 14377
rect 18061 14365 18095 14399
rect 18199 14365 18233 14399
rect 18429 14365 18463 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 20269 14365 20303 14399
rect 21097 14365 21131 14399
rect 21833 14365 21867 14399
rect 22201 14365 22235 14399
rect 22661 14365 22695 14399
rect 22845 14365 22879 14399
rect 22937 14365 22971 14399
rect 24869 14365 24903 14399
rect 25237 14365 25271 14399
rect 25605 14365 25639 14399
rect 25881 14365 25915 14399
rect 26433 14365 26467 14399
rect 26801 14365 26835 14399
rect 27353 14365 27387 14399
rect 27445 14365 27479 14399
rect 27629 14365 27663 14399
rect 27813 14365 27847 14399
rect 27997 14365 28031 14399
rect 28181 14365 28215 14399
rect 29745 14365 29779 14399
rect 30481 14365 30515 14399
rect 30574 14365 30608 14399
rect 30757 14365 30791 14399
rect 30987 14365 31021 14399
rect 4445 14297 4479 14331
rect 4537 14297 4571 14331
rect 6745 14297 6779 14331
rect 10793 14297 10827 14331
rect 14749 14297 14783 14331
rect 16589 14297 16623 14331
rect 27537 14297 27571 14331
rect 28089 14297 28123 14331
rect 30849 14297 30883 14331
rect 4813 14229 4847 14263
rect 6009 14229 6043 14263
rect 6653 14229 6687 14263
rect 8953 14229 8987 14263
rect 17325 14229 17359 14263
rect 20177 14229 20211 14263
rect 21189 14229 21223 14263
rect 22017 14229 22051 14263
rect 24685 14229 24719 14263
rect 29561 14229 29595 14263
rect 31125 14229 31159 14263
rect 4353 14025 4387 14059
rect 5181 14025 5215 14059
rect 5923 14025 5957 14059
rect 8677 14025 8711 14059
rect 9781 14025 9815 14059
rect 10149 14025 10183 14059
rect 12725 14025 12759 14059
rect 15485 14025 15519 14059
rect 15945 14025 15979 14059
rect 17233 14025 17267 14059
rect 20085 14025 20119 14059
rect 26617 14025 26651 14059
rect 27077 14025 27111 14059
rect 27721 14025 27755 14059
rect 32597 14025 32631 14059
rect 4813 13957 4847 13991
rect 5365 13957 5399 13991
rect 6009 13957 6043 13991
rect 8033 13957 8067 13991
rect 8217 13957 8251 13991
rect 9045 13957 9079 13991
rect 15117 13957 15151 13991
rect 17601 13957 17635 13991
rect 19717 13957 19751 13991
rect 19927 13957 19961 13991
rect 29009 13957 29043 13991
rect 29745 13957 29779 13991
rect 32137 13957 32171 13991
rect 2605 13889 2639 13923
rect 4629 13889 4663 13923
rect 4905 13889 4939 13923
rect 5089 13889 5123 13923
rect 5273 13889 5307 13923
rect 5549 13889 5583 13923
rect 5733 13889 5767 13923
rect 5825 13889 5859 13923
rect 6101 13889 6135 13923
rect 7297 13889 7331 13923
rect 7481 13889 7515 13923
rect 7573 13889 7607 13923
rect 7844 13911 7878 13945
rect 7941 13889 7975 13923
rect 8493 13889 8527 13923
rect 8769 13889 8803 13923
rect 9229 13889 9263 13923
rect 9505 13889 9539 13923
rect 9689 13889 9723 13923
rect 9965 13889 9999 13923
rect 10241 13889 10275 13923
rect 10333 13889 10367 13923
rect 10517 13889 10551 13923
rect 10609 13889 10643 13923
rect 10885 13889 10919 13923
rect 12357 13889 12391 13923
rect 12541 13889 12575 13923
rect 13185 13889 13219 13923
rect 13553 13889 13587 13923
rect 14105 13889 14139 13923
rect 14289 13889 14323 13923
rect 14657 13889 14691 13923
rect 15025 13889 15059 13923
rect 15301 13889 15335 13923
rect 15577 13889 15611 13923
rect 15761 13889 15795 13923
rect 17417 13889 17451 13923
rect 25053 13889 25087 13923
rect 25329 13889 25363 13923
rect 25513 13889 25547 13923
rect 26525 13889 26559 13923
rect 26709 13889 26743 13923
rect 26985 13889 27019 13923
rect 27169 13889 27203 13923
rect 27537 13889 27571 13923
rect 28181 13889 28215 13923
rect 28273 13889 28307 13923
rect 28365 13889 28399 13923
rect 28503 13889 28537 13923
rect 28912 13889 28946 13923
rect 29101 13889 29135 13923
rect 29284 13889 29318 13923
rect 29388 13889 29422 13923
rect 29476 13889 29510 13923
rect 29562 13889 29596 13923
rect 29837 13889 29871 13923
rect 29975 13889 30009 13923
rect 30665 13889 30699 13923
rect 32413 13889 32447 13923
rect 7113 13821 7147 13855
rect 8309 13821 8343 13855
rect 9321 13821 9355 13855
rect 10701 13821 10735 13855
rect 13001 13821 13035 13855
rect 13369 13821 13403 13855
rect 24961 13821 24995 13855
rect 27353 13821 27387 13855
rect 27997 13821 28031 13855
rect 28641 13821 28675 13855
rect 30757 13821 30791 13855
rect 32229 13821 32263 13855
rect 4445 13753 4479 13787
rect 8217 13753 8251 13787
rect 9413 13753 9447 13787
rect 13461 13753 13495 13787
rect 28733 13753 28767 13787
rect 30113 13753 30147 13787
rect 2868 13685 2902 13719
rect 11069 13685 11103 13719
rect 12541 13685 12575 13719
rect 15669 13685 15703 13719
rect 19892 13685 19926 13719
rect 32137 13685 32171 13719
rect 4905 13481 4939 13515
rect 5365 13481 5399 13515
rect 9413 13481 9447 13515
rect 15301 13481 15335 13515
rect 15761 13481 15795 13515
rect 16037 13481 16071 13515
rect 17877 13481 17911 13515
rect 18061 13481 18095 13515
rect 18705 13481 18739 13515
rect 18889 13481 18923 13515
rect 26249 13481 26283 13515
rect 26801 13481 26835 13515
rect 31677 13481 31711 13515
rect 33333 13481 33367 13515
rect 34161 13481 34195 13515
rect 34989 13481 35023 13515
rect 10425 13413 10459 13447
rect 33149 13413 33183 13447
rect 4353 13345 4387 13379
rect 12633 13345 12667 13379
rect 16129 13345 16163 13379
rect 19257 13345 19291 13379
rect 25697 13345 25731 13379
rect 25789 13345 25823 13379
rect 31861 13345 31895 13379
rect 33517 13345 33551 13379
rect 35173 13345 35207 13379
rect 4261 13277 4295 13311
rect 4813 13277 4847 13311
rect 4997 13277 5031 13311
rect 5273 13277 5307 13311
rect 5457 13277 5491 13311
rect 6377 13277 6411 13311
rect 6561 13277 6595 13311
rect 9321 13277 9355 13311
rect 9505 13277 9539 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 10793 13277 10827 13311
rect 10977 13277 11011 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 15761 13277 15795 13311
rect 16221 13277 16255 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 18245 13277 18279 13311
rect 19441 13277 19475 13311
rect 19533 13277 19567 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 20269 13277 20303 13311
rect 20362 13277 20396 13311
rect 20637 13277 20671 13311
rect 20775 13277 20809 13311
rect 21281 13277 21315 13311
rect 21465 13277 21499 13311
rect 21649 13277 21683 13311
rect 21833 13277 21867 13311
rect 22201 13277 22235 13311
rect 25513 13277 25547 13311
rect 25605 13277 25639 13311
rect 26249 13277 26283 13311
rect 26433 13277 26467 13311
rect 26801 13277 26835 13311
rect 26985 13277 27019 13311
rect 31953 13277 31987 13311
rect 33333 13277 33367 13311
rect 34161 13277 34195 13311
rect 34345 13277 34379 13311
rect 34989 13277 35023 13311
rect 35449 13277 35483 13311
rect 19073 13209 19107 13243
rect 20545 13209 20579 13243
rect 22109 13209 22143 13243
rect 31677 13209 31711 13243
rect 33609 13209 33643 13243
rect 4629 13141 4663 13175
rect 6469 13141 6503 13175
rect 15853 13141 15887 13175
rect 17509 13141 17543 13175
rect 18873 13141 18907 13175
rect 20913 13141 20947 13175
rect 25329 13141 25363 13175
rect 32137 13141 32171 13175
rect 34529 13141 34563 13175
rect 34805 13141 34839 13175
rect 5365 12937 5399 12971
rect 15301 12937 15335 12971
rect 15761 12937 15795 12971
rect 17233 12937 17267 12971
rect 18429 12937 18463 12971
rect 19809 12937 19843 12971
rect 20529 12937 20563 12971
rect 31217 12937 31251 12971
rect 5733 12869 5767 12903
rect 6469 12869 6503 12903
rect 8217 12869 8251 12903
rect 9137 12869 9171 12903
rect 17417 12869 17451 12903
rect 20729 12869 20763 12903
rect 27721 12869 27755 12903
rect 28273 12869 28307 12903
rect 5549 12801 5583 12835
rect 6377 12801 6411 12835
rect 6561 12801 6595 12835
rect 7021 12801 7055 12835
rect 8125 12801 8159 12835
rect 8309 12801 8343 12835
rect 8580 12801 8614 12835
rect 8677 12801 8711 12835
rect 8769 12801 8803 12835
rect 8897 12801 8931 12835
rect 9045 12801 9079 12835
rect 9321 12801 9355 12835
rect 10241 12801 10275 12835
rect 10517 12801 10551 12835
rect 10793 12801 10827 12835
rect 10977 12801 11011 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 15025 12801 15059 12835
rect 15209 12801 15243 12835
rect 15577 12801 15611 12835
rect 15669 12801 15703 12835
rect 15945 12801 15979 12835
rect 16129 12801 16163 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 17601 12801 17635 12835
rect 17693 12801 17727 12835
rect 17877 12801 17911 12835
rect 17969 12801 18003 12835
rect 18061 12801 18095 12835
rect 18245 12801 18279 12835
rect 19993 12801 20027 12835
rect 20177 12801 20211 12835
rect 22569 12801 22603 12835
rect 23581 12801 23615 12835
rect 23673 12801 23707 12835
rect 24225 12801 24259 12835
rect 25421 12801 25455 12835
rect 26157 12801 26191 12835
rect 26341 12801 26375 12835
rect 26525 12801 26559 12835
rect 26709 12801 26743 12835
rect 27077 12801 27111 12835
rect 27445 12801 27479 12835
rect 27813 12801 27847 12835
rect 27997 12801 28031 12835
rect 28089 12801 28123 12835
rect 28365 12801 28399 12835
rect 28457 12801 28491 12835
rect 29009 12801 29043 12835
rect 30573 12801 30607 12835
rect 30721 12801 30755 12835
rect 30849 12801 30883 12835
rect 30941 12801 30975 12835
rect 31038 12801 31072 12835
rect 7573 12733 7607 12767
rect 8033 12733 8067 12767
rect 10425 12733 10459 12767
rect 20269 12733 20303 12767
rect 24409 12733 24443 12767
rect 25145 12733 25179 12767
rect 25513 12733 25547 12767
rect 25973 12733 26007 12767
rect 7941 12665 7975 12699
rect 24685 12665 24719 12699
rect 25881 12665 25915 12699
rect 26709 12665 26743 12699
rect 28641 12665 28675 12699
rect 8401 12597 8435 12631
rect 9505 12597 9539 12631
rect 10057 12597 10091 12631
rect 10609 12597 10643 12631
rect 10977 12597 11011 12631
rect 11713 12597 11747 12631
rect 15025 12597 15059 12631
rect 15669 12597 15703 12631
rect 16865 12597 16899 12631
rect 18061 12597 18095 12631
rect 20361 12597 20395 12631
rect 20545 12597 20579 12631
rect 26157 12597 26191 12631
rect 27997 12597 28031 12631
rect 28825 12597 28859 12631
rect 3985 12393 4019 12427
rect 8769 12393 8803 12427
rect 13093 12393 13127 12427
rect 13737 12393 13771 12427
rect 14197 12393 14231 12427
rect 14749 12393 14783 12427
rect 15209 12393 15243 12427
rect 15669 12393 15703 12427
rect 16865 12393 16899 12427
rect 17325 12393 17359 12427
rect 18061 12393 18095 12427
rect 18521 12393 18555 12427
rect 18889 12393 18923 12427
rect 19257 12393 19291 12427
rect 20085 12393 20119 12427
rect 20269 12393 20303 12427
rect 21373 12393 21407 12427
rect 24409 12393 24443 12427
rect 27353 12393 27387 12427
rect 32505 12393 32539 12427
rect 33149 12393 33183 12427
rect 10517 12325 10551 12359
rect 14565 12325 14599 12359
rect 14841 12325 14875 12359
rect 19533 12325 19567 12359
rect 26433 12325 26467 12359
rect 5457 12257 5491 12291
rect 6837 12257 6871 12291
rect 9137 12257 9171 12291
rect 9597 12257 9631 12291
rect 9873 12257 9907 12291
rect 11345 12257 11379 12291
rect 12081 12257 12115 12291
rect 12173 12257 12207 12291
rect 15393 12257 15427 12291
rect 16957 12257 16991 12291
rect 18429 12257 18463 12291
rect 21189 12257 21223 12291
rect 22569 12257 22603 12291
rect 29101 12257 29135 12291
rect 33057 12257 33091 12291
rect 4445 12189 4479 12223
rect 4537 12189 4571 12223
rect 4813 12189 4847 12223
rect 6101 12189 6135 12223
rect 6377 12189 6411 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 8125 12189 8159 12223
rect 8401 12189 8435 12223
rect 8493 12189 8527 12223
rect 8585 12189 8619 12223
rect 9229 12189 9263 12223
rect 9965 12189 9999 12223
rect 10336 12189 10370 12223
rect 10793 12189 10827 12223
rect 10885 12189 10919 12223
rect 11161 12189 11195 12223
rect 11253 12189 11287 12223
rect 11529 12189 11563 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 12357 12189 12391 12223
rect 12817 12189 12851 12223
rect 13001 12189 13035 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14105 12189 14139 12223
rect 14381 12189 14415 12223
rect 14933 12189 14967 12223
rect 15485 12189 15519 12223
rect 16129 12189 16163 12223
rect 16222 12189 16256 12223
rect 16497 12189 16531 12223
rect 16594 12189 16628 12223
rect 17141 12189 17175 12223
rect 18245 12189 18279 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 19717 12189 19751 12223
rect 21373 12189 21407 12223
rect 23673 12189 23707 12223
rect 24041 12189 24075 12223
rect 24593 12189 24627 12223
rect 24869 12189 24903 12223
rect 26433 12189 26467 12223
rect 26617 12189 26651 12223
rect 27077 12189 27111 12223
rect 27169 12189 27203 12223
rect 27353 12189 27387 12223
rect 28917 12189 28951 12223
rect 32229 12189 32263 12223
rect 32413 12189 32447 12223
rect 32505 12189 32539 12223
rect 32965 12189 32999 12223
rect 33241 12189 33275 12223
rect 4077 12121 4111 12155
rect 4629 12121 4663 12155
rect 6193 12121 6227 12155
rect 7573 12121 7607 12155
rect 7941 12121 7975 12155
rect 8283 12121 8317 12155
rect 9505 12121 9539 12155
rect 10977 12121 11011 12155
rect 12909 12121 12943 12155
rect 13921 12121 13955 12155
rect 14657 12121 14691 12155
rect 15209 12121 15243 12155
rect 16405 12121 16439 12155
rect 16865 12121 16899 12155
rect 18521 12121 18555 12155
rect 18873 12121 18907 12155
rect 19073 12121 19107 12155
rect 20453 12121 20487 12155
rect 21097 12121 21131 12155
rect 22017 12121 22051 12155
rect 22201 12121 22235 12155
rect 22385 12121 22419 12155
rect 23397 12121 23431 12155
rect 23765 12121 23799 12155
rect 23857 12121 23891 12155
rect 27629 12121 27663 12155
rect 28365 12121 28399 12155
rect 4261 12053 4295 12087
rect 4905 12053 4939 12087
rect 5273 12053 5307 12087
rect 5365 12053 5399 12087
rect 6561 12053 6595 12087
rect 8953 12053 8987 12087
rect 10333 12053 10367 12087
rect 10609 12053 10643 12087
rect 11713 12053 11747 12087
rect 12541 12053 12575 12087
rect 13553 12053 13587 12087
rect 13721 12053 13755 12087
rect 16773 12053 16807 12087
rect 18705 12053 18739 12087
rect 20253 12053 20287 12087
rect 21557 12053 21591 12087
rect 23489 12053 23523 12087
rect 24777 12053 24811 12087
rect 26893 12053 26927 12087
rect 28733 12053 28767 12087
rect 32689 12053 32723 12087
rect 32781 12053 32815 12087
rect 4629 11849 4663 11883
rect 4721 11849 4755 11883
rect 5181 11849 5215 11883
rect 6193 11849 6227 11883
rect 7665 11849 7699 11883
rect 7757 11849 7791 11883
rect 10701 11849 10735 11883
rect 11529 11849 11563 11883
rect 12449 11849 12483 11883
rect 14841 11849 14875 11883
rect 27353 11849 27387 11883
rect 31677 11849 31711 11883
rect 35357 11849 35391 11883
rect 3157 11781 3191 11815
rect 7297 11781 7331 11815
rect 15025 11781 15059 11815
rect 15577 11781 15611 11815
rect 18337 11781 18371 11815
rect 18429 11781 18463 11815
rect 20545 11781 20579 11815
rect 20761 11781 20795 11815
rect 23029 11781 23063 11815
rect 28523 11781 28557 11815
rect 28641 11781 28675 11815
rect 28733 11781 28767 11815
rect 31309 11781 31343 11815
rect 32321 11781 32355 11815
rect 34897 11781 34931 11815
rect 4905 11713 4939 11747
rect 4997 11713 5031 11747
rect 5733 11713 5767 11747
rect 5825 11713 5859 11747
rect 7573 11713 7607 11747
rect 8217 11713 8251 11747
rect 8401 11713 8435 11747
rect 9321 11713 9355 11747
rect 10333 11713 10367 11747
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 10977 11713 11011 11747
rect 11529 11713 11563 11747
rect 12357 11713 12391 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 15209 11713 15243 11747
rect 15761 11713 15795 11747
rect 18153 11713 18187 11747
rect 18613 11713 18647 11747
rect 18797 11713 18831 11747
rect 18889 11713 18923 11747
rect 21189 11713 21223 11747
rect 21465 11713 21499 11747
rect 22845 11713 22879 11747
rect 23765 11713 23799 11747
rect 24041 11713 24075 11747
rect 24961 11713 24995 11747
rect 25237 11713 25271 11747
rect 25789 11713 25823 11747
rect 26709 11713 26743 11747
rect 26985 11713 27019 11747
rect 27629 11713 27663 11747
rect 28273 11713 28307 11747
rect 28825 11713 28859 11747
rect 29009 11713 29043 11747
rect 29101 11713 29135 11747
rect 29193 11713 29227 11747
rect 31033 11713 31067 11747
rect 31126 11713 31160 11747
rect 31401 11713 31435 11747
rect 31539 11713 31573 11747
rect 32597 11713 32631 11747
rect 33149 11713 33183 11747
rect 33307 11713 33341 11747
rect 33425 11713 33459 11747
rect 33517 11713 33551 11747
rect 33609 11713 33643 11747
rect 33885 11713 33919 11747
rect 33977 11713 34011 11747
rect 35173 11713 35207 11747
rect 2881 11645 2915 11679
rect 4721 11645 4755 11679
rect 5457 11645 5491 11679
rect 5917 11645 5951 11679
rect 6469 11645 6503 11679
rect 8493 11645 8527 11679
rect 9413 11645 9447 11679
rect 9505 11645 9539 11679
rect 9597 11645 9631 11679
rect 11805 11645 11839 11679
rect 24685 11645 24719 11679
rect 25513 11645 25547 11679
rect 27169 11645 27203 11679
rect 27261 11645 27295 11679
rect 27537 11645 27571 11679
rect 28365 11645 28399 11679
rect 32413 11645 32447 11679
rect 34989 11645 35023 11679
rect 7941 11577 7975 11611
rect 8861 11577 8895 11611
rect 11621 11577 11655 11611
rect 12725 11577 12759 11611
rect 20913 11577 20947 11611
rect 24777 11577 24811 11611
rect 26065 11577 26099 11611
rect 29469 11577 29503 11611
rect 5457 11509 5491 11543
rect 5917 11509 5951 11543
rect 7389 11509 7423 11543
rect 8033 11509 8067 11543
rect 8953 11509 8987 11543
rect 9137 11509 9171 11543
rect 11069 11509 11103 11543
rect 15945 11509 15979 11543
rect 17969 11509 18003 11543
rect 20729 11509 20763 11543
rect 21281 11509 21315 11543
rect 21649 11509 21683 11543
rect 24225 11509 24259 11543
rect 29193 11509 29227 11543
rect 32505 11509 32539 11543
rect 32781 11509 32815 11543
rect 33793 11509 33827 11543
rect 33885 11509 33919 11543
rect 34253 11509 34287 11543
rect 34897 11509 34931 11543
rect 5273 11305 5307 11339
rect 5825 11305 5859 11339
rect 7481 11305 7515 11339
rect 12541 11305 12575 11339
rect 18153 11305 18187 11339
rect 19257 11305 19291 11339
rect 20545 11305 20579 11339
rect 21465 11305 21499 11339
rect 22477 11305 22511 11339
rect 22661 11305 22695 11339
rect 23029 11305 23063 11339
rect 23121 11305 23155 11339
rect 24777 11305 24811 11339
rect 25145 11305 25179 11339
rect 30389 11305 30423 11339
rect 30573 11305 30607 11339
rect 33517 11305 33551 11339
rect 33793 11305 33827 11339
rect 7297 11237 7331 11271
rect 19533 11237 19567 11271
rect 20361 11237 20395 11271
rect 22109 11237 22143 11271
rect 25237 11237 25271 11271
rect 29377 11237 29411 11271
rect 6193 11169 6227 11203
rect 8401 11169 8435 11203
rect 17509 11169 17543 11203
rect 19625 11169 19659 11203
rect 19993 11169 20027 11203
rect 20453 11169 20487 11203
rect 22385 11169 22419 11203
rect 25421 11169 25455 11203
rect 30665 11169 30699 11203
rect 33885 11169 33919 11203
rect 5089 11101 5123 11135
rect 5273 11101 5307 11135
rect 6009 11101 6043 11135
rect 6377 11101 6411 11135
rect 8125 11101 8159 11135
rect 8217 11101 8251 11135
rect 8493 11101 8527 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 13001 11101 13035 11135
rect 16312 11101 16346 11135
rect 16405 11101 16439 11135
rect 16497 11101 16531 11135
rect 16681 11101 16715 11135
rect 17141 11101 17175 11135
rect 17325 11101 17359 11135
rect 18061 11101 18095 11135
rect 18153 11101 18187 11135
rect 18337 11101 18371 11135
rect 19441 11101 19475 11135
rect 19717 11101 19751 11135
rect 19901 11101 19935 11135
rect 20177 11101 20211 11135
rect 20729 11101 20763 11135
rect 20821 11101 20855 11135
rect 21189 11101 21223 11135
rect 21281 11101 21315 11135
rect 21557 11101 21591 11135
rect 21741 11101 21775 11135
rect 22201 11101 22235 11135
rect 22477 11101 22511 11135
rect 23213 11101 23247 11135
rect 23489 11101 23523 11135
rect 24501 11101 24535 11135
rect 24961 11101 24995 11135
rect 25145 11101 25179 11135
rect 25697 11101 25731 11135
rect 25881 11101 25915 11135
rect 26893 11101 26927 11135
rect 27261 11101 27295 11135
rect 28089 11101 28123 11135
rect 28181 11101 28215 11135
rect 28365 11101 28399 11135
rect 28457 11101 28491 11135
rect 28549 11101 28583 11135
rect 28825 11101 28859 11135
rect 29009 11101 29043 11135
rect 29101 11101 29135 11135
rect 29193 11101 29227 11135
rect 30573 11101 30607 11135
rect 30849 11101 30883 11135
rect 32689 11101 32723 11135
rect 33701 11101 33735 11135
rect 33977 11101 34011 11135
rect 7465 11033 7499 11067
rect 7665 11033 7699 11067
rect 7941 11033 7975 11067
rect 16037 11033 16071 11067
rect 20959 11033 20993 11067
rect 21097 11033 21131 11067
rect 21925 11033 21959 11067
rect 22753 11033 22787 11067
rect 25789 11033 25823 11067
rect 32321 11033 32355 11067
rect 32505 11033 32539 11067
rect 13001 10965 13035 10999
rect 17877 10965 17911 10999
rect 21833 10965 21867 10999
rect 23397 10965 23431 10999
rect 28733 10965 28767 10999
rect 6101 10761 6135 10795
rect 8401 10761 8435 10795
rect 21097 10761 21131 10795
rect 27905 10761 27939 10795
rect 29285 10761 29319 10795
rect 32597 10761 32631 10795
rect 35173 10761 35207 10795
rect 5917 10693 5951 10727
rect 6377 10693 6411 10727
rect 10425 10693 10459 10727
rect 14473 10693 14507 10727
rect 15853 10693 15887 10727
rect 17141 10693 17175 10727
rect 21265 10693 21299 10727
rect 21465 10693 21499 10727
rect 23857 10693 23891 10727
rect 24317 10693 24351 10727
rect 28825 10693 28859 10727
rect 34345 10693 34379 10727
rect 34529 10693 34563 10727
rect 35633 10693 35667 10727
rect 6193 10625 6227 10659
rect 6561 10625 6595 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 6837 10625 6871 10659
rect 7021 10625 7055 10659
rect 7113 10625 7147 10659
rect 7665 10625 7699 10659
rect 7757 10625 7791 10659
rect 7941 10625 7975 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 8585 10625 8619 10659
rect 9689 10625 9723 10659
rect 9873 10625 9907 10659
rect 10241 10625 10275 10659
rect 10701 10625 10735 10659
rect 10793 10625 10827 10659
rect 10885 10625 10919 10659
rect 11069 10625 11103 10659
rect 12081 10625 12115 10659
rect 12725 10625 12759 10659
rect 13001 10625 13035 10659
rect 13185 10625 13219 10659
rect 13277 10625 13311 10659
rect 13461 10625 13495 10659
rect 13921 10625 13955 10659
rect 14105 10625 14139 10659
rect 14749 10625 14783 10659
rect 15117 10625 15151 10659
rect 15577 10625 15611 10659
rect 15669 10625 15703 10659
rect 16037 10625 16071 10659
rect 16865 10625 16899 10659
rect 19901 10625 19935 10659
rect 19993 10625 20027 10659
rect 20177 10625 20211 10659
rect 20269 10625 20303 10659
rect 23581 10625 23615 10659
rect 24225 10625 24259 10659
rect 24409 10625 24443 10659
rect 24593 10625 24627 10659
rect 25237 10625 25271 10659
rect 25421 10625 25455 10659
rect 25697 10625 25731 10659
rect 25881 10625 25915 10659
rect 25973 10625 26007 10659
rect 26249 10625 26283 10659
rect 26341 10625 26375 10659
rect 26709 10625 26743 10659
rect 27169 10625 27203 10659
rect 27445 10625 27479 10659
rect 28089 10625 28123 10659
rect 28365 10625 28399 10659
rect 28549 10625 28583 10659
rect 28641 10625 28675 10659
rect 28917 10625 28951 10659
rect 29033 10625 29067 10659
rect 29469 10625 29503 10659
rect 29653 10625 29687 10659
rect 32137 10625 32171 10659
rect 32413 10625 32447 10659
rect 34713 10625 34747 10659
rect 35357 10625 35391 10659
rect 35449 10625 35483 10659
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 11805 10557 11839 10591
rect 11989 10557 12023 10591
rect 12541 10557 12575 10591
rect 14013 10557 14047 10591
rect 16957 10557 16991 10591
rect 23765 10557 23799 10591
rect 25513 10557 25547 10591
rect 27261 10557 27295 10591
rect 28273 10557 28307 10591
rect 32229 10557 32263 10591
rect 6653 10489 6687 10523
rect 19717 10489 19751 10523
rect 25237 10489 25271 10523
rect 26433 10489 26467 10523
rect 28549 10489 28583 10523
rect 5917 10421 5951 10455
rect 7297 10421 7331 10455
rect 8217 10421 8251 10455
rect 8585 10421 8619 10455
rect 10517 10421 10551 10455
rect 12449 10421 12483 10455
rect 13553 10421 13587 10455
rect 16681 10421 16715 10455
rect 17141 10421 17175 10455
rect 21281 10421 21315 10455
rect 23397 10421 23431 10455
rect 23857 10421 23891 10455
rect 24041 10421 24075 10455
rect 26525 10421 26559 10455
rect 29193 10421 29227 10455
rect 32321 10421 32355 10455
rect 35633 10421 35667 10455
rect 6285 10217 6319 10251
rect 7021 10217 7055 10251
rect 7849 10217 7883 10251
rect 8585 10217 8619 10251
rect 9413 10217 9447 10251
rect 10057 10217 10091 10251
rect 11345 10217 11379 10251
rect 16037 10217 16071 10251
rect 16589 10217 16623 10251
rect 17509 10217 17543 10251
rect 17693 10217 17727 10251
rect 19809 10217 19843 10251
rect 20637 10217 20671 10251
rect 20821 10217 20855 10251
rect 22109 10217 22143 10251
rect 22201 10217 22235 10251
rect 22569 10217 22603 10251
rect 29101 10217 29135 10251
rect 31033 10217 31067 10251
rect 5549 10149 5583 10183
rect 16405 10149 16439 10183
rect 18797 10149 18831 10183
rect 18889 10149 18923 10183
rect 25973 10149 26007 10183
rect 28181 10149 28215 10183
rect 28733 10149 28767 10183
rect 3801 10081 3835 10115
rect 6377 10081 6411 10115
rect 6929 10081 6963 10115
rect 7389 10081 7423 10115
rect 7941 10081 7975 10115
rect 8677 10081 8711 10115
rect 9689 10081 9723 10115
rect 11069 10081 11103 10115
rect 12081 10081 12115 10115
rect 13001 10081 13035 10115
rect 13093 10081 13127 10115
rect 13369 10081 13403 10115
rect 16497 10081 16531 10115
rect 16957 10081 16991 10115
rect 17417 10081 17451 10115
rect 18521 10081 18555 10115
rect 20177 10081 20211 10115
rect 21097 10081 21131 10115
rect 24869 10081 24903 10115
rect 25329 10081 25363 10115
rect 25881 10081 25915 10115
rect 26433 10081 26467 10115
rect 27261 10081 27295 10115
rect 5914 10013 5948 10047
rect 7205 10013 7239 10047
rect 7665 10013 7699 10047
rect 8214 10013 8248 10047
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 9505 10013 9539 10047
rect 9781 10013 9815 10047
rect 10425 10013 10459 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 10793 10013 10827 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 11437 10013 11471 10047
rect 11621 10013 11655 10047
rect 11897 10013 11931 10047
rect 12357 10013 12391 10047
rect 12633 10013 12667 10047
rect 13461 10013 13495 10047
rect 14749 10013 14783 10047
rect 14933 10013 14967 10047
rect 16221 10013 16255 10047
rect 16773 10013 16807 10047
rect 17325 10013 17359 10047
rect 18705 10013 18739 10047
rect 18981 10013 19015 10047
rect 20085 10013 20119 10047
rect 20269 10013 20303 10047
rect 20361 10013 20395 10047
rect 20545 10013 20579 10047
rect 21465 10013 21499 10047
rect 21833 10013 21867 10047
rect 22017 10013 22051 10047
rect 22293 10013 22327 10047
rect 24777 10013 24811 10047
rect 25145 10013 25179 10047
rect 26157 10013 26191 10047
rect 26617 10013 26651 10047
rect 26985 10013 27019 10047
rect 27905 10013 27939 10047
rect 28929 10013 28963 10047
rect 29285 10013 29319 10047
rect 29653 10013 29687 10047
rect 29811 10013 29845 10047
rect 30113 10013 30147 10047
rect 30389 10013 30423 10047
rect 30757 10013 30791 10047
rect 31212 10013 31246 10047
rect 31309 10013 31343 10047
rect 31529 10013 31563 10047
rect 31677 10013 31711 10047
rect 4077 9945 4111 9979
rect 9137 9945 9171 9979
rect 12173 9945 12207 9979
rect 14657 9945 14691 9979
rect 21005 9945 21039 9979
rect 21281 9945 21315 9979
rect 28475 9945 28509 9979
rect 29929 9945 29963 9979
rect 30021 9945 30055 9979
rect 31401 9945 31435 9979
rect 5733 9877 5767 9911
rect 5917 9877 5951 9911
rect 7481 9877 7515 9911
rect 8033 9877 8067 9911
rect 8217 9877 8251 9911
rect 9051 9877 9085 9911
rect 12541 9877 12575 9911
rect 13277 9877 13311 9911
rect 13645 9877 13679 9911
rect 14841 9877 14875 9911
rect 20805 9877 20839 9911
rect 30297 9877 30331 9911
rect 10793 9673 10827 9707
rect 13461 9673 13495 9707
rect 14381 9673 14415 9707
rect 33517 9673 33551 9707
rect 34897 9673 34931 9707
rect 6837 9605 6871 9639
rect 13737 9605 13771 9639
rect 13829 9605 13863 9639
rect 19257 9605 19291 9639
rect 20453 9605 20487 9639
rect 28089 9605 28123 9639
rect 34529 9605 34563 9639
rect 6740 9537 6774 9571
rect 6929 9537 6963 9571
rect 7112 9537 7146 9571
rect 7205 9537 7239 9571
rect 10149 9537 10183 9571
rect 10241 9537 10275 9571
rect 10425 9537 10459 9571
rect 10885 9537 10919 9571
rect 11713 9537 11747 9571
rect 13645 9537 13679 9571
rect 13967 9537 14001 9571
rect 14322 9537 14356 9571
rect 14749 9537 14783 9571
rect 15393 9537 15427 9571
rect 15577 9537 15611 9571
rect 15761 9537 15795 9571
rect 15945 9537 15979 9571
rect 16221 9537 16255 9571
rect 18061 9537 18095 9571
rect 18226 9537 18260 9571
rect 18337 9537 18371 9571
rect 18429 9537 18463 9571
rect 18797 9537 18831 9571
rect 18889 9543 18923 9577
rect 19533 9537 19567 9571
rect 19625 9537 19659 9571
rect 19717 9537 19751 9571
rect 19993 9537 20027 9571
rect 20269 9537 20303 9571
rect 22477 9537 22511 9571
rect 22569 9537 22603 9571
rect 22937 9537 22971 9571
rect 23305 9537 23339 9571
rect 23397 9537 23431 9571
rect 23581 9537 23615 9571
rect 24317 9537 24351 9571
rect 24409 9537 24443 9571
rect 24593 9537 24627 9571
rect 25789 9537 25823 9571
rect 26065 9537 26099 9571
rect 26341 9537 26375 9571
rect 26617 9537 26651 9571
rect 27169 9537 27203 9571
rect 27721 9537 27755 9571
rect 27997 9537 28031 9571
rect 28549 9537 28583 9571
rect 28641 9537 28675 9571
rect 29193 9537 29227 9571
rect 29653 9537 29687 9571
rect 30113 9537 30147 9571
rect 32873 9537 32907 9571
rect 33031 9537 33065 9571
rect 33149 9537 33183 9571
rect 33241 9537 33275 9571
rect 33333 9537 33367 9571
rect 33609 9537 33643 9571
rect 34253 9537 34287 9571
rect 34346 9537 34380 9571
rect 34621 9537 34655 9571
rect 34718 9537 34752 9571
rect 4445 9469 4479 9503
rect 4721 9469 4755 9503
rect 10609 9469 10643 9503
rect 11621 9469 11655 9503
rect 14105 9469 14139 9503
rect 14841 9469 14875 9503
rect 15669 9469 15703 9503
rect 25697 9469 25731 9503
rect 27353 9469 27387 9503
rect 29009 9469 29043 9503
rect 6193 9401 6227 9435
rect 6561 9401 6595 9435
rect 12081 9401 12115 9435
rect 14197 9401 14231 9435
rect 16129 9401 16163 9435
rect 20085 9401 20119 9435
rect 22661 9401 22695 9435
rect 23581 9401 23615 9435
rect 26341 9401 26375 9435
rect 29377 9401 29411 9435
rect 33793 9401 33827 9435
rect 15209 9333 15243 9367
rect 17877 9333 17911 9367
rect 18521 9333 18555 9367
rect 18705 9333 18739 9367
rect 19809 9333 19843 9367
rect 22201 9333 22235 9367
rect 22753 9333 22787 9367
rect 24133 9333 24167 9367
rect 24593 9333 24627 9367
rect 28825 9333 28859 9367
rect 29561 9333 29595 9367
rect 30297 9333 30331 9367
rect 6285 9129 6319 9163
rect 6837 9129 6871 9163
rect 7297 9129 7331 9163
rect 18153 9129 18187 9163
rect 18613 9129 18647 9163
rect 21097 9129 21131 9163
rect 21465 9129 21499 9163
rect 21557 9129 21591 9163
rect 21925 9129 21959 9163
rect 22661 9129 22695 9163
rect 22845 9129 22879 9163
rect 24409 9129 24443 9163
rect 25053 9129 25087 9163
rect 25421 9129 25455 9163
rect 27721 9129 27755 9163
rect 31401 9129 31435 9163
rect 32781 9129 32815 9163
rect 17509 9061 17543 9095
rect 17601 9061 17635 9095
rect 24777 9061 24811 9095
rect 25881 9061 25915 9095
rect 26801 9061 26835 9095
rect 26985 9061 27019 9095
rect 27077 9061 27111 9095
rect 28641 9061 28675 9095
rect 30481 9061 30515 9095
rect 33517 9061 33551 9095
rect 8493 8993 8527 9027
rect 14749 8993 14783 9027
rect 17233 8993 17267 9027
rect 18245 8993 18279 9027
rect 18705 8993 18739 9027
rect 21649 8993 21683 9027
rect 25697 8993 25731 9027
rect 26893 8993 26927 9027
rect 32045 8993 32079 9027
rect 4537 8925 4571 8959
rect 7205 8925 7239 8959
rect 7573 8925 7607 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 9689 8925 9723 8959
rect 9965 8925 9999 8959
rect 10425 8925 10459 8959
rect 11161 8925 11195 8959
rect 11713 8925 11747 8959
rect 12817 8925 12851 8959
rect 14933 8925 14967 8959
rect 15117 8925 15151 8959
rect 17417 8925 17451 8959
rect 17693 8925 17727 8959
rect 18153 8925 18187 8959
rect 18429 8925 18463 8959
rect 21005 8925 21039 8959
rect 21281 8925 21315 8959
rect 21557 8925 21591 8959
rect 24593 8925 24627 8959
rect 24685 8925 24719 8959
rect 24869 8925 24903 8959
rect 25237 8925 25271 8959
rect 25513 8925 25547 8959
rect 27445 8925 27479 8959
rect 27905 8925 27939 8959
rect 28273 8925 28307 8959
rect 28457 8925 28491 8959
rect 29009 8925 29043 8959
rect 29561 8925 29595 8959
rect 30297 8925 30331 8959
rect 31585 8925 31619 8959
rect 31677 8925 31711 8959
rect 31769 8925 31803 8959
rect 4813 8857 4847 8891
rect 7021 8857 7055 8891
rect 7297 8857 7331 8891
rect 7481 8857 7515 8891
rect 8493 8857 8527 8891
rect 10333 8857 10367 8891
rect 12081 8857 12115 8891
rect 14473 8857 14507 8891
rect 18889 8857 18923 8891
rect 19073 8857 19107 8891
rect 22829 8857 22863 8891
rect 23029 8857 23063 8891
rect 26157 8857 26191 8891
rect 27997 8857 28031 8891
rect 28089 8857 28123 8891
rect 30113 8857 30147 8891
rect 31907 8857 31941 8891
rect 33517 8857 33551 8891
rect 9781 8789 9815 8823
rect 10149 8789 10183 8823
rect 14105 8789 14139 8823
rect 14565 8789 14599 8823
rect 15117 8789 15151 8823
rect 28917 8789 28951 8823
rect 29745 8789 29779 8823
rect 30021 8789 30055 8823
rect 32965 8789 32999 8823
rect 33057 8789 33091 8823
rect 5549 8585 5583 8619
rect 9045 8585 9079 8619
rect 17969 8585 18003 8619
rect 18705 8585 18739 8619
rect 22753 8585 22787 8619
rect 24777 8585 24811 8619
rect 27077 8585 27111 8619
rect 28181 8585 28215 8619
rect 29101 8585 29135 8619
rect 33609 8585 33643 8619
rect 34345 8585 34379 8619
rect 34989 8585 35023 8619
rect 12449 8517 12483 8551
rect 13369 8517 13403 8551
rect 22201 8517 22235 8551
rect 25789 8517 25823 8551
rect 29745 8517 29779 8551
rect 30297 8517 30331 8551
rect 30389 8517 30423 8551
rect 35081 8517 35115 8551
rect 5273 8449 5307 8483
rect 6837 8449 6871 8483
rect 8309 8449 8343 8483
rect 8677 8449 8711 8483
rect 9413 8449 9447 8483
rect 10057 8449 10091 8483
rect 10333 8449 10367 8483
rect 10977 8449 11011 8483
rect 13093 8449 13127 8483
rect 16037 8449 16071 8483
rect 16221 8449 16255 8483
rect 16773 8449 16807 8483
rect 16957 8459 16991 8493
rect 21971 8483 22005 8517
rect 17325 8449 17359 8483
rect 17417 8449 17451 8483
rect 17785 8449 17819 8483
rect 18153 8449 18187 8483
rect 18337 8449 18371 8483
rect 18521 8449 18555 8483
rect 19257 8449 19291 8483
rect 19349 8449 19383 8483
rect 19441 8449 19475 8483
rect 19625 8449 19659 8483
rect 20085 8449 20119 8483
rect 20545 8449 20579 8483
rect 20821 8449 20855 8483
rect 20913 8449 20947 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 22293 8449 22327 8483
rect 22477 8449 22511 8483
rect 22569 8449 22603 8483
rect 23765 8449 23799 8483
rect 23949 8449 23983 8483
rect 24221 8449 24255 8483
rect 24593 8449 24627 8483
rect 24685 8449 24719 8483
rect 24869 8449 24903 8483
rect 26617 8449 26651 8483
rect 27813 8449 27847 8483
rect 27905 8449 27939 8483
rect 29285 8449 29319 8483
rect 30205 8449 30239 8483
rect 30941 8449 30975 8483
rect 31033 8449 31067 8483
rect 31125 8449 31159 8483
rect 32689 8449 32723 8483
rect 33057 8449 33091 8483
rect 33425 8449 33459 8483
rect 33609 8449 33643 8483
rect 34161 8449 34195 8483
rect 34805 8449 34839 8483
rect 5549 8381 5583 8415
rect 6929 8381 6963 8415
rect 7021 8381 7055 8415
rect 7849 8381 7883 8415
rect 9505 8381 9539 8415
rect 9597 8381 9631 8415
rect 10885 8381 10919 8415
rect 11621 8381 11655 8415
rect 14841 8381 14875 8415
rect 18245 8381 18279 8415
rect 21189 8381 21223 8415
rect 24317 8373 24351 8407
rect 26157 8381 26191 8415
rect 26709 8381 26743 8415
rect 27353 8381 27387 8415
rect 28457 8381 28491 8415
rect 29469 8381 29503 8415
rect 29837 8381 29871 8415
rect 31493 8381 31527 8415
rect 31677 8381 31711 8415
rect 5365 8313 5399 8347
rect 6469 8313 6503 8347
rect 10149 8313 10183 8347
rect 10241 8313 10275 8347
rect 10517 8313 10551 8347
rect 17049 8313 17083 8347
rect 17509 8313 17543 8347
rect 17601 8313 17635 8347
rect 18981 8313 19015 8347
rect 20269 8313 20303 8347
rect 20361 8313 20395 8347
rect 21281 8313 21315 8347
rect 21649 8313 21683 8347
rect 24409 8313 24443 8347
rect 24501 8313 24535 8347
rect 29009 8313 29043 8347
rect 32873 8313 32907 8347
rect 34069 8313 34103 8347
rect 34621 8313 34655 8347
rect 10701 8245 10735 8279
rect 16129 8245 16163 8279
rect 16865 8245 16899 8279
rect 20453 8245 20487 8279
rect 21833 8245 21867 8279
rect 22017 8245 22051 8279
rect 22293 8245 22327 8279
rect 24133 8245 24167 8279
rect 26249 8245 26283 8279
rect 27445 8245 27479 8279
rect 28549 8245 28583 8279
rect 28641 8245 28675 8279
rect 7113 8041 7147 8075
rect 9229 8041 9263 8075
rect 9689 8041 9723 8075
rect 9965 8041 9999 8075
rect 10517 8041 10551 8075
rect 11253 8041 11287 8075
rect 13461 8041 13495 8075
rect 16589 8041 16623 8075
rect 17325 8041 17359 8075
rect 18889 8041 18923 8075
rect 19257 8041 19291 8075
rect 21005 8041 21039 8075
rect 21373 8041 21407 8075
rect 26801 8041 26835 8075
rect 27169 8041 27203 8075
rect 28549 8041 28583 8075
rect 28917 8041 28951 8075
rect 8125 7973 8159 8007
rect 15393 7973 15427 8007
rect 25053 7973 25087 8007
rect 26341 7973 26375 8007
rect 26709 7973 26743 8007
rect 29101 7973 29135 8007
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 7297 7905 7331 7939
rect 8217 7905 8251 7939
rect 8585 7905 8619 7939
rect 16037 7905 16071 7939
rect 26893 7905 26927 7939
rect 28273 7905 28307 7939
rect 34069 7905 34103 7939
rect 6561 7837 6595 7871
rect 7389 7837 7423 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 8401 7837 8435 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 10149 7837 10183 7871
rect 10425 7837 10459 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 11161 7837 11195 7871
rect 11345 7837 11379 7871
rect 11437 7837 11471 7871
rect 11713 7837 11747 7871
rect 14657 7837 14691 7871
rect 14750 7837 14784 7871
rect 15122 7837 15156 7871
rect 16221 7837 16255 7871
rect 17693 7837 17727 7871
rect 19533 7837 19567 7871
rect 19625 7837 19659 7871
rect 19717 7837 19751 7871
rect 19901 7837 19935 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 21741 7837 21775 7871
rect 24869 7837 24903 7871
rect 27629 7837 27663 7871
rect 27905 7837 27939 7871
rect 28181 7837 28215 7871
rect 29745 7837 29779 7871
rect 29837 7837 29871 7871
rect 30113 7837 30147 7871
rect 30389 7837 30423 7871
rect 30573 7837 30607 7871
rect 31033 7837 31067 7871
rect 31861 7837 31895 7871
rect 32045 7837 32079 7871
rect 32597 7837 32631 7871
rect 33057 7837 33091 7871
rect 33517 7837 33551 7871
rect 33609 7837 33643 7871
rect 34253 7837 34287 7871
rect 34805 7837 34839 7871
rect 34989 7837 35023 7871
rect 11989 7769 12023 7803
rect 14933 7769 14967 7803
rect 15025 7769 15059 7803
rect 15853 7769 15887 7803
rect 17509 7769 17543 7803
rect 19073 7769 19107 7803
rect 28390 7769 28424 7803
rect 29377 7769 29411 7803
rect 29561 7769 29595 7803
rect 33977 7769 34011 7803
rect 34437 7769 34471 7803
rect 9505 7701 9539 7735
rect 10333 7701 10367 7735
rect 11621 7701 11655 7735
rect 15301 7701 15335 7735
rect 15761 7701 15795 7735
rect 16589 7701 16623 7735
rect 16773 7701 16807 7735
rect 18705 7701 18739 7735
rect 18873 7701 18907 7735
rect 21557 7701 21591 7735
rect 27445 7701 27479 7735
rect 30665 7701 30699 7735
rect 31493 7701 31527 7735
rect 11621 7497 11655 7531
rect 11989 7497 12023 7531
rect 13277 7497 13311 7531
rect 14013 7497 14047 7531
rect 15025 7497 15059 7531
rect 22201 7497 22235 7531
rect 25421 7497 25455 7531
rect 25605 7497 25639 7531
rect 25881 7497 25915 7531
rect 27077 7497 27111 7531
rect 28089 7497 28123 7531
rect 29009 7497 29043 7531
rect 30113 7497 30147 7531
rect 30573 7497 30607 7531
rect 35357 7497 35391 7531
rect 11529 7429 11563 7463
rect 11897 7429 11931 7463
rect 13461 7429 13495 7463
rect 18981 7429 19015 7463
rect 20729 7429 20763 7463
rect 21465 7429 21499 7463
rect 21833 7429 21867 7463
rect 22017 7429 22051 7463
rect 22109 7429 22143 7463
rect 23213 7429 23247 7463
rect 24777 7429 24811 7463
rect 27997 7429 28031 7463
rect 29193 7429 29227 7463
rect 30941 7429 30975 7463
rect 31033 7429 31067 7463
rect 33885 7429 33919 7463
rect 20499 7395 20533 7429
rect 12173 7361 12207 7395
rect 12265 7361 12299 7395
rect 12434 7361 12468 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 13185 7361 13219 7395
rect 13829 7361 13863 7395
rect 14105 7361 14139 7395
rect 14381 7361 14415 7395
rect 16865 7361 16899 7395
rect 17141 7361 17175 7395
rect 17325 7361 17359 7395
rect 19257 7361 19291 7395
rect 19349 7361 19383 7395
rect 19441 7361 19475 7395
rect 19625 7361 19659 7395
rect 19993 7361 20027 7395
rect 21373 7361 21407 7395
rect 23029 7361 23063 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 24409 7361 24443 7395
rect 24501 7361 24535 7395
rect 24869 7361 24903 7395
rect 24961 7361 24995 7395
rect 25145 7361 25179 7395
rect 25237 7361 25271 7395
rect 25513 7361 25547 7395
rect 26617 7361 26651 7395
rect 27261 7361 27295 7395
rect 27629 7361 27663 7395
rect 28641 7361 28675 7395
rect 29285 7361 29319 7395
rect 29653 7361 29687 7395
rect 30021 7361 30055 7395
rect 30205 7361 30239 7395
rect 30757 7361 30791 7395
rect 31401 7361 31435 7395
rect 31493 7361 31527 7395
rect 31953 7361 31987 7395
rect 14197 7293 14231 7327
rect 14565 7293 14599 7327
rect 15117 7293 15151 7327
rect 15209 7293 15243 7327
rect 19717 7293 19751 7327
rect 19901 7293 19935 7327
rect 20085 7293 20119 7327
rect 20177 7293 20211 7327
rect 26157 7293 26191 7327
rect 26709 7293 26743 7327
rect 27721 7293 27755 7327
rect 28825 7293 28859 7327
rect 29377 7293 29411 7327
rect 33609 7293 33643 7327
rect 11713 7225 11747 7259
rect 14657 7225 14691 7259
rect 16957 7225 16991 7259
rect 17049 7225 17083 7259
rect 20361 7225 20395 7259
rect 28457 7225 28491 7259
rect 11805 7157 11839 7191
rect 12633 7157 12667 7191
rect 12817 7157 12851 7191
rect 13461 7157 13495 7191
rect 16681 7157 16715 7191
rect 20545 7157 20579 7191
rect 22385 7157 22419 7191
rect 26249 7157 26283 7191
rect 27261 7157 27295 7191
rect 15466 6953 15500 6987
rect 21189 6953 21223 6987
rect 21373 6953 21407 6987
rect 22385 6953 22419 6987
rect 22661 6953 22695 6987
rect 23397 6953 23431 6987
rect 26157 6953 26191 6987
rect 27169 6953 27203 6987
rect 32492 6953 32526 6987
rect 33977 6953 34011 6987
rect 24869 6885 24903 6919
rect 25329 6885 25363 6919
rect 26249 6885 26283 6919
rect 28733 6885 28767 6919
rect 29009 6885 29043 6919
rect 13185 6817 13219 6851
rect 13829 6817 13863 6851
rect 15209 6817 15243 6851
rect 17233 6817 17267 6851
rect 22753 6817 22787 6851
rect 25605 6817 25639 6851
rect 26065 6817 26099 6851
rect 29285 6817 29319 6851
rect 29653 6817 29687 6851
rect 30021 6817 30055 6851
rect 30824 6817 30858 6851
rect 31033 6817 31067 6851
rect 31309 6817 31343 6851
rect 32229 6817 32263 6851
rect 11437 6749 11471 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 13737 6749 13771 6783
rect 17601 6749 17635 6783
rect 17785 6749 17819 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 22845 6749 22879 6783
rect 22937 6749 22971 6783
rect 23121 6749 23155 6783
rect 24041 6749 24075 6783
rect 24593 6749 24627 6783
rect 24777 6749 24811 6783
rect 24869 6749 24903 6783
rect 26617 6749 26651 6783
rect 26709 6749 26743 6783
rect 27077 6749 27111 6783
rect 27353 6749 27387 6783
rect 27629 6749 27663 6783
rect 28365 6749 28399 6783
rect 29837 6749 29871 6783
rect 30205 6749 30239 6783
rect 30389 6749 30423 6783
rect 11713 6681 11747 6715
rect 19257 6681 19291 6715
rect 21341 6681 21375 6715
rect 21557 6681 21591 6715
rect 23581 6681 23615 6715
rect 23673 6681 23707 6715
rect 23857 6681 23891 6715
rect 25697 6681 25731 6715
rect 28457 6681 28491 6715
rect 28549 6681 28583 6715
rect 30113 6681 30147 6715
rect 13369 6613 13403 6647
rect 17693 6613 17727 6647
rect 19533 6613 19567 6647
rect 19809 6613 19843 6647
rect 23213 6613 23247 6647
rect 23381 6613 23415 6647
rect 25145 6613 25179 6647
rect 28181 6613 28215 6647
rect 28825 6613 28859 6647
rect 30665 6613 30699 6647
rect 30941 6613 30975 6647
rect 11621 6409 11655 6443
rect 30205 6409 30239 6443
rect 33885 6409 33919 6443
rect 13369 6341 13403 6375
rect 15117 6341 15151 6375
rect 17601 6341 17635 6375
rect 20085 6341 20119 6375
rect 20545 6341 20579 6375
rect 25421 6341 25455 6375
rect 26801 6341 26835 6375
rect 27629 6341 27663 6375
rect 27813 6341 27847 6375
rect 28181 6341 28215 6375
rect 28733 6341 28767 6375
rect 11805 6273 11839 6307
rect 11989 6273 12023 6307
rect 12081 6273 12115 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16037 6273 16071 6307
rect 16129 6273 16163 6307
rect 17049 6273 17083 6307
rect 17325 6273 17359 6307
rect 19625 6273 19659 6307
rect 20177 6273 20211 6307
rect 20361 6273 20395 6307
rect 25237 6273 25271 6307
rect 25789 6273 25823 6307
rect 27445 6273 27479 6307
rect 27997 6273 28031 6307
rect 28457 6273 28491 6307
rect 32137 6273 32171 6307
rect 12173 6205 12207 6239
rect 13093 6205 13127 6239
rect 19349 6205 19383 6239
rect 19717 6205 19751 6239
rect 26065 6205 26099 6239
rect 26433 6205 26467 6239
rect 27077 6205 27111 6239
rect 27169 6205 27203 6239
rect 32413 6205 32447 6239
rect 12817 6069 12851 6103
rect 15577 6069 15611 6103
rect 16773 6069 16807 6103
rect 19441 6069 19475 6103
rect 19625 6069 19659 6103
rect 25697 6069 25731 6103
rect 26525 6069 26559 6103
rect 26663 6069 26697 6103
rect 10412 5865 10446 5899
rect 11989 5865 12023 5899
rect 13093 5865 13127 5899
rect 16957 5865 16991 5899
rect 19441 5865 19475 5899
rect 23765 5865 23799 5899
rect 29561 5865 29595 5899
rect 33885 5865 33919 5899
rect 25329 5797 25363 5831
rect 10149 5729 10183 5763
rect 12449 5729 12483 5763
rect 12541 5729 12575 5763
rect 13277 5729 13311 5763
rect 14565 5729 14599 5763
rect 14749 5729 14783 5763
rect 15485 5729 15519 5763
rect 31309 5729 31343 5763
rect 32137 5729 32171 5763
rect 13185 5661 13219 5695
rect 13829 5661 13863 5695
rect 15209 5661 15243 5695
rect 18429 5661 18463 5695
rect 18705 5661 18739 5695
rect 18889 5661 18923 5695
rect 18981 5661 19015 5695
rect 19257 5661 19291 5695
rect 19901 5661 19935 5695
rect 20545 5661 20579 5695
rect 20637 5661 20671 5695
rect 20913 5661 20947 5695
rect 21189 5661 21223 5695
rect 21281 5661 21315 5695
rect 21741 5661 21775 5695
rect 22017 5661 22051 5695
rect 22109 5661 22143 5695
rect 22661 5661 22695 5695
rect 23029 5661 23063 5695
rect 23305 5661 23339 5695
rect 23397 5661 23431 5695
rect 23949 5661 23983 5695
rect 24685 5661 24719 5695
rect 24869 5661 24903 5695
rect 24961 5661 24995 5695
rect 25053 5661 25087 5695
rect 25513 5661 25547 5695
rect 12357 5593 12391 5627
rect 21097 5593 21131 5627
rect 21925 5593 21959 5627
rect 23213 5593 23247 5627
rect 31033 5593 31067 5627
rect 32413 5593 32447 5627
rect 11897 5525 11931 5559
rect 14105 5525 14139 5559
rect 14473 5525 14507 5559
rect 17785 5525 17819 5559
rect 18521 5525 18555 5559
rect 20729 5525 20763 5559
rect 21465 5525 21499 5559
rect 22293 5525 22327 5559
rect 22477 5525 22511 5559
rect 23581 5525 23615 5559
rect 25237 5525 25271 5559
rect 12265 5321 12299 5355
rect 12633 5321 12667 5355
rect 19533 5321 19567 5355
rect 14105 5253 14139 5287
rect 24317 5253 24351 5287
rect 12173 5185 12207 5219
rect 14381 5185 14415 5219
rect 15209 5185 15243 5219
rect 15761 5185 15795 5219
rect 17233 5185 17267 5219
rect 17417 5185 17451 5219
rect 17509 5185 17543 5219
rect 17693 5185 17727 5219
rect 19625 5185 19659 5219
rect 21833 5185 21867 5219
rect 24133 5185 24167 5219
rect 24409 5185 24443 5219
rect 24501 5185 24535 5219
rect 24869 5185 24903 5219
rect 12357 5117 12391 5151
rect 15301 5117 15335 5151
rect 15393 5117 15427 5151
rect 16313 5117 16347 5151
rect 17325 5117 17359 5151
rect 17785 5117 17819 5151
rect 18061 5117 18095 5151
rect 19901 5117 19935 5151
rect 21649 5117 21683 5151
rect 22109 5117 22143 5151
rect 23857 5117 23891 5151
rect 25145 5117 25179 5151
rect 24685 5049 24719 5083
rect 11805 4981 11839 5015
rect 14841 4981 14875 5015
rect 17049 4981 17083 5015
rect 26617 4981 26651 5015
rect 20085 4777 20119 4811
rect 20361 4777 20395 4811
rect 23857 4777 23891 4811
rect 26801 4777 26835 4811
rect 17969 4709 18003 4743
rect 14381 4641 14415 4675
rect 16221 4641 16255 4675
rect 16497 4641 16531 4675
rect 22109 4641 22143 4675
rect 25053 4641 25087 4675
rect 25329 4641 25363 4675
rect 11253 4573 11287 4607
rect 13369 4573 13403 4607
rect 18705 4573 18739 4607
rect 19257 4573 19291 4607
rect 19901 4573 19935 4607
rect 20269 4573 20303 4607
rect 20545 4573 20579 4607
rect 20729 4573 20763 4607
rect 20913 4573 20947 4607
rect 11529 4505 11563 4539
rect 14657 4505 14691 4539
rect 20637 4505 20671 4539
rect 22385 4505 22419 4539
rect 13001 4437 13035 4471
rect 13921 4437 13955 4471
rect 16129 4437 16163 4471
rect 18153 4437 18187 4471
rect 11989 4233 12023 4267
rect 14933 4233 14967 4267
rect 19901 4233 19935 4267
rect 16037 4165 16071 4199
rect 16681 4165 16715 4199
rect 17509 4165 17543 4199
rect 18061 4165 18095 4199
rect 26985 4165 27019 4199
rect 27169 4165 27203 4199
rect 2053 4097 2087 4131
rect 14473 4097 14507 4131
rect 15025 4097 15059 4131
rect 16129 4097 16163 4131
rect 17417 4097 17451 4131
rect 17693 4097 17727 4131
rect 20177 4097 20211 4131
rect 20269 4097 20303 4131
rect 23305 4097 23339 4131
rect 25145 4097 25179 4131
rect 26801 4097 26835 4131
rect 27353 4097 27387 4131
rect 11345 4029 11379 4063
rect 12633 4029 12667 4063
rect 14197 4029 14231 4063
rect 15209 4029 15243 4063
rect 16221 4029 16255 4063
rect 17325 4029 17359 4063
rect 17785 4029 17819 4063
rect 19809 4029 19843 4063
rect 19901 4029 19935 4063
rect 23581 4029 23615 4063
rect 25053 4029 25087 4063
rect 26433 4029 26467 4063
rect 1869 3961 1903 3995
rect 14565 3961 14599 3995
rect 20085 3961 20119 3995
rect 25513 3961 25547 3995
rect 25881 3961 25915 3995
rect 10701 3893 10735 3927
rect 12725 3893 12759 3927
rect 15669 3893 15703 3927
rect 17693 3893 17727 3927
rect 20361 3893 20395 3927
rect 25605 3893 25639 3927
rect 26709 3893 26743 3927
rect 16957 3689 16991 3723
rect 17785 3689 17819 3723
rect 26157 3689 26191 3723
rect 36001 3689 36035 3723
rect 11161 3553 11195 3587
rect 13185 3553 13219 3587
rect 13829 3553 13863 3587
rect 14565 3553 14599 3587
rect 14749 3553 14783 3587
rect 15209 3553 15243 3587
rect 24409 3553 24443 3587
rect 24685 3553 24719 3587
rect 26801 3553 26835 3587
rect 10977 3485 11011 3519
rect 11069 3485 11103 3519
rect 11437 3485 11471 3519
rect 17601 3485 17635 3519
rect 17969 3485 18003 3519
rect 18061 3485 18095 3519
rect 18153 3485 18187 3519
rect 18705 3485 18739 3519
rect 18889 3485 18923 3519
rect 19257 3485 19291 3519
rect 19441 3485 19475 3519
rect 19625 3485 19659 3519
rect 27353 3485 27387 3519
rect 11713 3417 11747 3451
rect 13277 3417 13311 3451
rect 14473 3417 14507 3451
rect 15485 3417 15519 3451
rect 17785 3417 17819 3451
rect 18981 3417 19015 3451
rect 26985 3417 27019 3451
rect 36093 3417 36127 3451
rect 10609 3349 10643 3383
rect 14105 3349 14139 3383
rect 17049 3349 17083 3383
rect 19717 3349 19751 3383
rect 26249 3349 26283 3383
rect 11897 3145 11931 3179
rect 12265 3145 12299 3179
rect 24409 3145 24443 3179
rect 9873 3077 9907 3111
rect 13185 3077 13219 3111
rect 17141 3077 17175 3111
rect 25881 3077 25915 3111
rect 9597 3009 9631 3043
rect 12357 3009 12391 3043
rect 12909 3009 12943 3043
rect 14749 3009 14783 3043
rect 16865 3009 16899 3043
rect 18705 3009 18739 3043
rect 23949 3009 23983 3043
rect 24041 3009 24075 3043
rect 26157 3009 26191 3043
rect 11345 2941 11379 2975
rect 12449 2941 12483 2975
rect 15025 2941 15059 2975
rect 16497 2941 16531 2975
rect 18981 2941 19015 2975
rect 20453 2941 20487 2975
rect 14657 2805 14691 2839
rect 18613 2805 18647 2839
rect 23765 2805 23799 2839
rect 14657 2601 14691 2635
rect 18705 2601 18739 2635
rect 19257 2601 19291 2635
rect 18429 2533 18463 2567
rect 15209 2465 15243 2499
rect 16681 2465 16715 2499
rect 16957 2465 16991 2499
rect 19809 2465 19843 2499
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 13001 2397 13035 2431
rect 13645 2397 13679 2431
rect 14289 2397 14323 2431
rect 15577 2397 15611 2431
rect 16221 2397 16255 2431
rect 18521 2397 18555 2431
rect 24685 2397 24719 2431
rect 24869 2397 24903 2431
rect 25237 2397 25271 2431
rect 24777 2329 24811 2363
rect 11805 2261 11839 2295
rect 12541 2261 12575 2295
rect 13185 2261 13219 2295
rect 13829 2261 13863 2295
rect 14473 2261 14507 2295
rect 15761 2261 15795 2295
rect 16405 2261 16439 2295
rect 25421 2261 25455 2295
<< metal1 >>
rect 1104 37562 36524 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 36524 37562
rect 1104 37488 36524 37510
rect 22278 37380 22284 37392
rect 12820 37352 22284 37380
rect 7009 37315 7067 37321
rect 7009 37281 7021 37315
rect 7055 37312 7067 37315
rect 7558 37312 7564 37324
rect 7055 37284 7564 37312
rect 7055 37281 7067 37284
rect 7009 37275 7067 37281
rect 7558 37272 7564 37284
rect 7616 37312 7622 37324
rect 8113 37315 8171 37321
rect 8113 37312 8125 37315
rect 7616 37284 8125 37312
rect 7616 37272 7622 37284
rect 8113 37281 8125 37284
rect 8159 37312 8171 37315
rect 9582 37312 9588 37324
rect 8159 37284 9588 37312
rect 8159 37281 8171 37284
rect 8113 37275 8171 37281
rect 9582 37272 9588 37284
rect 9640 37312 9646 37324
rect 12820 37321 12848 37352
rect 22278 37340 22284 37352
rect 22336 37340 22342 37392
rect 10229 37315 10287 37321
rect 10229 37312 10241 37315
rect 9640 37284 10241 37312
rect 9640 37272 9646 37284
rect 10229 37281 10241 37284
rect 10275 37312 10287 37315
rect 11241 37315 11299 37321
rect 11241 37312 11253 37315
rect 10275 37284 11253 37312
rect 10275 37281 10287 37284
rect 10229 37275 10287 37281
rect 11241 37281 11253 37284
rect 11287 37312 11299 37315
rect 12805 37315 12863 37321
rect 12805 37312 12817 37315
rect 11287 37284 12817 37312
rect 11287 37281 11299 37284
rect 11241 37275 11299 37281
rect 12805 37281 12817 37284
rect 12851 37281 12863 37315
rect 12805 37275 12863 37281
rect 17218 37272 17224 37324
rect 17276 37272 17282 37324
rect 17497 37315 17555 37321
rect 17497 37281 17509 37315
rect 17543 37312 17555 37315
rect 18138 37312 18144 37324
rect 17543 37284 18144 37312
rect 17543 37281 17555 37284
rect 17497 37275 17555 37281
rect 18138 37272 18144 37284
rect 18196 37272 18202 37324
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 5868 37216 6837 37244
rect 5868 37204 5874 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 6825 37207 6883 37213
rect 7929 37247 7987 37253
rect 7929 37213 7941 37247
rect 7975 37244 7987 37247
rect 8386 37244 8392 37256
rect 7975 37216 8392 37244
rect 7975 37213 7987 37216
rect 7929 37207 7987 37213
rect 8386 37204 8392 37216
rect 8444 37204 8450 37256
rect 10045 37247 10103 37253
rect 8956 37216 9674 37244
rect 6733 37179 6791 37185
rect 6733 37145 6745 37179
rect 6779 37176 6791 37179
rect 8294 37176 8300 37188
rect 6779 37148 8300 37176
rect 6779 37145 6791 37148
rect 6733 37139 6791 37145
rect 8294 37136 8300 37148
rect 8352 37136 8358 37188
rect 4430 37068 4436 37120
rect 4488 37108 4494 37120
rect 6365 37111 6423 37117
rect 6365 37108 6377 37111
rect 4488 37080 6377 37108
rect 4488 37068 4494 37080
rect 6365 37077 6377 37080
rect 6411 37077 6423 37111
rect 6365 37071 6423 37077
rect 7466 37068 7472 37120
rect 7524 37068 7530 37120
rect 7837 37111 7895 37117
rect 7837 37077 7849 37111
rect 7883 37108 7895 37111
rect 8956 37108 8984 37216
rect 9646 37176 9674 37216
rect 10045 37213 10057 37247
rect 10091 37244 10103 37247
rect 10962 37244 10968 37256
rect 10091 37216 10968 37244
rect 10091 37213 10103 37216
rect 10045 37207 10103 37213
rect 10962 37204 10968 37216
rect 11020 37204 11026 37256
rect 11057 37247 11115 37253
rect 11057 37213 11069 37247
rect 11103 37244 11115 37247
rect 11606 37244 11612 37256
rect 11103 37216 11612 37244
rect 11103 37213 11115 37216
rect 11057 37207 11115 37213
rect 11606 37204 11612 37216
rect 11664 37204 11670 37256
rect 12250 37204 12256 37256
rect 12308 37244 12314 37256
rect 12621 37247 12679 37253
rect 12621 37244 12633 37247
rect 12308 37216 12633 37244
rect 12308 37204 12314 37216
rect 12621 37213 12633 37216
rect 12667 37213 12679 37247
rect 12621 37207 12679 37213
rect 17034 37204 17040 37256
rect 17092 37244 17098 37256
rect 17129 37247 17187 37253
rect 17129 37244 17141 37247
rect 17092 37216 17141 37244
rect 17092 37204 17098 37216
rect 17129 37213 17141 37216
rect 17175 37213 17187 37247
rect 17129 37207 17187 37213
rect 10778 37176 10784 37188
rect 9646 37148 10784 37176
rect 10778 37136 10784 37148
rect 10836 37136 10842 37188
rect 7883 37080 8984 37108
rect 7883 37077 7895 37080
rect 7837 37071 7895 37077
rect 9030 37068 9036 37120
rect 9088 37108 9094 37120
rect 9585 37111 9643 37117
rect 9585 37108 9597 37111
rect 9088 37080 9597 37108
rect 9088 37068 9094 37080
rect 9585 37077 9597 37080
rect 9631 37077 9643 37111
rect 9585 37071 9643 37077
rect 9953 37111 10011 37117
rect 9953 37077 9965 37111
rect 9999 37108 10011 37111
rect 10042 37108 10048 37120
rect 9999 37080 10048 37108
rect 9999 37077 10011 37080
rect 9953 37071 10011 37077
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 10594 37068 10600 37120
rect 10652 37068 10658 37120
rect 10870 37068 10876 37120
rect 10928 37108 10934 37120
rect 10965 37111 11023 37117
rect 10965 37108 10977 37111
rect 10928 37080 10977 37108
rect 10928 37068 10934 37080
rect 10965 37077 10977 37080
rect 11011 37077 11023 37111
rect 10965 37071 11023 37077
rect 11882 37068 11888 37120
rect 11940 37108 11946 37120
rect 12161 37111 12219 37117
rect 12161 37108 12173 37111
rect 11940 37080 12173 37108
rect 11940 37068 11946 37080
rect 12161 37077 12173 37080
rect 12207 37077 12219 37111
rect 12161 37071 12219 37077
rect 12342 37068 12348 37120
rect 12400 37108 12406 37120
rect 12529 37111 12587 37117
rect 12529 37108 12541 37111
rect 12400 37080 12541 37108
rect 12400 37068 12406 37080
rect 12529 37077 12541 37080
rect 12575 37077 12587 37111
rect 12529 37071 12587 37077
rect 1104 37018 36524 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 36524 37018
rect 1104 36944 36524 36966
rect 9674 36904 9680 36916
rect 8680 36876 9680 36904
rect 4430 36796 4436 36848
rect 4488 36796 4494 36848
rect 7374 36836 7380 36848
rect 5658 36808 7380 36836
rect 7374 36796 7380 36808
rect 7432 36796 7438 36848
rect 8680 36845 8708 36876
rect 9674 36864 9680 36876
rect 9732 36864 9738 36916
rect 13814 36904 13820 36916
rect 12268 36876 13820 36904
rect 8665 36839 8723 36845
rect 8665 36805 8677 36839
rect 8711 36805 8723 36839
rect 10781 36839 10839 36845
rect 8665 36799 8723 36805
rect 8772 36808 9522 36836
rect 5810 36728 5816 36780
rect 5868 36768 5874 36780
rect 6181 36771 6239 36777
rect 6181 36768 6193 36771
rect 5868 36740 6193 36768
rect 5868 36728 5874 36740
rect 6181 36737 6193 36740
rect 6227 36737 6239 36771
rect 6181 36731 6239 36737
rect 8018 36728 8024 36780
rect 8076 36768 8082 36780
rect 8772 36768 8800 36808
rect 10781 36805 10793 36839
rect 10827 36836 10839 36839
rect 10962 36836 10968 36848
rect 10827 36808 10968 36836
rect 10827 36805 10839 36808
rect 10781 36799 10839 36805
rect 10962 36796 10968 36808
rect 11020 36796 11026 36848
rect 11882 36796 11888 36848
rect 11940 36796 11946 36848
rect 12158 36796 12164 36848
rect 12216 36836 12222 36848
rect 12268 36836 12296 36876
rect 13814 36864 13820 36876
rect 13872 36904 13878 36916
rect 26602 36904 26608 36916
rect 13872 36876 14320 36904
rect 13872 36864 13878 36876
rect 14292 36836 14320 36876
rect 20272 36876 22094 36904
rect 14734 36836 14740 36848
rect 12216 36808 12374 36836
rect 14292 36808 14740 36836
rect 12216 36796 12222 36808
rect 14734 36796 14740 36808
rect 14792 36796 14798 36848
rect 16942 36796 16948 36848
rect 17000 36836 17006 36848
rect 19886 36836 19892 36848
rect 17000 36808 19892 36836
rect 17000 36796 17006 36808
rect 8076 36740 8800 36768
rect 8076 36728 8082 36740
rect 17402 36728 17408 36780
rect 17460 36728 17466 36780
rect 18138 36728 18144 36780
rect 18196 36728 18202 36780
rect 18708 36777 18736 36808
rect 19886 36796 19892 36808
rect 19944 36836 19950 36848
rect 20162 36836 20168 36848
rect 19944 36808 20168 36836
rect 19944 36796 19950 36808
rect 20162 36796 20168 36808
rect 20220 36796 20226 36848
rect 20272 36836 20300 36876
rect 20346 36836 20352 36848
rect 20272 36808 20352 36836
rect 20346 36796 20352 36808
rect 20404 36796 20410 36848
rect 22066 36836 22094 36876
rect 23492 36876 25360 36904
rect 23492 36836 23520 36876
rect 25332 36836 25360 36876
rect 25608 36876 26608 36904
rect 25608 36836 25636 36876
rect 26602 36864 26608 36876
rect 26660 36864 26666 36916
rect 22066 36808 23598 36836
rect 25332 36808 25714 36836
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36737 18751 36771
rect 18693 36731 18751 36737
rect 19153 36771 19211 36777
rect 19153 36737 19165 36771
rect 19199 36768 19211 36771
rect 19518 36768 19524 36780
rect 19199 36740 19524 36768
rect 19199 36737 19211 36740
rect 19153 36731 19211 36737
rect 19518 36728 19524 36740
rect 19576 36728 19582 36780
rect 4157 36703 4215 36709
rect 4157 36669 4169 36703
rect 4203 36669 4215 36703
rect 4157 36663 4215 36669
rect 6641 36703 6699 36709
rect 6641 36669 6653 36703
rect 6687 36669 6699 36703
rect 6641 36663 6699 36669
rect 4172 36564 4200 36663
rect 5534 36564 5540 36576
rect 4172 36536 5540 36564
rect 5534 36524 5540 36536
rect 5592 36564 5598 36576
rect 6454 36564 6460 36576
rect 5592 36536 6460 36564
rect 5592 36524 5598 36536
rect 6454 36524 6460 36536
rect 6512 36564 6518 36576
rect 6656 36564 6684 36663
rect 6914 36660 6920 36712
rect 6972 36660 6978 36712
rect 8754 36660 8760 36712
rect 8812 36660 8818 36712
rect 9030 36660 9036 36712
rect 9088 36660 9094 36712
rect 10686 36660 10692 36712
rect 10744 36700 10750 36712
rect 11609 36703 11667 36709
rect 11609 36700 11621 36703
rect 10744 36672 11621 36700
rect 10744 36660 10750 36672
rect 11609 36669 11621 36672
rect 11655 36669 11667 36703
rect 11609 36663 11667 36669
rect 6512 36536 6684 36564
rect 6512 36524 6518 36536
rect 8294 36524 8300 36576
rect 8352 36564 8358 36576
rect 9214 36564 9220 36576
rect 8352 36536 9220 36564
rect 8352 36524 8358 36536
rect 9214 36524 9220 36536
rect 9272 36524 9278 36576
rect 11624 36564 11652 36663
rect 12250 36660 12256 36712
rect 12308 36700 12314 36712
rect 13633 36703 13691 36709
rect 13633 36700 13645 36703
rect 12308 36672 13645 36700
rect 12308 36660 12314 36672
rect 13633 36669 13645 36672
rect 13679 36669 13691 36703
rect 13633 36663 13691 36669
rect 14001 36703 14059 36709
rect 14001 36669 14013 36703
rect 14047 36669 14059 36703
rect 14001 36663 14059 36669
rect 14016 36576 14044 36663
rect 14274 36660 14280 36712
rect 14332 36660 14338 36712
rect 15010 36660 15016 36712
rect 15068 36700 15074 36712
rect 15749 36703 15807 36709
rect 15749 36700 15761 36703
rect 15068 36672 15761 36700
rect 15068 36660 15074 36672
rect 15749 36669 15761 36672
rect 15795 36700 15807 36703
rect 17034 36700 17040 36712
rect 15795 36672 17040 36700
rect 15795 36669 15807 36672
rect 15749 36663 15807 36669
rect 17034 36660 17040 36672
rect 17092 36660 17098 36712
rect 17494 36660 17500 36712
rect 17552 36660 17558 36712
rect 18230 36660 18236 36712
rect 18288 36660 18294 36712
rect 19334 36660 19340 36712
rect 19392 36700 19398 36712
rect 19429 36703 19487 36709
rect 19429 36700 19441 36703
rect 19392 36672 19441 36700
rect 19392 36660 19398 36672
rect 19429 36669 19441 36672
rect 19475 36669 19487 36703
rect 19429 36663 19487 36669
rect 19613 36703 19671 36709
rect 19613 36669 19625 36703
rect 19659 36669 19671 36703
rect 19613 36663 19671 36669
rect 19889 36703 19947 36709
rect 19889 36669 19901 36703
rect 19935 36700 19947 36703
rect 19978 36700 19984 36712
rect 19935 36672 19984 36700
rect 19935 36669 19947 36672
rect 19889 36663 19947 36669
rect 17773 36635 17831 36641
rect 17773 36632 17785 36635
rect 15304 36604 17785 36632
rect 13998 36564 14004 36576
rect 11624 36536 14004 36564
rect 13998 36524 14004 36536
rect 14056 36524 14062 36576
rect 14642 36524 14648 36576
rect 14700 36564 14706 36576
rect 15304 36564 15332 36604
rect 17773 36601 17785 36604
rect 17819 36601 17831 36635
rect 17773 36595 17831 36601
rect 14700 36536 15332 36564
rect 14700 36524 14706 36536
rect 16574 36524 16580 36576
rect 16632 36564 16638 36576
rect 17037 36567 17095 36573
rect 17037 36564 17049 36567
rect 16632 36536 17049 36564
rect 16632 36524 16638 36536
rect 17037 36533 17049 36536
rect 17083 36533 17095 36567
rect 19628 36564 19656 36663
rect 19978 36660 19984 36672
rect 20036 36660 20042 36712
rect 20254 36660 20260 36712
rect 20312 36700 20318 36712
rect 21637 36703 21695 36709
rect 21637 36700 21649 36703
rect 20312 36672 21649 36700
rect 20312 36660 20318 36672
rect 21637 36669 21649 36672
rect 21683 36669 21695 36703
rect 21637 36663 21695 36669
rect 22833 36703 22891 36709
rect 22833 36669 22845 36703
rect 22879 36669 22891 36703
rect 22833 36663 22891 36669
rect 23109 36703 23167 36709
rect 23109 36669 23121 36703
rect 23155 36700 23167 36703
rect 23198 36700 23204 36712
rect 23155 36672 23204 36700
rect 23155 36669 23167 36672
rect 23109 36663 23167 36669
rect 22848 36564 22876 36663
rect 23198 36660 23204 36672
rect 23256 36660 23262 36712
rect 24578 36660 24584 36712
rect 24636 36700 24642 36712
rect 24857 36703 24915 36709
rect 24857 36700 24869 36703
rect 24636 36672 24869 36700
rect 24636 36660 24642 36672
rect 24857 36669 24869 36672
rect 24903 36669 24915 36703
rect 24857 36663 24915 36669
rect 24946 36660 24952 36712
rect 25004 36660 25010 36712
rect 25222 36660 25228 36712
rect 25280 36660 25286 36712
rect 23106 36564 23112 36576
rect 19628 36536 23112 36564
rect 17037 36527 17095 36533
rect 23106 36524 23112 36536
rect 23164 36524 23170 36576
rect 25958 36524 25964 36576
rect 26016 36564 26022 36576
rect 26697 36567 26755 36573
rect 26697 36564 26709 36567
rect 26016 36536 26709 36564
rect 26016 36524 26022 36536
rect 26697 36533 26709 36536
rect 26743 36533 26755 36567
rect 26697 36527 26755 36533
rect 1104 36474 36524 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 36524 36474
rect 1104 36400 36524 36422
rect 6914 36320 6920 36372
rect 6972 36360 6978 36372
rect 8941 36363 8999 36369
rect 8941 36360 8953 36363
rect 6972 36332 8953 36360
rect 6972 36320 6978 36332
rect 8941 36329 8953 36332
rect 8987 36329 8999 36363
rect 13446 36360 13452 36372
rect 8941 36323 8999 36329
rect 13188 36332 13452 36360
rect 8754 36252 8760 36304
rect 8812 36292 8818 36304
rect 8812 36264 10364 36292
rect 8812 36252 8818 36264
rect 6454 36184 6460 36236
rect 6512 36184 6518 36236
rect 6733 36227 6791 36233
rect 6733 36193 6745 36227
rect 6779 36224 6791 36227
rect 7466 36224 7472 36236
rect 6779 36196 7472 36224
rect 6779 36193 6791 36196
rect 6733 36187 6791 36193
rect 7466 36184 7472 36196
rect 7524 36184 7530 36236
rect 8386 36184 8392 36236
rect 8444 36224 8450 36236
rect 8481 36227 8539 36233
rect 8481 36224 8493 36227
rect 8444 36196 8493 36224
rect 8444 36184 8450 36196
rect 8481 36193 8493 36196
rect 8527 36193 8539 36227
rect 8481 36187 8539 36193
rect 9582 36184 9588 36236
rect 9640 36184 9646 36236
rect 9401 36159 9459 36165
rect 9401 36125 9413 36159
rect 9447 36156 9459 36159
rect 9674 36156 9680 36168
rect 9447 36128 9680 36156
rect 9447 36125 9459 36128
rect 9401 36119 9459 36125
rect 9674 36116 9680 36128
rect 9732 36116 9738 36168
rect 10336 36165 10364 36264
rect 11698 36252 11704 36304
rect 11756 36292 11762 36304
rect 11756 36264 12388 36292
rect 11756 36252 11762 36264
rect 10594 36184 10600 36236
rect 10652 36184 10658 36236
rect 12360 36233 12388 36264
rect 13188 36233 13216 36332
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 14734 36320 14740 36372
rect 14792 36360 14798 36372
rect 14792 36332 16436 36360
rect 14792 36320 14798 36332
rect 13262 36252 13268 36304
rect 13320 36252 13326 36304
rect 13998 36252 14004 36304
rect 14056 36292 14062 36304
rect 14056 36264 15148 36292
rect 14056 36252 14062 36264
rect 12345 36227 12403 36233
rect 12345 36193 12357 36227
rect 12391 36193 12403 36227
rect 12345 36187 12403 36193
rect 13173 36227 13231 36233
rect 13173 36193 13185 36227
rect 13219 36193 13231 36227
rect 13280 36224 13308 36252
rect 13280 36196 14872 36224
rect 13173 36187 13231 36193
rect 10321 36159 10379 36165
rect 10321 36125 10333 36159
rect 10367 36125 10379 36159
rect 12158 36156 12164 36168
rect 11730 36128 12164 36156
rect 10321 36119 10379 36125
rect 8018 36088 8024 36100
rect 7958 36060 8024 36088
rect 8018 36048 8024 36060
rect 8076 36048 8082 36100
rect 9309 36091 9367 36097
rect 9309 36057 9321 36091
rect 9355 36088 9367 36091
rect 9766 36088 9772 36100
rect 9355 36060 9772 36088
rect 9355 36057 9367 36060
rect 9309 36051 9367 36057
rect 9766 36048 9772 36060
rect 9824 36048 9830 36100
rect 10336 36088 10364 36119
rect 12158 36116 12164 36128
rect 12216 36116 12222 36168
rect 12618 36116 12624 36168
rect 12676 36156 12682 36168
rect 13265 36159 13323 36165
rect 13265 36156 13277 36159
rect 12676 36128 13277 36156
rect 12676 36116 12682 36128
rect 13265 36125 13277 36128
rect 13311 36125 13323 36159
rect 13265 36119 13323 36125
rect 14642 36116 14648 36168
rect 14700 36116 14706 36168
rect 14734 36116 14740 36168
rect 14792 36116 14798 36168
rect 14844 36156 14872 36196
rect 14918 36184 14924 36236
rect 14976 36184 14982 36236
rect 15120 36233 15148 36264
rect 15105 36227 15163 36233
rect 15105 36193 15117 36227
rect 15151 36193 15163 36227
rect 15105 36187 15163 36193
rect 15010 36156 15016 36168
rect 14844 36128 15016 36156
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 16408 36156 16436 36332
rect 17494 36320 17500 36372
rect 17552 36360 17558 36372
rect 18141 36363 18199 36369
rect 18141 36360 18153 36363
rect 17552 36332 18153 36360
rect 17552 36320 17558 36332
rect 18141 36329 18153 36332
rect 18187 36329 18199 36363
rect 18141 36323 18199 36329
rect 19978 36320 19984 36372
rect 20036 36320 20042 36372
rect 25133 36363 25191 36369
rect 22066 36332 25084 36360
rect 18230 36292 18236 36304
rect 17972 36264 18236 36292
rect 17972 36233 18000 36264
rect 18230 36252 18236 36264
rect 18288 36292 18294 36304
rect 19429 36295 19487 36301
rect 19429 36292 19441 36295
rect 18288 36264 19441 36292
rect 18288 36252 18294 36264
rect 19429 36261 19441 36264
rect 19475 36261 19487 36295
rect 19705 36295 19763 36301
rect 19705 36292 19717 36295
rect 19429 36255 19487 36261
rect 19536 36264 19717 36292
rect 19536 36233 19564 36264
rect 19705 36261 19717 36264
rect 19751 36261 19763 36295
rect 19705 36255 19763 36261
rect 17957 36227 18015 36233
rect 17957 36193 17969 36227
rect 18003 36193 18015 36227
rect 17957 36187 18015 36193
rect 19521 36227 19579 36233
rect 19521 36193 19533 36227
rect 19567 36193 19579 36227
rect 19521 36187 19579 36193
rect 19610 36184 19616 36236
rect 19668 36184 19674 36236
rect 20625 36227 20683 36233
rect 20625 36224 20637 36227
rect 19996 36196 20637 36224
rect 16482 36156 16488 36168
rect 16408 36128 16488 36156
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 17034 36116 17040 36168
rect 17092 36156 17098 36168
rect 17129 36159 17187 36165
rect 17129 36156 17141 36159
rect 17092 36128 17141 36156
rect 17092 36116 17098 36128
rect 17129 36125 17141 36128
rect 17175 36125 17187 36159
rect 17129 36119 17187 36125
rect 17310 36116 17316 36168
rect 17368 36116 17374 36168
rect 17865 36159 17923 36165
rect 17865 36125 17877 36159
rect 17911 36156 17923 36159
rect 18138 36156 18144 36168
rect 17911 36128 18144 36156
rect 17911 36125 17923 36128
rect 17865 36119 17923 36125
rect 18138 36116 18144 36128
rect 18196 36116 18202 36168
rect 19242 36116 19248 36168
rect 19300 36116 19306 36168
rect 19334 36116 19340 36168
rect 19392 36116 19398 36168
rect 19702 36116 19708 36168
rect 19760 36156 19766 36168
rect 19797 36159 19855 36165
rect 19797 36156 19809 36159
rect 19760 36128 19809 36156
rect 19760 36116 19766 36128
rect 19797 36125 19809 36128
rect 19843 36125 19855 36159
rect 19797 36119 19855 36125
rect 19886 36116 19892 36168
rect 19944 36116 19950 36168
rect 10594 36088 10600 36100
rect 10336 36060 10600 36088
rect 10594 36048 10600 36060
rect 10652 36048 10658 36100
rect 15286 36088 15292 36100
rect 13648 36060 15292 36088
rect 7374 35980 7380 36032
rect 7432 36020 7438 36032
rect 8036 36020 8064 36048
rect 13648 36029 13676 36060
rect 15286 36048 15292 36060
rect 15344 36048 15350 36100
rect 15378 36048 15384 36100
rect 15436 36048 15442 36100
rect 16758 36048 16764 36100
rect 16816 36088 16822 36100
rect 19996 36088 20024 36196
rect 20625 36193 20637 36196
rect 20671 36224 20683 36227
rect 20990 36224 20996 36236
rect 20671 36196 20996 36224
rect 20671 36193 20683 36196
rect 20625 36187 20683 36193
rect 20990 36184 20996 36196
rect 21048 36224 21054 36236
rect 22066 36224 22094 36332
rect 21048 36196 22094 36224
rect 21048 36184 21054 36196
rect 23106 36184 23112 36236
rect 23164 36224 23170 36236
rect 23385 36227 23443 36233
rect 23385 36224 23397 36227
rect 23164 36196 23397 36224
rect 23164 36184 23170 36196
rect 23385 36193 23397 36196
rect 23431 36224 23443 36227
rect 24946 36224 24952 36236
rect 23431 36196 24952 36224
rect 23431 36193 23443 36196
rect 23385 36187 23443 36193
rect 24946 36184 24952 36196
rect 25004 36184 25010 36236
rect 25056 36224 25084 36332
rect 25133 36329 25145 36363
rect 25179 36360 25191 36363
rect 25222 36360 25228 36372
rect 25179 36332 25228 36360
rect 25179 36329 25191 36332
rect 25133 36323 25191 36329
rect 25222 36320 25228 36332
rect 25280 36320 25286 36372
rect 25682 36224 25688 36236
rect 25056 36196 25688 36224
rect 25682 36184 25688 36196
rect 25740 36184 25746 36236
rect 25958 36184 25964 36236
rect 26016 36224 26022 36236
rect 26016 36196 26556 36224
rect 26016 36184 26022 36196
rect 20346 36116 20352 36168
rect 20404 36156 20410 36168
rect 24029 36159 24087 36165
rect 20404 36128 22034 36156
rect 20404 36116 20410 36128
rect 24029 36125 24041 36159
rect 24075 36125 24087 36159
rect 24029 36119 24087 36125
rect 16816 36060 20024 36088
rect 16816 36048 16822 36060
rect 23106 36048 23112 36100
rect 23164 36048 23170 36100
rect 24044 36088 24072 36119
rect 24210 36116 24216 36168
rect 24268 36156 24274 36168
rect 24578 36156 24584 36168
rect 24268 36128 24584 36156
rect 24268 36116 24274 36128
rect 24578 36116 24584 36128
rect 24636 36116 24642 36168
rect 25498 36116 25504 36168
rect 25556 36156 25562 36168
rect 25593 36159 25651 36165
rect 25593 36156 25605 36159
rect 25556 36128 25605 36156
rect 25556 36116 25562 36128
rect 25593 36125 25605 36128
rect 25639 36125 25651 36159
rect 25593 36119 25651 36125
rect 24118 36088 24124 36100
rect 24044 36060 24124 36088
rect 24118 36048 24124 36060
rect 24176 36088 24182 36100
rect 24397 36091 24455 36097
rect 24397 36088 24409 36091
rect 24176 36060 24409 36088
rect 24176 36048 24182 36060
rect 24397 36057 24409 36060
rect 24443 36057 24455 36091
rect 25976 36088 26004 36184
rect 26053 36159 26111 36165
rect 26053 36125 26065 36159
rect 26099 36125 26111 36159
rect 26053 36119 26111 36125
rect 24397 36051 24455 36057
rect 25516 36060 26004 36088
rect 26068 36088 26096 36119
rect 26234 36116 26240 36168
rect 26292 36116 26298 36168
rect 26326 36116 26332 36168
rect 26384 36116 26390 36168
rect 26528 36165 26556 36196
rect 26513 36159 26571 36165
rect 26513 36125 26525 36159
rect 26559 36125 26571 36159
rect 26513 36119 26571 36125
rect 26421 36091 26479 36097
rect 26421 36088 26433 36091
rect 26068 36060 26433 36088
rect 7432 35992 8064 36020
rect 13633 36023 13691 36029
rect 7432 35980 7438 35992
rect 13633 35989 13645 36023
rect 13679 35989 13691 36023
rect 13633 35983 13691 35989
rect 14366 35980 14372 36032
rect 14424 36020 14430 36032
rect 14461 36023 14519 36029
rect 14461 36020 14473 36023
rect 14424 35992 14473 36020
rect 14424 35980 14430 35992
rect 14461 35989 14473 35992
rect 14507 35989 14519 36023
rect 14461 35983 14519 35989
rect 16850 35980 16856 36032
rect 16908 35980 16914 36032
rect 17221 36023 17279 36029
rect 17221 35989 17233 36023
rect 17267 36020 17279 36023
rect 17497 36023 17555 36029
rect 17497 36020 17509 36023
rect 17267 35992 17509 36020
rect 17267 35989 17279 35992
rect 17221 35983 17279 35989
rect 17497 35989 17509 35992
rect 17543 35989 17555 36023
rect 17497 35983 17555 35989
rect 19886 35980 19892 36032
rect 19944 36020 19950 36032
rect 20349 36023 20407 36029
rect 20349 36020 20361 36023
rect 19944 35992 20361 36020
rect 19944 35980 19950 35992
rect 20349 35989 20361 35992
rect 20395 35989 20407 36023
rect 20349 35983 20407 35989
rect 20438 35980 20444 36032
rect 20496 35980 20502 36032
rect 21637 36023 21695 36029
rect 21637 35989 21649 36023
rect 21683 36020 21695 36023
rect 22094 36020 22100 36032
rect 21683 35992 22100 36020
rect 21683 35989 21695 35992
rect 21637 35983 21695 35989
rect 22094 35980 22100 35992
rect 22152 35980 22158 36032
rect 24213 36023 24271 36029
rect 24213 35989 24225 36023
rect 24259 36020 24271 36023
rect 24670 36020 24676 36032
rect 24259 35992 24676 36020
rect 24259 35989 24271 35992
rect 24213 35983 24271 35989
rect 24670 35980 24676 35992
rect 24728 35980 24734 36032
rect 24765 36023 24823 36029
rect 24765 35989 24777 36023
rect 24811 36020 24823 36023
rect 24854 36020 24860 36032
rect 24811 35992 24860 36020
rect 24811 35989 24823 35992
rect 24765 35983 24823 35989
rect 24854 35980 24860 35992
rect 24912 35980 24918 36032
rect 25314 35980 25320 36032
rect 25372 36020 25378 36032
rect 25516 36029 25544 36060
rect 26421 36057 26433 36060
rect 26467 36057 26479 36091
rect 26421 36051 26479 36057
rect 25501 36023 25559 36029
rect 25501 36020 25513 36023
rect 25372 35992 25513 36020
rect 25372 35980 25378 35992
rect 25501 35989 25513 35992
rect 25547 35989 25559 36023
rect 25501 35983 25559 35989
rect 26142 35980 26148 36032
rect 26200 35980 26206 36032
rect 1104 35930 36524 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 36524 35930
rect 1104 35856 36524 35878
rect 7374 35776 7380 35828
rect 7432 35816 7438 35828
rect 9585 35819 9643 35825
rect 7432 35788 7972 35816
rect 7432 35776 7438 35788
rect 7944 35760 7972 35788
rect 9585 35785 9597 35819
rect 9631 35816 9643 35819
rect 12894 35816 12900 35828
rect 9631 35788 12900 35816
rect 9631 35785 9643 35788
rect 9585 35779 9643 35785
rect 12894 35776 12900 35788
rect 12952 35776 12958 35828
rect 12989 35819 13047 35825
rect 12989 35785 13001 35819
rect 13035 35816 13047 35819
rect 13035 35788 13124 35816
rect 13035 35785 13047 35788
rect 12989 35779 13047 35785
rect 7926 35748 7932 35760
rect 7866 35720 7932 35748
rect 7926 35708 7932 35720
rect 7984 35708 7990 35760
rect 13096 35748 13124 35788
rect 13170 35776 13176 35828
rect 13228 35816 13234 35828
rect 13725 35819 13783 35825
rect 13725 35816 13737 35819
rect 13228 35788 13737 35816
rect 13228 35776 13234 35788
rect 13725 35785 13737 35788
rect 13771 35816 13783 35819
rect 15013 35819 15071 35825
rect 13771 35788 14504 35816
rect 13771 35785 13783 35788
rect 13725 35779 13783 35785
rect 13630 35748 13636 35760
rect 13096 35720 13636 35748
rect 13630 35708 13636 35720
rect 13688 35748 13694 35760
rect 13688 35720 14412 35748
rect 13688 35708 13694 35720
rect 9214 35640 9220 35692
rect 9272 35680 9278 35692
rect 9490 35680 9496 35692
rect 9272 35652 9496 35680
rect 9272 35640 9278 35652
rect 9490 35640 9496 35652
rect 9548 35640 9554 35692
rect 9766 35640 9772 35692
rect 9824 35680 9830 35692
rect 9861 35683 9919 35689
rect 9861 35680 9873 35683
rect 9824 35652 9873 35680
rect 9824 35640 9830 35652
rect 9861 35649 9873 35652
rect 9907 35649 9919 35683
rect 9861 35643 9919 35649
rect 12158 35640 12164 35692
rect 12216 35680 12222 35692
rect 12437 35683 12495 35689
rect 12437 35680 12449 35683
rect 12216 35652 12449 35680
rect 12216 35640 12222 35652
rect 12437 35649 12449 35652
rect 12483 35649 12495 35683
rect 12437 35643 12495 35649
rect 12526 35640 12532 35692
rect 12584 35680 12590 35692
rect 12621 35683 12679 35689
rect 12621 35680 12633 35683
rect 12584 35652 12633 35680
rect 12584 35640 12590 35652
rect 12621 35649 12633 35652
rect 12667 35649 12679 35683
rect 12621 35643 12679 35649
rect 12711 35683 12769 35689
rect 12711 35649 12723 35683
rect 12757 35649 12769 35683
rect 12711 35643 12769 35649
rect 12897 35683 12955 35689
rect 12897 35649 12909 35683
rect 12943 35680 12955 35683
rect 12986 35680 12992 35692
rect 12943 35652 12992 35680
rect 12943 35649 12955 35652
rect 12897 35643 12955 35649
rect 5534 35572 5540 35624
rect 5592 35612 5598 35624
rect 6365 35615 6423 35621
rect 6365 35612 6377 35615
rect 5592 35584 6377 35612
rect 5592 35572 5598 35584
rect 6365 35581 6377 35584
rect 6411 35581 6423 35615
rect 6365 35575 6423 35581
rect 6641 35615 6699 35621
rect 6641 35581 6653 35615
rect 6687 35612 6699 35615
rect 7006 35612 7012 35624
rect 6687 35584 7012 35612
rect 6687 35581 6699 35584
rect 6641 35575 6699 35581
rect 7006 35572 7012 35584
rect 7064 35572 7070 35624
rect 7098 35572 7104 35624
rect 7156 35612 7162 35624
rect 8389 35615 8447 35621
rect 8389 35612 8401 35615
rect 7156 35584 8401 35612
rect 7156 35572 7162 35584
rect 8389 35581 8401 35584
rect 8435 35581 8447 35615
rect 8389 35575 8447 35581
rect 9306 35572 9312 35624
rect 9364 35572 9370 35624
rect 9950 35572 9956 35624
rect 10008 35572 10014 35624
rect 12250 35572 12256 35624
rect 12308 35612 12314 35624
rect 12723 35612 12751 35643
rect 12986 35640 12992 35652
rect 13044 35640 13050 35692
rect 14384 35689 14412 35720
rect 14476 35689 14504 35788
rect 15013 35785 15025 35819
rect 15059 35816 15071 35819
rect 15378 35816 15384 35828
rect 15059 35788 15384 35816
rect 15059 35785 15071 35788
rect 15013 35779 15071 35785
rect 15378 35776 15384 35788
rect 15436 35776 15442 35828
rect 17957 35819 18015 35825
rect 17957 35785 17969 35819
rect 18003 35816 18015 35819
rect 18046 35816 18052 35828
rect 18003 35788 18052 35816
rect 18003 35785 18015 35788
rect 17957 35779 18015 35785
rect 18046 35776 18052 35788
rect 18104 35776 18110 35828
rect 19242 35776 19248 35828
rect 19300 35816 19306 35828
rect 19429 35819 19487 35825
rect 19429 35816 19441 35819
rect 19300 35788 19441 35816
rect 19300 35776 19306 35788
rect 19429 35785 19441 35788
rect 19475 35785 19487 35819
rect 19429 35779 19487 35785
rect 20165 35819 20223 35825
rect 20165 35785 20177 35819
rect 20211 35816 20223 35819
rect 20438 35816 20444 35828
rect 20211 35788 20444 35816
rect 20211 35785 20223 35788
rect 20165 35779 20223 35785
rect 20438 35776 20444 35788
rect 20496 35776 20502 35828
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 23106 35816 23112 35828
rect 22511 35788 23112 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 23106 35776 23112 35788
rect 23164 35776 23170 35828
rect 23198 35776 23204 35828
rect 23256 35776 23262 35828
rect 23569 35819 23627 35825
rect 23569 35785 23581 35819
rect 23615 35785 23627 35819
rect 23569 35779 23627 35785
rect 14550 35708 14556 35760
rect 14608 35748 14614 35760
rect 14918 35748 14924 35760
rect 14608 35720 14924 35748
rect 14608 35708 14614 35720
rect 14918 35708 14924 35720
rect 14976 35748 14982 35760
rect 16209 35751 16267 35757
rect 16209 35748 16221 35751
rect 14976 35720 16221 35748
rect 14976 35708 14982 35720
rect 16209 35717 16221 35720
rect 16255 35748 16267 35751
rect 16758 35748 16764 35760
rect 16255 35720 16764 35748
rect 16255 35717 16267 35720
rect 16209 35711 16267 35717
rect 16758 35708 16764 35720
rect 16816 35708 16822 35760
rect 17405 35751 17463 35757
rect 17405 35717 17417 35751
rect 17451 35748 17463 35751
rect 18141 35751 18199 35757
rect 18141 35748 18153 35751
rect 17451 35720 18153 35748
rect 17451 35717 17463 35720
rect 17405 35711 17463 35717
rect 18141 35717 18153 35720
rect 18187 35717 18199 35751
rect 18141 35711 18199 35717
rect 18230 35708 18236 35760
rect 18288 35748 18294 35760
rect 20714 35748 20720 35760
rect 18288 35720 20720 35748
rect 18288 35708 18294 35720
rect 20714 35708 20720 35720
rect 20772 35708 20778 35760
rect 21634 35708 21640 35760
rect 21692 35748 21698 35760
rect 22833 35751 22891 35757
rect 21692 35720 22692 35748
rect 21692 35708 21698 35720
rect 13173 35683 13231 35689
rect 13173 35680 13185 35683
rect 13096 35652 13185 35680
rect 12308 35584 12751 35612
rect 12308 35572 12314 35584
rect 10226 35504 10232 35556
rect 10284 35504 10290 35556
rect 12723 35544 12751 35584
rect 13096 35544 13124 35652
rect 13173 35649 13185 35652
rect 13219 35680 13231 35683
rect 14277 35683 14335 35689
rect 14277 35680 14289 35683
rect 13219 35652 14289 35680
rect 13219 35649 13231 35652
rect 13173 35643 13231 35649
rect 13722 35612 13728 35624
rect 13188 35584 13728 35612
rect 13188 35553 13216 35584
rect 13722 35572 13728 35584
rect 13780 35572 13786 35624
rect 13832 35621 13860 35652
rect 14277 35649 14289 35652
rect 14323 35649 14335 35683
rect 14277 35643 14335 35649
rect 14369 35683 14427 35689
rect 14369 35649 14381 35683
rect 14415 35649 14427 35683
rect 14369 35643 14427 35649
rect 14461 35683 14519 35689
rect 14461 35649 14473 35683
rect 14507 35649 14519 35683
rect 14461 35643 14519 35649
rect 14734 35640 14740 35692
rect 14792 35680 14798 35692
rect 15194 35680 15200 35692
rect 14792 35652 15200 35680
rect 14792 35640 14798 35652
rect 15194 35640 15200 35652
rect 15252 35640 15258 35692
rect 15286 35640 15292 35692
rect 15344 35680 15350 35692
rect 15565 35683 15623 35689
rect 15565 35680 15577 35683
rect 15344 35652 15577 35680
rect 15344 35640 15350 35652
rect 15565 35649 15577 35652
rect 15611 35649 15623 35683
rect 15565 35643 15623 35649
rect 15749 35683 15807 35689
rect 15749 35649 15761 35683
rect 15795 35680 15807 35683
rect 15841 35683 15899 35689
rect 15841 35680 15853 35683
rect 15795 35652 15853 35680
rect 15795 35649 15807 35652
rect 15749 35643 15807 35649
rect 15841 35649 15853 35652
rect 15887 35649 15899 35683
rect 15841 35643 15899 35649
rect 15930 35640 15936 35692
rect 15988 35680 15994 35692
rect 16025 35683 16083 35689
rect 16025 35680 16037 35683
rect 15988 35652 16037 35680
rect 15988 35640 15994 35652
rect 16025 35649 16037 35652
rect 16071 35649 16083 35683
rect 16025 35643 16083 35649
rect 16669 35683 16727 35689
rect 16669 35649 16681 35683
rect 16715 35680 16727 35683
rect 16850 35680 16856 35692
rect 16715 35652 16856 35680
rect 16715 35649 16727 35652
rect 16669 35643 16727 35649
rect 13817 35615 13875 35621
rect 13817 35581 13829 35615
rect 13863 35581 13875 35615
rect 13817 35575 13875 35581
rect 14182 35572 14188 35624
rect 14240 35572 14246 35624
rect 15381 35615 15439 35621
rect 15381 35581 15393 35615
rect 15427 35581 15439 35615
rect 15381 35575 15439 35581
rect 15473 35615 15531 35621
rect 15473 35581 15485 35615
rect 15519 35612 15531 35615
rect 15654 35612 15660 35624
rect 15519 35584 15660 35612
rect 15519 35581 15531 35584
rect 15473 35575 15531 35581
rect 12723 35516 13124 35544
rect 13173 35547 13231 35553
rect 13173 35513 13185 35547
rect 13219 35513 13231 35547
rect 13173 35507 13231 35513
rect 13265 35547 13323 35553
rect 13265 35513 13277 35547
rect 13311 35544 13323 35547
rect 13446 35544 13452 35556
rect 13311 35516 13452 35544
rect 13311 35513 13323 35516
rect 13265 35507 13323 35513
rect 13446 35504 13452 35516
rect 13504 35504 13510 35556
rect 15396 35544 15424 35575
rect 15654 35572 15660 35584
rect 15712 35572 15718 35624
rect 16040 35612 16068 35643
rect 16684 35612 16712 35643
rect 16850 35640 16856 35652
rect 16908 35640 16914 35692
rect 17034 35640 17040 35692
rect 17092 35640 17098 35692
rect 17129 35683 17187 35689
rect 17129 35649 17141 35683
rect 17175 35680 17187 35683
rect 17218 35680 17224 35692
rect 17175 35652 17224 35680
rect 17175 35649 17187 35652
rect 17129 35643 17187 35649
rect 17218 35640 17224 35652
rect 17276 35680 17282 35692
rect 17770 35680 17776 35692
rect 17276 35652 17776 35680
rect 17276 35640 17282 35652
rect 17770 35640 17776 35652
rect 17828 35640 17834 35692
rect 17862 35640 17868 35692
rect 17920 35640 17926 35692
rect 19153 35683 19211 35689
rect 19153 35649 19165 35683
rect 19199 35680 19211 35683
rect 19334 35680 19340 35692
rect 19199 35652 19340 35680
rect 19199 35649 19211 35652
rect 19153 35643 19211 35649
rect 19334 35640 19340 35652
rect 19392 35640 19398 35692
rect 19610 35640 19616 35692
rect 19668 35680 19674 35692
rect 19889 35683 19947 35689
rect 19889 35680 19901 35683
rect 19668 35652 19901 35680
rect 19668 35640 19674 35652
rect 19889 35649 19901 35652
rect 19935 35649 19947 35683
rect 19889 35643 19947 35649
rect 20070 35640 20076 35692
rect 20128 35680 20134 35692
rect 20533 35683 20591 35689
rect 20533 35680 20545 35683
rect 20128 35652 20545 35680
rect 20128 35640 20134 35652
rect 20533 35649 20545 35652
rect 20579 35649 20591 35683
rect 21269 35683 21327 35689
rect 20533 35643 20591 35649
rect 20732 35652 21220 35680
rect 16040 35584 16712 35612
rect 19702 35572 19708 35624
rect 19760 35612 19766 35624
rect 19797 35615 19855 35621
rect 19797 35612 19809 35615
rect 19760 35584 19809 35612
rect 19760 35572 19766 35584
rect 19797 35581 19809 35584
rect 19843 35581 19855 35615
rect 19797 35575 19855 35581
rect 20622 35572 20628 35624
rect 20680 35572 20686 35624
rect 16574 35544 16580 35556
rect 15396 35516 16580 35544
rect 16574 35504 16580 35516
rect 16632 35504 16638 35556
rect 18141 35547 18199 35553
rect 18141 35513 18153 35547
rect 18187 35544 18199 35547
rect 20732 35544 20760 35652
rect 21192 35621 21220 35652
rect 21269 35649 21281 35683
rect 21315 35680 21327 35683
rect 21450 35682 21456 35692
rect 21376 35680 21456 35682
rect 21315 35654 21456 35680
rect 21315 35652 21404 35654
rect 21315 35649 21327 35652
rect 21269 35643 21327 35649
rect 21450 35640 21456 35654
rect 21508 35640 21514 35692
rect 21928 35689 21956 35720
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21560 35652 21833 35680
rect 20809 35615 20867 35621
rect 20809 35581 20821 35615
rect 20855 35581 20867 35615
rect 20809 35575 20867 35581
rect 21177 35615 21235 35621
rect 21177 35581 21189 35615
rect 21223 35581 21235 35615
rect 21177 35575 21235 35581
rect 18187 35516 20760 35544
rect 18187 35513 18199 35516
rect 18141 35507 18199 35513
rect 12713 35479 12771 35485
rect 12713 35445 12725 35479
rect 12759 35476 12771 35479
rect 12802 35476 12808 35488
rect 12759 35448 12808 35476
rect 12759 35445 12771 35448
rect 12713 35439 12771 35445
rect 12802 35436 12808 35448
rect 12860 35436 12866 35488
rect 14182 35436 14188 35488
rect 14240 35476 14246 35488
rect 14645 35479 14703 35485
rect 14645 35476 14657 35479
rect 14240 35448 14657 35476
rect 14240 35436 14246 35448
rect 14645 35445 14657 35448
rect 14691 35445 14703 35479
rect 14645 35439 14703 35445
rect 16850 35436 16856 35488
rect 16908 35436 16914 35488
rect 16945 35479 17003 35485
rect 16945 35445 16957 35479
rect 16991 35476 17003 35479
rect 17218 35476 17224 35488
rect 16991 35448 17224 35476
rect 16991 35445 17003 35448
rect 16945 35439 17003 35445
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 18322 35436 18328 35488
rect 18380 35476 18386 35488
rect 19061 35479 19119 35485
rect 19061 35476 19073 35479
rect 18380 35448 19073 35476
rect 18380 35436 18386 35448
rect 19061 35445 19073 35448
rect 19107 35445 19119 35479
rect 19061 35439 19119 35445
rect 19886 35436 19892 35488
rect 19944 35476 19950 35488
rect 20073 35479 20131 35485
rect 20073 35476 20085 35479
rect 19944 35448 20085 35476
rect 19944 35436 19950 35448
rect 20073 35445 20085 35448
rect 20119 35445 20131 35479
rect 20824 35476 20852 35575
rect 21192 35544 21220 35575
rect 21358 35572 21364 35624
rect 21416 35612 21422 35624
rect 21560 35612 21588 35652
rect 21821 35649 21833 35652
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 21914 35683 21972 35689
rect 21914 35649 21926 35683
rect 21960 35649 21972 35683
rect 21914 35643 21972 35649
rect 22051 35683 22109 35689
rect 22051 35649 22063 35683
rect 22097 35649 22109 35683
rect 22051 35643 22109 35649
rect 21416 35584 21588 35612
rect 21637 35615 21695 35621
rect 21416 35572 21422 35584
rect 21637 35581 21649 35615
rect 21683 35612 21695 35615
rect 22066 35612 22094 35643
rect 22186 35640 22192 35692
rect 22244 35640 22250 35692
rect 22327 35683 22385 35689
rect 22327 35649 22339 35683
rect 22373 35680 22385 35683
rect 22462 35680 22468 35692
rect 22373 35652 22468 35680
rect 22373 35649 22385 35652
rect 22327 35643 22385 35649
rect 22462 35640 22468 35652
rect 22520 35640 22526 35692
rect 22554 35640 22560 35692
rect 22612 35640 22618 35692
rect 22664 35689 22692 35720
rect 22833 35717 22845 35751
rect 22879 35748 22891 35751
rect 23584 35748 23612 35779
rect 23658 35776 23664 35828
rect 23716 35816 23722 35828
rect 24210 35816 24216 35828
rect 23716 35788 24216 35816
rect 23716 35776 23722 35788
rect 24210 35776 24216 35788
rect 24268 35816 24274 35828
rect 24305 35819 24363 35825
rect 24305 35816 24317 35819
rect 24268 35788 24317 35816
rect 24268 35776 24274 35788
rect 24305 35785 24317 35788
rect 24351 35785 24363 35819
rect 24305 35779 24363 35785
rect 24673 35819 24731 35825
rect 24673 35785 24685 35819
rect 24719 35816 24731 35819
rect 24762 35816 24768 35828
rect 24719 35788 24768 35816
rect 24719 35785 24731 35788
rect 24673 35779 24731 35785
rect 24762 35776 24768 35788
rect 24820 35816 24826 35828
rect 25885 35819 25943 35825
rect 25885 35816 25897 35819
rect 24820 35788 25897 35816
rect 24820 35776 24826 35788
rect 25885 35785 25897 35788
rect 25931 35785 25943 35819
rect 25885 35779 25943 35785
rect 26234 35776 26240 35828
rect 26292 35816 26298 35828
rect 26513 35819 26571 35825
rect 26513 35816 26525 35819
rect 26292 35788 26525 35816
rect 26292 35776 26298 35788
rect 26513 35785 26525 35788
rect 26559 35785 26571 35819
rect 26513 35779 26571 35785
rect 22879 35720 23612 35748
rect 23952 35720 24532 35748
rect 22879 35717 22891 35720
rect 22833 35711 22891 35717
rect 23952 35692 23980 35720
rect 22650 35683 22708 35689
rect 22650 35649 22662 35683
rect 22696 35649 22708 35683
rect 22650 35643 22708 35649
rect 22922 35640 22928 35692
rect 22980 35640 22986 35692
rect 23014 35640 23020 35692
rect 23072 35689 23078 35692
rect 23072 35680 23080 35689
rect 23293 35683 23351 35689
rect 23072 35652 23117 35680
rect 23072 35643 23080 35652
rect 23293 35649 23305 35683
rect 23339 35649 23351 35683
rect 23293 35643 23351 35649
rect 23477 35683 23535 35689
rect 23477 35649 23489 35683
rect 23523 35649 23535 35683
rect 23477 35643 23535 35649
rect 23072 35640 23078 35643
rect 21683 35584 22094 35612
rect 22204 35612 22232 35640
rect 23308 35612 23336 35643
rect 22204 35584 23336 35612
rect 21683 35581 21695 35584
rect 21637 35575 21695 35581
rect 22646 35544 22652 35556
rect 21192 35516 22652 35544
rect 22646 35504 22652 35516
rect 22704 35504 22710 35556
rect 23492 35544 23520 35643
rect 23934 35640 23940 35692
rect 23992 35640 23998 35692
rect 24118 35640 24124 35692
rect 24176 35680 24182 35692
rect 24504 35689 24532 35720
rect 24854 35708 24860 35760
rect 24912 35748 24918 35760
rect 25685 35751 25743 35757
rect 25685 35748 25697 35751
rect 24912 35720 25697 35748
rect 24912 35708 24918 35720
rect 25685 35717 25697 35720
rect 25731 35717 25743 35751
rect 25685 35711 25743 35717
rect 24213 35683 24271 35689
rect 24213 35680 24225 35683
rect 24176 35652 24225 35680
rect 24176 35640 24182 35652
rect 24213 35649 24225 35652
rect 24259 35649 24271 35683
rect 24213 35643 24271 35649
rect 24489 35683 24547 35689
rect 24489 35649 24501 35683
rect 24535 35649 24547 35683
rect 24489 35643 24547 35649
rect 24670 35640 24676 35692
rect 24728 35680 24734 35692
rect 24765 35683 24823 35689
rect 24765 35680 24777 35683
rect 24728 35652 24777 35680
rect 24728 35640 24734 35652
rect 24765 35649 24777 35652
rect 24811 35649 24823 35683
rect 24872 35680 24900 35708
rect 24949 35683 25007 35689
rect 24949 35680 24961 35683
rect 24872 35652 24961 35680
rect 24765 35643 24823 35649
rect 24949 35649 24961 35652
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 25038 35640 25044 35692
rect 25096 35640 25102 35692
rect 25317 35683 25375 35689
rect 25317 35680 25329 35683
rect 25240 35652 25329 35680
rect 24029 35615 24087 35621
rect 24029 35581 24041 35615
rect 24075 35612 24087 35615
rect 24857 35615 24915 35621
rect 24857 35612 24869 35615
rect 24075 35584 24869 35612
rect 24075 35581 24087 35584
rect 24029 35575 24087 35581
rect 24857 35581 24869 35584
rect 24903 35581 24915 35615
rect 24857 35575 24915 35581
rect 25130 35572 25136 35624
rect 25188 35612 25194 35624
rect 25240 35612 25268 35652
rect 25317 35649 25329 35652
rect 25363 35649 25375 35683
rect 25317 35643 25375 35649
rect 25406 35640 25412 35692
rect 25464 35680 25470 35692
rect 26145 35683 26203 35689
rect 26145 35680 26157 35683
rect 25464 35652 26157 35680
rect 25464 35640 25470 35652
rect 26145 35649 26157 35652
rect 26191 35649 26203 35683
rect 26145 35643 26203 35649
rect 26326 35640 26332 35692
rect 26384 35640 26390 35692
rect 26344 35612 26372 35640
rect 25188 35584 25268 35612
rect 25332 35584 26372 35612
rect 25188 35572 25194 35584
rect 22740 35516 23520 35544
rect 22094 35476 22100 35488
rect 20824 35448 22100 35476
rect 20073 35439 20131 35445
rect 22094 35436 22100 35448
rect 22152 35436 22158 35488
rect 22186 35436 22192 35488
rect 22244 35476 22250 35488
rect 22740 35476 22768 35516
rect 24118 35504 24124 35556
rect 24176 35544 24182 35556
rect 25332 35544 25360 35584
rect 26053 35547 26111 35553
rect 26053 35544 26065 35547
rect 24176 35516 25360 35544
rect 25424 35516 26065 35544
rect 24176 35504 24182 35516
rect 22244 35448 22768 35476
rect 22244 35436 22250 35448
rect 23106 35436 23112 35488
rect 23164 35476 23170 35488
rect 25424 35485 25452 35516
rect 26053 35513 26065 35516
rect 26099 35544 26111 35547
rect 26510 35544 26516 35556
rect 26099 35516 26516 35544
rect 26099 35513 26111 35516
rect 26053 35507 26111 35513
rect 26510 35504 26516 35516
rect 26568 35504 26574 35556
rect 23385 35479 23443 35485
rect 23385 35476 23397 35479
rect 23164 35448 23397 35476
rect 23164 35436 23170 35448
rect 23385 35445 23397 35448
rect 23431 35445 23443 35479
rect 23385 35439 23443 35445
rect 25409 35479 25467 35485
rect 25409 35445 25421 35479
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 25590 35436 25596 35488
rect 25648 35436 25654 35488
rect 25869 35479 25927 35485
rect 25869 35445 25881 35479
rect 25915 35476 25927 35479
rect 26142 35476 26148 35488
rect 25915 35448 26148 35476
rect 25915 35445 25927 35448
rect 25869 35439 25927 35445
rect 26142 35436 26148 35448
rect 26200 35436 26206 35488
rect 1104 35386 36524 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 36524 35386
rect 1104 35312 36524 35334
rect 7006 35232 7012 35284
rect 7064 35232 7070 35284
rect 9306 35232 9312 35284
rect 9364 35232 9370 35284
rect 9861 35275 9919 35281
rect 9861 35241 9873 35275
rect 9907 35272 9919 35275
rect 9950 35272 9956 35284
rect 9907 35244 9956 35272
rect 9907 35241 9919 35244
rect 9861 35235 9919 35241
rect 9950 35232 9956 35244
rect 10008 35232 10014 35284
rect 12526 35232 12532 35284
rect 12584 35272 12590 35284
rect 12621 35275 12679 35281
rect 12621 35272 12633 35275
rect 12584 35244 12633 35272
rect 12584 35232 12590 35244
rect 12621 35241 12633 35244
rect 12667 35272 12679 35275
rect 12710 35272 12716 35284
rect 12667 35244 12716 35272
rect 12667 35241 12679 35244
rect 12621 35235 12679 35241
rect 12710 35232 12716 35244
rect 12768 35232 12774 35284
rect 12805 35275 12863 35281
rect 12805 35241 12817 35275
rect 12851 35272 12863 35275
rect 12986 35272 12992 35284
rect 12851 35244 12992 35272
rect 12851 35241 12863 35244
rect 12805 35235 12863 35241
rect 12986 35232 12992 35244
rect 13044 35232 13050 35284
rect 13449 35275 13507 35281
rect 13449 35272 13461 35275
rect 13096 35244 13461 35272
rect 10042 35164 10048 35216
rect 10100 35204 10106 35216
rect 10100 35176 12848 35204
rect 10100 35164 10106 35176
rect 4893 35139 4951 35145
rect 4893 35105 4905 35139
rect 4939 35136 4951 35139
rect 5534 35136 5540 35148
rect 4939 35108 5540 35136
rect 4939 35105 4951 35108
rect 4893 35099 4951 35105
rect 5534 35096 5540 35108
rect 5592 35096 5598 35148
rect 6546 35096 6552 35148
rect 6604 35136 6610 35148
rect 6917 35139 6975 35145
rect 6917 35136 6929 35139
rect 6604 35108 6929 35136
rect 6604 35096 6610 35108
rect 6917 35105 6929 35108
rect 6963 35105 6975 35139
rect 6917 35099 6975 35105
rect 7098 35096 7104 35148
rect 7156 35136 7162 35148
rect 7469 35139 7527 35145
rect 7469 35136 7481 35139
rect 7156 35108 7481 35136
rect 7156 35096 7162 35108
rect 7469 35105 7481 35108
rect 7515 35105 7527 35139
rect 7469 35099 7527 35105
rect 7558 35096 7564 35148
rect 7616 35096 7622 35148
rect 11425 35139 11483 35145
rect 11425 35105 11437 35139
rect 11471 35136 11483 35139
rect 11514 35136 11520 35148
rect 11471 35108 11520 35136
rect 11471 35105 11483 35108
rect 11425 35099 11483 35105
rect 11514 35096 11520 35108
rect 11572 35096 11578 35148
rect 11606 35096 11612 35148
rect 11664 35136 11670 35148
rect 12250 35136 12256 35148
rect 11664 35108 12256 35136
rect 11664 35096 11670 35108
rect 12250 35096 12256 35108
rect 12308 35136 12314 35148
rect 12529 35139 12587 35145
rect 12529 35136 12541 35139
rect 12308 35108 12541 35136
rect 12308 35096 12314 35108
rect 12529 35105 12541 35108
rect 12575 35105 12587 35139
rect 12529 35099 12587 35105
rect 9214 35028 9220 35080
rect 9272 35028 9278 35080
rect 9398 35028 9404 35080
rect 9456 35028 9462 35080
rect 9677 35071 9735 35077
rect 9677 35037 9689 35071
rect 9723 35037 9735 35071
rect 9677 35031 9735 35037
rect 9861 35071 9919 35077
rect 9861 35037 9873 35071
rect 9907 35068 9919 35071
rect 9950 35068 9956 35080
rect 9907 35040 9956 35068
rect 9907 35037 9919 35040
rect 9861 35031 9919 35037
rect 5169 35003 5227 35009
rect 5169 34969 5181 35003
rect 5215 35000 5227 35003
rect 5442 35000 5448 35012
rect 5215 34972 5448 35000
rect 5215 34969 5227 34972
rect 5169 34963 5227 34969
rect 5442 34960 5448 34972
rect 5500 34960 5506 35012
rect 7926 35000 7932 35012
rect 6394 34972 7932 35000
rect 7926 34960 7932 34972
rect 7984 34960 7990 35012
rect 9692 35000 9720 35031
rect 9950 35028 9956 35040
rect 10008 35028 10014 35080
rect 10137 35071 10195 35077
rect 10137 35037 10149 35071
rect 10183 35068 10195 35071
rect 10226 35068 10232 35080
rect 10183 35040 10232 35068
rect 10183 35037 10195 35040
rect 10137 35031 10195 35037
rect 10226 35028 10232 35040
rect 10284 35028 10290 35080
rect 11333 35071 11391 35077
rect 11333 35037 11345 35071
rect 11379 35068 11391 35071
rect 12342 35068 12348 35080
rect 11379 35040 12348 35068
rect 11379 35037 11391 35040
rect 11333 35031 11391 35037
rect 10042 35000 10048 35012
rect 9692 34972 10048 35000
rect 10042 34960 10048 34972
rect 10100 34960 10106 35012
rect 7377 34935 7435 34941
rect 7377 34901 7389 34935
rect 7423 34932 7435 34935
rect 11348 34932 11376 35031
rect 12342 35028 12348 35040
rect 12400 35028 12406 35080
rect 12618 35028 12624 35080
rect 12676 35028 12682 35080
rect 12713 35071 12771 35077
rect 12713 35037 12725 35071
rect 12759 35037 12771 35071
rect 12713 35031 12771 35037
rect 12434 34960 12440 35012
rect 12492 35000 12498 35012
rect 12728 35000 12756 35031
rect 12492 34972 12756 35000
rect 12820 35000 12848 35176
rect 13096 35136 13124 35244
rect 13449 35241 13461 35244
rect 13495 35241 13507 35275
rect 13449 35235 13507 35241
rect 14182 35232 14188 35284
rect 14240 35232 14246 35284
rect 14274 35232 14280 35284
rect 14332 35272 14338 35284
rect 14553 35275 14611 35281
rect 14553 35272 14565 35275
rect 14332 35244 14565 35272
rect 14332 35232 14338 35244
rect 14553 35241 14565 35244
rect 14599 35241 14611 35275
rect 14553 35235 14611 35241
rect 20070 35232 20076 35284
rect 20128 35232 20134 35284
rect 21729 35275 21787 35281
rect 21729 35241 21741 35275
rect 21775 35272 21787 35275
rect 22554 35272 22560 35284
rect 21775 35244 22560 35272
rect 21775 35241 21787 35244
rect 21729 35235 21787 35241
rect 22554 35232 22560 35244
rect 22612 35232 22618 35284
rect 22646 35232 22652 35284
rect 22704 35232 22710 35284
rect 22741 35275 22799 35281
rect 22741 35241 22753 35275
rect 22787 35272 22799 35275
rect 23934 35272 23940 35284
rect 22787 35244 23940 35272
rect 22787 35241 22799 35244
rect 22741 35235 22799 35241
rect 23934 35232 23940 35244
rect 23992 35232 23998 35284
rect 25038 35232 25044 35284
rect 25096 35272 25102 35284
rect 25225 35275 25283 35281
rect 25225 35272 25237 35275
rect 25096 35244 25237 35272
rect 25096 35232 25102 35244
rect 25225 35241 25237 35244
rect 25271 35241 25283 35275
rect 25225 35235 25283 35241
rect 25498 35232 25504 35284
rect 25556 35232 25562 35284
rect 26053 35275 26111 35281
rect 26053 35241 26065 35275
rect 26099 35272 26111 35275
rect 26329 35275 26387 35281
rect 26329 35272 26341 35275
rect 26099 35244 26341 35272
rect 26099 35241 26111 35244
rect 26053 35235 26111 35241
rect 26329 35241 26341 35244
rect 26375 35241 26387 35275
rect 26329 35235 26387 35241
rect 26510 35232 26516 35284
rect 26568 35272 26574 35284
rect 26973 35275 27031 35281
rect 26973 35272 26985 35275
rect 26568 35244 26985 35272
rect 26568 35232 26574 35244
rect 26973 35241 26985 35244
rect 27019 35241 27031 35275
rect 26973 35235 27031 35241
rect 13265 35207 13323 35213
rect 13265 35173 13277 35207
rect 13311 35173 13323 35207
rect 13265 35167 13323 35173
rect 13004 35108 13124 35136
rect 13280 35136 13308 35167
rect 14734 35164 14740 35216
rect 14792 35204 14798 35216
rect 14792 35176 20024 35204
rect 14792 35164 14798 35176
rect 13280 35108 13676 35136
rect 13004 35080 13032 35108
rect 12986 35028 12992 35080
rect 13044 35028 13050 35080
rect 13648 35077 13676 35108
rect 13722 35096 13728 35148
rect 13780 35136 13786 35148
rect 14093 35139 14151 35145
rect 14093 35136 14105 35139
rect 13780 35108 14105 35136
rect 13780 35096 13786 35108
rect 14093 35105 14105 35108
rect 14139 35105 14151 35139
rect 14093 35099 14151 35105
rect 16761 35139 16819 35145
rect 16761 35105 16773 35139
rect 16807 35105 16819 35139
rect 16761 35099 16819 35105
rect 17037 35139 17095 35145
rect 17037 35105 17049 35139
rect 17083 35136 17095 35139
rect 17402 35136 17408 35148
rect 17083 35108 17408 35136
rect 17083 35105 17095 35108
rect 17037 35099 17095 35105
rect 13357 35071 13415 35077
rect 13357 35068 13369 35071
rect 13096 35040 13369 35068
rect 13096 35009 13124 35040
rect 13357 35037 13369 35040
rect 13403 35037 13415 35071
rect 13357 35031 13415 35037
rect 13633 35071 13691 35077
rect 13633 35037 13645 35071
rect 13679 35037 13691 35071
rect 13998 35068 14004 35080
rect 13633 35031 13691 35037
rect 13740 35040 14004 35068
rect 13081 35003 13139 35009
rect 13081 35000 13093 35003
rect 12820 34972 13093 35000
rect 12492 34960 12498 34972
rect 13081 34969 13093 34972
rect 13127 34969 13139 35003
rect 13081 34963 13139 34969
rect 13265 35003 13323 35009
rect 13265 34969 13277 35003
rect 13311 35000 13323 35003
rect 13740 35000 13768 35040
rect 13998 35028 14004 35040
rect 14056 35028 14062 35080
rect 14366 35028 14372 35080
rect 14424 35028 14430 35080
rect 15930 35028 15936 35080
rect 15988 35068 15994 35080
rect 16669 35071 16727 35077
rect 16669 35068 16681 35071
rect 15988 35040 16681 35068
rect 15988 35028 15994 35040
rect 16669 35037 16681 35040
rect 16715 35037 16727 35071
rect 16776 35068 16804 35099
rect 17402 35096 17408 35108
rect 17460 35136 17466 35148
rect 17460 35108 18276 35136
rect 17460 35096 17466 35108
rect 17310 35068 17316 35080
rect 16776 35040 17316 35068
rect 16669 35031 16727 35037
rect 17310 35028 17316 35040
rect 17368 35028 17374 35080
rect 17862 35028 17868 35080
rect 17920 35028 17926 35080
rect 18138 35028 18144 35080
rect 18196 35028 18202 35080
rect 18248 35077 18276 35108
rect 19886 35096 19892 35148
rect 19944 35096 19950 35148
rect 19996 35136 20024 35176
rect 21450 35164 21456 35216
rect 21508 35204 21514 35216
rect 23017 35207 23075 35213
rect 23017 35204 23029 35207
rect 21508 35176 22094 35204
rect 21508 35164 21514 35176
rect 22066 35136 22094 35176
rect 22572 35176 23029 35204
rect 22572 35136 22600 35176
rect 23017 35173 23029 35176
rect 23063 35173 23075 35207
rect 26142 35204 26148 35216
rect 23017 35167 23075 35173
rect 25240 35176 26148 35204
rect 19996 35108 21772 35136
rect 22066 35108 22600 35136
rect 18233 35071 18291 35077
rect 18233 35037 18245 35071
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 18322 35028 18328 35080
rect 18380 35028 18386 35080
rect 18506 35028 18512 35080
rect 18564 35028 18570 35080
rect 18598 35028 18604 35080
rect 18656 35028 18662 35080
rect 19334 35028 19340 35080
rect 19392 35068 19398 35080
rect 21744 35077 21772 35108
rect 19797 35071 19855 35077
rect 19797 35068 19809 35071
rect 19392 35040 19809 35068
rect 19392 35028 19398 35040
rect 19797 35037 19809 35040
rect 19843 35037 19855 35071
rect 19797 35031 19855 35037
rect 21735 35071 21793 35077
rect 21735 35037 21747 35071
rect 21781 35037 21793 35071
rect 21735 35031 21793 35037
rect 21910 35028 21916 35080
rect 21968 35028 21974 35080
rect 22002 35028 22008 35080
rect 22060 35068 22066 35080
rect 22572 35077 22600 35108
rect 22833 35139 22891 35145
rect 22833 35105 22845 35139
rect 22879 35136 22891 35139
rect 22879 35108 23152 35136
rect 22879 35105 22891 35108
rect 22833 35099 22891 35105
rect 23124 35080 23152 35108
rect 22281 35071 22339 35077
rect 22281 35068 22293 35071
rect 22060 35040 22293 35068
rect 22060 35028 22066 35040
rect 22281 35037 22293 35040
rect 22327 35037 22339 35071
rect 22281 35031 22339 35037
rect 22557 35071 22615 35077
rect 22557 35037 22569 35071
rect 22603 35037 22615 35071
rect 22557 35031 22615 35037
rect 22925 35071 22983 35077
rect 22925 35037 22937 35071
rect 22971 35037 22983 35071
rect 22925 35031 22983 35037
rect 13311 34972 13768 35000
rect 13817 35003 13875 35009
rect 13311 34969 13323 34972
rect 13265 34963 13323 34969
rect 13817 34969 13829 35003
rect 13863 35000 13875 35003
rect 21358 35000 21364 35012
rect 13863 34972 21364 35000
rect 13863 34969 13875 34972
rect 13817 34963 13875 34969
rect 21358 34960 21364 34972
rect 21416 34960 21422 35012
rect 21542 34960 21548 35012
rect 21600 35000 21606 35012
rect 22020 35000 22048 35028
rect 21600 34972 22048 35000
rect 22097 35003 22155 35009
rect 21600 34960 21606 34972
rect 22097 34969 22109 35003
rect 22143 35000 22155 35003
rect 22186 35000 22192 35012
rect 22143 34972 22192 35000
rect 22143 34969 22155 34972
rect 22097 34963 22155 34969
rect 22186 34960 22192 34972
rect 22244 34960 22250 35012
rect 22465 35003 22523 35009
rect 22465 34969 22477 35003
rect 22511 35000 22523 35003
rect 22940 35000 22968 35031
rect 23106 35028 23112 35080
rect 23164 35028 23170 35080
rect 24762 35028 24768 35080
rect 24820 35028 24826 35080
rect 24854 35028 24860 35080
rect 24912 35028 24918 35080
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35068 25099 35071
rect 25240 35068 25268 35176
rect 26142 35164 26148 35176
rect 26200 35164 26206 35216
rect 26528 35176 27108 35204
rect 25332 35108 25544 35136
rect 25332 35077 25360 35108
rect 25087 35040 25268 35068
rect 25317 35071 25375 35077
rect 25087 35037 25099 35040
rect 25041 35031 25099 35037
rect 25317 35037 25329 35071
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 25424 35000 25452 35031
rect 22511 34972 22968 35000
rect 23768 34972 25452 35000
rect 22511 34969 22523 34972
rect 22465 34963 22523 34969
rect 7423 34904 11376 34932
rect 7423 34901 7435 34904
rect 7377 34895 7435 34901
rect 11698 34892 11704 34944
rect 11756 34892 11762 34944
rect 11790 34892 11796 34944
rect 11848 34932 11854 34944
rect 12253 34935 12311 34941
rect 12253 34932 12265 34935
rect 11848 34904 12265 34932
rect 11848 34892 11854 34904
rect 12253 34901 12265 34904
rect 12299 34932 12311 34935
rect 12710 34932 12716 34944
rect 12299 34904 12716 34932
rect 12299 34901 12311 34904
rect 12253 34895 12311 34901
rect 12710 34892 12716 34904
rect 12768 34892 12774 34944
rect 12894 34892 12900 34944
rect 12952 34932 12958 34944
rect 20622 34932 20628 34944
rect 12952 34904 20628 34932
rect 12952 34892 12958 34904
rect 20622 34892 20628 34904
rect 20680 34892 20686 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 23768 34932 23796 34972
rect 20772 34904 23796 34932
rect 20772 34892 20778 34904
rect 23842 34892 23848 34944
rect 23900 34932 23906 34944
rect 25516 34932 25544 35108
rect 25590 35096 25596 35148
rect 25648 35096 25654 35148
rect 26234 35028 26240 35080
rect 26292 35068 26298 35080
rect 26528 35077 26556 35176
rect 26786 35096 26792 35148
rect 26844 35096 26850 35148
rect 26513 35071 26571 35077
rect 26513 35068 26525 35071
rect 26292 35040 26525 35068
rect 26292 35028 26298 35040
rect 26513 35037 26525 35040
rect 26559 35037 26571 35071
rect 26513 35031 26571 35037
rect 26697 35071 26755 35077
rect 26697 35037 26709 35071
rect 26743 35068 26755 35071
rect 26804 35068 26832 35096
rect 27080 35077 27108 35176
rect 26743 35040 26832 35068
rect 27065 35071 27123 35077
rect 26743 35037 26755 35040
rect 26697 35031 26755 35037
rect 27065 35037 27077 35071
rect 27111 35037 27123 35071
rect 27065 35031 27123 35037
rect 25866 34960 25872 35012
rect 25924 34960 25930 35012
rect 26085 35003 26143 35009
rect 26085 34969 26097 35003
rect 26131 35000 26143 35003
rect 26789 35003 26847 35009
rect 26789 35000 26801 35003
rect 26131 34972 26801 35000
rect 26131 34969 26143 34972
rect 26085 34963 26143 34969
rect 26789 34969 26801 34972
rect 26835 34969 26847 35003
rect 26789 34963 26847 34969
rect 23900 34904 25544 34932
rect 23900 34892 23906 34904
rect 26234 34892 26240 34944
rect 26292 34892 26298 34944
rect 1104 34842 36524 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 36524 34842
rect 1104 34768 36524 34790
rect 5442 34688 5448 34740
rect 5500 34728 5506 34740
rect 6365 34731 6423 34737
rect 6365 34728 6377 34731
rect 5500 34700 6377 34728
rect 5500 34688 5506 34700
rect 6365 34697 6377 34700
rect 6411 34697 6423 34731
rect 6365 34691 6423 34697
rect 6546 34688 6552 34740
rect 6604 34728 6610 34740
rect 6825 34731 6883 34737
rect 6825 34728 6837 34731
rect 6604 34700 6837 34728
rect 6604 34688 6610 34700
rect 6825 34697 6837 34700
rect 6871 34697 6883 34731
rect 6825 34691 6883 34697
rect 9125 34731 9183 34737
rect 9125 34697 9137 34731
rect 9171 34728 9183 34731
rect 9214 34728 9220 34740
rect 9171 34700 9220 34728
rect 9171 34697 9183 34700
rect 9125 34691 9183 34697
rect 9214 34688 9220 34700
rect 9272 34728 9278 34740
rect 9585 34731 9643 34737
rect 9585 34728 9597 34731
rect 9272 34700 9597 34728
rect 9272 34688 9278 34700
rect 9585 34697 9597 34700
rect 9631 34697 9643 34731
rect 9585 34691 9643 34697
rect 11514 34688 11520 34740
rect 11572 34688 11578 34740
rect 12894 34728 12900 34740
rect 12406 34700 12900 34728
rect 9398 34660 9404 34672
rect 9232 34632 9404 34660
rect 6733 34595 6791 34601
rect 6733 34561 6745 34595
rect 6779 34592 6791 34595
rect 8294 34592 8300 34604
rect 6779 34564 8300 34592
rect 6779 34561 6791 34564
rect 6733 34555 6791 34561
rect 8294 34552 8300 34564
rect 8352 34552 8358 34604
rect 9232 34601 9260 34632
rect 9398 34620 9404 34632
rect 9456 34660 9462 34672
rect 10137 34663 10195 34669
rect 10137 34660 10149 34663
rect 9456 34632 10149 34660
rect 9456 34620 9462 34632
rect 10137 34629 10149 34632
rect 10183 34629 10195 34663
rect 10137 34623 10195 34629
rect 11698 34620 11704 34672
rect 11756 34660 11762 34672
rect 12406 34660 12434 34700
rect 12894 34688 12900 34700
rect 12952 34688 12958 34740
rect 12986 34688 12992 34740
rect 13044 34688 13050 34740
rect 14458 34688 14464 34740
rect 14516 34728 14522 34740
rect 16850 34728 16856 34740
rect 14516 34700 16856 34728
rect 14516 34688 14522 34700
rect 16850 34688 16856 34700
rect 16908 34688 16914 34740
rect 18598 34728 18604 34740
rect 18524 34700 18604 34728
rect 11756 34632 12434 34660
rect 11756 34620 11762 34632
rect 12710 34620 12716 34672
rect 12768 34660 12774 34672
rect 17954 34660 17960 34672
rect 12768 34632 13032 34660
rect 12768 34620 12774 34632
rect 9217 34595 9275 34601
rect 9217 34561 9229 34595
rect 9263 34561 9275 34595
rect 9217 34555 9275 34561
rect 9766 34552 9772 34604
rect 9824 34592 9830 34604
rect 9953 34595 10011 34601
rect 9953 34592 9965 34595
rect 9824 34564 9965 34592
rect 9824 34552 9830 34564
rect 9953 34561 9965 34564
rect 9999 34592 10011 34595
rect 10045 34595 10103 34601
rect 10045 34592 10057 34595
rect 9999 34564 10057 34592
rect 9999 34561 10011 34564
rect 9953 34555 10011 34561
rect 10045 34561 10057 34564
rect 10091 34561 10103 34595
rect 10045 34555 10103 34561
rect 10226 34552 10232 34604
rect 10284 34552 10290 34604
rect 11790 34592 11796 34604
rect 10796 34564 11796 34592
rect 7009 34527 7067 34533
rect 7009 34493 7021 34527
rect 7055 34524 7067 34527
rect 7558 34524 7564 34536
rect 7055 34496 7564 34524
rect 7055 34493 7067 34496
rect 7009 34487 7067 34493
rect 7558 34484 7564 34496
rect 7616 34484 7622 34536
rect 8389 34527 8447 34533
rect 8389 34493 8401 34527
rect 8435 34524 8447 34527
rect 9401 34527 9459 34533
rect 8435 34496 8800 34524
rect 8435 34493 8447 34496
rect 8389 34487 8447 34493
rect 8662 34416 8668 34468
rect 8720 34416 8726 34468
rect 8772 34465 8800 34496
rect 9401 34493 9413 34527
rect 9447 34524 9459 34527
rect 9490 34524 9496 34536
rect 9447 34496 9496 34524
rect 9447 34493 9459 34496
rect 9401 34487 9459 34493
rect 9490 34484 9496 34496
rect 9548 34484 9554 34536
rect 9861 34527 9919 34533
rect 9861 34493 9873 34527
rect 9907 34524 9919 34527
rect 10502 34524 10508 34536
rect 9907 34496 10508 34524
rect 9907 34493 9919 34496
rect 9861 34487 9919 34493
rect 10060 34468 10088 34496
rect 10502 34484 10508 34496
rect 10560 34484 10566 34536
rect 8757 34459 8815 34465
rect 8757 34425 8769 34459
rect 8803 34425 8815 34459
rect 8757 34419 8815 34425
rect 10042 34416 10048 34468
rect 10100 34416 10106 34468
rect 9950 34348 9956 34400
rect 10008 34388 10014 34400
rect 10796 34388 10824 34564
rect 11790 34552 11796 34564
rect 11848 34552 11854 34604
rect 11882 34552 11888 34604
rect 11940 34552 11946 34604
rect 12342 34552 12348 34604
rect 12400 34552 12406 34604
rect 12802 34552 12808 34604
rect 12860 34552 12866 34604
rect 13004 34601 13032 34632
rect 15028 34632 15884 34660
rect 15028 34604 15056 34632
rect 12989 34595 13047 34601
rect 12989 34561 13001 34595
rect 13035 34561 13047 34595
rect 12989 34555 13047 34561
rect 15010 34552 15016 34604
rect 15068 34552 15074 34604
rect 15856 34601 15884 34632
rect 17144 34632 17960 34660
rect 15197 34595 15255 34601
rect 15197 34561 15209 34595
rect 15243 34561 15255 34595
rect 15197 34555 15255 34561
rect 15841 34595 15899 34601
rect 15841 34561 15853 34595
rect 15887 34561 15899 34595
rect 15841 34555 15899 34561
rect 11054 34484 11060 34536
rect 11112 34524 11118 34536
rect 11977 34527 12035 34533
rect 11977 34524 11989 34527
rect 11112 34496 11989 34524
rect 11112 34484 11118 34496
rect 11977 34493 11989 34496
rect 12023 34493 12035 34527
rect 11977 34487 12035 34493
rect 12069 34527 12127 34533
rect 12069 34493 12081 34527
rect 12115 34493 12127 34527
rect 12069 34487 12127 34493
rect 12437 34527 12495 34533
rect 12437 34493 12449 34527
rect 12483 34493 12495 34527
rect 12437 34487 12495 34493
rect 14921 34527 14979 34533
rect 14921 34493 14933 34527
rect 14967 34493 14979 34527
rect 15212 34524 15240 34555
rect 16758 34552 16764 34604
rect 16816 34552 16822 34604
rect 16945 34595 17003 34601
rect 16945 34561 16957 34595
rect 16991 34592 17003 34595
rect 17144 34592 17172 34632
rect 17954 34620 17960 34632
rect 18012 34660 18018 34672
rect 18524 34660 18552 34700
rect 18598 34688 18604 34700
rect 18656 34728 18662 34740
rect 18966 34728 18972 34740
rect 18656 34700 18972 34728
rect 18656 34688 18662 34700
rect 18966 34688 18972 34700
rect 19024 34688 19030 34740
rect 19242 34688 19248 34740
rect 19300 34688 19306 34740
rect 19610 34688 19616 34740
rect 19668 34728 19674 34740
rect 19978 34728 19984 34740
rect 19668 34700 19984 34728
rect 19668 34688 19674 34700
rect 19978 34688 19984 34700
rect 20036 34728 20042 34740
rect 22186 34728 22192 34740
rect 20036 34700 22192 34728
rect 20036 34688 20042 34700
rect 22186 34688 22192 34700
rect 22244 34688 22250 34740
rect 25866 34728 25872 34740
rect 22572 34700 25872 34728
rect 19260 34660 19288 34688
rect 18012 34632 18552 34660
rect 18012 34620 18018 34632
rect 16991 34564 17172 34592
rect 16991 34561 17003 34564
rect 16945 34555 17003 34561
rect 17218 34552 17224 34604
rect 17276 34592 17282 34604
rect 18524 34601 18552 34632
rect 18708 34632 19288 34660
rect 18708 34601 18736 34632
rect 21726 34620 21732 34672
rect 21784 34660 21790 34672
rect 21910 34660 21916 34672
rect 21784 34632 21916 34660
rect 21784 34620 21790 34632
rect 21910 34620 21916 34632
rect 21968 34660 21974 34672
rect 22572 34660 22600 34700
rect 25866 34688 25872 34700
rect 25924 34688 25930 34740
rect 21968 34632 22600 34660
rect 22649 34663 22707 34669
rect 21968 34620 21974 34632
rect 22649 34629 22661 34663
rect 22695 34660 22707 34663
rect 22695 34632 25912 34660
rect 22695 34629 22707 34632
rect 22649 34623 22707 34629
rect 17681 34595 17739 34601
rect 17681 34592 17693 34595
rect 17276 34564 17693 34592
rect 17276 34552 17282 34564
rect 17681 34561 17693 34564
rect 17727 34561 17739 34595
rect 17681 34555 17739 34561
rect 18417 34595 18475 34601
rect 18417 34561 18429 34595
rect 18463 34561 18475 34595
rect 18417 34555 18475 34561
rect 18509 34595 18567 34601
rect 18509 34561 18521 34595
rect 18555 34561 18567 34595
rect 18509 34555 18567 34561
rect 18693 34595 18751 34601
rect 18693 34561 18705 34595
rect 18739 34561 18751 34595
rect 18693 34555 18751 34561
rect 15749 34527 15807 34533
rect 15749 34524 15761 34527
rect 15212 34496 15761 34524
rect 14921 34487 14979 34493
rect 15749 34493 15761 34496
rect 15795 34524 15807 34527
rect 16853 34527 16911 34533
rect 16853 34524 16865 34527
rect 15795 34496 16865 34524
rect 15795 34493 15807 34496
rect 15749 34487 15807 34493
rect 16853 34493 16865 34496
rect 16899 34493 16911 34527
rect 16853 34487 16911 34493
rect 10870 34416 10876 34468
rect 10928 34456 10934 34468
rect 12084 34456 12112 34487
rect 12452 34456 12480 34487
rect 10928 34428 12480 34456
rect 10928 34416 10934 34428
rect 12526 34416 12532 34468
rect 12584 34456 12590 34468
rect 12713 34459 12771 34465
rect 12713 34456 12725 34459
rect 12584 34428 12725 34456
rect 12584 34416 12590 34428
rect 12713 34425 12725 34428
rect 12759 34425 12771 34459
rect 12713 34419 12771 34425
rect 14826 34416 14832 34468
rect 14884 34456 14890 34468
rect 14936 34456 14964 34487
rect 17310 34484 17316 34536
rect 17368 34524 17374 34536
rect 17589 34527 17647 34533
rect 17589 34524 17601 34527
rect 17368 34496 17601 34524
rect 17368 34484 17374 34496
rect 17589 34493 17601 34496
rect 17635 34493 17647 34527
rect 17589 34487 17647 34493
rect 18049 34527 18107 34533
rect 18049 34493 18061 34527
rect 18095 34524 18107 34527
rect 18138 34524 18144 34536
rect 18095 34496 18144 34524
rect 18095 34493 18107 34496
rect 18049 34487 18107 34493
rect 18138 34484 18144 34496
rect 18196 34524 18202 34536
rect 18432 34524 18460 34555
rect 18782 34552 18788 34604
rect 18840 34592 18846 34604
rect 18877 34595 18935 34601
rect 18877 34592 18889 34595
rect 18840 34564 18889 34592
rect 18840 34552 18846 34564
rect 18877 34561 18889 34564
rect 18923 34561 18935 34595
rect 18877 34555 18935 34561
rect 18966 34552 18972 34604
rect 19024 34552 19030 34604
rect 19058 34552 19064 34604
rect 19116 34592 19122 34604
rect 21542 34592 21548 34604
rect 19116 34564 21548 34592
rect 19116 34552 19122 34564
rect 21542 34552 21548 34564
rect 21600 34552 21606 34604
rect 22186 34552 22192 34604
rect 22244 34552 22250 34604
rect 22281 34595 22339 34601
rect 22281 34561 22293 34595
rect 22327 34561 22339 34595
rect 22281 34555 22339 34561
rect 19245 34527 19303 34533
rect 19245 34524 19257 34527
rect 18196 34496 19257 34524
rect 18196 34484 18202 34496
rect 19245 34493 19257 34496
rect 19291 34493 19303 34527
rect 19245 34487 19303 34493
rect 22002 34484 22008 34536
rect 22060 34524 22066 34536
rect 22296 34524 22324 34555
rect 22462 34552 22468 34604
rect 22520 34592 22526 34604
rect 22830 34592 22836 34604
rect 22520 34564 22836 34592
rect 22520 34552 22526 34564
rect 22830 34552 22836 34564
rect 22888 34552 22894 34604
rect 23198 34552 23204 34604
rect 23256 34552 23262 34604
rect 23293 34595 23351 34601
rect 23293 34561 23305 34595
rect 23339 34561 23351 34595
rect 23293 34555 23351 34561
rect 23308 34524 23336 34555
rect 23474 34552 23480 34604
rect 23532 34552 23538 34604
rect 25884 34601 25912 34632
rect 26326 34620 26332 34672
rect 26384 34660 26390 34672
rect 26384 34632 26556 34660
rect 26384 34620 26390 34632
rect 25593 34595 25651 34601
rect 25593 34561 25605 34595
rect 25639 34561 25651 34595
rect 25593 34555 25651 34561
rect 25869 34595 25927 34601
rect 25869 34561 25881 34595
rect 25915 34561 25927 34595
rect 25869 34555 25927 34561
rect 25961 34595 26019 34601
rect 25961 34561 25973 34595
rect 26007 34592 26019 34595
rect 26234 34592 26240 34604
rect 26007 34564 26240 34592
rect 26007 34561 26019 34564
rect 25961 34555 26019 34561
rect 25130 34524 25136 34536
rect 22060 34496 25136 34524
rect 22060 34484 22066 34496
rect 25130 34484 25136 34496
rect 25188 34484 25194 34536
rect 25608 34524 25636 34555
rect 26234 34552 26240 34564
rect 26292 34552 26298 34604
rect 26414 34595 26472 34601
rect 26414 34592 26426 34595
rect 26344 34564 26426 34592
rect 26344 34524 26372 34564
rect 26414 34561 26426 34564
rect 26460 34561 26472 34595
rect 26414 34555 26472 34561
rect 26528 34533 26556 34632
rect 25608 34496 26372 34524
rect 14884 34428 15700 34456
rect 14884 34416 14890 34428
rect 10008 34360 10824 34388
rect 10008 34348 10014 34360
rect 11882 34348 11888 34400
rect 11940 34388 11946 34400
rect 12345 34391 12403 34397
rect 12345 34388 12357 34391
rect 11940 34360 12357 34388
rect 11940 34348 11946 34360
rect 12345 34357 12357 34360
rect 12391 34357 12403 34391
rect 12345 34351 12403 34357
rect 12618 34348 12624 34400
rect 12676 34388 12682 34400
rect 13354 34388 13360 34400
rect 12676 34360 13360 34388
rect 12676 34348 12682 34360
rect 13354 34348 13360 34360
rect 13412 34348 13418 34400
rect 15378 34348 15384 34400
rect 15436 34348 15442 34400
rect 15470 34348 15476 34400
rect 15528 34348 15534 34400
rect 15672 34397 15700 34428
rect 18598 34416 18604 34468
rect 18656 34456 18662 34468
rect 19061 34459 19119 34465
rect 19061 34456 19073 34459
rect 18656 34428 19073 34456
rect 18656 34416 18662 34428
rect 19061 34425 19073 34428
rect 19107 34425 19119 34459
rect 19061 34419 19119 34425
rect 19150 34416 19156 34468
rect 19208 34456 19214 34468
rect 25608 34456 25636 34496
rect 19208 34428 25636 34456
rect 19208 34416 19214 34428
rect 25682 34416 25688 34468
rect 25740 34416 25746 34468
rect 26344 34456 26372 34496
rect 26513 34527 26571 34533
rect 26513 34493 26525 34527
rect 26559 34493 26571 34527
rect 26513 34487 26571 34493
rect 26786 34484 26792 34536
rect 26844 34484 26850 34536
rect 27522 34456 27528 34468
rect 26344 34428 27528 34456
rect 27522 34416 27528 34428
rect 27580 34416 27586 34468
rect 15657 34391 15715 34397
rect 15657 34357 15669 34391
rect 15703 34357 15715 34391
rect 15657 34351 15715 34357
rect 18233 34391 18291 34397
rect 18233 34357 18245 34391
rect 18279 34388 18291 34391
rect 18414 34388 18420 34400
rect 18279 34360 18420 34388
rect 18279 34357 18291 34360
rect 18233 34351 18291 34357
rect 18414 34348 18420 34360
rect 18472 34348 18478 34400
rect 23658 34348 23664 34400
rect 23716 34348 23722 34400
rect 26050 34348 26056 34400
rect 26108 34388 26114 34400
rect 26145 34391 26203 34397
rect 26145 34388 26157 34391
rect 26108 34360 26157 34388
rect 26108 34348 26114 34360
rect 26145 34357 26157 34360
rect 26191 34357 26203 34391
rect 26145 34351 26203 34357
rect 1104 34298 36524 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 36524 34298
rect 1104 34224 36524 34246
rect 10045 34187 10103 34193
rect 10045 34153 10057 34187
rect 10091 34184 10103 34187
rect 10226 34184 10232 34196
rect 10091 34156 10232 34184
rect 10091 34153 10103 34156
rect 10045 34147 10103 34153
rect 10226 34144 10232 34156
rect 10284 34144 10290 34196
rect 11517 34187 11575 34193
rect 11517 34153 11529 34187
rect 11563 34184 11575 34187
rect 12434 34184 12440 34196
rect 11563 34156 12440 34184
rect 11563 34153 11575 34156
rect 11517 34147 11575 34153
rect 12434 34144 12440 34156
rect 12492 34144 12498 34196
rect 16040 34156 16252 34184
rect 8938 34116 8944 34128
rect 8772 34088 8944 34116
rect 5534 34008 5540 34060
rect 5592 34048 5598 34060
rect 6362 34048 6368 34060
rect 5592 34020 6368 34048
rect 5592 34008 5598 34020
rect 6362 34008 6368 34020
rect 6420 34048 6426 34060
rect 6733 34051 6791 34057
rect 6733 34048 6745 34051
rect 6420 34020 6745 34048
rect 6420 34008 6426 34020
rect 6733 34017 6745 34020
rect 6779 34017 6791 34051
rect 6733 34011 6791 34017
rect 8662 34008 8668 34060
rect 8720 34048 8726 34060
rect 8772 34057 8800 34088
rect 8938 34076 8944 34088
rect 8996 34076 9002 34128
rect 10870 34076 10876 34128
rect 10928 34116 10934 34128
rect 10928 34088 11192 34116
rect 10928 34076 10934 34088
rect 8757 34051 8815 34057
rect 8757 34048 8769 34051
rect 8720 34020 8769 34048
rect 8720 34008 8726 34020
rect 8757 34017 8769 34020
rect 8803 34017 8815 34051
rect 8757 34011 8815 34017
rect 9490 34008 9496 34060
rect 9548 34048 9554 34060
rect 11164 34057 11192 34088
rect 10229 34051 10287 34057
rect 10229 34048 10241 34051
rect 9548 34020 10241 34048
rect 9548 34008 9554 34020
rect 10229 34017 10241 34020
rect 10275 34017 10287 34051
rect 10229 34011 10287 34017
rect 11149 34051 11207 34057
rect 11149 34017 11161 34051
rect 11195 34017 11207 34051
rect 11149 34011 11207 34017
rect 11977 34051 12035 34057
rect 11977 34017 11989 34051
rect 12023 34048 12035 34051
rect 15381 34051 15439 34057
rect 12023 34020 15332 34048
rect 12023 34017 12035 34020
rect 11977 34011 12035 34017
rect 8846 33940 8852 33992
rect 8904 33980 8910 33992
rect 8941 33983 8999 33989
rect 8941 33980 8953 33983
rect 8904 33952 8953 33980
rect 8904 33940 8910 33952
rect 8941 33949 8953 33952
rect 8987 33949 8999 33983
rect 8941 33943 8999 33949
rect 9401 33983 9459 33989
rect 9401 33949 9413 33983
rect 9447 33949 9459 33983
rect 9401 33943 9459 33949
rect 9886 33983 9944 33989
rect 9886 33949 9898 33983
rect 9932 33980 9944 33983
rect 10042 33980 10048 33992
rect 9932 33952 10048 33980
rect 9932 33949 9944 33952
rect 9886 33943 9944 33949
rect 7006 33872 7012 33924
rect 7064 33872 7070 33924
rect 9416 33912 9444 33943
rect 10042 33940 10048 33952
rect 10100 33940 10106 33992
rect 10134 33940 10140 33992
rect 10192 33940 10198 33992
rect 10778 33940 10784 33992
rect 10836 33980 10842 33992
rect 10873 33983 10931 33989
rect 10873 33980 10885 33983
rect 10836 33952 10885 33980
rect 10836 33940 10842 33952
rect 10873 33949 10885 33952
rect 10919 33949 10931 33983
rect 11606 33980 11612 33992
rect 10873 33943 10931 33949
rect 11164 33952 11612 33980
rect 10796 33912 10824 33940
rect 8234 33884 9168 33912
rect 9416 33884 10824 33912
rect 7926 33804 7932 33856
rect 7984 33844 7990 33856
rect 8312 33844 8340 33884
rect 9140 33853 9168 33884
rect 7984 33816 8340 33844
rect 9125 33847 9183 33853
rect 7984 33804 7990 33816
rect 9125 33813 9137 33847
rect 9171 33813 9183 33847
rect 9125 33807 9183 33813
rect 9674 33804 9680 33856
rect 9732 33804 9738 33856
rect 9766 33804 9772 33856
rect 9824 33804 9830 33856
rect 10226 33804 10232 33856
rect 10284 33844 10290 33856
rect 11164 33844 11192 33952
rect 11606 33940 11612 33952
rect 11664 33940 11670 33992
rect 11882 33940 11888 33992
rect 11940 33940 11946 33992
rect 12066 33940 12072 33992
rect 12124 33940 12130 33992
rect 14185 33983 14243 33989
rect 14185 33949 14197 33983
rect 14231 33980 14243 33983
rect 14645 33983 14703 33989
rect 14645 33980 14657 33983
rect 14231 33952 14657 33980
rect 14231 33949 14243 33952
rect 14185 33943 14243 33949
rect 14645 33949 14657 33952
rect 14691 33949 14703 33983
rect 14645 33943 14703 33949
rect 14734 33940 14740 33992
rect 14792 33980 14798 33992
rect 14829 33983 14887 33989
rect 14829 33980 14841 33983
rect 14792 33952 14841 33980
rect 14792 33940 14798 33952
rect 14829 33949 14841 33952
rect 14875 33949 14887 33983
rect 14829 33943 14887 33949
rect 14918 33940 14924 33992
rect 14976 33940 14982 33992
rect 15013 33983 15071 33989
rect 15013 33949 15025 33983
rect 15059 33980 15071 33983
rect 15102 33980 15108 33992
rect 15059 33952 15108 33980
rect 15059 33949 15071 33952
rect 15013 33943 15071 33949
rect 15102 33940 15108 33952
rect 15160 33940 15166 33992
rect 15194 33940 15200 33992
rect 15252 33940 15258 33992
rect 15304 33980 15332 34020
rect 15381 34017 15393 34051
rect 15427 34048 15439 34051
rect 16040 34048 16068 34156
rect 15427 34020 16068 34048
rect 16224 34048 16252 34156
rect 17218 34144 17224 34196
rect 17276 34184 17282 34196
rect 17276 34156 17908 34184
rect 17276 34144 17282 34156
rect 17880 34116 17908 34156
rect 17954 34144 17960 34196
rect 18012 34144 18018 34196
rect 18322 34144 18328 34196
rect 18380 34184 18386 34196
rect 19058 34184 19064 34196
rect 18380 34156 19064 34184
rect 18380 34144 18386 34156
rect 19058 34144 19064 34156
rect 19116 34144 19122 34196
rect 19702 34184 19708 34196
rect 19306 34156 19708 34184
rect 19306 34116 19334 34156
rect 19702 34144 19708 34156
rect 19760 34184 19766 34196
rect 20806 34184 20812 34196
rect 19760 34156 20812 34184
rect 19760 34144 19766 34156
rect 20806 34144 20812 34156
rect 20864 34144 20870 34196
rect 23109 34187 23167 34193
rect 23109 34153 23121 34187
rect 23155 34184 23167 34187
rect 23198 34184 23204 34196
rect 23155 34156 23204 34184
rect 23155 34153 23167 34156
rect 23109 34147 23167 34153
rect 23198 34144 23204 34156
rect 23256 34144 23262 34196
rect 27522 34144 27528 34196
rect 27580 34144 27586 34196
rect 17880 34088 19334 34116
rect 20548 34088 20944 34116
rect 17221 34051 17279 34057
rect 17221 34048 17233 34051
rect 16224 34020 17233 34048
rect 15427 34017 15439 34020
rect 15381 34011 15439 34017
rect 17221 34017 17233 34020
rect 17267 34017 17279 34051
rect 17221 34011 17279 34017
rect 17497 34051 17555 34057
rect 17497 34017 17509 34051
rect 17543 34048 17555 34051
rect 18322 34048 18328 34060
rect 17543 34020 18328 34048
rect 17543 34017 17555 34020
rect 17497 34011 17555 34017
rect 18322 34008 18328 34020
rect 18380 34008 18386 34060
rect 15304 33952 15976 33980
rect 11330 33872 11336 33924
rect 11388 33921 11394 33924
rect 11388 33915 11416 33921
rect 11404 33912 11416 33915
rect 11974 33912 11980 33924
rect 11404 33884 11980 33912
rect 11404 33881 11416 33884
rect 11388 33875 11416 33881
rect 11388 33872 11394 33875
rect 11974 33872 11980 33884
rect 12032 33912 12038 33924
rect 12342 33912 12348 33924
rect 12032 33884 12348 33912
rect 12032 33872 12038 33884
rect 12342 33872 12348 33884
rect 12400 33872 12406 33924
rect 13354 33872 13360 33924
rect 13412 33912 13418 33924
rect 14369 33915 14427 33921
rect 14369 33912 14381 33915
rect 13412 33884 14381 33912
rect 13412 33872 13418 33884
rect 14369 33881 14381 33884
rect 14415 33881 14427 33915
rect 14369 33875 14427 33881
rect 10284 33816 11192 33844
rect 10284 33804 10290 33816
rect 11238 33804 11244 33856
rect 11296 33804 11302 33856
rect 14384 33844 14412 33875
rect 14550 33872 14556 33924
rect 14608 33872 14614 33924
rect 15473 33915 15531 33921
rect 15473 33912 15485 33915
rect 15212 33884 15485 33912
rect 15212 33844 15240 33884
rect 15473 33881 15485 33884
rect 15519 33912 15531 33915
rect 15838 33912 15844 33924
rect 15519 33884 15844 33912
rect 15519 33881 15531 33884
rect 15473 33875 15531 33881
rect 15838 33872 15844 33884
rect 15896 33872 15902 33924
rect 14384 33816 15240 33844
rect 15948 33844 15976 33952
rect 17586 33940 17592 33992
rect 17644 33940 17650 33992
rect 17770 33940 17776 33992
rect 17828 33940 17834 33992
rect 18414 33940 18420 33992
rect 18472 33940 18478 33992
rect 18506 33940 18512 33992
rect 18564 33980 18570 33992
rect 18800 33989 18828 34088
rect 19058 34008 19064 34060
rect 19116 34048 19122 34060
rect 19245 34051 19303 34057
rect 19245 34048 19257 34051
rect 19116 34020 19257 34048
rect 19116 34008 19122 34020
rect 19245 34017 19257 34020
rect 19291 34048 19303 34051
rect 20548 34048 20576 34088
rect 19291 34020 20576 34048
rect 20916 34048 20944 34088
rect 21174 34076 21180 34128
rect 21232 34116 21238 34128
rect 21634 34116 21640 34128
rect 21232 34088 21640 34116
rect 21232 34076 21238 34088
rect 21634 34076 21640 34088
rect 21692 34076 21698 34128
rect 23014 34116 23020 34128
rect 22066 34088 23020 34116
rect 22066 34048 22094 34088
rect 23014 34076 23020 34088
rect 23072 34116 23078 34128
rect 24946 34116 24952 34128
rect 23072 34088 24952 34116
rect 23072 34076 23078 34088
rect 20916 34020 22094 34048
rect 19291 34017 19303 34020
rect 19245 34011 19303 34017
rect 22462 34008 22468 34060
rect 22520 34048 22526 34060
rect 22649 34051 22707 34057
rect 22649 34048 22661 34051
rect 22520 34020 22661 34048
rect 22520 34008 22526 34020
rect 22649 34017 22661 34020
rect 22695 34017 22707 34051
rect 22649 34011 22707 34017
rect 18785 33983 18843 33989
rect 18564 33952 18609 33980
rect 18564 33940 18570 33952
rect 18785 33949 18797 33983
rect 18831 33949 18843 33983
rect 18785 33943 18843 33949
rect 18882 33983 18940 33989
rect 18882 33949 18894 33983
rect 18928 33949 18940 33983
rect 18882 33943 18940 33949
rect 16482 33872 16488 33924
rect 16540 33872 16546 33924
rect 18693 33915 18751 33921
rect 18693 33912 18705 33915
rect 16868 33884 18705 33912
rect 16868 33844 16896 33884
rect 18693 33881 18705 33884
rect 18739 33881 18751 33915
rect 18693 33875 18751 33881
rect 18892 33912 18920 33943
rect 20806 33940 20812 33992
rect 20864 33980 20870 33992
rect 21269 33983 21327 33989
rect 21269 33980 21281 33983
rect 20864 33952 21281 33980
rect 20864 33940 20870 33952
rect 21269 33949 21281 33952
rect 21315 33949 21327 33983
rect 21269 33943 21327 33949
rect 21726 33940 21732 33992
rect 21784 33980 21790 33992
rect 21821 33983 21879 33989
rect 21821 33980 21833 33983
rect 21784 33952 21833 33980
rect 21784 33940 21790 33952
rect 21821 33949 21833 33952
rect 21867 33949 21879 33983
rect 21821 33943 21879 33949
rect 21910 33940 21916 33992
rect 21968 33940 21974 33992
rect 22554 33940 22560 33992
rect 22612 33980 22618 33992
rect 23492 33989 23520 34088
rect 24946 34076 24952 34088
rect 25004 34116 25010 34128
rect 25004 34088 25820 34116
rect 25004 34076 25010 34088
rect 25792 34057 25820 34088
rect 25777 34051 25835 34057
rect 25777 34017 25789 34051
rect 25823 34017 25835 34051
rect 25777 34011 25835 34017
rect 26050 34008 26056 34060
rect 26108 34008 26114 34060
rect 22741 33983 22799 33989
rect 22741 33980 22753 33983
rect 22612 33952 22753 33980
rect 22612 33940 22618 33952
rect 22741 33949 22753 33952
rect 22787 33949 22799 33983
rect 22741 33943 22799 33949
rect 23477 33983 23535 33989
rect 23477 33949 23489 33983
rect 23523 33949 23535 33983
rect 23477 33943 23535 33949
rect 19426 33912 19432 33924
rect 18892 33884 19432 33912
rect 15948 33816 16896 33844
rect 17494 33804 17500 33856
rect 17552 33844 17558 33856
rect 18892 33844 18920 33884
rect 19426 33872 19432 33884
rect 19484 33872 19490 33924
rect 19528 33915 19586 33921
rect 19528 33881 19540 33915
rect 19574 33912 19586 33915
rect 19794 33912 19800 33924
rect 19574 33884 19800 33912
rect 19574 33881 19586 33884
rect 19528 33875 19586 33881
rect 19794 33872 19800 33884
rect 19852 33872 19858 33924
rect 20254 33872 20260 33924
rect 20312 33872 20318 33924
rect 21542 33872 21548 33924
rect 21600 33912 21606 33924
rect 21928 33912 21956 33940
rect 21600 33884 21956 33912
rect 21600 33872 21606 33884
rect 24118 33872 24124 33924
rect 24176 33872 24182 33924
rect 26602 33872 26608 33924
rect 26660 33872 26666 33924
rect 17552 33816 18920 33844
rect 19061 33847 19119 33853
rect 17552 33804 17558 33816
rect 19061 33813 19073 33847
rect 19107 33844 19119 33847
rect 19334 33844 19340 33856
rect 19107 33816 19340 33844
rect 19107 33813 19119 33816
rect 19061 33807 19119 33813
rect 19334 33804 19340 33816
rect 19392 33804 19398 33856
rect 22186 33804 22192 33856
rect 22244 33844 22250 33856
rect 23566 33844 23572 33856
rect 22244 33816 23572 33844
rect 22244 33804 22250 33816
rect 23566 33804 23572 33816
rect 23624 33844 23630 33856
rect 23842 33844 23848 33856
rect 23624 33816 23848 33844
rect 23624 33804 23630 33816
rect 23842 33804 23848 33816
rect 23900 33804 23906 33856
rect 24026 33804 24032 33856
rect 24084 33804 24090 33856
rect 1104 33754 36524 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 36524 33754
rect 1104 33680 36524 33702
rect 7006 33600 7012 33652
rect 7064 33640 7070 33652
rect 8849 33643 8907 33649
rect 8849 33640 8861 33643
rect 7064 33612 8861 33640
rect 7064 33600 7070 33612
rect 8849 33609 8861 33612
rect 8895 33609 8907 33643
rect 8849 33603 8907 33609
rect 9585 33643 9643 33649
rect 9585 33609 9597 33643
rect 9631 33640 9643 33643
rect 9766 33640 9772 33652
rect 9631 33612 9772 33640
rect 9631 33609 9643 33612
rect 9585 33603 9643 33609
rect 9766 33600 9772 33612
rect 9824 33600 9830 33652
rect 11054 33600 11060 33652
rect 11112 33640 11118 33652
rect 11717 33643 11775 33649
rect 11717 33640 11729 33643
rect 11112 33612 11729 33640
rect 11112 33600 11118 33612
rect 11717 33609 11729 33612
rect 11763 33609 11775 33643
rect 11717 33603 11775 33609
rect 11885 33643 11943 33649
rect 11885 33609 11897 33643
rect 11931 33640 11943 33643
rect 12066 33640 12072 33652
rect 11931 33612 12072 33640
rect 11931 33609 11943 33612
rect 11885 33603 11943 33609
rect 12066 33600 12072 33612
rect 12124 33600 12130 33652
rect 13648 33612 14780 33640
rect 7926 33572 7932 33584
rect 7866 33544 7932 33572
rect 7926 33532 7932 33544
rect 7984 33532 7990 33584
rect 9490 33532 9496 33584
rect 9548 33572 9554 33584
rect 9953 33575 10011 33581
rect 9953 33572 9965 33575
rect 9548 33544 9965 33572
rect 9548 33532 9554 33544
rect 9953 33541 9965 33544
rect 9999 33541 10011 33575
rect 9953 33535 10011 33541
rect 10137 33575 10195 33581
rect 10137 33541 10149 33575
rect 10183 33572 10195 33575
rect 10870 33572 10876 33584
rect 10183 33544 10876 33572
rect 10183 33541 10195 33544
rect 10137 33535 10195 33541
rect 10870 33532 10876 33544
rect 10928 33572 10934 33584
rect 10928 33544 11468 33572
rect 10928 33532 10934 33544
rect 6362 33464 6368 33516
rect 6420 33464 6426 33516
rect 8478 33464 8484 33516
rect 8536 33464 8542 33516
rect 8662 33464 8668 33516
rect 8720 33464 8726 33516
rect 8757 33507 8815 33513
rect 8757 33473 8769 33507
rect 8803 33473 8815 33507
rect 8757 33467 8815 33473
rect 8941 33507 8999 33513
rect 8941 33473 8953 33507
rect 8987 33473 8999 33507
rect 8941 33467 8999 33473
rect 9769 33507 9827 33513
rect 9769 33473 9781 33507
rect 9815 33473 9827 33507
rect 9769 33467 9827 33473
rect 9861 33507 9919 33513
rect 9861 33473 9873 33507
rect 9907 33504 9919 33507
rect 9907 33476 10364 33504
rect 9907 33473 9919 33476
rect 9861 33467 9919 33473
rect 6641 33439 6699 33445
rect 6641 33405 6653 33439
rect 6687 33436 6699 33439
rect 7006 33436 7012 33448
rect 6687 33408 7012 33436
rect 6687 33405 6699 33408
rect 6641 33399 6699 33405
rect 7006 33396 7012 33408
rect 7064 33396 7070 33448
rect 7834 33396 7840 33448
rect 7892 33436 7898 33448
rect 8389 33439 8447 33445
rect 8389 33436 8401 33439
rect 7892 33408 8401 33436
rect 7892 33396 7898 33408
rect 8389 33405 8401 33408
rect 8435 33405 8447 33439
rect 8389 33399 8447 33405
rect 8573 33439 8631 33445
rect 8573 33405 8585 33439
rect 8619 33436 8631 33439
rect 8772 33436 8800 33467
rect 8619 33408 8800 33436
rect 8619 33405 8631 33408
rect 8573 33399 8631 33405
rect 8956 33300 8984 33467
rect 9784 33436 9812 33467
rect 10226 33436 10232 33448
rect 9784 33408 10232 33436
rect 10226 33396 10232 33408
rect 10284 33396 10290 33448
rect 10336 33368 10364 33476
rect 11054 33464 11060 33516
rect 11112 33464 11118 33516
rect 11149 33507 11207 33513
rect 11149 33473 11161 33507
rect 11195 33504 11207 33507
rect 11195 33476 11284 33504
rect 11195 33473 11207 33476
rect 11149 33467 11207 33473
rect 11146 33368 11152 33380
rect 10336 33340 11152 33368
rect 11146 33328 11152 33340
rect 11204 33328 11210 33380
rect 10962 33300 10968 33312
rect 8956 33272 10968 33300
rect 10962 33260 10968 33272
rect 11020 33260 11026 33312
rect 11256 33300 11284 33476
rect 11330 33464 11336 33516
rect 11388 33464 11394 33516
rect 11440 33436 11468 33544
rect 11514 33532 11520 33584
rect 11572 33572 11578 33584
rect 12253 33575 12311 33581
rect 11572 33544 12020 33572
rect 11572 33532 11578 33544
rect 11992 33513 12020 33544
rect 12253 33541 12265 33575
rect 12299 33572 12311 33575
rect 12618 33572 12624 33584
rect 12299 33544 12624 33572
rect 12299 33541 12311 33544
rect 12253 33535 12311 33541
rect 12618 33532 12624 33544
rect 12676 33532 12682 33584
rect 13648 33572 13676 33612
rect 13570 33544 13676 33572
rect 13722 33532 13728 33584
rect 13780 33572 13786 33584
rect 13780 33544 14320 33572
rect 13780 33532 13786 33544
rect 11977 33507 12035 33513
rect 11977 33473 11989 33507
rect 12023 33504 12035 33507
rect 12342 33504 12348 33516
rect 12023 33476 12348 33504
rect 12023 33473 12035 33476
rect 11977 33467 12035 33473
rect 12342 33464 12348 33476
rect 12400 33464 12406 33516
rect 14292 33513 14320 33544
rect 14277 33507 14335 33513
rect 14277 33473 14289 33507
rect 14323 33473 14335 33507
rect 14277 33467 14335 33473
rect 14550 33464 14556 33516
rect 14608 33504 14614 33516
rect 14645 33507 14703 33513
rect 14645 33504 14657 33507
rect 14608 33476 14657 33504
rect 14608 33464 14614 33476
rect 14645 33473 14657 33476
rect 14691 33473 14703 33507
rect 14752 33504 14780 33612
rect 14826 33600 14832 33652
rect 14884 33600 14890 33652
rect 15102 33600 15108 33652
rect 15160 33600 15166 33652
rect 16758 33600 16764 33652
rect 16816 33640 16822 33652
rect 16945 33643 17003 33649
rect 16945 33640 16957 33643
rect 16816 33612 16957 33640
rect 16816 33600 16822 33612
rect 16945 33609 16957 33612
rect 16991 33609 17003 33643
rect 16945 33603 17003 33609
rect 17034 33600 17040 33652
rect 17092 33640 17098 33652
rect 17770 33640 17776 33652
rect 17092 33612 17776 33640
rect 17092 33600 17098 33612
rect 17770 33600 17776 33612
rect 17828 33600 17834 33652
rect 18506 33600 18512 33652
rect 18564 33640 18570 33652
rect 22002 33640 22008 33652
rect 18564 33612 22008 33640
rect 18564 33600 18570 33612
rect 15378 33532 15384 33584
rect 15436 33572 15442 33584
rect 15565 33575 15623 33581
rect 15565 33572 15577 33575
rect 15436 33544 15577 33572
rect 15436 33532 15442 33544
rect 15565 33541 15577 33544
rect 15611 33572 15623 33575
rect 18598 33572 18604 33584
rect 15611 33544 18604 33572
rect 15611 33541 15623 33544
rect 15565 33535 15623 33541
rect 18598 33532 18604 33544
rect 18656 33532 18662 33584
rect 20898 33532 20904 33584
rect 20956 33572 20962 33584
rect 21542 33572 21548 33584
rect 20956 33544 21548 33572
rect 20956 33532 20962 33544
rect 16022 33504 16028 33516
rect 14752 33476 16028 33504
rect 14645 33467 14703 33473
rect 16022 33464 16028 33476
rect 16080 33464 16086 33516
rect 16853 33507 16911 33513
rect 16853 33473 16865 33507
rect 16899 33504 16911 33507
rect 16942 33504 16948 33516
rect 16899 33476 16948 33504
rect 16899 33473 16911 33476
rect 16853 33467 16911 33473
rect 16942 33464 16948 33476
rect 17000 33464 17006 33516
rect 17037 33507 17095 33513
rect 17037 33473 17049 33507
rect 17083 33504 17095 33507
rect 17586 33504 17592 33516
rect 17083 33476 17592 33504
rect 17083 33473 17095 33476
rect 17037 33467 17095 33473
rect 12069 33439 12127 33445
rect 12069 33436 12081 33439
rect 11440 33408 12081 33436
rect 12069 33405 12081 33408
rect 12115 33405 12127 33439
rect 12069 33399 12127 33405
rect 13998 33396 14004 33448
rect 14056 33396 14062 33448
rect 14461 33439 14519 33445
rect 14461 33405 14473 33439
rect 14507 33436 14519 33439
rect 14507 33408 14688 33436
rect 14507 33405 14519 33408
rect 14461 33399 14519 33405
rect 14660 33380 14688 33408
rect 15194 33396 15200 33448
rect 15252 33436 15258 33448
rect 15252 33408 15608 33436
rect 15252 33396 15258 33408
rect 15580 33380 15608 33408
rect 15838 33396 15844 33448
rect 15896 33436 15902 33448
rect 17052 33436 17080 33467
rect 17586 33464 17592 33476
rect 17644 33464 17650 33516
rect 21376 33513 21404 33544
rect 21542 33532 21548 33544
rect 21600 33532 21606 33584
rect 21177 33507 21235 33513
rect 21177 33473 21189 33507
rect 21223 33473 21235 33507
rect 21177 33467 21235 33473
rect 21361 33507 21419 33513
rect 21361 33473 21373 33507
rect 21407 33473 21419 33507
rect 21361 33467 21419 33473
rect 21637 33507 21695 33513
rect 21637 33473 21649 33507
rect 21683 33473 21695 33507
rect 21744 33504 21772 33612
rect 22002 33600 22008 33612
rect 22060 33600 22066 33652
rect 23017 33643 23075 33649
rect 23017 33609 23029 33643
rect 23063 33640 23075 33643
rect 23474 33640 23480 33652
rect 23063 33612 23480 33640
rect 23063 33609 23075 33612
rect 23017 33603 23075 33609
rect 23474 33600 23480 33612
rect 23532 33600 23538 33652
rect 21910 33532 21916 33584
rect 21968 33572 21974 33584
rect 22741 33575 22799 33581
rect 22741 33572 22753 33575
rect 21968 33544 22753 33572
rect 21968 33532 21974 33544
rect 22741 33541 22753 33544
rect 22787 33572 22799 33575
rect 23385 33575 23443 33581
rect 22787 33544 22968 33572
rect 22787 33541 22799 33544
rect 22741 33535 22799 33541
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 21744 33476 21833 33504
rect 21637 33467 21695 33473
rect 21821 33473 21833 33476
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 22097 33507 22155 33513
rect 22097 33473 22109 33507
rect 22143 33473 22155 33507
rect 22097 33467 22155 33473
rect 15896 33408 17080 33436
rect 15896 33396 15902 33408
rect 11333 33371 11391 33377
rect 11333 33337 11345 33371
rect 11379 33368 11391 33371
rect 11882 33368 11888 33380
rect 11379 33340 11888 33368
rect 11379 33337 11391 33340
rect 11333 33331 11391 33337
rect 11882 33328 11888 33340
rect 11940 33328 11946 33380
rect 14642 33328 14648 33380
rect 14700 33328 14706 33380
rect 15289 33371 15347 33377
rect 15289 33337 15301 33371
rect 15335 33368 15347 33371
rect 15470 33368 15476 33380
rect 15335 33340 15476 33368
rect 15335 33337 15347 33340
rect 15289 33331 15347 33337
rect 15470 33328 15476 33340
rect 15528 33328 15534 33380
rect 15562 33328 15568 33380
rect 15620 33368 15626 33380
rect 16114 33368 16120 33380
rect 15620 33340 16120 33368
rect 15620 33328 15626 33340
rect 16114 33328 16120 33340
rect 16172 33368 16178 33380
rect 21192 33368 21220 33467
rect 21652 33436 21680 33467
rect 21726 33436 21732 33448
rect 21652 33408 21732 33436
rect 21726 33396 21732 33408
rect 21784 33436 21790 33448
rect 22112 33436 22140 33467
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 22465 33507 22523 33513
rect 22465 33504 22477 33507
rect 22428 33476 22477 33504
rect 22428 33464 22434 33476
rect 22465 33473 22477 33476
rect 22511 33473 22523 33507
rect 22465 33467 22523 33473
rect 22646 33464 22652 33516
rect 22704 33464 22710 33516
rect 22830 33464 22836 33516
rect 22888 33464 22894 33516
rect 22738 33436 22744 33448
rect 21784 33408 22744 33436
rect 21784 33396 21790 33408
rect 22738 33396 22744 33408
rect 22796 33396 22802 33448
rect 22940 33436 22968 33544
rect 23385 33541 23397 33575
rect 23431 33572 23443 33575
rect 23658 33572 23664 33584
rect 23431 33544 23664 33572
rect 23431 33541 23443 33544
rect 23385 33535 23443 33541
rect 23658 33532 23664 33544
rect 23716 33532 23722 33584
rect 24670 33572 24676 33584
rect 24610 33544 24676 33572
rect 24670 33532 24676 33544
rect 24728 33532 24734 33584
rect 25130 33532 25136 33584
rect 25188 33572 25194 33584
rect 25225 33575 25283 33581
rect 25225 33572 25237 33575
rect 25188 33544 25237 33572
rect 25188 33532 25194 33544
rect 25225 33541 25237 33544
rect 25271 33541 25283 33575
rect 25225 33535 25283 33541
rect 25409 33575 25467 33581
rect 25409 33541 25421 33575
rect 25455 33572 25467 33575
rect 25682 33572 25688 33584
rect 25455 33544 25688 33572
rect 25455 33541 25467 33544
rect 25409 33535 25467 33541
rect 25682 33532 25688 33544
rect 25740 33532 25746 33584
rect 23014 33464 23020 33516
rect 23072 33504 23078 33516
rect 23109 33507 23167 33513
rect 23109 33504 23121 33507
rect 23072 33476 23121 33504
rect 23072 33464 23078 33476
rect 23109 33473 23121 33476
rect 23155 33473 23167 33507
rect 23109 33467 23167 33473
rect 25038 33464 25044 33516
rect 25096 33464 25102 33516
rect 24394 33436 24400 33448
rect 22940 33408 24400 33436
rect 24394 33396 24400 33408
rect 24452 33436 24458 33448
rect 24857 33439 24915 33445
rect 24857 33436 24869 33439
rect 24452 33408 24869 33436
rect 24452 33396 24458 33408
rect 24857 33405 24869 33408
rect 24903 33436 24915 33439
rect 25682 33436 25688 33448
rect 24903 33408 25688 33436
rect 24903 33405 24915 33408
rect 24857 33399 24915 33405
rect 25682 33396 25688 33408
rect 25740 33396 25746 33448
rect 16172 33340 21128 33368
rect 21192 33340 21680 33368
rect 16172 33328 16178 33340
rect 11701 33303 11759 33309
rect 11701 33300 11713 33303
rect 11256 33272 11713 33300
rect 11701 33269 11713 33272
rect 11747 33300 11759 33303
rect 11790 33300 11796 33312
rect 11747 33272 11796 33300
rect 11747 33269 11759 33272
rect 11701 33263 11759 33269
rect 11790 33260 11796 33272
rect 11848 33260 11854 33312
rect 14918 33260 14924 33312
rect 14976 33300 14982 33312
rect 15654 33300 15660 33312
rect 14976 33272 15660 33300
rect 14976 33260 14982 33272
rect 15654 33260 15660 33272
rect 15712 33300 15718 33312
rect 18138 33300 18144 33312
rect 15712 33272 18144 33300
rect 15712 33260 15718 33272
rect 18138 33260 18144 33272
rect 18196 33300 18202 33312
rect 20898 33300 20904 33312
rect 18196 33272 20904 33300
rect 18196 33260 18202 33272
rect 20898 33260 20904 33272
rect 20956 33300 20962 33312
rect 20993 33303 21051 33309
rect 20993 33300 21005 33303
rect 20956 33272 21005 33300
rect 20956 33260 20962 33272
rect 20993 33269 21005 33272
rect 21039 33269 21051 33303
rect 21100 33300 21128 33340
rect 21545 33303 21603 33309
rect 21545 33300 21557 33303
rect 21100 33272 21557 33300
rect 20993 33263 21051 33269
rect 21545 33269 21557 33272
rect 21591 33269 21603 33303
rect 21652 33300 21680 33340
rect 21818 33328 21824 33380
rect 21876 33368 21882 33380
rect 22097 33371 22155 33377
rect 22097 33368 22109 33371
rect 21876 33340 22109 33368
rect 21876 33328 21882 33340
rect 22097 33337 22109 33340
rect 22143 33337 22155 33371
rect 22097 33331 22155 33337
rect 22186 33300 22192 33312
rect 21652 33272 22192 33300
rect 21545 33263 21603 33269
rect 22186 33260 22192 33272
rect 22244 33260 22250 33312
rect 22738 33260 22744 33312
rect 22796 33300 22802 33312
rect 25038 33300 25044 33312
rect 22796 33272 25044 33300
rect 22796 33260 22802 33272
rect 25038 33260 25044 33272
rect 25096 33260 25102 33312
rect 1104 33210 36524 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 36524 33210
rect 1104 33136 36524 33158
rect 7006 33056 7012 33108
rect 7064 33056 7070 33108
rect 9674 33056 9680 33108
rect 9732 33096 9738 33108
rect 10686 33096 10692 33108
rect 9732 33068 10692 33096
rect 9732 33056 9738 33068
rect 10686 33056 10692 33068
rect 10744 33056 10750 33108
rect 10870 33056 10876 33108
rect 10928 33056 10934 33108
rect 11054 33056 11060 33108
rect 11112 33096 11118 33108
rect 11149 33099 11207 33105
rect 11149 33096 11161 33099
rect 11112 33068 11161 33096
rect 11112 33056 11118 33068
rect 11149 33065 11161 33068
rect 11195 33065 11207 33099
rect 11149 33059 11207 33065
rect 11238 33056 11244 33108
rect 11296 33056 11302 33108
rect 13449 33099 13507 33105
rect 13449 33065 13461 33099
rect 13495 33096 13507 33099
rect 13998 33096 14004 33108
rect 13495 33068 14004 33096
rect 13495 33065 13507 33068
rect 13449 33059 13507 33065
rect 13998 33056 14004 33068
rect 14056 33056 14062 33108
rect 18322 33096 18328 33108
rect 14936 33068 18328 33096
rect 8294 33028 8300 33040
rect 7668 33000 8300 33028
rect 7668 32969 7696 33000
rect 8294 32988 8300 33000
rect 8352 33028 8358 33040
rect 8478 33028 8484 33040
rect 8352 33000 8484 33028
rect 8352 32988 8358 33000
rect 8478 32988 8484 33000
rect 8536 33028 8542 33040
rect 14936 33028 14964 33068
rect 18322 33056 18328 33068
rect 18380 33056 18386 33108
rect 18782 33096 18788 33108
rect 18708 33068 18788 33096
rect 8536 33000 14964 33028
rect 8536 32988 8542 33000
rect 7653 32963 7711 32969
rect 7653 32929 7665 32963
rect 7699 32929 7711 32963
rect 7653 32923 7711 32929
rect 10888 32932 11468 32960
rect 10888 32904 10916 32932
rect 7469 32895 7527 32901
rect 7469 32861 7481 32895
rect 7515 32892 7527 32895
rect 7834 32892 7840 32904
rect 7515 32864 7840 32892
rect 7515 32861 7527 32864
rect 7469 32855 7527 32861
rect 7834 32852 7840 32864
rect 7892 32852 7898 32904
rect 10781 32895 10839 32901
rect 10781 32861 10793 32895
rect 10827 32861 10839 32895
rect 10781 32855 10839 32861
rect 10796 32824 10824 32855
rect 10870 32852 10876 32904
rect 10928 32852 10934 32904
rect 11440 32901 11468 32932
rect 12618 32920 12624 32972
rect 12676 32960 12682 32972
rect 13280 32969 13308 33000
rect 15010 32988 15016 33040
rect 15068 33028 15074 33040
rect 18506 33028 18512 33040
rect 15068 33000 15700 33028
rect 15068 32988 15074 33000
rect 13173 32963 13231 32969
rect 13173 32960 13185 32963
rect 12676 32932 13185 32960
rect 12676 32920 12682 32932
rect 13173 32929 13185 32932
rect 13219 32929 13231 32963
rect 13173 32923 13231 32929
rect 13265 32963 13323 32969
rect 13265 32929 13277 32963
rect 13311 32929 13323 32963
rect 15289 32963 15347 32969
rect 13265 32923 13323 32929
rect 14292 32932 15240 32960
rect 11241 32895 11299 32901
rect 11241 32861 11253 32895
rect 11287 32861 11299 32895
rect 11241 32855 11299 32861
rect 11425 32895 11483 32901
rect 11425 32861 11437 32895
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 11054 32824 11060 32836
rect 10796 32796 11060 32824
rect 11054 32784 11060 32796
rect 11112 32824 11118 32836
rect 11256 32824 11284 32855
rect 11112 32796 11284 32824
rect 12805 32827 12863 32833
rect 11112 32784 11118 32796
rect 12805 32793 12817 32827
rect 12851 32824 12863 32827
rect 14292 32824 14320 32932
rect 14369 32895 14427 32901
rect 14369 32861 14381 32895
rect 14415 32861 14427 32895
rect 14369 32855 14427 32861
rect 12851 32796 14320 32824
rect 12851 32793 12863 32796
rect 12805 32787 12863 32793
rect 7377 32759 7435 32765
rect 7377 32725 7389 32759
rect 7423 32756 7435 32759
rect 9122 32756 9128 32768
rect 7423 32728 9128 32756
rect 7423 32725 7435 32728
rect 7377 32719 7435 32725
rect 9122 32716 9128 32728
rect 9180 32716 9186 32768
rect 14384 32756 14412 32855
rect 14550 32852 14556 32904
rect 14608 32852 14614 32904
rect 14645 32895 14703 32901
rect 14645 32861 14657 32895
rect 14691 32861 14703 32895
rect 14645 32855 14703 32861
rect 14461 32827 14519 32833
rect 14461 32793 14473 32827
rect 14507 32824 14519 32827
rect 14660 32824 14688 32855
rect 14826 32852 14832 32904
rect 14884 32852 14890 32904
rect 14921 32895 14979 32901
rect 14921 32861 14933 32895
rect 14967 32892 14979 32895
rect 15010 32892 15016 32904
rect 14967 32864 15016 32892
rect 14967 32861 14979 32864
rect 14921 32855 14979 32861
rect 15010 32852 15016 32864
rect 15068 32852 15074 32904
rect 15105 32895 15163 32901
rect 15105 32861 15117 32895
rect 15151 32861 15163 32895
rect 15212 32892 15240 32932
rect 15289 32929 15301 32963
rect 15335 32960 15347 32963
rect 15562 32960 15568 32972
rect 15335 32932 15568 32960
rect 15335 32929 15347 32932
rect 15289 32923 15347 32929
rect 15562 32920 15568 32932
rect 15620 32920 15626 32972
rect 15212 32864 15332 32892
rect 15105 32855 15163 32861
rect 14507 32796 14688 32824
rect 14737 32827 14795 32833
rect 14507 32793 14519 32796
rect 14461 32787 14519 32793
rect 14737 32793 14749 32827
rect 14783 32824 14795 32827
rect 15120 32824 15148 32855
rect 15194 32824 15200 32836
rect 14783 32796 15200 32824
rect 14783 32793 14795 32796
rect 14737 32787 14795 32793
rect 15194 32784 15200 32796
rect 15252 32784 15258 32836
rect 15304 32824 15332 32864
rect 15378 32852 15384 32904
rect 15436 32852 15442 32904
rect 15470 32852 15476 32904
rect 15528 32852 15534 32904
rect 15672 32901 15700 33000
rect 17788 33000 18512 33028
rect 15657 32895 15715 32901
rect 15657 32861 15669 32895
rect 15703 32861 15715 32895
rect 15657 32855 15715 32861
rect 16574 32824 16580 32836
rect 15304 32796 16580 32824
rect 16574 32784 16580 32796
rect 16632 32784 16638 32836
rect 14642 32756 14648 32768
rect 14384 32728 14648 32756
rect 14642 32716 14648 32728
rect 14700 32716 14706 32768
rect 15102 32716 15108 32768
rect 15160 32756 15166 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 15160 32728 15577 32756
rect 15160 32716 15166 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 15565 32719 15623 32725
rect 15654 32716 15660 32768
rect 15712 32756 15718 32768
rect 17788 32756 17816 33000
rect 18506 32988 18512 33000
rect 18564 32988 18570 33040
rect 17954 32920 17960 32972
rect 18012 32960 18018 32972
rect 18708 32969 18736 33068
rect 18782 33056 18788 33068
rect 18840 33096 18846 33108
rect 21174 33096 21180 33108
rect 18840 33068 21180 33096
rect 18840 33056 18846 33068
rect 21174 33056 21180 33068
rect 21232 33096 21238 33108
rect 21726 33096 21732 33108
rect 21232 33068 21732 33096
rect 21232 33056 21238 33068
rect 21726 33056 21732 33068
rect 21784 33056 21790 33108
rect 22462 33056 22468 33108
rect 22520 33056 22526 33108
rect 18877 33031 18935 33037
rect 18877 32997 18889 33031
rect 18923 33028 18935 33031
rect 19426 33028 19432 33040
rect 18923 33000 19432 33028
rect 18923 32997 18935 33000
rect 18877 32991 18935 32997
rect 19426 32988 19432 33000
rect 19484 32988 19490 33040
rect 18693 32963 18751 32969
rect 18693 32960 18705 32963
rect 18012 32932 18705 32960
rect 18012 32920 18018 32932
rect 18693 32929 18705 32932
rect 18739 32929 18751 32963
rect 18693 32923 18751 32929
rect 18782 32920 18788 32972
rect 18840 32960 18846 32972
rect 19150 32960 19156 32972
rect 18840 32932 19156 32960
rect 18840 32920 18846 32932
rect 19150 32920 19156 32932
rect 19208 32960 19214 32972
rect 20165 32963 20223 32969
rect 20165 32960 20177 32963
rect 19208 32932 20177 32960
rect 19208 32920 19214 32932
rect 20165 32929 20177 32932
rect 20211 32960 20223 32963
rect 20211 32932 22094 32960
rect 20211 32929 20223 32932
rect 20165 32923 20223 32929
rect 17862 32852 17868 32904
rect 17920 32852 17926 32904
rect 18046 32852 18052 32904
rect 18104 32852 18110 32904
rect 18138 32852 18144 32904
rect 18196 32852 18202 32904
rect 18233 32895 18291 32901
rect 18233 32861 18245 32895
rect 18279 32861 18291 32895
rect 18233 32855 18291 32861
rect 15712 32728 17816 32756
rect 15712 32716 15718 32728
rect 18138 32716 18144 32768
rect 18196 32756 18202 32768
rect 18248 32756 18276 32855
rect 18414 32852 18420 32904
rect 18472 32852 18478 32904
rect 18966 32852 18972 32904
rect 19024 32852 19030 32904
rect 22066 32892 22094 32932
rect 22738 32920 22744 32972
rect 22796 32960 22802 32972
rect 23017 32963 23075 32969
rect 23017 32960 23029 32963
rect 22796 32932 23029 32960
rect 22796 32920 22802 32932
rect 23017 32929 23029 32932
rect 23063 32929 23075 32963
rect 24670 32960 24676 32972
rect 23017 32923 23075 32929
rect 23768 32932 24676 32960
rect 23477 32895 23535 32901
rect 23477 32892 23489 32895
rect 22066 32864 23489 32892
rect 23477 32861 23489 32864
rect 23523 32892 23535 32895
rect 23566 32892 23572 32904
rect 23523 32864 23572 32892
rect 23523 32861 23535 32864
rect 23477 32855 23535 32861
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 18690 32784 18696 32836
rect 18748 32784 18754 32836
rect 20441 32827 20499 32833
rect 20441 32793 20453 32827
rect 20487 32824 20499 32827
rect 20530 32824 20536 32836
rect 20487 32796 20536 32824
rect 20487 32793 20499 32796
rect 20441 32787 20499 32793
rect 20530 32784 20536 32796
rect 20588 32784 20594 32836
rect 23768 32824 23796 32932
rect 24670 32920 24676 32932
rect 24728 32920 24734 32972
rect 25130 32920 25136 32972
rect 25188 32960 25194 32972
rect 25225 32963 25283 32969
rect 25225 32960 25237 32963
rect 25188 32932 25237 32960
rect 25188 32920 25194 32932
rect 25225 32929 25237 32932
rect 25271 32929 25283 32963
rect 25225 32923 25283 32929
rect 27617 32963 27675 32969
rect 27617 32929 27629 32963
rect 27663 32960 27675 32963
rect 29549 32963 29607 32969
rect 29549 32960 29561 32963
rect 27663 32932 29561 32960
rect 27663 32929 27675 32932
rect 27617 32923 27675 32929
rect 29549 32929 29561 32932
rect 29595 32960 29607 32963
rect 30190 32960 30196 32972
rect 29595 32932 30196 32960
rect 29595 32929 29607 32932
rect 29549 32923 29607 32929
rect 30190 32920 30196 32932
rect 30248 32920 30254 32972
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24397 32895 24455 32901
rect 24397 32892 24409 32895
rect 23900 32864 24409 32892
rect 23900 32852 23906 32864
rect 24397 32861 24409 32864
rect 24443 32861 24455 32895
rect 24397 32855 24455 32861
rect 28810 32852 28816 32904
rect 28868 32892 28874 32904
rect 29181 32895 29239 32901
rect 29181 32892 29193 32895
rect 28868 32864 29193 32892
rect 28868 32852 28874 32864
rect 29181 32861 29193 32864
rect 29227 32861 29239 32895
rect 29181 32855 29239 32861
rect 29914 32852 29920 32904
rect 29972 32852 29978 32904
rect 20824 32796 20930 32824
rect 21744 32796 23796 32824
rect 20824 32768 20852 32796
rect 18196 32728 18276 32756
rect 18196 32716 18202 32728
rect 18598 32716 18604 32768
rect 18656 32716 18662 32768
rect 18874 32716 18880 32768
rect 18932 32756 18938 32768
rect 20714 32756 20720 32768
rect 18932 32728 20720 32756
rect 18932 32716 18938 32728
rect 20714 32716 20720 32728
rect 20772 32716 20778 32768
rect 20806 32716 20812 32768
rect 20864 32756 20870 32768
rect 21744 32756 21772 32796
rect 24210 32784 24216 32836
rect 24268 32784 24274 32836
rect 24302 32784 24308 32836
rect 24360 32824 24366 32836
rect 25041 32827 25099 32833
rect 25041 32824 25053 32827
rect 24360 32796 25053 32824
rect 24360 32784 24366 32796
rect 25041 32793 25053 32796
rect 25087 32793 25099 32827
rect 25041 32787 25099 32793
rect 25593 32827 25651 32833
rect 25593 32793 25605 32827
rect 25639 32824 25651 32827
rect 25958 32824 25964 32836
rect 25639 32796 25964 32824
rect 25639 32793 25651 32796
rect 25593 32787 25651 32793
rect 25958 32784 25964 32796
rect 26016 32784 26022 32836
rect 26602 32784 26608 32836
rect 26660 32784 26666 32836
rect 27338 32784 27344 32836
rect 27396 32784 27402 32836
rect 30834 32784 30840 32836
rect 30892 32784 30898 32836
rect 20864 32728 21772 32756
rect 20864 32716 20870 32728
rect 21818 32716 21824 32768
rect 21876 32756 21882 32768
rect 21913 32759 21971 32765
rect 21913 32756 21925 32759
rect 21876 32728 21925 32756
rect 21876 32716 21882 32728
rect 21913 32725 21925 32728
rect 21959 32725 21971 32759
rect 21913 32719 21971 32725
rect 22554 32716 22560 32768
rect 22612 32756 22618 32768
rect 22833 32759 22891 32765
rect 22833 32756 22845 32759
rect 22612 32728 22845 32756
rect 22612 32716 22618 32728
rect 22833 32725 22845 32728
rect 22879 32725 22891 32759
rect 22833 32719 22891 32725
rect 22925 32759 22983 32765
rect 22925 32725 22937 32759
rect 22971 32756 22983 32759
rect 24489 32759 24547 32765
rect 24489 32756 24501 32759
rect 22971 32728 24501 32756
rect 22971 32725 22983 32728
rect 22925 32719 22983 32725
rect 24489 32725 24501 32728
rect 24535 32725 24547 32759
rect 24489 32719 24547 32725
rect 24673 32759 24731 32765
rect 24673 32725 24685 32759
rect 24719 32756 24731 32759
rect 24854 32756 24860 32768
rect 24719 32728 24860 32756
rect 24719 32725 24731 32728
rect 24673 32719 24731 32725
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 25133 32759 25191 32765
rect 25133 32725 25145 32759
rect 25179 32756 25191 32759
rect 25498 32756 25504 32768
rect 25179 32728 25504 32756
rect 25179 32725 25191 32728
rect 25133 32719 25191 32725
rect 25498 32716 25504 32728
rect 25556 32716 25562 32768
rect 28166 32716 28172 32768
rect 28224 32756 28230 32768
rect 28629 32759 28687 32765
rect 28629 32756 28641 32759
rect 28224 32728 28641 32756
rect 28224 32716 28230 32728
rect 28629 32725 28641 32728
rect 28675 32725 28687 32759
rect 28629 32719 28687 32725
rect 30006 32716 30012 32768
rect 30064 32756 30070 32768
rect 30650 32756 30656 32768
rect 30064 32728 30656 32756
rect 30064 32716 30070 32728
rect 30650 32716 30656 32728
rect 30708 32756 30714 32768
rect 31343 32759 31401 32765
rect 31343 32756 31355 32759
rect 30708 32728 31355 32756
rect 30708 32716 30714 32728
rect 31343 32725 31355 32728
rect 31389 32725 31401 32759
rect 31343 32719 31401 32725
rect 1104 32666 36524 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 36524 32666
rect 1104 32592 36524 32614
rect 6546 32512 6552 32564
rect 6604 32552 6610 32564
rect 8478 32552 8484 32564
rect 6604 32524 8484 32552
rect 6604 32512 6610 32524
rect 8478 32512 8484 32524
rect 8536 32512 8542 32564
rect 8846 32512 8852 32564
rect 8904 32552 8910 32564
rect 8904 32524 11008 32552
rect 8904 32512 8910 32524
rect 2682 32444 2688 32496
rect 2740 32484 2746 32496
rect 5077 32487 5135 32493
rect 5077 32484 5089 32487
rect 2740 32456 5089 32484
rect 2740 32444 2746 32456
rect 5077 32453 5089 32456
rect 5123 32453 5135 32487
rect 5077 32447 5135 32453
rect 7282 32444 7288 32496
rect 7340 32444 7346 32496
rect 7926 32444 7932 32496
rect 7984 32484 7990 32496
rect 8389 32487 8447 32493
rect 8389 32484 8401 32487
rect 7984 32456 8401 32484
rect 7984 32444 7990 32456
rect 8389 32453 8401 32456
rect 8435 32484 8447 32487
rect 10318 32484 10324 32496
rect 8435 32456 10324 32484
rect 8435 32453 8447 32456
rect 8389 32447 8447 32453
rect 10318 32444 10324 32456
rect 10376 32444 10382 32496
rect 10980 32484 11008 32524
rect 11054 32512 11060 32564
rect 11112 32512 11118 32564
rect 11790 32512 11796 32564
rect 11848 32552 11854 32564
rect 11885 32555 11943 32561
rect 11885 32552 11897 32555
rect 11848 32524 11897 32552
rect 11848 32512 11854 32524
rect 11885 32521 11897 32524
rect 11931 32521 11943 32555
rect 11885 32515 11943 32521
rect 12529 32555 12587 32561
rect 12529 32521 12541 32555
rect 12575 32552 12587 32555
rect 14734 32552 14740 32564
rect 12575 32524 14740 32552
rect 12575 32521 12587 32524
rect 12529 32515 12587 32521
rect 14734 32512 14740 32524
rect 14792 32512 14798 32564
rect 15197 32555 15255 32561
rect 15197 32552 15209 32555
rect 14936 32524 15209 32552
rect 13814 32484 13820 32496
rect 10980 32456 13820 32484
rect 13814 32444 13820 32456
rect 13872 32444 13878 32496
rect 14642 32444 14648 32496
rect 14700 32484 14706 32496
rect 14936 32493 14964 32524
rect 15197 32521 15209 32524
rect 15243 32521 15255 32555
rect 15197 32515 15255 32521
rect 17310 32512 17316 32564
rect 17368 32552 17374 32564
rect 17497 32555 17555 32561
rect 17497 32552 17509 32555
rect 17368 32524 17509 32552
rect 17368 32512 17374 32524
rect 17497 32521 17509 32524
rect 17543 32521 17555 32555
rect 17497 32515 17555 32521
rect 18414 32512 18420 32564
rect 18472 32552 18478 32564
rect 18690 32552 18696 32564
rect 18472 32524 18696 32552
rect 18472 32512 18478 32524
rect 18690 32512 18696 32524
rect 18748 32552 18754 32564
rect 19981 32555 20039 32561
rect 19981 32552 19993 32555
rect 18748 32524 19993 32552
rect 18748 32512 18754 32524
rect 19981 32521 19993 32524
rect 20027 32521 20039 32555
rect 19981 32515 20039 32521
rect 20530 32512 20536 32564
rect 20588 32512 20594 32564
rect 21634 32552 21640 32564
rect 20640 32524 21640 32552
rect 14829 32487 14887 32493
rect 14829 32484 14841 32487
rect 14700 32456 14841 32484
rect 14700 32444 14706 32456
rect 14829 32453 14841 32456
rect 14875 32453 14887 32487
rect 14829 32447 14887 32453
rect 14921 32487 14979 32493
rect 14921 32453 14933 32487
rect 14967 32453 14979 32487
rect 14921 32447 14979 32453
rect 15378 32444 15384 32496
rect 15436 32484 15442 32496
rect 15436 32456 15688 32484
rect 15436 32444 15442 32456
rect 4890 32376 4896 32428
rect 4948 32376 4954 32428
rect 5169 32419 5227 32425
rect 5169 32385 5181 32419
rect 5215 32416 5227 32419
rect 5350 32416 5356 32428
rect 5215 32388 5356 32416
rect 5215 32385 5227 32388
rect 5169 32379 5227 32385
rect 5350 32376 5356 32388
rect 5408 32376 5414 32428
rect 8202 32376 8208 32428
rect 8260 32416 8266 32428
rect 8941 32419 8999 32425
rect 8941 32416 8953 32419
rect 8260 32388 8953 32416
rect 8260 32376 8266 32388
rect 8941 32385 8953 32388
rect 8987 32385 8999 32419
rect 8941 32379 8999 32385
rect 9398 32376 9404 32428
rect 9456 32376 9462 32428
rect 9582 32376 9588 32428
rect 9640 32376 9646 32428
rect 10134 32376 10140 32428
rect 10192 32416 10198 32428
rect 10597 32419 10655 32425
rect 10597 32416 10609 32419
rect 10192 32388 10609 32416
rect 10192 32376 10198 32388
rect 10597 32385 10609 32388
rect 10643 32385 10655 32419
rect 10597 32379 10655 32385
rect 10873 32419 10931 32425
rect 10873 32385 10885 32419
rect 10919 32416 10931 32419
rect 11054 32416 11060 32428
rect 10919 32388 11060 32416
rect 10919 32385 10931 32388
rect 10873 32379 10931 32385
rect 11054 32376 11060 32388
rect 11112 32376 11118 32428
rect 11149 32419 11207 32425
rect 11149 32385 11161 32419
rect 11195 32416 11207 32419
rect 11238 32416 11244 32428
rect 11195 32388 11244 32416
rect 11195 32385 11207 32388
rect 11149 32379 11207 32385
rect 11238 32376 11244 32388
rect 11296 32376 11302 32428
rect 11514 32376 11520 32428
rect 11572 32376 11578 32428
rect 11698 32376 11704 32428
rect 11756 32416 11762 32428
rect 12161 32419 12219 32425
rect 12161 32416 12173 32419
rect 11756 32388 12173 32416
rect 11756 32376 11762 32388
rect 12161 32385 12173 32388
rect 12207 32385 12219 32419
rect 12161 32379 12219 32385
rect 12989 32419 13047 32425
rect 12989 32385 13001 32419
rect 13035 32416 13047 32419
rect 13170 32416 13176 32428
rect 13035 32388 13176 32416
rect 13035 32385 13047 32388
rect 12989 32379 13047 32385
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 14734 32376 14740 32428
rect 14792 32376 14798 32428
rect 15102 32376 15108 32428
rect 15160 32376 15166 32428
rect 15194 32376 15200 32428
rect 15252 32416 15258 32428
rect 15660 32425 15688 32456
rect 15746 32444 15752 32496
rect 15804 32484 15810 32496
rect 18782 32484 18788 32496
rect 15804 32456 15976 32484
rect 15804 32444 15810 32456
rect 15473 32419 15531 32425
rect 15473 32416 15485 32419
rect 15252 32388 15485 32416
rect 15252 32376 15258 32388
rect 15473 32385 15485 32388
rect 15519 32385 15531 32419
rect 15473 32379 15531 32385
rect 15565 32419 15623 32425
rect 15565 32385 15577 32419
rect 15611 32385 15623 32419
rect 15565 32379 15623 32385
rect 15657 32419 15715 32425
rect 15657 32385 15669 32419
rect 15703 32385 15715 32419
rect 15657 32379 15715 32385
rect 6365 32351 6423 32357
rect 6365 32317 6377 32351
rect 6411 32317 6423 32351
rect 6365 32311 6423 32317
rect 6641 32351 6699 32357
rect 6641 32317 6653 32351
rect 6687 32348 6699 32351
rect 7098 32348 7104 32360
rect 6687 32320 7104 32348
rect 6687 32317 6699 32320
rect 6641 32311 6699 32317
rect 4709 32215 4767 32221
rect 4709 32181 4721 32215
rect 4755 32212 4767 32215
rect 5534 32212 5540 32224
rect 4755 32184 5540 32212
rect 4755 32181 4767 32184
rect 4709 32175 4767 32181
rect 5534 32172 5540 32184
rect 5592 32172 5598 32224
rect 6380 32212 6408 32311
rect 7098 32308 7104 32320
rect 7156 32308 7162 32360
rect 9033 32351 9091 32357
rect 9033 32317 9045 32351
rect 9079 32348 9091 32351
rect 9493 32351 9551 32357
rect 9493 32348 9505 32351
rect 9079 32320 9505 32348
rect 9079 32317 9091 32320
rect 9033 32311 9091 32317
rect 9493 32317 9505 32320
rect 9539 32317 9551 32351
rect 9493 32311 9551 32317
rect 10318 32308 10324 32360
rect 10376 32348 10382 32360
rect 10689 32351 10747 32357
rect 10689 32348 10701 32351
rect 10376 32320 10701 32348
rect 10376 32308 10382 32320
rect 10689 32317 10701 32320
rect 10735 32317 10747 32351
rect 11716 32348 11744 32376
rect 10689 32311 10747 32317
rect 10796 32320 11744 32348
rect 9306 32240 9312 32292
rect 9364 32240 9370 32292
rect 9674 32240 9680 32292
rect 9732 32280 9738 32292
rect 10796 32280 10824 32320
rect 11974 32308 11980 32360
rect 12032 32348 12038 32360
rect 12069 32351 12127 32357
rect 12069 32348 12081 32351
rect 12032 32320 12081 32348
rect 12032 32308 12038 32320
rect 12069 32317 12081 32320
rect 12115 32317 12127 32351
rect 12805 32351 12863 32357
rect 12805 32348 12817 32351
rect 12069 32311 12127 32317
rect 12406 32320 12817 32348
rect 11241 32283 11299 32289
rect 11241 32280 11253 32283
rect 9732 32252 10824 32280
rect 10888 32252 11253 32280
rect 9732 32240 9738 32252
rect 7190 32212 7196 32224
rect 6380 32184 7196 32212
rect 7190 32172 7196 32184
rect 7248 32172 7254 32224
rect 10410 32172 10416 32224
rect 10468 32212 10474 32224
rect 10888 32221 10916 32252
rect 11241 32249 11253 32252
rect 11287 32249 11299 32283
rect 11241 32243 11299 32249
rect 11330 32240 11336 32292
rect 11388 32280 11394 32292
rect 12406 32280 12434 32320
rect 12805 32317 12817 32320
rect 12851 32317 12863 32351
rect 12805 32311 12863 32317
rect 12894 32308 12900 32360
rect 12952 32308 12958 32360
rect 13081 32351 13139 32357
rect 13081 32317 13093 32351
rect 13127 32317 13139 32351
rect 15580 32348 15608 32379
rect 15838 32376 15844 32428
rect 15896 32376 15902 32428
rect 15948 32425 15976 32456
rect 17696 32456 18184 32484
rect 15933 32419 15991 32425
rect 15933 32385 15945 32419
rect 15979 32385 15991 32419
rect 15933 32379 15991 32385
rect 15948 32348 15976 32379
rect 16114 32376 16120 32428
rect 16172 32376 16178 32428
rect 16666 32376 16672 32428
rect 16724 32376 16730 32428
rect 16850 32376 16856 32428
rect 16908 32416 16914 32428
rect 17696 32425 17724 32456
rect 17129 32419 17187 32425
rect 17129 32416 17141 32419
rect 16908 32388 17141 32416
rect 16908 32376 16914 32388
rect 17129 32385 17141 32388
rect 17175 32385 17187 32419
rect 17129 32379 17187 32385
rect 17313 32419 17371 32425
rect 17313 32385 17325 32419
rect 17359 32385 17371 32419
rect 17313 32379 17371 32385
rect 17681 32419 17739 32425
rect 17681 32385 17693 32419
rect 17727 32385 17739 32419
rect 17681 32379 17739 32385
rect 16298 32348 16304 32360
rect 15580 32320 16304 32348
rect 13081 32311 13139 32317
rect 11388 32252 12434 32280
rect 13096 32280 13124 32311
rect 16298 32308 16304 32320
rect 16356 32308 16362 32360
rect 16942 32308 16948 32360
rect 17000 32308 17006 32360
rect 17328 32348 17356 32379
rect 17770 32376 17776 32428
rect 17828 32376 17834 32428
rect 17957 32419 18015 32425
rect 17957 32385 17969 32419
rect 18003 32385 18015 32419
rect 17957 32379 18015 32385
rect 17865 32351 17923 32357
rect 17865 32348 17877 32351
rect 17328 32320 17877 32348
rect 17865 32317 17877 32320
rect 17911 32317 17923 32351
rect 17865 32311 17923 32317
rect 14553 32283 14611 32289
rect 14553 32280 14565 32283
rect 13096 32252 14565 32280
rect 11388 32240 11394 32252
rect 14553 32249 14565 32252
rect 14599 32249 14611 32283
rect 16853 32283 16911 32289
rect 14553 32243 14611 32249
rect 15304 32252 15516 32280
rect 10873 32215 10931 32221
rect 10873 32212 10885 32215
rect 10468 32184 10885 32212
rect 10468 32172 10474 32184
rect 10873 32181 10885 32184
rect 10919 32181 10931 32215
rect 10873 32175 10931 32181
rect 11146 32172 11152 32224
rect 11204 32212 11210 32224
rect 11517 32215 11575 32221
rect 11517 32212 11529 32215
rect 11204 32184 11529 32212
rect 11204 32172 11210 32184
rect 11517 32181 11529 32184
rect 11563 32181 11575 32215
rect 11517 32175 11575 32181
rect 12526 32172 12532 32224
rect 12584 32212 12590 32224
rect 12621 32215 12679 32221
rect 12621 32212 12633 32215
rect 12584 32184 12633 32212
rect 12584 32172 12590 32184
rect 12621 32181 12633 32184
rect 12667 32181 12679 32215
rect 12621 32175 12679 32181
rect 13170 32172 13176 32224
rect 13228 32212 13234 32224
rect 15304 32212 15332 32252
rect 13228 32184 15332 32212
rect 13228 32172 13234 32184
rect 15378 32172 15384 32224
rect 15436 32172 15442 32224
rect 15488 32212 15516 32252
rect 16853 32249 16865 32283
rect 16899 32280 16911 32283
rect 16899 32252 17724 32280
rect 16899 32249 16911 32252
rect 16853 32243 16911 32249
rect 15654 32212 15660 32224
rect 15488 32184 15660 32212
rect 15654 32172 15660 32184
rect 15712 32172 15718 32224
rect 15746 32172 15752 32224
rect 15804 32212 15810 32224
rect 15841 32215 15899 32221
rect 15841 32212 15853 32215
rect 15804 32184 15853 32212
rect 15804 32172 15810 32184
rect 15841 32181 15853 32184
rect 15887 32181 15899 32215
rect 15841 32175 15899 32181
rect 16114 32172 16120 32224
rect 16172 32172 16178 32224
rect 16758 32172 16764 32224
rect 16816 32172 16822 32224
rect 17313 32215 17371 32221
rect 17313 32181 17325 32215
rect 17359 32212 17371 32215
rect 17586 32212 17592 32224
rect 17359 32184 17592 32212
rect 17359 32181 17371 32184
rect 17313 32175 17371 32181
rect 17586 32172 17592 32184
rect 17644 32172 17650 32224
rect 17696 32212 17724 32252
rect 17770 32240 17776 32292
rect 17828 32280 17834 32292
rect 17972 32280 18000 32379
rect 18156 32348 18184 32456
rect 18248 32456 18788 32484
rect 18248 32425 18276 32456
rect 18782 32444 18788 32456
rect 18840 32444 18846 32496
rect 20438 32484 20444 32496
rect 19734 32456 20444 32484
rect 20438 32444 20444 32456
rect 20496 32444 20502 32496
rect 18233 32419 18291 32425
rect 18233 32385 18245 32419
rect 18279 32385 18291 32419
rect 20640 32416 20668 32524
rect 21634 32512 21640 32524
rect 21692 32512 21698 32564
rect 21726 32512 21732 32564
rect 21784 32552 21790 32564
rect 22557 32555 22615 32561
rect 21784 32524 22094 32552
rect 21784 32512 21790 32524
rect 22066 32484 22094 32524
rect 22557 32521 22569 32555
rect 22603 32552 22615 32555
rect 22646 32552 22652 32564
rect 22603 32524 22652 32552
rect 22603 32521 22615 32524
rect 22557 32515 22615 32521
rect 22646 32512 22652 32524
rect 22704 32512 22710 32564
rect 24946 32552 24952 32564
rect 23492 32524 24952 32552
rect 23492 32493 23520 32524
rect 24946 32512 24952 32524
rect 25004 32512 25010 32564
rect 25317 32555 25375 32561
rect 25317 32521 25329 32555
rect 25363 32552 25375 32555
rect 27338 32552 27344 32564
rect 25363 32524 27344 32552
rect 25363 32521 25375 32524
rect 25317 32515 25375 32521
rect 27338 32512 27344 32524
rect 27396 32512 27402 32564
rect 30926 32552 30932 32564
rect 29012 32524 30932 32552
rect 23477 32487 23535 32493
rect 22066 32456 22784 32484
rect 18233 32379 18291 32385
rect 20088 32388 20668 32416
rect 20717 32419 20775 32425
rect 20088 32348 20116 32388
rect 20717 32385 20729 32419
rect 20763 32416 20775 32419
rect 20806 32416 20812 32428
rect 20763 32388 20812 32416
rect 20763 32385 20775 32388
rect 20717 32379 20775 32385
rect 20806 32376 20812 32388
rect 20864 32376 20870 32428
rect 20898 32376 20904 32428
rect 20956 32376 20962 32428
rect 21634 32376 21640 32428
rect 21692 32416 21698 32428
rect 21692 32388 21956 32416
rect 21692 32376 21698 32388
rect 20993 32351 21051 32357
rect 20993 32348 21005 32351
rect 18156 32320 20116 32348
rect 20548 32320 21005 32348
rect 17828 32252 18000 32280
rect 17828 32240 17834 32252
rect 20070 32240 20076 32292
rect 20128 32280 20134 32292
rect 20548 32280 20576 32320
rect 20993 32317 21005 32320
rect 21039 32348 21051 32351
rect 21726 32348 21732 32360
rect 21039 32320 21732 32348
rect 21039 32317 21051 32320
rect 20993 32311 21051 32317
rect 21726 32308 21732 32320
rect 21784 32308 21790 32360
rect 21821 32351 21879 32357
rect 21821 32317 21833 32351
rect 21867 32317 21879 32351
rect 21821 32311 21879 32317
rect 21836 32280 21864 32311
rect 20128 32252 20576 32280
rect 20640 32252 21864 32280
rect 21928 32280 21956 32388
rect 22002 32376 22008 32428
rect 22060 32376 22066 32428
rect 22094 32376 22100 32428
rect 22152 32376 22158 32428
rect 22186 32376 22192 32428
rect 22244 32376 22250 32428
rect 22756 32425 22784 32456
rect 23477 32453 23489 32487
rect 23523 32453 23535 32487
rect 23477 32447 23535 32453
rect 24673 32487 24731 32493
rect 24673 32453 24685 32487
rect 24719 32484 24731 32487
rect 28902 32484 28908 32496
rect 24719 32456 25636 32484
rect 28474 32456 28908 32484
rect 24719 32453 24731 32456
rect 24673 32447 24731 32453
rect 22741 32419 22799 32425
rect 22741 32385 22753 32419
rect 22787 32385 22799 32419
rect 22741 32379 22799 32385
rect 23014 32376 23020 32428
rect 23072 32376 23078 32428
rect 24210 32376 24216 32428
rect 24268 32376 24274 32428
rect 24394 32376 24400 32428
rect 24452 32376 24458 32428
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32385 24547 32419
rect 24489 32379 24547 32385
rect 22020 32348 22048 32376
rect 22020 32320 22416 32348
rect 22388 32289 22416 32320
rect 22646 32308 22652 32360
rect 22704 32348 22710 32360
rect 24026 32348 24032 32360
rect 22704 32320 24032 32348
rect 22704 32308 22710 32320
rect 24026 32308 24032 32320
rect 24084 32348 24090 32360
rect 24504 32348 24532 32379
rect 24578 32376 24584 32428
rect 24636 32416 24642 32428
rect 24949 32419 25007 32425
rect 24949 32416 24961 32419
rect 24636 32388 24961 32416
rect 24636 32376 24642 32388
rect 24949 32385 24961 32388
rect 24995 32416 25007 32419
rect 25038 32416 25044 32428
rect 24995 32388 25044 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 25038 32376 25044 32388
rect 25096 32376 25102 32428
rect 25406 32376 25412 32428
rect 25464 32376 25470 32428
rect 25608 32425 25636 32456
rect 28902 32444 28908 32456
rect 28960 32484 28966 32496
rect 29012 32484 29040 32524
rect 30926 32512 30932 32524
rect 30984 32552 30990 32564
rect 33318 32552 33324 32564
rect 30984 32524 33324 32552
rect 30984 32512 30990 32524
rect 28960 32456 29118 32484
rect 28960 32444 28966 32456
rect 30190 32444 30196 32496
rect 30248 32484 30254 32496
rect 32784 32484 32812 32524
rect 33318 32512 33324 32524
rect 33376 32512 33382 32564
rect 30248 32456 32168 32484
rect 32784 32456 32890 32484
rect 30248 32444 30254 32456
rect 25593 32419 25651 32425
rect 25593 32385 25605 32419
rect 25639 32385 25651 32419
rect 25593 32379 25651 32385
rect 25682 32376 25688 32428
rect 25740 32376 25746 32428
rect 25958 32376 25964 32428
rect 26016 32376 26022 32428
rect 30576 32425 30604 32456
rect 30561 32419 30619 32425
rect 30561 32385 30573 32419
rect 30607 32385 30619 32419
rect 30561 32379 30619 32385
rect 30650 32376 30656 32428
rect 30708 32376 30714 32428
rect 31110 32376 31116 32428
rect 31168 32376 31174 32428
rect 31294 32376 31300 32428
rect 31352 32376 31358 32428
rect 31478 32376 31484 32428
rect 31536 32376 31542 32428
rect 32140 32425 32168 32456
rect 32125 32419 32183 32425
rect 32125 32385 32137 32419
rect 32171 32385 32183 32419
rect 32125 32379 32183 32385
rect 24084 32320 24532 32348
rect 24084 32308 24090 32320
rect 24854 32308 24860 32360
rect 24912 32308 24918 32360
rect 25774 32308 25780 32360
rect 25832 32348 25838 32360
rect 26973 32351 27031 32357
rect 26973 32348 26985 32351
rect 25832 32320 26985 32348
rect 25832 32308 25838 32320
rect 26973 32317 26985 32320
rect 27019 32317 27031 32351
rect 26973 32311 27031 32317
rect 27246 32308 27252 32360
rect 27304 32308 27310 32360
rect 29086 32308 29092 32360
rect 29144 32348 29150 32360
rect 30285 32351 30343 32357
rect 30285 32348 30297 32351
rect 29144 32320 30297 32348
rect 29144 32308 29150 32320
rect 30285 32317 30297 32320
rect 30331 32317 30343 32351
rect 30929 32351 30987 32357
rect 30929 32348 30941 32351
rect 30285 32311 30343 32317
rect 30576 32320 30941 32348
rect 30576 32292 30604 32320
rect 30929 32317 30941 32320
rect 30975 32317 30987 32351
rect 32140 32348 32168 32379
rect 32306 32348 32312 32360
rect 32140 32320 32312 32348
rect 30929 32311 30987 32317
rect 32306 32308 32312 32320
rect 32364 32308 32370 32360
rect 32490 32308 32496 32360
rect 32548 32308 32554 32360
rect 33919 32351 33977 32357
rect 33919 32317 33931 32351
rect 33965 32348 33977 32351
rect 34422 32348 34428 32360
rect 33965 32320 34428 32348
rect 33965 32317 33977 32320
rect 33919 32311 33977 32317
rect 34422 32308 34428 32320
rect 34480 32348 34486 32360
rect 34609 32351 34667 32357
rect 34609 32348 34621 32351
rect 34480 32320 34621 32348
rect 34480 32308 34486 32320
rect 34609 32317 34621 32320
rect 34655 32317 34667 32351
rect 34609 32311 34667 32317
rect 22373 32283 22431 32289
rect 21928 32252 22094 32280
rect 20128 32240 20134 32252
rect 20640 32224 20668 32252
rect 18138 32212 18144 32224
rect 17696 32184 18144 32212
rect 18138 32172 18144 32184
rect 18196 32172 18202 32224
rect 18496 32215 18554 32221
rect 18496 32181 18508 32215
rect 18542 32212 18554 32215
rect 18598 32212 18604 32224
rect 18542 32184 18604 32212
rect 18542 32181 18554 32184
rect 18496 32175 18554 32181
rect 18598 32172 18604 32184
rect 18656 32172 18662 32224
rect 19518 32172 19524 32224
rect 19576 32212 19582 32224
rect 20622 32212 20628 32224
rect 19576 32184 20628 32212
rect 19576 32172 19582 32184
rect 20622 32172 20628 32184
rect 20680 32172 20686 32224
rect 21450 32172 21456 32224
rect 21508 32212 21514 32224
rect 21913 32215 21971 32221
rect 21913 32212 21925 32215
rect 21508 32184 21925 32212
rect 21508 32172 21514 32184
rect 21913 32181 21925 32184
rect 21959 32181 21971 32215
rect 22066 32212 22094 32252
rect 22373 32249 22385 32283
rect 22419 32249 22431 32283
rect 24118 32280 24124 32292
rect 22373 32243 22431 32249
rect 22480 32252 24124 32280
rect 22480 32212 22508 32252
rect 24118 32240 24124 32252
rect 24176 32240 24182 32292
rect 24394 32240 24400 32292
rect 24452 32280 24458 32292
rect 26053 32283 26111 32289
rect 26053 32280 26065 32283
rect 24452 32252 26065 32280
rect 24452 32240 24458 32252
rect 26053 32249 26065 32252
rect 26099 32249 26111 32283
rect 28810 32280 28816 32292
rect 26053 32243 26111 32249
rect 28276 32252 28816 32280
rect 22066 32184 22508 32212
rect 22925 32215 22983 32221
rect 21913 32175 21971 32181
rect 22925 32181 22937 32215
rect 22971 32212 22983 32215
rect 23198 32212 23204 32224
rect 22971 32184 23204 32212
rect 22971 32181 22983 32184
rect 22925 32175 22983 32181
rect 23198 32172 23204 32184
rect 23256 32212 23262 32224
rect 25409 32215 25467 32221
rect 25409 32212 25421 32215
rect 23256 32184 25421 32212
rect 23256 32172 23262 32184
rect 25409 32181 25421 32184
rect 25455 32181 25467 32215
rect 25409 32175 25467 32181
rect 25498 32172 25504 32224
rect 25556 32212 25562 32224
rect 25777 32215 25835 32221
rect 25777 32212 25789 32215
rect 25556 32184 25789 32212
rect 25556 32172 25562 32184
rect 25777 32181 25789 32184
rect 25823 32181 25835 32215
rect 25777 32175 25835 32181
rect 26234 32172 26240 32224
rect 26292 32212 26298 32224
rect 28276 32212 28304 32252
rect 28810 32240 28816 32252
rect 28868 32240 28874 32292
rect 30558 32240 30564 32292
rect 30616 32240 30622 32292
rect 26292 32184 28304 32212
rect 26292 32172 26298 32184
rect 28718 32172 28724 32224
rect 28776 32172 28782 32224
rect 28994 32172 29000 32224
rect 29052 32212 29058 32224
rect 31294 32212 31300 32224
rect 29052 32184 31300 32212
rect 29052 32172 29058 32184
rect 31294 32172 31300 32184
rect 31352 32172 31358 32224
rect 34054 32172 34060 32224
rect 34112 32172 34118 32224
rect 1104 32122 36524 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 36524 32122
rect 1104 32048 36524 32070
rect 4890 31968 4896 32020
rect 4948 32008 4954 32020
rect 4948 31980 7052 32008
rect 4948 31968 4954 31980
rect 6365 31943 6423 31949
rect 6365 31909 6377 31943
rect 6411 31940 6423 31943
rect 6914 31940 6920 31952
rect 6411 31912 6920 31940
rect 6411 31909 6423 31912
rect 6365 31903 6423 31909
rect 6914 31900 6920 31912
rect 6972 31900 6978 31952
rect 7024 31940 7052 31980
rect 7098 31968 7104 32020
rect 7156 31968 7162 32020
rect 7208 31980 8984 32008
rect 7208 31940 7236 31980
rect 7926 31940 7932 31952
rect 7024 31912 7236 31940
rect 7576 31912 7932 31940
rect 5534 31832 5540 31884
rect 5592 31832 5598 31884
rect 5813 31875 5871 31881
rect 5813 31841 5825 31875
rect 5859 31872 5871 31875
rect 7190 31872 7196 31884
rect 5859 31844 7196 31872
rect 5859 31841 5871 31844
rect 5813 31835 5871 31841
rect 7190 31832 7196 31844
rect 7248 31832 7254 31884
rect 7576 31881 7604 31912
rect 7926 31900 7932 31912
rect 7984 31900 7990 31952
rect 8956 31949 8984 31980
rect 9490 31968 9496 32020
rect 9548 31968 9554 32020
rect 9582 31968 9588 32020
rect 9640 31968 9646 32020
rect 10042 31968 10048 32020
rect 10100 32008 10106 32020
rect 10413 32011 10471 32017
rect 10413 32008 10425 32011
rect 10100 31980 10425 32008
rect 10100 31968 10106 31980
rect 10413 31977 10425 31980
rect 10459 32008 10471 32011
rect 10778 32008 10784 32020
rect 10459 31980 10784 32008
rect 10459 31977 10471 31980
rect 10413 31971 10471 31977
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 11149 32011 11207 32017
rect 11149 31977 11161 32011
rect 11195 32008 11207 32011
rect 11330 32008 11336 32020
rect 11195 31980 11336 32008
rect 11195 31977 11207 31980
rect 11149 31971 11207 31977
rect 11330 31968 11336 31980
rect 11388 31968 11394 32020
rect 11974 31968 11980 32020
rect 12032 31968 12038 32020
rect 12332 32011 12390 32017
rect 12332 31977 12344 32011
rect 12378 32008 12390 32011
rect 12526 32008 12532 32020
rect 12378 31980 12532 32008
rect 12378 31977 12390 31980
rect 12332 31971 12390 31977
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 13817 32011 13875 32017
rect 13817 31977 13829 32011
rect 13863 32008 13875 32011
rect 14642 32008 14648 32020
rect 13863 31980 14648 32008
rect 13863 31977 13875 31980
rect 13817 31971 13875 31977
rect 14642 31968 14648 31980
rect 14700 31968 14706 32020
rect 15378 31968 15384 32020
rect 15436 31968 15442 32020
rect 15948 31980 16712 32008
rect 8941 31943 8999 31949
rect 8941 31909 8953 31943
rect 8987 31940 8999 31943
rect 9674 31940 9680 31952
rect 8987 31912 9680 31940
rect 8987 31909 8999 31912
rect 8941 31903 8999 31909
rect 9674 31900 9680 31912
rect 9732 31900 9738 31952
rect 15948 31949 15976 31980
rect 10597 31943 10655 31949
rect 10597 31909 10609 31943
rect 10643 31940 10655 31943
rect 15933 31943 15991 31949
rect 10643 31912 11560 31940
rect 10643 31909 10655 31912
rect 10597 31903 10655 31909
rect 7561 31875 7619 31881
rect 7561 31841 7573 31875
rect 7607 31841 7619 31875
rect 7561 31835 7619 31841
rect 7745 31875 7803 31881
rect 7745 31841 7757 31875
rect 7791 31872 7803 31875
rect 8294 31872 8300 31884
rect 7791 31844 8300 31872
rect 7791 31841 7803 31844
rect 7745 31835 7803 31841
rect 2682 31764 2688 31816
rect 2740 31804 2746 31816
rect 3789 31807 3847 31813
rect 3789 31804 3801 31807
rect 2740 31776 3801 31804
rect 2740 31764 2746 31776
rect 3789 31773 3801 31776
rect 3835 31773 3847 31807
rect 3789 31767 3847 31773
rect 5828 31776 6500 31804
rect 4062 31696 4068 31748
rect 4120 31736 4126 31748
rect 4120 31708 4370 31736
rect 4120 31696 4126 31708
rect 5258 31696 5264 31748
rect 5316 31736 5322 31748
rect 5828 31736 5856 31776
rect 5316 31708 5856 31736
rect 6472 31736 6500 31776
rect 6546 31764 6552 31816
rect 6604 31764 6610 31816
rect 6733 31807 6791 31813
rect 6733 31804 6745 31807
rect 6656 31776 6745 31804
rect 6656 31736 6684 31776
rect 6733 31773 6745 31776
rect 6779 31773 6791 31807
rect 6733 31767 6791 31773
rect 6825 31807 6883 31813
rect 6825 31773 6837 31807
rect 6871 31804 6883 31807
rect 7760 31804 7788 31835
rect 8294 31832 8300 31844
rect 8352 31832 8358 31884
rect 8389 31875 8447 31881
rect 8389 31841 8401 31875
rect 8435 31872 8447 31875
rect 8478 31872 8484 31884
rect 8435 31844 8484 31872
rect 8435 31841 8447 31844
rect 8389 31835 8447 31841
rect 8478 31832 8484 31844
rect 8536 31832 8542 31884
rect 6871 31776 7788 31804
rect 8113 31807 8171 31813
rect 6871 31773 6883 31776
rect 6825 31767 6883 31773
rect 8113 31773 8125 31807
rect 8159 31804 8171 31807
rect 8202 31804 8208 31816
rect 8159 31776 8208 31804
rect 8159 31773 8171 31776
rect 8113 31767 8171 31773
rect 6472 31708 6684 31736
rect 5316 31696 5322 31708
rect 5350 31628 5356 31680
rect 5408 31668 5414 31680
rect 6840 31668 6868 31767
rect 8202 31764 8208 31776
rect 8260 31804 8266 31816
rect 8573 31807 8631 31813
rect 8573 31804 8585 31807
rect 8260 31776 8585 31804
rect 8260 31764 8266 31776
rect 8573 31773 8585 31776
rect 8619 31773 8631 31807
rect 8573 31767 8631 31773
rect 8665 31807 8723 31813
rect 8665 31773 8677 31807
rect 8711 31804 8723 31807
rect 9953 31807 10011 31813
rect 9953 31804 9965 31807
rect 8711 31776 9965 31804
rect 8711 31773 8723 31776
rect 8665 31767 8723 31773
rect 9953 31773 9965 31776
rect 9999 31804 10011 31807
rect 10318 31804 10324 31816
rect 9999 31776 10324 31804
rect 9999 31773 10011 31776
rect 9953 31767 10011 31773
rect 10318 31764 10324 31776
rect 10376 31764 10382 31816
rect 10410 31764 10416 31816
rect 10468 31764 10474 31816
rect 10612 31804 10640 31903
rect 11532 31884 11560 31912
rect 15933 31909 15945 31943
rect 15979 31909 15991 31943
rect 15933 31903 15991 31909
rect 16298 31900 16304 31952
rect 16356 31900 16362 31952
rect 16684 31940 16712 31980
rect 16758 31968 16764 32020
rect 16816 32008 16822 32020
rect 17957 32011 18015 32017
rect 17957 32008 17969 32011
rect 16816 31980 17969 32008
rect 16816 31968 16822 31980
rect 17957 31977 17969 31980
rect 18003 31977 18015 32011
rect 17957 31971 18015 31977
rect 18049 32011 18107 32017
rect 18049 31977 18061 32011
rect 18095 32008 18107 32011
rect 18785 32011 18843 32017
rect 18785 32008 18797 32011
rect 18095 31980 18797 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18785 31977 18797 31980
rect 18831 32008 18843 32011
rect 18966 32008 18972 32020
rect 18831 31980 18972 32008
rect 18831 31977 18843 31980
rect 18785 31971 18843 31977
rect 18966 31968 18972 31980
rect 19024 31968 19030 32020
rect 19058 31968 19064 32020
rect 19116 32008 19122 32020
rect 19116 31980 20484 32008
rect 19116 31968 19122 31980
rect 16850 31940 16856 31952
rect 16684 31912 16856 31940
rect 10796 31844 11100 31872
rect 10796 31813 10824 31844
rect 10689 31807 10747 31813
rect 10689 31804 10701 31807
rect 10612 31776 10701 31804
rect 10689 31773 10701 31776
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 10781 31807 10839 31813
rect 10781 31773 10793 31807
rect 10827 31773 10839 31807
rect 10781 31767 10839 31773
rect 10965 31807 11023 31813
rect 10965 31773 10977 31807
rect 11011 31773 11023 31807
rect 11072 31804 11100 31844
rect 11146 31832 11152 31884
rect 11204 31872 11210 31884
rect 11333 31875 11391 31881
rect 11333 31872 11345 31875
rect 11204 31844 11345 31872
rect 11204 31832 11210 31844
rect 11333 31841 11345 31844
rect 11379 31841 11391 31875
rect 11333 31835 11391 31841
rect 11514 31832 11520 31884
rect 11572 31832 11578 31884
rect 14550 31832 14556 31884
rect 14608 31872 14614 31884
rect 14608 31844 15240 31872
rect 14608 31832 14614 31844
rect 11606 31804 11612 31816
rect 11072 31776 11612 31804
rect 10965 31767 11023 31773
rect 9309 31739 9367 31745
rect 9309 31736 9321 31739
rect 8680 31708 9321 31736
rect 5408 31640 6868 31668
rect 7469 31671 7527 31677
rect 5408 31628 5414 31640
rect 7469 31637 7481 31671
rect 7515 31668 7527 31671
rect 8018 31668 8024 31680
rect 7515 31640 8024 31668
rect 7515 31637 7527 31640
rect 7469 31631 7527 31637
rect 8018 31628 8024 31640
rect 8076 31628 8082 31680
rect 8680 31677 8708 31708
rect 9309 31705 9321 31708
rect 9355 31705 9367 31739
rect 9309 31699 9367 31705
rect 9769 31739 9827 31745
rect 9769 31705 9781 31739
rect 9815 31736 9827 31739
rect 10042 31736 10048 31748
rect 9815 31708 10048 31736
rect 9815 31705 9827 31708
rect 9769 31699 9827 31705
rect 10042 31696 10048 31708
rect 10100 31696 10106 31748
rect 10134 31696 10140 31748
rect 10192 31696 10198 31748
rect 10980 31736 11008 31767
rect 11606 31764 11612 31776
rect 11664 31764 11670 31816
rect 12066 31764 12072 31816
rect 12124 31764 12130 31816
rect 13814 31804 13820 31816
rect 13478 31776 13820 31804
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 13998 31764 14004 31816
rect 14056 31804 14062 31816
rect 15010 31804 15016 31816
rect 14056 31776 15016 31804
rect 14056 31764 14062 31776
rect 15010 31764 15016 31776
rect 15068 31764 15074 31816
rect 15212 31813 15240 31844
rect 15856 31844 16574 31872
rect 15197 31807 15255 31813
rect 15197 31773 15209 31807
rect 15243 31804 15255 31807
rect 15286 31804 15292 31816
rect 15243 31776 15292 31804
rect 15243 31773 15255 31776
rect 15197 31767 15255 31773
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 15746 31764 15752 31816
rect 15804 31804 15810 31816
rect 15856 31813 15884 31844
rect 15841 31807 15899 31813
rect 15841 31804 15853 31807
rect 15804 31776 15853 31804
rect 15804 31764 15810 31776
rect 15841 31773 15853 31776
rect 15887 31773 15899 31807
rect 15841 31767 15899 31773
rect 16025 31807 16083 31813
rect 16025 31773 16037 31807
rect 16071 31773 16083 31807
rect 16025 31767 16083 31773
rect 11054 31736 11060 31748
rect 10980 31708 11060 31736
rect 11054 31696 11060 31708
rect 11112 31696 11118 31748
rect 13832 31736 13860 31764
rect 15102 31736 15108 31748
rect 13832 31708 15108 31736
rect 15102 31696 15108 31708
rect 15160 31696 15166 31748
rect 16040 31736 16068 31767
rect 16114 31764 16120 31816
rect 16172 31764 16178 31816
rect 16546 31813 16574 31844
rect 16666 31832 16672 31884
rect 16724 31832 16730 31884
rect 16776 31881 16804 31912
rect 16850 31900 16856 31912
rect 16908 31900 16914 31952
rect 17589 31943 17647 31949
rect 17589 31909 17601 31943
rect 17635 31940 17647 31943
rect 17678 31940 17684 31952
rect 17635 31912 17684 31940
rect 17635 31909 17647 31912
rect 17589 31903 17647 31909
rect 16761 31875 16819 31881
rect 16761 31841 16773 31875
rect 16807 31841 16819 31875
rect 17604 31872 17632 31903
rect 17678 31900 17684 31912
rect 17736 31900 17742 31952
rect 17862 31900 17868 31952
rect 17920 31940 17926 31952
rect 18417 31943 18475 31949
rect 18417 31940 18429 31943
rect 17920 31912 18429 31940
rect 17920 31900 17926 31912
rect 18417 31909 18429 31912
rect 18463 31909 18475 31943
rect 18417 31903 18475 31909
rect 16761 31835 16819 31841
rect 17052 31844 17632 31872
rect 17788 31844 18368 31872
rect 16531 31807 16589 31813
rect 16531 31773 16543 31807
rect 16577 31773 16589 31807
rect 16531 31767 16589 31773
rect 16684 31736 16712 31832
rect 16850 31764 16856 31816
rect 16908 31804 16914 31816
rect 17052 31813 17080 31844
rect 17037 31807 17095 31813
rect 17037 31804 17049 31807
rect 16908 31776 17049 31804
rect 16908 31764 16914 31776
rect 17037 31773 17049 31776
rect 17083 31773 17095 31807
rect 17037 31767 17095 31773
rect 17126 31764 17132 31816
rect 17184 31764 17190 31816
rect 17310 31764 17316 31816
rect 17368 31804 17374 31816
rect 17405 31807 17463 31813
rect 17405 31804 17417 31807
rect 17368 31776 17417 31804
rect 17368 31764 17374 31776
rect 17405 31773 17417 31776
rect 17451 31773 17463 31807
rect 17405 31767 17463 31773
rect 17586 31764 17592 31816
rect 17644 31804 17650 31816
rect 17788 31804 17816 31844
rect 17644 31776 17816 31804
rect 17865 31807 17923 31813
rect 17644 31764 17650 31776
rect 17865 31773 17877 31807
rect 17911 31804 17923 31807
rect 17954 31804 17960 31816
rect 17911 31776 17960 31804
rect 17911 31773 17923 31776
rect 17865 31767 17923 31773
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18340 31813 18368 31844
rect 18874 31832 18880 31884
rect 18932 31832 18938 31884
rect 18187 31807 18245 31813
rect 18187 31804 18199 31807
rect 18165 31776 18199 31804
rect 18187 31773 18199 31776
rect 18233 31773 18245 31807
rect 18187 31767 18245 31773
rect 18325 31807 18383 31813
rect 18325 31773 18337 31807
rect 18371 31804 18383 31807
rect 18601 31807 18659 31813
rect 18601 31804 18613 31807
rect 18371 31776 18613 31804
rect 18371 31773 18383 31776
rect 18325 31767 18383 31773
rect 18601 31773 18613 31776
rect 18647 31773 18659 31807
rect 18984 31804 19012 31968
rect 19242 31900 19248 31952
rect 19300 31900 19306 31952
rect 19260 31872 19288 31900
rect 19996 31872 20208 31880
rect 20349 31875 20407 31881
rect 20349 31872 20361 31875
rect 19260 31852 20361 31872
rect 19260 31844 20024 31852
rect 20180 31844 20361 31852
rect 19444 31813 19472 31844
rect 20349 31841 20361 31844
rect 20395 31841 20407 31875
rect 20349 31835 20407 31841
rect 19245 31807 19303 31813
rect 19245 31804 19257 31807
rect 18984 31776 19257 31804
rect 18601 31767 18659 31773
rect 19245 31773 19257 31776
rect 19291 31773 19303 31807
rect 19245 31767 19303 31773
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31773 19487 31807
rect 19429 31767 19487 31773
rect 15580 31708 15976 31736
rect 16040 31708 16712 31736
rect 17144 31736 17172 31764
rect 17770 31736 17776 31748
rect 17144 31708 17776 31736
rect 8665 31671 8723 31677
rect 8665 31637 8677 31671
rect 8711 31637 8723 31671
rect 8665 31631 8723 31637
rect 8754 31628 8760 31680
rect 8812 31668 8818 31680
rect 9122 31668 9128 31680
rect 8812 31640 9128 31668
rect 8812 31628 8818 31640
rect 9122 31628 9128 31640
rect 9180 31628 9186 31680
rect 9214 31628 9220 31680
rect 9272 31628 9278 31680
rect 9398 31628 9404 31680
rect 9456 31668 9462 31680
rect 11882 31668 11888 31680
rect 9456 31640 11888 31668
rect 9456 31628 9462 31640
rect 11882 31628 11888 31640
rect 11940 31628 11946 31680
rect 14734 31628 14740 31680
rect 14792 31668 14798 31680
rect 15580 31668 15608 31708
rect 14792 31640 15608 31668
rect 14792 31628 14798 31640
rect 15654 31628 15660 31680
rect 15712 31628 15718 31680
rect 15948 31668 15976 31708
rect 17770 31696 17776 31708
rect 17828 31696 17834 31748
rect 18202 31736 18230 31767
rect 19518 31764 19524 31816
rect 19576 31804 19582 31816
rect 19613 31807 19671 31813
rect 19613 31804 19625 31807
rect 19576 31776 19625 31804
rect 19576 31764 19582 31776
rect 19613 31773 19625 31776
rect 19659 31773 19671 31807
rect 19613 31767 19671 31773
rect 19705 31807 19763 31813
rect 19705 31773 19717 31807
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 18874 31736 18880 31748
rect 18202 31708 18880 31736
rect 18874 31696 18880 31708
rect 18932 31696 18938 31748
rect 17494 31668 17500 31680
rect 15948 31640 17500 31668
rect 17494 31628 17500 31640
rect 17552 31628 17558 31680
rect 19334 31628 19340 31680
rect 19392 31668 19398 31680
rect 19720 31668 19748 31767
rect 19978 31764 19984 31816
rect 20036 31764 20042 31816
rect 20070 31764 20076 31816
rect 20128 31764 20134 31816
rect 20456 31813 20484 31980
rect 20806 31968 20812 32020
rect 20864 31968 20870 32020
rect 22646 31968 22652 32020
rect 22704 32008 22710 32020
rect 22741 32011 22799 32017
rect 22741 32008 22753 32011
rect 22704 31980 22753 32008
rect 22704 31968 22710 31980
rect 22741 31977 22753 31980
rect 22787 31977 22799 32011
rect 22741 31971 22799 31977
rect 22830 31968 22836 32020
rect 22888 32008 22894 32020
rect 23842 32008 23848 32020
rect 22888 31980 23848 32008
rect 22888 31968 22894 31980
rect 23842 31968 23848 31980
rect 23900 31968 23906 32020
rect 23934 31968 23940 32020
rect 23992 32008 23998 32020
rect 24397 32011 24455 32017
rect 24397 32008 24409 32011
rect 23992 31980 24409 32008
rect 23992 31968 23998 31980
rect 24397 31977 24409 31980
rect 24443 31977 24455 32011
rect 24397 31971 24455 31977
rect 24762 31968 24768 32020
rect 24820 32008 24826 32020
rect 25133 32011 25191 32017
rect 25133 32008 25145 32011
rect 24820 31980 25145 32008
rect 24820 31968 24826 31980
rect 25133 31977 25145 31980
rect 25179 31977 25191 32011
rect 25133 31971 25191 31977
rect 27246 31968 27252 32020
rect 27304 32008 27310 32020
rect 27433 32011 27491 32017
rect 27433 32008 27445 32011
rect 27304 31980 27445 32008
rect 27304 31968 27310 31980
rect 27433 31977 27445 31980
rect 27479 31977 27491 32011
rect 27433 31971 27491 31977
rect 27522 31968 27528 32020
rect 27580 32008 27586 32020
rect 28445 32011 28503 32017
rect 28445 32008 28457 32011
rect 27580 31980 28457 32008
rect 27580 31968 27586 31980
rect 28445 31977 28457 31980
rect 28491 31977 28503 32011
rect 28445 31971 28503 31977
rect 28994 31968 29000 32020
rect 29052 31968 29058 32020
rect 30561 32011 30619 32017
rect 30561 32008 30573 32011
rect 29196 31980 30573 32008
rect 20622 31900 20628 31952
rect 20680 31940 20686 31952
rect 22097 31943 22155 31949
rect 22097 31940 22109 31943
rect 20680 31912 22109 31940
rect 20680 31900 20686 31912
rect 22097 31909 22109 31912
rect 22143 31909 22155 31943
rect 22097 31903 22155 31909
rect 22186 31900 22192 31952
rect 22244 31900 22250 31952
rect 22370 31900 22376 31952
rect 22428 31940 22434 31952
rect 23109 31943 23167 31949
rect 23109 31940 23121 31943
rect 22428 31912 23121 31940
rect 22428 31900 22434 31912
rect 23109 31909 23121 31912
rect 23155 31909 23167 31943
rect 24029 31943 24087 31949
rect 24029 31940 24041 31943
rect 23109 31903 23167 31909
rect 23216 31912 24041 31940
rect 22204 31872 22232 31900
rect 22830 31872 22836 31884
rect 21192 31844 22232 31872
rect 22296 31844 22836 31872
rect 20257 31807 20315 31813
rect 20257 31804 20269 31807
rect 20235 31776 20269 31804
rect 20257 31773 20269 31776
rect 20303 31773 20315 31807
rect 20257 31767 20315 31773
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31773 20499 31807
rect 20441 31767 20499 31773
rect 19886 31696 19892 31748
rect 19944 31736 19950 31748
rect 20272 31736 20300 31767
rect 20990 31764 20996 31816
rect 21048 31764 21054 31816
rect 21192 31813 21220 31844
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31773 21235 31807
rect 21177 31767 21235 31773
rect 21358 31764 21364 31816
rect 21416 31764 21422 31816
rect 21450 31764 21456 31816
rect 21508 31764 21514 31816
rect 21634 31764 21640 31816
rect 21692 31764 21698 31816
rect 22296 31813 22324 31844
rect 22830 31832 22836 31844
rect 22888 31872 22894 31884
rect 23216 31872 23244 31912
rect 24029 31909 24041 31912
rect 24075 31909 24087 31943
rect 24029 31903 24087 31909
rect 24121 31943 24179 31949
rect 24121 31909 24133 31943
rect 24167 31940 24179 31943
rect 24949 31943 25007 31949
rect 24949 31940 24961 31943
rect 24167 31912 24961 31940
rect 24167 31909 24179 31912
rect 24121 31903 24179 31909
rect 24949 31909 24961 31912
rect 24995 31940 25007 31943
rect 25406 31940 25412 31952
rect 24995 31912 25412 31940
rect 24995 31909 25007 31912
rect 24949 31903 25007 31909
rect 25406 31900 25412 31912
rect 25464 31900 25470 31952
rect 28258 31940 28264 31952
rect 28092 31912 28264 31940
rect 22888 31844 23244 31872
rect 22888 31832 22894 31844
rect 23934 31832 23940 31884
rect 23992 31832 23998 31884
rect 25774 31872 25780 31884
rect 24044 31844 25780 31872
rect 22281 31807 22339 31813
rect 22281 31773 22293 31807
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 22462 31764 22468 31816
rect 22520 31764 22526 31816
rect 22738 31764 22744 31816
rect 22796 31764 22802 31816
rect 23017 31807 23075 31813
rect 23017 31773 23029 31807
rect 23063 31804 23075 31807
rect 23106 31804 23112 31816
rect 23063 31776 23112 31804
rect 23063 31773 23075 31776
rect 23017 31767 23075 31773
rect 23106 31764 23112 31776
rect 23164 31764 23170 31816
rect 23198 31764 23204 31816
rect 23256 31764 23262 31816
rect 23566 31764 23572 31816
rect 23624 31804 23630 31816
rect 24044 31804 24072 31844
rect 25774 31832 25780 31844
rect 25832 31832 25838 31884
rect 28092 31881 28120 31912
rect 28258 31900 28264 31912
rect 28316 31900 28322 31952
rect 28077 31875 28135 31881
rect 28077 31841 28089 31875
rect 28123 31841 28135 31875
rect 28442 31872 28448 31884
rect 28077 31835 28135 31841
rect 28276 31844 28448 31872
rect 23624 31776 24072 31804
rect 24213 31807 24271 31813
rect 23624 31764 23630 31776
rect 24213 31773 24225 31807
rect 24259 31804 24271 31807
rect 24302 31804 24308 31816
rect 24259 31776 24308 31804
rect 24259 31773 24271 31776
rect 24213 31767 24271 31773
rect 24302 31764 24308 31776
rect 24360 31764 24366 31816
rect 24581 31807 24639 31813
rect 24581 31773 24593 31807
rect 24627 31804 24639 31807
rect 24627 31776 24808 31804
rect 24627 31773 24639 31776
rect 24581 31767 24639 31773
rect 19944 31708 20300 31736
rect 19944 31696 19950 31708
rect 21082 31696 21088 31748
rect 21140 31696 21146 31748
rect 21542 31696 21548 31748
rect 21600 31736 21606 31748
rect 21600 31708 22094 31736
rect 21600 31696 21606 31708
rect 19797 31671 19855 31677
rect 19797 31668 19809 31671
rect 19392 31640 19809 31668
rect 19392 31628 19398 31640
rect 19797 31637 19809 31640
rect 19843 31637 19855 31671
rect 19797 31631 19855 31637
rect 19978 31628 19984 31680
rect 20036 31668 20042 31680
rect 21821 31671 21879 31677
rect 21821 31668 21833 31671
rect 20036 31640 21833 31668
rect 20036 31628 20042 31640
rect 21821 31637 21833 31640
rect 21867 31637 21879 31671
rect 22066 31668 22094 31708
rect 22740 31677 22768 31764
rect 22922 31696 22928 31748
rect 22980 31696 22986 31748
rect 24780 31736 24808 31776
rect 24854 31764 24860 31816
rect 24912 31764 24918 31816
rect 27614 31764 27620 31816
rect 27672 31764 27678 31816
rect 25317 31739 25375 31745
rect 25317 31736 25329 31739
rect 24780 31708 25329 31736
rect 25317 31705 25329 31708
rect 25363 31736 25375 31739
rect 25498 31736 25504 31748
rect 25363 31708 25504 31736
rect 25363 31705 25375 31708
rect 25317 31699 25375 31705
rect 25498 31696 25504 31708
rect 25556 31696 25562 31748
rect 27709 31739 27767 31745
rect 27709 31705 27721 31739
rect 27755 31705 27767 31739
rect 27709 31699 27767 31705
rect 22557 31671 22615 31677
rect 22557 31668 22569 31671
rect 22066 31640 22569 31668
rect 21821 31631 21879 31637
rect 22557 31637 22569 31640
rect 22603 31637 22615 31671
rect 22557 31631 22615 31637
rect 22725 31671 22783 31677
rect 22725 31637 22737 31671
rect 22771 31637 22783 31671
rect 22725 31631 22783 31637
rect 24394 31628 24400 31680
rect 24452 31668 24458 31680
rect 24762 31668 24768 31680
rect 24452 31640 24768 31668
rect 24452 31628 24458 31640
rect 24762 31628 24768 31640
rect 24820 31628 24826 31680
rect 24854 31628 24860 31680
rect 24912 31668 24918 31680
rect 25107 31671 25165 31677
rect 25107 31668 25119 31671
rect 24912 31640 25119 31668
rect 24912 31628 24918 31640
rect 25107 31637 25119 31640
rect 25153 31637 25165 31671
rect 27724 31668 27752 31699
rect 27798 31696 27804 31748
rect 27856 31696 27862 31748
rect 27939 31739 27997 31745
rect 27939 31705 27951 31739
rect 27985 31736 27997 31739
rect 28276 31736 28304 31844
rect 28442 31832 28448 31844
rect 28500 31832 28506 31884
rect 29089 31875 29147 31881
rect 29089 31841 29101 31875
rect 29135 31841 29147 31875
rect 29089 31835 29147 31841
rect 28721 31807 28779 31813
rect 27985 31708 28304 31736
rect 28399 31773 28457 31779
rect 28399 31739 28411 31773
rect 28445 31770 28457 31773
rect 28534 31770 28540 31782
rect 28445 31742 28540 31770
rect 28445 31739 28457 31742
rect 28399 31733 28457 31739
rect 28534 31730 28540 31742
rect 28592 31730 28598 31782
rect 28721 31773 28733 31807
rect 28767 31804 28779 31807
rect 28767 31776 29040 31804
rect 28767 31773 28779 31776
rect 28721 31767 28779 31773
rect 28629 31739 28687 31745
rect 27985 31705 27997 31708
rect 27939 31699 27997 31705
rect 28629 31705 28641 31739
rect 28675 31705 28687 31739
rect 28629 31699 28687 31705
rect 28074 31668 28080 31680
rect 27724 31640 28080 31668
rect 25107 31631 25165 31637
rect 28074 31628 28080 31640
rect 28132 31668 28138 31680
rect 28261 31671 28319 31677
rect 28261 31668 28273 31671
rect 28132 31640 28273 31668
rect 28132 31628 28138 31640
rect 28261 31637 28273 31640
rect 28307 31637 28319 31671
rect 28261 31631 28319 31637
rect 28442 31628 28448 31680
rect 28500 31668 28506 31680
rect 28644 31668 28672 31699
rect 28500 31640 28672 31668
rect 29012 31668 29040 31776
rect 29104 31736 29132 31835
rect 29196 31813 29224 31980
rect 30561 31977 30573 31980
rect 30607 32008 30619 32011
rect 30742 32008 30748 32020
rect 30607 31980 30748 32008
rect 30607 31977 30619 31980
rect 30561 31971 30619 31977
rect 30742 31968 30748 31980
rect 30800 32008 30806 32020
rect 31478 32008 31484 32020
rect 30800 31980 31484 32008
rect 30800 31968 30806 31980
rect 31478 31968 31484 31980
rect 31536 31968 31542 32020
rect 29365 31943 29423 31949
rect 29365 31909 29377 31943
rect 29411 31940 29423 31943
rect 30650 31940 30656 31952
rect 29411 31912 30656 31940
rect 29411 31909 29423 31912
rect 29365 31903 29423 31909
rect 30650 31900 30656 31912
rect 30708 31900 30714 31952
rect 29730 31832 29736 31884
rect 29788 31872 29794 31884
rect 30190 31872 30196 31884
rect 29788 31844 30196 31872
rect 29788 31832 29794 31844
rect 30190 31832 30196 31844
rect 30248 31872 30254 31884
rect 30285 31875 30343 31881
rect 30285 31872 30297 31875
rect 30248 31844 30297 31872
rect 30248 31832 30254 31844
rect 30285 31841 30297 31844
rect 30331 31841 30343 31875
rect 30285 31835 30343 31841
rect 31386 31832 31392 31884
rect 31444 31872 31450 31884
rect 32033 31875 32091 31881
rect 32033 31872 32045 31875
rect 31444 31844 32045 31872
rect 31444 31832 31450 31844
rect 32033 31841 32045 31844
rect 32079 31841 32091 31875
rect 32033 31835 32091 31841
rect 32306 31832 32312 31884
rect 32364 31872 32370 31884
rect 32769 31875 32827 31881
rect 32769 31872 32781 31875
rect 32364 31844 32781 31872
rect 32364 31832 32370 31844
rect 32769 31841 32781 31844
rect 32815 31841 32827 31875
rect 32769 31835 32827 31841
rect 33045 31875 33103 31881
rect 33045 31841 33057 31875
rect 33091 31872 33103 31875
rect 33410 31872 33416 31884
rect 33091 31844 33416 31872
rect 33091 31841 33103 31844
rect 33045 31835 33103 31841
rect 33410 31832 33416 31844
rect 33468 31832 33474 31884
rect 34514 31832 34520 31884
rect 34572 31872 34578 31884
rect 35253 31875 35311 31881
rect 35253 31872 35265 31875
rect 34572 31844 35265 31872
rect 34572 31832 34578 31844
rect 35253 31841 35265 31844
rect 35299 31841 35311 31875
rect 35253 31835 35311 31841
rect 29181 31807 29239 31813
rect 29181 31773 29193 31807
rect 29227 31773 29239 31807
rect 29181 31767 29239 31773
rect 29546 31764 29552 31816
rect 29604 31764 29610 31816
rect 29656 31776 30788 31804
rect 29656 31736 29684 31776
rect 29104 31708 29684 31736
rect 30006 31668 30012 31680
rect 29012 31640 30012 31668
rect 28500 31628 28506 31640
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 30098 31628 30104 31680
rect 30156 31668 30162 31680
rect 30558 31668 30564 31680
rect 30156 31640 30564 31668
rect 30156 31628 30162 31640
rect 30558 31628 30564 31640
rect 30616 31628 30622 31680
rect 30760 31668 30788 31776
rect 30926 31764 30932 31816
rect 30984 31764 30990 31816
rect 32582 31764 32588 31816
rect 32640 31804 32646 31816
rect 32677 31807 32735 31813
rect 32677 31804 32689 31807
rect 32640 31776 32689 31804
rect 32640 31764 32646 31776
rect 32677 31773 32689 31776
rect 32723 31773 32735 31807
rect 32677 31767 32735 31773
rect 34330 31736 34336 31748
rect 34270 31708 34336 31736
rect 34330 31696 34336 31708
rect 34388 31696 34394 31748
rect 31110 31668 31116 31680
rect 30760 31640 31116 31668
rect 31110 31628 31116 31640
rect 31168 31628 31174 31680
rect 32398 31628 32404 31680
rect 32456 31668 32462 31680
rect 32493 31671 32551 31677
rect 32493 31668 32505 31671
rect 32456 31640 32505 31668
rect 32456 31628 32462 31640
rect 32493 31637 32505 31640
rect 32539 31668 32551 31671
rect 33962 31668 33968 31680
rect 32539 31640 33968 31668
rect 32539 31637 32551 31640
rect 32493 31631 32551 31637
rect 33962 31628 33968 31640
rect 34020 31628 34026 31680
rect 34698 31628 34704 31680
rect 34756 31628 34762 31680
rect 1104 31578 36524 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 36524 31578
rect 1104 31504 36524 31526
rect 5261 31467 5319 31473
rect 5261 31433 5273 31467
rect 5307 31464 5319 31467
rect 6730 31464 6736 31476
rect 5307 31436 6736 31464
rect 5307 31433 5319 31436
rect 5261 31427 5319 31433
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 7561 31467 7619 31473
rect 7561 31433 7573 31467
rect 7607 31464 7619 31467
rect 9490 31464 9496 31476
rect 7607 31436 9496 31464
rect 7607 31433 7619 31436
rect 7561 31427 7619 31433
rect 9490 31424 9496 31436
rect 9548 31424 9554 31476
rect 9861 31467 9919 31473
rect 9861 31433 9873 31467
rect 9907 31464 9919 31467
rect 11149 31467 11207 31473
rect 9907 31436 10180 31464
rect 9907 31433 9919 31436
rect 9861 31427 9919 31433
rect 10152 31408 10180 31436
rect 11149 31433 11161 31467
rect 11195 31464 11207 31467
rect 11195 31436 11652 31464
rect 11195 31433 11207 31436
rect 11149 31427 11207 31433
rect 11624 31408 11652 31436
rect 11882 31424 11888 31476
rect 11940 31424 11946 31476
rect 14734 31464 14740 31476
rect 12406 31436 13308 31464
rect 5350 31396 5356 31408
rect 5092 31368 5356 31396
rect 5092 31269 5120 31368
rect 5350 31356 5356 31368
rect 5408 31356 5414 31408
rect 6362 31396 6368 31408
rect 6104 31368 6368 31396
rect 6104 31337 6132 31368
rect 6362 31356 6368 31368
rect 6420 31396 6426 31408
rect 6457 31399 6515 31405
rect 6457 31396 6469 31399
rect 6420 31368 6469 31396
rect 6420 31356 6426 31368
rect 6457 31365 6469 31368
rect 6503 31365 6515 31399
rect 6457 31359 6515 31365
rect 7190 31356 7196 31408
rect 7248 31396 7254 31408
rect 8021 31399 8079 31405
rect 8021 31396 8033 31399
rect 7248 31368 8033 31396
rect 7248 31356 7254 31368
rect 8021 31365 8033 31368
rect 8067 31365 8079 31399
rect 8021 31359 8079 31365
rect 9677 31399 9735 31405
rect 9677 31365 9689 31399
rect 9723 31365 9735 31399
rect 9677 31359 9735 31365
rect 6089 31331 6147 31337
rect 6089 31297 6101 31331
rect 6135 31297 6147 31331
rect 6089 31291 6147 31297
rect 7285 31331 7343 31337
rect 7285 31297 7297 31331
rect 7331 31328 7343 31331
rect 7650 31328 7656 31340
rect 7331 31300 7656 31328
rect 7331 31297 7343 31300
rect 7285 31291 7343 31297
rect 7650 31288 7656 31300
rect 7708 31288 7714 31340
rect 7745 31331 7803 31337
rect 7745 31297 7757 31331
rect 7791 31297 7803 31331
rect 7745 31291 7803 31297
rect 7929 31331 7987 31337
rect 7929 31297 7941 31331
rect 7975 31328 7987 31331
rect 8202 31328 8208 31340
rect 7975 31300 8208 31328
rect 7975 31297 7987 31300
rect 7929 31291 7987 31297
rect 5077 31263 5135 31269
rect 5077 31229 5089 31263
rect 5123 31229 5135 31263
rect 5077 31223 5135 31229
rect 5169 31263 5227 31269
rect 5169 31229 5181 31263
rect 5215 31229 5227 31263
rect 5169 31223 5227 31229
rect 3694 31152 3700 31204
rect 3752 31192 3758 31204
rect 5184 31192 5212 31223
rect 3752 31164 5212 31192
rect 7760 31192 7788 31291
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 9214 31288 9220 31340
rect 9272 31288 9278 31340
rect 9306 31288 9312 31340
rect 9364 31328 9370 31340
rect 9493 31331 9551 31337
rect 9493 31328 9505 31331
rect 9364 31300 9505 31328
rect 9364 31288 9370 31300
rect 9493 31297 9505 31300
rect 9539 31297 9551 31331
rect 9493 31291 9551 31297
rect 8938 31220 8944 31272
rect 8996 31260 9002 31272
rect 9401 31263 9459 31269
rect 9401 31260 9413 31263
rect 8996 31232 9413 31260
rect 8996 31220 9002 31232
rect 9401 31229 9413 31232
rect 9447 31260 9459 31263
rect 9692 31260 9720 31359
rect 10134 31356 10140 31408
rect 10192 31356 10198 31408
rect 10778 31356 10784 31408
rect 10836 31356 10842 31408
rect 11330 31396 11336 31408
rect 10980 31368 11336 31396
rect 9950 31288 9956 31340
rect 10008 31288 10014 31340
rect 10321 31331 10379 31337
rect 10321 31297 10333 31331
rect 10367 31328 10379 31331
rect 10502 31328 10508 31340
rect 10367 31300 10508 31328
rect 10367 31297 10379 31300
rect 10321 31291 10379 31297
rect 10502 31288 10508 31300
rect 10560 31328 10566 31340
rect 10980 31337 11008 31368
rect 11330 31356 11336 31368
rect 11388 31356 11394 31408
rect 11514 31356 11520 31408
rect 11572 31356 11578 31408
rect 11606 31356 11612 31408
rect 11664 31396 11670 31408
rect 11701 31399 11759 31405
rect 11701 31396 11713 31399
rect 11664 31368 11713 31396
rect 11664 31356 11670 31368
rect 11701 31365 11713 31368
rect 11747 31365 11759 31399
rect 11701 31359 11759 31365
rect 10965 31331 11023 31337
rect 10965 31328 10977 31331
rect 10560 31300 10977 31328
rect 10560 31288 10566 31300
rect 10965 31297 10977 31300
rect 11011 31297 11023 31331
rect 10965 31291 11023 31297
rect 11054 31288 11060 31340
rect 11112 31328 11118 31340
rect 11238 31328 11244 31340
rect 11112 31300 11244 31328
rect 11112 31288 11118 31300
rect 11238 31288 11244 31300
rect 11296 31328 11302 31340
rect 11793 31331 11851 31337
rect 11793 31328 11805 31331
rect 11296 31300 11805 31328
rect 11296 31288 11302 31300
rect 11793 31297 11805 31300
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 11882 31288 11888 31340
rect 11940 31288 11946 31340
rect 12066 31288 12072 31340
rect 12124 31288 12130 31340
rect 9447 31232 9720 31260
rect 10229 31263 10287 31269
rect 9447 31229 9459 31232
rect 9401 31223 9459 31229
rect 10229 31229 10241 31263
rect 10275 31229 10287 31263
rect 12406 31260 12434 31436
rect 13280 31405 13308 31436
rect 13464 31436 14740 31464
rect 13265 31399 13323 31405
rect 13265 31365 13277 31399
rect 13311 31365 13323 31399
rect 13265 31359 13323 31365
rect 13081 31331 13139 31337
rect 13081 31297 13093 31331
rect 13127 31328 13139 31331
rect 13170 31328 13176 31340
rect 13127 31300 13176 31328
rect 13127 31297 13139 31300
rect 13081 31291 13139 31297
rect 13170 31288 13176 31300
rect 13228 31288 13234 31340
rect 13464 31337 13492 31436
rect 14734 31424 14740 31436
rect 14792 31424 14798 31476
rect 15657 31467 15715 31473
rect 15657 31433 15669 31467
rect 15703 31464 15715 31467
rect 15838 31464 15844 31476
rect 15703 31436 15844 31464
rect 15703 31433 15715 31436
rect 15657 31427 15715 31433
rect 15838 31424 15844 31436
rect 15896 31424 15902 31476
rect 16022 31424 16028 31476
rect 16080 31464 16086 31476
rect 17310 31464 17316 31476
rect 16080 31436 17316 31464
rect 16080 31424 16086 31436
rect 17310 31424 17316 31436
rect 17368 31424 17374 31476
rect 18874 31424 18880 31476
rect 18932 31424 18938 31476
rect 19426 31424 19432 31476
rect 19484 31424 19490 31476
rect 19613 31467 19671 31473
rect 19613 31433 19625 31467
rect 19659 31464 19671 31467
rect 19886 31464 19892 31476
rect 19659 31436 19892 31464
rect 19659 31433 19671 31436
rect 19613 31427 19671 31433
rect 19886 31424 19892 31436
rect 19944 31424 19950 31476
rect 20714 31424 20720 31476
rect 20772 31464 20778 31476
rect 24210 31464 24216 31476
rect 20772 31436 24216 31464
rect 20772 31424 20778 31436
rect 24210 31424 24216 31436
rect 24268 31424 24274 31476
rect 24673 31467 24731 31473
rect 24673 31464 24685 31467
rect 24504 31436 24685 31464
rect 13998 31396 14004 31408
rect 13648 31368 14004 31396
rect 13357 31331 13415 31337
rect 13357 31297 13369 31331
rect 13403 31297 13415 31331
rect 13357 31291 13415 31297
rect 13449 31331 13507 31337
rect 13449 31297 13461 31331
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 10229 31223 10287 31229
rect 10704 31232 12434 31260
rect 13372 31260 13400 31291
rect 13648 31260 13676 31368
rect 13998 31356 14004 31368
rect 14056 31356 14062 31408
rect 15286 31356 15292 31408
rect 15344 31396 15350 31408
rect 15344 31368 15792 31396
rect 15344 31356 15350 31368
rect 13722 31288 13728 31340
rect 13780 31288 13786 31340
rect 15102 31288 15108 31340
rect 15160 31288 15166 31340
rect 15764 31337 15792 31368
rect 17678 31356 17684 31408
rect 17736 31356 17742 31408
rect 18138 31356 18144 31408
rect 18196 31356 18202 31408
rect 18598 31396 18604 31408
rect 18432 31368 18604 31396
rect 15565 31331 15623 31337
rect 15565 31328 15577 31331
rect 15488 31300 15577 31328
rect 13372 31232 13676 31260
rect 14001 31263 14059 31269
rect 8478 31192 8484 31204
rect 7760 31164 8484 31192
rect 3752 31152 3758 31164
rect 8478 31152 8484 31164
rect 8536 31152 8542 31204
rect 9306 31152 9312 31204
rect 9364 31152 9370 31204
rect 9677 31195 9735 31201
rect 9677 31161 9689 31195
rect 9723 31192 9735 31195
rect 10244 31192 10272 31223
rect 10704 31201 10732 31232
rect 14001 31229 14013 31263
rect 14047 31260 14059 31263
rect 14550 31260 14556 31272
rect 14047 31232 14556 31260
rect 14047 31229 14059 31232
rect 14001 31223 14059 31229
rect 14550 31220 14556 31232
rect 14608 31220 14614 31272
rect 15010 31220 15016 31272
rect 15068 31260 15074 31272
rect 15488 31269 15516 31300
rect 15565 31297 15577 31300
rect 15611 31297 15623 31331
rect 15565 31291 15623 31297
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31328 15807 31331
rect 16850 31328 16856 31340
rect 15795 31300 16856 31328
rect 15795 31297 15807 31300
rect 15749 31291 15807 31297
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 18432 31337 18460 31368
rect 18598 31356 18604 31368
rect 18656 31396 18662 31408
rect 19150 31396 19156 31408
rect 18656 31368 19156 31396
rect 18656 31356 18662 31368
rect 19150 31356 19156 31368
rect 19208 31356 19214 31408
rect 19978 31396 19984 31408
rect 19260 31368 19984 31396
rect 18417 31331 18475 31337
rect 18417 31297 18429 31331
rect 18463 31297 18475 31331
rect 18417 31291 18475 31297
rect 18693 31331 18751 31337
rect 18693 31297 18705 31331
rect 18739 31328 18751 31331
rect 19260 31328 19288 31368
rect 18739 31300 19288 31328
rect 18739 31297 18751 31300
rect 18693 31291 18751 31297
rect 19334 31288 19340 31340
rect 19392 31288 19398 31340
rect 19426 31288 19432 31340
rect 19484 31288 19490 31340
rect 19720 31337 19748 31368
rect 19978 31356 19984 31368
rect 20036 31396 20042 31408
rect 20036 31368 21956 31396
rect 20036 31356 20042 31368
rect 19521 31331 19579 31337
rect 19521 31297 19533 31331
rect 19567 31297 19579 31331
rect 19521 31291 19579 31297
rect 19705 31331 19763 31337
rect 19705 31297 19717 31331
rect 19751 31297 19763 31331
rect 19705 31291 19763 31297
rect 15473 31263 15531 31269
rect 15473 31260 15485 31263
rect 15068 31232 15485 31260
rect 15068 31220 15074 31232
rect 15473 31229 15485 31232
rect 15519 31229 15531 31263
rect 17678 31260 17684 31272
rect 15473 31223 15531 31229
rect 15580 31232 17684 31260
rect 9723 31164 10272 31192
rect 10689 31195 10747 31201
rect 9723 31161 9735 31164
rect 9677 31155 9735 31161
rect 10689 31161 10701 31195
rect 10735 31161 10747 31195
rect 10689 31155 10747 31161
rect 11793 31195 11851 31201
rect 11793 31161 11805 31195
rect 11839 31192 11851 31195
rect 12894 31192 12900 31204
rect 11839 31164 12900 31192
rect 11839 31161 11851 31164
rect 11793 31155 11851 31161
rect 12894 31152 12900 31164
rect 12952 31152 12958 31204
rect 15102 31152 15108 31204
rect 15160 31192 15166 31204
rect 15580 31192 15608 31232
rect 17678 31220 17684 31232
rect 17736 31220 17742 31272
rect 18046 31220 18052 31272
rect 18104 31260 18110 31272
rect 18509 31263 18567 31269
rect 18509 31260 18521 31263
rect 18104 31232 18521 31260
rect 18104 31220 18110 31232
rect 18509 31229 18521 31232
rect 18555 31229 18567 31263
rect 18509 31223 18567 31229
rect 19153 31263 19211 31269
rect 19153 31229 19165 31263
rect 19199 31260 19211 31263
rect 19242 31260 19248 31272
rect 19199 31232 19248 31260
rect 19199 31229 19211 31232
rect 19153 31223 19211 31229
rect 15160 31164 15608 31192
rect 18524 31192 18552 31223
rect 19242 31220 19248 31232
rect 19300 31220 19306 31272
rect 18690 31192 18696 31204
rect 18524 31164 18696 31192
rect 15160 31152 15166 31164
rect 18690 31152 18696 31164
rect 18748 31192 18754 31204
rect 19536 31192 19564 31291
rect 19886 31288 19892 31340
rect 19944 31328 19950 31340
rect 20364 31337 20392 31368
rect 20073 31331 20131 31337
rect 20073 31328 20085 31331
rect 19944 31300 20085 31328
rect 19944 31288 19950 31300
rect 20073 31297 20085 31300
rect 20119 31297 20131 31331
rect 20073 31291 20131 31297
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31297 20315 31331
rect 20257 31291 20315 31297
rect 20349 31331 20407 31337
rect 20349 31297 20361 31331
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 20272 31260 20300 31291
rect 20548 31260 20576 31291
rect 20806 31288 20812 31340
rect 20864 31328 20870 31340
rect 21269 31331 21327 31337
rect 20864 31300 21220 31328
rect 20864 31288 20870 31300
rect 21085 31263 21143 31269
rect 21085 31260 21097 31263
rect 20272 31232 21097 31260
rect 21085 31229 21097 31232
rect 21131 31229 21143 31263
rect 21192 31260 21220 31300
rect 21269 31297 21281 31331
rect 21315 31328 21327 31331
rect 21358 31328 21364 31340
rect 21315 31300 21364 31328
rect 21315 31297 21327 31300
rect 21269 31291 21327 31297
rect 21358 31288 21364 31300
rect 21416 31288 21422 31340
rect 21450 31288 21456 31340
rect 21508 31288 21514 31340
rect 21542 31260 21548 31272
rect 21192 31232 21548 31260
rect 21085 31223 21143 31229
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 21928 31269 21956 31368
rect 22094 31356 22100 31408
rect 22152 31396 22158 31408
rect 22557 31399 22615 31405
rect 22557 31396 22569 31399
rect 22152 31368 22569 31396
rect 22152 31356 22158 31368
rect 22557 31365 22569 31368
rect 22603 31365 22615 31399
rect 22557 31359 22615 31365
rect 23842 31356 23848 31408
rect 23900 31356 23906 31408
rect 24118 31356 24124 31408
rect 24176 31396 24182 31408
rect 24504 31396 24532 31436
rect 24673 31433 24685 31436
rect 24719 31433 24731 31467
rect 24673 31427 24731 31433
rect 24762 31424 24768 31476
rect 24820 31464 24826 31476
rect 28353 31467 28411 31473
rect 24820 31436 28304 31464
rect 24820 31424 24826 31436
rect 24176 31368 24532 31396
rect 24176 31356 24182 31368
rect 24578 31356 24584 31408
rect 24636 31356 24642 31408
rect 27356 31405 27384 31436
rect 27341 31399 27399 31405
rect 27341 31365 27353 31399
rect 27387 31365 27399 31399
rect 27341 31359 27399 31365
rect 27617 31399 27675 31405
rect 27617 31365 27629 31399
rect 27663 31396 27675 31399
rect 27663 31368 27844 31396
rect 27663 31365 27675 31368
rect 27617 31359 27675 31365
rect 22005 31331 22063 31337
rect 22005 31297 22017 31331
rect 22051 31297 22063 31331
rect 22462 31328 22468 31340
rect 22005 31291 22063 31297
rect 22388 31300 22468 31328
rect 21913 31263 21971 31269
rect 21913 31229 21925 31263
rect 21959 31229 21971 31263
rect 21913 31223 21971 31229
rect 18748 31164 19564 31192
rect 18748 31152 18754 31164
rect 20070 31152 20076 31204
rect 20128 31192 20134 31204
rect 22020 31192 22048 31291
rect 22388 31269 22416 31300
rect 22462 31288 22468 31300
rect 22520 31288 22526 31340
rect 22649 31331 22707 31337
rect 22649 31297 22661 31331
rect 22695 31328 22707 31331
rect 22830 31328 22836 31340
rect 22695 31300 22836 31328
rect 22695 31297 22707 31300
rect 22649 31291 22707 31297
rect 22830 31288 22836 31300
rect 22888 31288 22894 31340
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31328 23719 31331
rect 24210 31328 24216 31340
rect 23707 31300 24216 31328
rect 23707 31297 23719 31300
rect 23661 31291 23719 31297
rect 24210 31288 24216 31300
rect 24268 31288 24274 31340
rect 24394 31288 24400 31340
rect 24452 31328 24458 31340
rect 24673 31331 24731 31337
rect 24673 31328 24685 31331
rect 24452 31300 24685 31328
rect 24452 31288 24458 31300
rect 24673 31297 24685 31300
rect 24719 31297 24731 31331
rect 24673 31291 24731 31297
rect 24854 31288 24860 31340
rect 24912 31288 24918 31340
rect 25869 31331 25927 31337
rect 25869 31297 25881 31331
rect 25915 31328 25927 31331
rect 26142 31328 26148 31340
rect 25915 31300 26148 31328
rect 25915 31297 25927 31300
rect 25869 31291 25927 31297
rect 26142 31288 26148 31300
rect 26200 31288 26206 31340
rect 27816 31337 27844 31368
rect 27982 31356 27988 31408
rect 28040 31356 28046 31408
rect 28074 31356 28080 31408
rect 28132 31356 28138 31408
rect 28276 31396 28304 31436
rect 28353 31433 28365 31467
rect 28399 31464 28411 31467
rect 29086 31464 29092 31476
rect 28399 31436 29092 31464
rect 28399 31433 28411 31436
rect 28353 31427 28411 31433
rect 29086 31424 29092 31436
rect 29144 31424 29150 31476
rect 30834 31464 30840 31476
rect 29472 31436 29868 31464
rect 29472 31396 29500 31436
rect 29730 31396 29736 31408
rect 28276 31368 29500 31396
rect 29564 31368 29736 31396
rect 27525 31331 27583 31337
rect 27525 31297 27537 31331
rect 27571 31297 27583 31331
rect 27525 31291 27583 31297
rect 27709 31331 27767 31337
rect 27709 31297 27721 31331
rect 27755 31297 27767 31331
rect 27709 31291 27767 31297
rect 27801 31331 27859 31337
rect 27801 31297 27813 31331
rect 27847 31297 27859 31331
rect 27801 31291 27859 31297
rect 28169 31331 28227 31337
rect 28169 31297 28181 31331
rect 28215 31328 28227 31331
rect 28350 31328 28356 31340
rect 28215 31300 28356 31328
rect 28215 31297 28227 31300
rect 28169 31291 28227 31297
rect 22373 31263 22431 31269
rect 22373 31229 22385 31263
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 22554 31220 22560 31272
rect 22612 31260 22618 31272
rect 23477 31263 23535 31269
rect 23477 31260 23489 31263
rect 22612 31232 23489 31260
rect 22612 31220 22618 31232
rect 23477 31229 23489 31232
rect 23523 31260 23535 31263
rect 25590 31260 25596 31272
rect 23523 31232 25596 31260
rect 23523 31229 23535 31232
rect 23477 31223 23535 31229
rect 25590 31220 25596 31232
rect 25648 31220 25654 31272
rect 25682 31220 25688 31272
rect 25740 31220 25746 31272
rect 20128 31164 22048 31192
rect 20128 31152 20134 31164
rect 5534 31084 5540 31136
rect 5592 31124 5598 31136
rect 5629 31127 5687 31133
rect 5629 31124 5641 31127
rect 5592 31096 5641 31124
rect 5592 31084 5598 31096
rect 5629 31093 5641 31096
rect 5675 31093 5687 31127
rect 5629 31087 5687 31093
rect 9030 31084 9036 31136
rect 9088 31084 9094 31136
rect 9214 31084 9220 31136
rect 9272 31124 9278 31136
rect 9950 31124 9956 31136
rect 9272 31096 9956 31124
rect 9272 31084 9278 31096
rect 9950 31084 9956 31096
rect 10008 31084 10014 31136
rect 13633 31127 13691 31133
rect 13633 31093 13645 31127
rect 13679 31124 13691 31127
rect 14182 31124 14188 31136
rect 13679 31096 14188 31124
rect 13679 31093 13691 31096
rect 13633 31087 13691 31093
rect 14182 31084 14188 31096
rect 14240 31084 14246 31136
rect 16666 31084 16672 31136
rect 16724 31084 16730 31136
rect 16758 31084 16764 31136
rect 16816 31124 16822 31136
rect 19889 31127 19947 31133
rect 19889 31124 19901 31127
rect 16816 31096 19901 31124
rect 16816 31084 16822 31096
rect 19889 31093 19901 31096
rect 19935 31093 19947 31127
rect 19889 31087 19947 31093
rect 20993 31127 21051 31133
rect 20993 31093 21005 31127
rect 21039 31124 21051 31127
rect 21266 31124 21272 31136
rect 21039 31096 21272 31124
rect 21039 31093 21051 31096
rect 20993 31087 21051 31093
rect 21266 31084 21272 31096
rect 21324 31084 21330 31136
rect 21450 31084 21456 31136
rect 21508 31124 21514 31136
rect 22572 31124 22600 31220
rect 21508 31096 22600 31124
rect 21508 31084 21514 31096
rect 25958 31084 25964 31136
rect 26016 31124 26022 31136
rect 26053 31127 26111 31133
rect 26053 31124 26065 31127
rect 26016 31096 26065 31124
rect 26016 31084 26022 31096
rect 26053 31093 26065 31096
rect 26099 31093 26111 31127
rect 26053 31087 26111 31093
rect 26602 31084 26608 31136
rect 26660 31124 26666 31136
rect 26970 31124 26976 31136
rect 26660 31096 26976 31124
rect 26660 31084 26666 31096
rect 26970 31084 26976 31096
rect 27028 31124 27034 31136
rect 27065 31127 27123 31133
rect 27065 31124 27077 31127
rect 27028 31096 27077 31124
rect 27028 31084 27034 31096
rect 27065 31093 27077 31096
rect 27111 31093 27123 31127
rect 27540 31124 27568 31291
rect 27614 31220 27620 31272
rect 27672 31260 27678 31272
rect 27724 31260 27752 31291
rect 28350 31288 28356 31300
rect 28408 31328 28414 31340
rect 28408 31300 28672 31328
rect 28408 31288 28414 31300
rect 27672 31232 27844 31260
rect 27672 31220 27678 31232
rect 27816 31192 27844 31232
rect 28258 31220 28264 31272
rect 28316 31260 28322 31272
rect 28445 31263 28503 31269
rect 28445 31260 28457 31263
rect 28316 31232 28457 31260
rect 28316 31220 28322 31232
rect 28445 31229 28457 31232
rect 28491 31229 28503 31263
rect 28644 31260 28672 31300
rect 28718 31288 28724 31340
rect 28776 31328 28782 31340
rect 28997 31331 29055 31337
rect 28997 31328 29009 31331
rect 28776 31300 29009 31328
rect 28776 31288 28782 31300
rect 28997 31297 29009 31300
rect 29043 31297 29055 31331
rect 28997 31291 29055 31297
rect 29178 31288 29184 31340
rect 29236 31288 29242 31340
rect 28810 31260 28816 31272
rect 28644 31232 28816 31260
rect 28445 31223 28503 31229
rect 28810 31220 28816 31232
rect 28868 31220 28874 31272
rect 29454 31220 29460 31272
rect 29512 31260 29518 31272
rect 29564 31269 29592 31368
rect 29730 31356 29736 31368
rect 29788 31356 29794 31408
rect 29840 31396 29868 31436
rect 30208 31436 30840 31464
rect 30208 31396 30236 31436
rect 30834 31424 30840 31436
rect 30892 31424 30898 31476
rect 32309 31467 32367 31473
rect 32309 31433 32321 31467
rect 32355 31464 32367 31467
rect 32490 31464 32496 31476
rect 32355 31436 32496 31464
rect 32355 31433 32367 31436
rect 32309 31427 32367 31433
rect 32490 31424 32496 31436
rect 32548 31424 32554 31476
rect 33410 31424 33416 31476
rect 33468 31464 33474 31476
rect 33505 31467 33563 31473
rect 33505 31464 33517 31467
rect 33468 31436 33517 31464
rect 33468 31424 33474 31436
rect 33505 31433 33517 31436
rect 33551 31433 33563 31467
rect 33505 31427 33563 31433
rect 33873 31467 33931 31473
rect 33873 31433 33885 31467
rect 33919 31464 33931 31467
rect 34698 31464 34704 31476
rect 33919 31436 34704 31464
rect 33919 31433 33931 31436
rect 33873 31427 33931 31433
rect 34698 31424 34704 31436
rect 34756 31424 34762 31476
rect 32585 31399 32643 31405
rect 29840 31368 30314 31396
rect 32585 31365 32597 31399
rect 32631 31396 32643 31399
rect 34054 31396 34060 31408
rect 32631 31368 34060 31396
rect 32631 31365 32643 31368
rect 32585 31359 32643 31365
rect 34054 31356 34060 31368
rect 34112 31356 34118 31408
rect 34422 31356 34428 31408
rect 34480 31356 34486 31408
rect 31941 31331 31999 31337
rect 31941 31297 31953 31331
rect 31987 31297 31999 31331
rect 31941 31291 31999 31297
rect 29549 31263 29607 31269
rect 29549 31260 29561 31263
rect 29512 31232 29561 31260
rect 29512 31220 29518 31232
rect 29549 31229 29561 31232
rect 29595 31229 29607 31263
rect 29549 31223 29607 31229
rect 29822 31220 29828 31272
rect 29880 31220 29886 31272
rect 30834 31220 30840 31272
rect 30892 31260 30898 31272
rect 31956 31260 31984 31291
rect 32398 31288 32404 31340
rect 32456 31328 32462 31340
rect 32493 31331 32551 31337
rect 32493 31328 32505 31331
rect 32456 31300 32505 31328
rect 32456 31288 32462 31300
rect 32493 31297 32505 31300
rect 32539 31297 32551 31331
rect 32493 31291 32551 31297
rect 32674 31288 32680 31340
rect 32732 31288 32738 31340
rect 32861 31331 32919 31337
rect 32861 31297 32873 31331
rect 32907 31328 32919 31331
rect 33042 31328 33048 31340
rect 32907 31300 33048 31328
rect 32907 31297 32919 31300
rect 32861 31291 32919 31297
rect 33042 31288 33048 31300
rect 33100 31288 33106 31340
rect 33689 31331 33747 31337
rect 33689 31297 33701 31331
rect 33735 31328 33747 31331
rect 33870 31328 33876 31340
rect 33735 31300 33876 31328
rect 33735 31297 33747 31300
rect 33689 31291 33747 31297
rect 33870 31288 33876 31300
rect 33928 31288 33934 31340
rect 33962 31288 33968 31340
rect 34020 31288 34026 31340
rect 34241 31331 34299 31337
rect 34241 31297 34253 31331
rect 34287 31328 34299 31331
rect 34514 31328 34520 31340
rect 34287 31300 34520 31328
rect 34287 31297 34299 31300
rect 34241 31291 34299 31297
rect 34514 31288 34520 31300
rect 34572 31288 34578 31340
rect 34146 31260 34152 31272
rect 30892 31232 34152 31260
rect 30892 31220 30898 31232
rect 34146 31220 34152 31232
rect 34204 31220 34210 31272
rect 29086 31192 29092 31204
rect 27816 31164 29092 31192
rect 29086 31152 29092 31164
rect 29144 31152 29150 31204
rect 31110 31152 31116 31204
rect 31168 31192 31174 31204
rect 34057 31195 34115 31201
rect 34057 31192 34069 31195
rect 31168 31164 34069 31192
rect 31168 31152 31174 31164
rect 34057 31161 34069 31164
rect 34103 31161 34115 31195
rect 34057 31155 34115 31161
rect 27614 31124 27620 31136
rect 27540 31096 27620 31124
rect 27065 31087 27123 31093
rect 27614 31084 27620 31096
rect 27672 31084 27678 31136
rect 27706 31084 27712 31136
rect 27764 31124 27770 31136
rect 29365 31127 29423 31133
rect 29365 31124 29377 31127
rect 27764 31096 29377 31124
rect 27764 31084 27770 31096
rect 29365 31093 29377 31096
rect 29411 31124 29423 31127
rect 30190 31124 30196 31136
rect 29411 31096 30196 31124
rect 29411 31093 29423 31096
rect 29365 31087 29423 31093
rect 30190 31084 30196 31096
rect 30248 31084 30254 31136
rect 31294 31084 31300 31136
rect 31352 31124 31358 31136
rect 31662 31124 31668 31136
rect 31352 31096 31668 31124
rect 31352 31084 31358 31096
rect 31662 31084 31668 31096
rect 31720 31084 31726 31136
rect 33318 31084 33324 31136
rect 33376 31124 33382 31136
rect 34422 31124 34428 31136
rect 33376 31096 34428 31124
rect 33376 31084 33382 31096
rect 34422 31084 34428 31096
rect 34480 31084 34486 31136
rect 1104 31034 36524 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 36524 31034
rect 1104 30960 36524 30982
rect 8938 30880 8944 30932
rect 8996 30920 9002 30932
rect 8996 30892 9260 30920
rect 8996 30880 9002 30892
rect 8386 30812 8392 30864
rect 8444 30852 8450 30864
rect 8570 30852 8576 30864
rect 8444 30824 8576 30852
rect 8444 30812 8450 30824
rect 8570 30812 8576 30824
rect 8628 30852 8634 30864
rect 9122 30852 9128 30864
rect 8628 30824 9128 30852
rect 8628 30812 8634 30824
rect 9122 30812 9128 30824
rect 9180 30812 9186 30864
rect 9232 30852 9260 30892
rect 9306 30880 9312 30932
rect 9364 30920 9370 30932
rect 9401 30923 9459 30929
rect 9401 30920 9413 30923
rect 9364 30892 9413 30920
rect 9364 30880 9370 30892
rect 9401 30889 9413 30892
rect 9447 30889 9459 30923
rect 10962 30920 10968 30932
rect 9401 30883 9459 30889
rect 9692 30892 10968 30920
rect 9585 30855 9643 30861
rect 9585 30852 9597 30855
rect 9232 30824 9597 30852
rect 9585 30821 9597 30824
rect 9631 30821 9643 30855
rect 9585 30815 9643 30821
rect 6914 30744 6920 30796
rect 6972 30744 6978 30796
rect 9692 30784 9720 30892
rect 10962 30880 10968 30892
rect 11020 30880 11026 30932
rect 11698 30880 11704 30932
rect 11756 30920 11762 30932
rect 11882 30920 11888 30932
rect 11756 30892 11888 30920
rect 11756 30880 11762 30892
rect 11882 30880 11888 30892
rect 11940 30920 11946 30932
rect 14458 30920 14464 30932
rect 11940 30892 14464 30920
rect 11940 30880 11946 30892
rect 14458 30880 14464 30892
rect 14516 30880 14522 30932
rect 14550 30880 14556 30932
rect 14608 30880 14614 30932
rect 16853 30923 16911 30929
rect 16853 30889 16865 30923
rect 16899 30920 16911 30923
rect 16899 30892 16988 30920
rect 16899 30889 16911 30892
rect 16853 30883 16911 30889
rect 9953 30855 10011 30861
rect 9953 30821 9965 30855
rect 9999 30852 10011 30855
rect 10778 30852 10784 30864
rect 9999 30824 10784 30852
rect 9999 30821 10011 30824
rect 9953 30815 10011 30821
rect 10778 30812 10784 30824
rect 10836 30812 10842 30864
rect 12066 30812 12072 30864
rect 12124 30852 12130 30864
rect 16960 30852 16988 30892
rect 17034 30880 17040 30932
rect 17092 30920 17098 30932
rect 17405 30923 17463 30929
rect 17405 30920 17417 30923
rect 17092 30892 17417 30920
rect 17092 30880 17098 30892
rect 17405 30889 17417 30892
rect 17451 30889 17463 30923
rect 17405 30883 17463 30889
rect 17678 30880 17684 30932
rect 17736 30920 17742 30932
rect 17773 30923 17831 30929
rect 17773 30920 17785 30923
rect 17736 30892 17785 30920
rect 17736 30880 17742 30892
rect 17773 30889 17785 30892
rect 17819 30889 17831 30923
rect 17773 30883 17831 30889
rect 17862 30880 17868 30932
rect 17920 30920 17926 30932
rect 17920 30892 20944 30920
rect 17920 30880 17926 30892
rect 18230 30852 18236 30864
rect 12124 30824 16896 30852
rect 16960 30824 18236 30852
rect 12124 30812 12130 30824
rect 8588 30756 9720 30784
rect 5166 30676 5172 30728
rect 5224 30676 5230 30728
rect 7190 30676 7196 30728
rect 7248 30716 7254 30728
rect 8588 30725 8616 30756
rect 10042 30744 10048 30796
rect 10100 30744 10106 30796
rect 14550 30744 14556 30796
rect 14608 30784 14614 30796
rect 16761 30787 16819 30793
rect 16761 30784 16773 30787
rect 14608 30756 16773 30784
rect 14608 30744 14614 30756
rect 16761 30753 16773 30756
rect 16807 30753 16819 30787
rect 16868 30784 16896 30824
rect 18230 30812 18236 30824
rect 18288 30812 18294 30864
rect 20806 30852 20812 30864
rect 20548 30824 20812 30852
rect 20548 30784 20576 30824
rect 20806 30812 20812 30824
rect 20864 30812 20870 30864
rect 20916 30852 20944 30892
rect 20990 30880 20996 30932
rect 21048 30880 21054 30932
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21177 30923 21235 30929
rect 21177 30920 21189 30923
rect 21140 30892 21189 30920
rect 21140 30880 21146 30892
rect 21177 30889 21189 30892
rect 21223 30889 21235 30923
rect 21177 30883 21235 30889
rect 22278 30880 22284 30932
rect 22336 30920 22342 30932
rect 22833 30923 22891 30929
rect 22833 30920 22845 30923
rect 22336 30892 22845 30920
rect 22336 30880 22342 30892
rect 22833 30889 22845 30892
rect 22879 30889 22891 30923
rect 22833 30883 22891 30889
rect 24854 30880 24860 30932
rect 24912 30920 24918 30932
rect 25133 30923 25191 30929
rect 25133 30920 25145 30923
rect 24912 30892 25145 30920
rect 24912 30880 24918 30892
rect 25133 30889 25145 30892
rect 25179 30889 25191 30923
rect 25133 30883 25191 30889
rect 28810 30880 28816 30932
rect 28868 30920 28874 30932
rect 29641 30923 29699 30929
rect 28868 30892 29500 30920
rect 28868 30880 28874 30892
rect 21450 30852 21456 30864
rect 20916 30824 21456 30852
rect 21450 30812 21456 30824
rect 21508 30812 21514 30864
rect 23477 30855 23535 30861
rect 23477 30821 23489 30855
rect 23523 30852 23535 30855
rect 23566 30852 23572 30864
rect 23523 30824 23572 30852
rect 23523 30821 23535 30824
rect 23477 30815 23535 30821
rect 23566 30812 23572 30824
rect 23624 30812 23630 30864
rect 27798 30812 27804 30864
rect 27856 30852 27862 30864
rect 27985 30855 28043 30861
rect 27985 30852 27997 30855
rect 27856 30824 27997 30852
rect 27856 30812 27862 30824
rect 27985 30821 27997 30824
rect 28031 30852 28043 30855
rect 29270 30852 29276 30864
rect 28031 30824 29276 30852
rect 28031 30821 28043 30824
rect 27985 30815 28043 30821
rect 29270 30812 29276 30824
rect 29328 30812 29334 30864
rect 29365 30855 29423 30861
rect 29365 30821 29377 30855
rect 29411 30821 29423 30855
rect 29472 30852 29500 30892
rect 29641 30889 29653 30923
rect 29687 30920 29699 30923
rect 29914 30920 29920 30932
rect 29687 30892 29920 30920
rect 29687 30889 29699 30892
rect 29641 30883 29699 30889
rect 29914 30880 29920 30892
rect 29972 30880 29978 30932
rect 30926 30880 30932 30932
rect 30984 30920 30990 30932
rect 34330 30920 34336 30932
rect 30984 30892 34336 30920
rect 30984 30880 30990 30892
rect 34330 30880 34336 30892
rect 34388 30880 34394 30932
rect 29733 30855 29791 30861
rect 29733 30852 29745 30855
rect 29472 30824 29745 30852
rect 29365 30815 29423 30821
rect 29733 30821 29745 30824
rect 29779 30852 29791 30855
rect 31018 30852 31024 30864
rect 29779 30824 31024 30852
rect 29779 30821 29791 30824
rect 29733 30815 29791 30821
rect 16868 30756 20576 30784
rect 20640 30756 21312 30784
rect 16761 30747 16819 30753
rect 8573 30719 8631 30725
rect 8573 30716 8585 30719
rect 7248 30688 8585 30716
rect 7248 30676 7254 30688
rect 8573 30685 8585 30688
rect 8619 30685 8631 30719
rect 8573 30679 8631 30685
rect 8941 30719 8999 30725
rect 8941 30685 8953 30719
rect 8987 30685 8999 30719
rect 8941 30679 8999 30685
rect 9033 30719 9091 30725
rect 9033 30685 9045 30719
rect 9079 30685 9091 30719
rect 9033 30679 9091 30685
rect 4062 30608 4068 30660
rect 4120 30648 4126 30660
rect 5626 30648 5632 30660
rect 4120 30620 5632 30648
rect 4120 30608 4126 30620
rect 5626 30608 5632 30620
rect 5684 30648 5690 30660
rect 7653 30651 7711 30657
rect 5684 30620 5750 30648
rect 5684 30608 5690 30620
rect 7653 30617 7665 30651
rect 7699 30617 7711 30651
rect 7653 30611 7711 30617
rect 7098 30540 7104 30592
rect 7156 30580 7162 30592
rect 7282 30580 7288 30592
rect 7156 30552 7288 30580
rect 7156 30540 7162 30552
rect 7282 30540 7288 30552
rect 7340 30580 7346 30592
rect 7377 30583 7435 30589
rect 7377 30580 7389 30583
rect 7340 30552 7389 30580
rect 7340 30540 7346 30552
rect 7377 30549 7389 30552
rect 7423 30549 7435 30583
rect 7668 30580 7696 30611
rect 7834 30608 7840 30660
rect 7892 30608 7898 30660
rect 8202 30608 8208 30660
rect 8260 30648 8266 30660
rect 8956 30648 8984 30679
rect 8260 30620 8984 30648
rect 9048 30648 9076 30679
rect 9122 30676 9128 30728
rect 9180 30716 9186 30728
rect 9217 30719 9275 30725
rect 9217 30716 9229 30719
rect 9180 30688 9229 30716
rect 9180 30676 9186 30688
rect 9217 30685 9229 30688
rect 9263 30685 9275 30719
rect 9582 30716 9588 30728
rect 9217 30679 9275 30685
rect 9497 30688 9588 30716
rect 9497 30648 9525 30688
rect 9582 30676 9588 30688
rect 9640 30676 9646 30728
rect 9766 30676 9772 30728
rect 9824 30676 9830 30728
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30685 9919 30719
rect 10060 30715 10088 30744
rect 9861 30679 9919 30685
rect 10045 30709 10103 30715
rect 9048 30620 9525 30648
rect 8260 30608 8266 30620
rect 9674 30608 9680 30660
rect 9732 30648 9738 30660
rect 9876 30648 9904 30679
rect 10045 30675 10057 30709
rect 10091 30675 10103 30709
rect 11146 30676 11152 30728
rect 11204 30676 11210 30728
rect 14182 30676 14188 30728
rect 14240 30676 14246 30728
rect 14369 30719 14427 30725
rect 14369 30685 14381 30719
rect 14415 30716 14427 30719
rect 15654 30716 15660 30728
rect 14415 30688 15660 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 15654 30676 15660 30688
rect 15712 30676 15718 30728
rect 16666 30676 16672 30728
rect 16724 30716 16730 30728
rect 17126 30716 17132 30728
rect 16724 30688 17132 30716
rect 16724 30676 16730 30688
rect 17126 30676 17132 30688
rect 17184 30716 17190 30728
rect 17224 30719 17282 30725
rect 17224 30716 17236 30719
rect 17184 30688 17236 30716
rect 17184 30676 17190 30688
rect 17224 30685 17236 30688
rect 17270 30685 17282 30719
rect 17224 30679 17282 30685
rect 17310 30676 17316 30728
rect 17368 30716 17374 30728
rect 20640 30725 20668 30756
rect 21284 30728 21312 30756
rect 21358 30744 21364 30796
rect 21416 30784 21422 30796
rect 22922 30784 22928 30796
rect 21416 30756 22928 30784
rect 21416 30744 21422 30756
rect 22922 30744 22928 30756
rect 22980 30744 22986 30796
rect 25041 30787 25099 30793
rect 25041 30784 25053 30787
rect 24688 30756 25053 30784
rect 24688 30728 24716 30756
rect 25041 30753 25053 30756
rect 25087 30753 25099 30787
rect 25041 30747 25099 30753
rect 25593 30787 25651 30793
rect 25593 30753 25605 30787
rect 25639 30784 25651 30787
rect 25774 30784 25780 30796
rect 25639 30756 25780 30784
rect 25639 30753 25651 30756
rect 25593 30747 25651 30753
rect 25774 30744 25780 30756
rect 25832 30744 25838 30796
rect 25958 30744 25964 30796
rect 26016 30744 26022 30796
rect 26142 30744 26148 30796
rect 26200 30784 26206 30796
rect 26200 30756 27936 30784
rect 26200 30744 26206 30756
rect 17681 30719 17739 30725
rect 17681 30716 17693 30719
rect 17368 30688 17693 30716
rect 17368 30676 17374 30688
rect 17681 30685 17693 30688
rect 17727 30685 17739 30719
rect 17681 30679 17739 30685
rect 20625 30719 20683 30725
rect 20625 30685 20637 30719
rect 20671 30685 20683 30719
rect 21085 30719 21143 30725
rect 21085 30716 21097 30719
rect 20625 30679 20683 30685
rect 20824 30688 21097 30716
rect 10045 30669 10103 30675
rect 9950 30648 9956 30660
rect 9732 30620 9956 30648
rect 9732 30608 9738 30620
rect 9950 30608 9956 30620
rect 10008 30608 10014 30660
rect 10318 30608 10324 30660
rect 10376 30648 10382 30660
rect 16758 30648 16764 30660
rect 10376 30620 16764 30648
rect 10376 30608 10382 30620
rect 16758 30608 16764 30620
rect 16816 30608 16822 30660
rect 16868 30620 17632 30648
rect 8846 30580 8852 30592
rect 7668 30552 8852 30580
rect 7377 30543 7435 30549
rect 8846 30540 8852 30552
rect 8904 30540 8910 30592
rect 11238 30540 11244 30592
rect 11296 30540 11302 30592
rect 13906 30540 13912 30592
rect 13964 30580 13970 30592
rect 16868 30580 16896 30620
rect 13964 30552 16896 30580
rect 17221 30583 17279 30589
rect 13964 30540 13970 30552
rect 17221 30549 17233 30583
rect 17267 30580 17279 30583
rect 17494 30580 17500 30592
rect 17267 30552 17500 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 17494 30540 17500 30552
rect 17552 30540 17558 30592
rect 17604 30580 17632 30620
rect 19886 30608 19892 30660
rect 19944 30648 19950 30660
rect 20824 30657 20852 30688
rect 21085 30685 21097 30688
rect 21131 30685 21143 30719
rect 21085 30679 21143 30685
rect 21266 30676 21272 30728
rect 21324 30676 21330 30728
rect 23106 30676 23112 30728
rect 23164 30676 23170 30728
rect 23198 30676 23204 30728
rect 23256 30716 23262 30728
rect 23293 30719 23351 30725
rect 23293 30716 23305 30719
rect 23256 30688 23305 30716
rect 23256 30676 23262 30688
rect 23293 30685 23305 30688
rect 23339 30685 23351 30719
rect 23293 30679 23351 30685
rect 23569 30719 23627 30725
rect 23569 30685 23581 30719
rect 23615 30685 23627 30719
rect 23569 30679 23627 30685
rect 20809 30651 20867 30657
rect 20809 30648 20821 30651
rect 19944 30620 20821 30648
rect 19944 30608 19950 30620
rect 20809 30617 20821 30620
rect 20855 30617 20867 30651
rect 20809 30611 20867 30617
rect 22922 30608 22928 30660
rect 22980 30648 22986 30660
rect 23584 30648 23612 30679
rect 24670 30676 24676 30728
rect 24728 30676 24734 30728
rect 24854 30676 24860 30728
rect 24912 30676 24918 30728
rect 25222 30676 25228 30728
rect 25280 30676 25286 30728
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30716 25375 30719
rect 25682 30716 25688 30728
rect 25363 30688 25688 30716
rect 25363 30685 25375 30688
rect 25317 30679 25375 30685
rect 22980 30620 23612 30648
rect 22980 30608 22986 30620
rect 23750 30608 23756 30660
rect 23808 30648 23814 30660
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 23808 30620 24593 30648
rect 23808 30608 23814 30620
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24872 30648 24900 30676
rect 25332 30648 25360 30679
rect 25682 30676 25688 30688
rect 25740 30676 25746 30728
rect 27706 30676 27712 30728
rect 27764 30676 27770 30728
rect 24872 30620 25360 30648
rect 24581 30611 24639 30617
rect 23014 30580 23020 30592
rect 17604 30552 23020 30580
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 23201 30583 23259 30589
rect 23201 30549 23213 30583
rect 23247 30580 23259 30583
rect 23658 30580 23664 30592
rect 23247 30552 23664 30580
rect 23247 30549 23259 30552
rect 23201 30543 23259 30549
rect 23658 30540 23664 30552
rect 23716 30540 23722 30592
rect 25700 30580 25728 30676
rect 26970 30608 26976 30660
rect 27028 30608 27034 30660
rect 27338 30580 27344 30592
rect 25700 30552 27344 30580
rect 27338 30540 27344 30552
rect 27396 30589 27402 30592
rect 27396 30583 27445 30589
rect 27396 30549 27399 30583
rect 27433 30549 27445 30583
rect 27908 30580 27936 30756
rect 28166 30744 28172 30796
rect 28224 30784 28230 30796
rect 28813 30787 28871 30793
rect 28813 30784 28825 30787
rect 28224 30756 28825 30784
rect 28224 30744 28230 30756
rect 28813 30753 28825 30756
rect 28859 30753 28871 30787
rect 29380 30784 29408 30815
rect 31018 30812 31024 30824
rect 31076 30852 31082 30864
rect 32490 30852 32496 30864
rect 31076 30824 32496 30852
rect 31076 30812 31082 30824
rect 32490 30812 32496 30824
rect 32548 30812 32554 30864
rect 29549 30787 29607 30793
rect 29549 30784 29561 30787
rect 29380 30756 29561 30784
rect 28813 30747 28871 30753
rect 29549 30753 29561 30756
rect 29595 30753 29607 30787
rect 30745 30787 30803 30793
rect 29549 30747 29607 30753
rect 29656 30756 29868 30784
rect 28074 30676 28080 30728
rect 28132 30716 28138 30728
rect 28721 30719 28779 30725
rect 28721 30716 28733 30719
rect 28132 30688 28733 30716
rect 28132 30676 28138 30688
rect 28721 30685 28733 30688
rect 28767 30685 28779 30719
rect 28721 30679 28779 30685
rect 29240 30719 29298 30725
rect 29240 30685 29252 30719
rect 29286 30716 29298 30719
rect 29656 30716 29684 30756
rect 29840 30725 29868 30756
rect 30745 30753 30757 30787
rect 30791 30784 30803 30787
rect 30834 30784 30840 30796
rect 30791 30756 30840 30784
rect 30791 30753 30803 30756
rect 30745 30747 30803 30753
rect 30834 30744 30840 30756
rect 30892 30744 30898 30796
rect 32306 30744 32312 30796
rect 32364 30784 32370 30796
rect 32585 30787 32643 30793
rect 32585 30784 32597 30787
rect 32364 30756 32597 30784
rect 32364 30744 32370 30756
rect 32585 30753 32597 30756
rect 32631 30753 32643 30787
rect 32585 30747 32643 30753
rect 29286 30688 29684 30716
rect 29825 30719 29883 30725
rect 29286 30685 29298 30688
rect 29240 30679 29298 30685
rect 29825 30685 29837 30719
rect 29871 30716 29883 30719
rect 30006 30716 30012 30728
rect 29871 30688 30012 30716
rect 29871 30685 29883 30688
rect 29825 30679 29883 30685
rect 30006 30676 30012 30688
rect 30064 30676 30070 30728
rect 30650 30676 30656 30728
rect 30708 30716 30714 30728
rect 30929 30719 30987 30725
rect 30929 30716 30941 30719
rect 30708 30688 30941 30716
rect 30708 30676 30714 30688
rect 30929 30685 30941 30688
rect 30975 30685 30987 30719
rect 30929 30679 30987 30685
rect 28169 30651 28227 30657
rect 28169 30617 28181 30651
rect 28215 30648 28227 30651
rect 29454 30648 29460 30660
rect 28215 30620 29460 30648
rect 28215 30617 28227 30620
rect 28169 30611 28227 30617
rect 29454 30608 29460 30620
rect 29512 30608 29518 30660
rect 29638 30608 29644 30660
rect 29696 30648 29702 30660
rect 29917 30651 29975 30657
rect 29917 30648 29929 30651
rect 29696 30620 29929 30648
rect 29696 30608 29702 30620
rect 29917 30617 29929 30620
rect 29963 30617 29975 30651
rect 29917 30611 29975 30617
rect 32858 30608 32864 30660
rect 32916 30608 32922 30660
rect 34422 30648 34428 30660
rect 34086 30620 34428 30648
rect 34422 30608 34428 30620
rect 34480 30608 34486 30660
rect 29181 30583 29239 30589
rect 29181 30580 29193 30583
rect 27908 30552 29193 30580
rect 27396 30543 27445 30549
rect 29181 30549 29193 30552
rect 29227 30580 29239 30583
rect 31018 30580 31024 30592
rect 29227 30552 31024 30580
rect 29227 30549 29239 30552
rect 29181 30543 29239 30549
rect 27396 30540 27402 30543
rect 31018 30540 31024 30552
rect 31076 30540 31082 30592
rect 31110 30540 31116 30592
rect 31168 30540 31174 30592
rect 33226 30540 33232 30592
rect 33284 30580 33290 30592
rect 34333 30583 34391 30589
rect 34333 30580 34345 30583
rect 33284 30552 34345 30580
rect 33284 30540 33290 30552
rect 34333 30549 34345 30552
rect 34379 30549 34391 30583
rect 34333 30543 34391 30549
rect 1104 30490 36524 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 36524 30490
rect 1104 30416 36524 30438
rect 5626 30336 5632 30388
rect 5684 30336 5690 30388
rect 8018 30336 8024 30388
rect 8076 30376 8082 30388
rect 8076 30348 8616 30376
rect 8076 30336 8082 30348
rect 3694 30268 3700 30320
rect 3752 30268 3758 30320
rect 4062 30268 4068 30320
rect 4120 30308 4126 30320
rect 5445 30311 5503 30317
rect 4120 30280 4278 30308
rect 4120 30268 4126 30280
rect 5445 30277 5457 30311
rect 5491 30308 5503 30311
rect 5534 30308 5540 30320
rect 5491 30280 5540 30308
rect 5491 30277 5503 30280
rect 5445 30271 5503 30277
rect 5534 30268 5540 30280
rect 5592 30268 5598 30320
rect 5644 30308 5672 30336
rect 7098 30308 7104 30320
rect 5644 30280 7104 30308
rect 7098 30268 7104 30280
rect 7156 30268 7162 30320
rect 8588 30308 8616 30348
rect 8754 30336 8760 30388
rect 8812 30376 8818 30388
rect 9125 30379 9183 30385
rect 8812 30348 9076 30376
rect 8812 30336 8818 30348
rect 9048 30308 9076 30348
rect 9125 30345 9137 30379
rect 9171 30376 9183 30379
rect 9214 30376 9220 30388
rect 9171 30348 9220 30376
rect 9171 30345 9183 30348
rect 9125 30339 9183 30345
rect 9214 30336 9220 30348
rect 9272 30336 9278 30388
rect 11146 30376 11152 30388
rect 9324 30348 11152 30376
rect 9324 30308 9352 30348
rect 11146 30336 11152 30348
rect 11204 30336 11210 30388
rect 14458 30336 14464 30388
rect 14516 30376 14522 30388
rect 19886 30376 19892 30388
rect 14516 30348 19892 30376
rect 14516 30336 14522 30348
rect 8220 30280 8524 30308
rect 8588 30280 8892 30308
rect 9048 30280 9352 30308
rect 5721 30243 5779 30249
rect 5721 30209 5733 30243
rect 5767 30240 5779 30243
rect 5810 30240 5816 30252
rect 5767 30212 5816 30240
rect 5767 30209 5779 30212
rect 5721 30203 5779 30209
rect 5810 30200 5816 30212
rect 5868 30240 5874 30252
rect 6270 30240 6276 30252
rect 5868 30212 6276 30240
rect 5868 30200 5874 30212
rect 6270 30200 6276 30212
rect 6328 30240 6334 30252
rect 8220 30249 8248 30280
rect 8496 30252 8524 30280
rect 8864 30252 8892 30280
rect 9398 30268 9404 30320
rect 9456 30308 9462 30320
rect 17972 30317 18000 30348
rect 19886 30336 19892 30348
rect 19944 30336 19950 30388
rect 20346 30336 20352 30388
rect 20404 30376 20410 30388
rect 23290 30376 23296 30388
rect 20404 30348 23296 30376
rect 20404 30336 20410 30348
rect 23290 30336 23296 30348
rect 23348 30336 23354 30388
rect 23658 30336 23664 30388
rect 23716 30376 23722 30388
rect 24762 30376 24768 30388
rect 23716 30348 24768 30376
rect 23716 30336 23722 30348
rect 24762 30336 24768 30348
rect 24820 30336 24826 30388
rect 28626 30376 28632 30388
rect 27264 30348 28632 30376
rect 17957 30311 18015 30317
rect 9456 30280 17908 30308
rect 9456 30268 9462 30280
rect 6365 30243 6423 30249
rect 6365 30240 6377 30243
rect 6328 30212 6377 30240
rect 6328 30200 6334 30212
rect 6365 30209 6377 30212
rect 6411 30209 6423 30243
rect 6365 30203 6423 30209
rect 8205 30243 8263 30249
rect 8205 30209 8217 30243
rect 8251 30209 8263 30243
rect 8205 30203 8263 30209
rect 8389 30243 8447 30249
rect 8389 30209 8401 30243
rect 8435 30209 8447 30243
rect 8389 30203 8447 30209
rect 6638 30132 6644 30184
rect 6696 30132 6702 30184
rect 6730 30132 6736 30184
rect 6788 30172 6794 30184
rect 6788 30144 8248 30172
rect 6788 30132 6794 30144
rect 8220 30113 8248 30144
rect 8294 30132 8300 30184
rect 8352 30172 8358 30184
rect 8404 30172 8432 30203
rect 8478 30200 8484 30252
rect 8536 30240 8542 30252
rect 8573 30243 8631 30249
rect 8573 30240 8585 30243
rect 8536 30212 8585 30240
rect 8536 30200 8542 30212
rect 8573 30209 8585 30212
rect 8619 30209 8631 30243
rect 8573 30203 8631 30209
rect 8757 30243 8815 30249
rect 8757 30209 8769 30243
rect 8803 30209 8815 30243
rect 8757 30203 8815 30209
rect 8772 30172 8800 30203
rect 8846 30200 8852 30252
rect 8904 30240 8910 30252
rect 9033 30243 9091 30249
rect 9033 30240 9045 30243
rect 8904 30212 9045 30240
rect 8904 30200 8910 30212
rect 9033 30209 9045 30212
rect 9079 30209 9091 30243
rect 9033 30203 9091 30209
rect 9217 30243 9275 30249
rect 9217 30209 9229 30243
rect 9263 30240 9275 30243
rect 9490 30240 9496 30252
rect 9263 30212 9496 30240
rect 9263 30209 9275 30212
rect 9217 30203 9275 30209
rect 9490 30200 9496 30212
rect 9548 30200 9554 30252
rect 9769 30243 9827 30249
rect 9769 30209 9781 30243
rect 9815 30209 9827 30243
rect 9769 30203 9827 30209
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30240 10011 30243
rect 10042 30240 10048 30252
rect 9999 30212 10048 30240
rect 9999 30209 10011 30212
rect 9953 30203 10011 30209
rect 9784 30172 9812 30203
rect 10042 30200 10048 30212
rect 10100 30240 10106 30252
rect 10870 30240 10876 30252
rect 10100 30212 10876 30240
rect 10100 30200 10106 30212
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 17880 30249 17908 30280
rect 17957 30277 17969 30311
rect 18003 30277 18015 30311
rect 17957 30271 18015 30277
rect 18782 30268 18788 30320
rect 18840 30308 18846 30320
rect 18877 30311 18935 30317
rect 18877 30308 18889 30311
rect 18840 30280 18889 30308
rect 18840 30268 18846 30280
rect 18877 30277 18889 30280
rect 18923 30277 18935 30311
rect 20254 30308 20260 30320
rect 20102 30280 20260 30308
rect 18877 30271 18935 30277
rect 20254 30268 20260 30280
rect 20312 30308 20318 30320
rect 20312 30280 24518 30308
rect 20312 30268 20318 30280
rect 26234 30268 26240 30320
rect 26292 30308 26298 30320
rect 26513 30311 26571 30317
rect 26513 30308 26525 30311
rect 26292 30280 26525 30308
rect 26292 30268 26298 30280
rect 26513 30277 26525 30280
rect 26559 30277 26571 30311
rect 26513 30271 26571 30277
rect 26602 30268 26608 30320
rect 26660 30308 26666 30320
rect 26697 30311 26755 30317
rect 26697 30308 26709 30311
rect 26660 30280 26709 30308
rect 26660 30268 26666 30280
rect 26697 30277 26709 30280
rect 26743 30308 26755 30311
rect 27264 30308 27292 30348
rect 28626 30336 28632 30348
rect 28684 30336 28690 30388
rect 29178 30376 29184 30388
rect 28736 30348 29184 30376
rect 27985 30311 28043 30317
rect 27985 30308 27997 30311
rect 26743 30280 27292 30308
rect 27356 30280 27997 30308
rect 26743 30277 26755 30280
rect 26697 30271 26755 30277
rect 27356 30252 27384 30280
rect 27985 30277 27997 30280
rect 28031 30277 28043 30311
rect 27985 30271 28043 30277
rect 28169 30311 28227 30317
rect 28169 30277 28181 30311
rect 28215 30308 28227 30311
rect 28736 30308 28764 30348
rect 29178 30336 29184 30348
rect 29236 30336 29242 30388
rect 29270 30336 29276 30388
rect 29328 30376 29334 30388
rect 29914 30376 29920 30388
rect 29328 30348 29920 30376
rect 29328 30336 29334 30348
rect 29914 30336 29920 30348
rect 29972 30336 29978 30388
rect 31021 30379 31079 30385
rect 31021 30345 31033 30379
rect 31067 30345 31079 30379
rect 31021 30339 31079 30345
rect 28215 30280 28764 30308
rect 28215 30277 28227 30280
rect 28169 30271 28227 30277
rect 29730 30268 29736 30320
rect 29788 30308 29794 30320
rect 29788 30280 30512 30308
rect 29788 30268 29794 30280
rect 17865 30243 17923 30249
rect 17865 30209 17877 30243
rect 17911 30240 17923 30243
rect 18138 30240 18144 30252
rect 17911 30212 18144 30240
rect 17911 30209 17923 30212
rect 17865 30203 17923 30209
rect 18138 30200 18144 30212
rect 18196 30200 18202 30252
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30240 18291 30243
rect 18506 30240 18512 30252
rect 18279 30212 18512 30240
rect 18279 30209 18291 30212
rect 18233 30203 18291 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 18598 30200 18604 30252
rect 18656 30200 18662 30252
rect 22922 30200 22928 30252
rect 22980 30200 22986 30252
rect 23017 30243 23075 30249
rect 23017 30209 23029 30243
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 8352 30144 17632 30172
rect 8352 30132 8358 30144
rect 8205 30107 8263 30113
rect 8205 30073 8217 30107
rect 8251 30073 8263 30107
rect 8205 30067 8263 30073
rect 9953 30107 10011 30113
rect 9953 30073 9965 30107
rect 9999 30073 10011 30107
rect 9953 30067 10011 30073
rect 8110 29996 8116 30048
rect 8168 29996 8174 30048
rect 8941 30039 8999 30045
rect 8941 30005 8953 30039
rect 8987 30036 8999 30039
rect 9122 30036 9128 30048
rect 8987 30008 9128 30036
rect 8987 30005 8999 30008
rect 8941 29999 8999 30005
rect 9122 29996 9128 30008
rect 9180 30036 9186 30048
rect 9490 30036 9496 30048
rect 9180 30008 9496 30036
rect 9180 29996 9186 30008
rect 9490 29996 9496 30008
rect 9548 29996 9554 30048
rect 9968 30036 9996 30067
rect 10134 30064 10140 30116
rect 10192 30104 10198 30116
rect 16942 30104 16948 30116
rect 10192 30076 16948 30104
rect 10192 30064 10198 30076
rect 16942 30064 16948 30076
rect 17000 30064 17006 30116
rect 17604 30104 17632 30144
rect 17678 30132 17684 30184
rect 17736 30172 17742 30184
rect 18414 30172 18420 30184
rect 17736 30144 18420 30172
rect 17736 30132 17742 30144
rect 18414 30132 18420 30144
rect 18472 30132 18478 30184
rect 19886 30172 19892 30184
rect 18708 30144 19892 30172
rect 17954 30104 17960 30116
rect 17604 30076 17960 30104
rect 17954 30064 17960 30076
rect 18012 30064 18018 30116
rect 18708 30104 18736 30144
rect 19886 30132 19892 30144
rect 19944 30132 19950 30184
rect 20625 30175 20683 30181
rect 20625 30172 20637 30175
rect 20088 30144 20637 30172
rect 18156 30076 18736 30104
rect 11790 30036 11796 30048
rect 9968 30008 11796 30036
rect 11790 29996 11796 30008
rect 11848 29996 11854 30048
rect 12710 29996 12716 30048
rect 12768 30036 12774 30048
rect 13170 30036 13176 30048
rect 12768 30008 13176 30036
rect 12768 29996 12774 30008
rect 13170 29996 13176 30008
rect 13228 30036 13234 30048
rect 13446 30036 13452 30048
rect 13228 30008 13452 30036
rect 13228 29996 13234 30008
rect 13446 29996 13452 30008
rect 13504 29996 13510 30048
rect 16960 30036 16988 30064
rect 18156 30036 18184 30076
rect 16960 30008 18184 30036
rect 18230 29996 18236 30048
rect 18288 30036 18294 30048
rect 20088 30036 20116 30144
rect 20625 30141 20637 30144
rect 20671 30172 20683 30175
rect 21174 30172 21180 30184
rect 20671 30144 21180 30172
rect 20671 30141 20683 30144
rect 20625 30135 20683 30141
rect 21174 30132 21180 30144
rect 21232 30132 21238 30184
rect 18288 30008 20116 30036
rect 23032 30036 23060 30203
rect 23198 30200 23204 30252
rect 23256 30240 23262 30252
rect 23293 30243 23351 30249
rect 23293 30240 23305 30243
rect 23256 30212 23305 30240
rect 23256 30200 23262 30212
rect 23293 30209 23305 30212
rect 23339 30209 23351 30243
rect 23293 30203 23351 30209
rect 23658 30200 23664 30252
rect 23716 30200 23722 30252
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30209 23903 30243
rect 23845 30203 23903 30209
rect 23474 30132 23480 30184
rect 23532 30172 23538 30184
rect 23753 30175 23811 30181
rect 23753 30172 23765 30175
rect 23532 30144 23765 30172
rect 23532 30132 23538 30144
rect 23753 30141 23765 30144
rect 23799 30141 23811 30175
rect 23753 30135 23811 30141
rect 23106 30064 23112 30116
rect 23164 30104 23170 30116
rect 23860 30104 23888 30203
rect 27338 30200 27344 30252
rect 27396 30200 27402 30252
rect 27522 30200 27528 30252
rect 27580 30240 27586 30252
rect 27801 30243 27859 30249
rect 27801 30240 27813 30243
rect 27580 30212 27813 30240
rect 27580 30200 27586 30212
rect 27801 30209 27813 30212
rect 27847 30240 27859 30243
rect 27847 30212 28488 30240
rect 27847 30209 27859 30212
rect 27801 30203 27859 30209
rect 24946 30132 24952 30184
rect 25004 30172 25010 30184
rect 25685 30175 25743 30181
rect 25685 30172 25697 30175
rect 25004 30144 25697 30172
rect 25004 30132 25010 30144
rect 25685 30141 25697 30144
rect 25731 30141 25743 30175
rect 25685 30135 25743 30141
rect 25961 30175 26019 30181
rect 25961 30141 25973 30175
rect 26007 30172 26019 30175
rect 26007 30144 28028 30172
rect 26007 30141 26019 30144
rect 25961 30135 26019 30141
rect 28000 30116 28028 30144
rect 28258 30132 28264 30184
rect 28316 30132 28322 30184
rect 28460 30172 28488 30212
rect 28534 30200 28540 30252
rect 28592 30240 28598 30252
rect 28902 30240 28908 30252
rect 28592 30212 28908 30240
rect 28592 30200 28598 30212
rect 28902 30200 28908 30212
rect 28960 30200 28966 30252
rect 30282 30200 30288 30252
rect 30340 30200 30346 30252
rect 30484 30249 30512 30280
rect 30742 30268 30748 30320
rect 30800 30268 30806 30320
rect 30377 30243 30435 30249
rect 30377 30209 30389 30243
rect 30423 30209 30435 30243
rect 30377 30203 30435 30209
rect 30470 30243 30528 30249
rect 30470 30209 30482 30243
rect 30516 30209 30528 30243
rect 30470 30203 30528 30209
rect 28994 30172 29000 30184
rect 28460 30144 29000 30172
rect 28994 30132 29000 30144
rect 29052 30132 29058 30184
rect 29362 30132 29368 30184
rect 29420 30172 29426 30184
rect 30009 30175 30067 30181
rect 30009 30172 30021 30175
rect 29420 30144 30021 30172
rect 29420 30132 29426 30144
rect 30009 30141 30021 30144
rect 30055 30141 30067 30175
rect 30392 30172 30420 30203
rect 30650 30200 30656 30252
rect 30708 30200 30714 30252
rect 30926 30249 30932 30252
rect 30883 30243 30932 30249
rect 30883 30209 30895 30243
rect 30929 30209 30932 30243
rect 30883 30203 30932 30209
rect 30926 30200 30932 30203
rect 30984 30200 30990 30252
rect 31036 30240 31064 30339
rect 32398 30336 32404 30388
rect 32456 30376 32462 30388
rect 32456 30348 32628 30376
rect 32456 30336 32462 30348
rect 31113 30311 31171 30317
rect 31113 30277 31125 30311
rect 31159 30308 31171 30311
rect 31386 30308 31392 30320
rect 31159 30280 31392 30308
rect 31159 30277 31171 30280
rect 31113 30271 31171 30277
rect 31386 30268 31392 30280
rect 31444 30268 31450 30320
rect 32214 30268 32220 30320
rect 32272 30308 32278 30320
rect 32600 30308 32628 30348
rect 32674 30336 32680 30388
rect 32732 30336 32738 30388
rect 32784 30348 33272 30376
rect 32784 30308 32812 30348
rect 32272 30280 32536 30308
rect 32600 30280 32812 30308
rect 32272 30268 32278 30280
rect 31297 30243 31355 30249
rect 31297 30240 31309 30243
rect 31036 30212 31309 30240
rect 31297 30209 31309 30212
rect 31343 30209 31355 30243
rect 31297 30203 31355 30209
rect 31478 30200 31484 30252
rect 31536 30200 31542 30252
rect 31573 30243 31631 30249
rect 31573 30209 31585 30243
rect 31619 30209 31631 30243
rect 31573 30203 31631 30209
rect 30558 30172 30564 30184
rect 30392 30144 30564 30172
rect 30009 30135 30067 30141
rect 30558 30132 30564 30144
rect 30616 30132 30622 30184
rect 31588 30172 31616 30203
rect 31754 30200 31760 30252
rect 31812 30200 31818 30252
rect 32122 30200 32128 30252
rect 32180 30200 32186 30252
rect 32306 30200 32312 30252
rect 32364 30200 32370 30252
rect 32398 30200 32404 30252
rect 32456 30200 32462 30252
rect 32508 30249 32536 30280
rect 32858 30268 32864 30320
rect 32916 30308 32922 30320
rect 33137 30311 33195 30317
rect 33137 30308 33149 30311
rect 32916 30280 33149 30308
rect 32916 30268 32922 30280
rect 33137 30277 33149 30280
rect 33183 30277 33195 30311
rect 33137 30271 33195 30277
rect 32493 30243 32551 30249
rect 32493 30209 32505 30243
rect 32539 30209 32551 30243
rect 32493 30203 32551 30209
rect 32766 30200 32772 30252
rect 32824 30200 32830 30252
rect 32950 30200 32956 30252
rect 33008 30200 33014 30252
rect 33244 30249 33272 30348
rect 34808 30348 35756 30376
rect 33594 30268 33600 30320
rect 33652 30308 33658 30320
rect 33781 30311 33839 30317
rect 33781 30308 33793 30311
rect 33652 30280 33793 30308
rect 33652 30268 33658 30280
rect 33781 30277 33793 30280
rect 33827 30308 33839 30311
rect 34808 30308 34836 30348
rect 33827 30280 34836 30308
rect 35728 30308 35756 30348
rect 36173 30311 36231 30317
rect 36173 30308 36185 30311
rect 35728 30280 36185 30308
rect 33827 30277 33839 30280
rect 33781 30271 33839 30277
rect 36173 30277 36185 30280
rect 36219 30277 36231 30311
rect 36173 30271 36231 30277
rect 33229 30243 33287 30249
rect 33229 30209 33241 30243
rect 33275 30209 33287 30243
rect 33229 30203 33287 30209
rect 33410 30200 33416 30252
rect 33468 30200 33474 30252
rect 33505 30243 33563 30249
rect 33505 30209 33517 30243
rect 33551 30209 33563 30243
rect 33505 30203 33563 30209
rect 33520 30172 33548 30203
rect 33686 30200 33692 30252
rect 33744 30200 33750 30252
rect 33873 30243 33931 30249
rect 33873 30240 33885 30243
rect 33796 30212 33885 30240
rect 31588 30144 33548 30172
rect 23164 30076 23888 30104
rect 26252 30076 27568 30104
rect 23164 30064 23170 30076
rect 23566 30036 23572 30048
rect 23032 30008 23572 30036
rect 18288 29996 18294 30008
rect 23566 29996 23572 30008
rect 23624 29996 23630 30048
rect 24210 29996 24216 30048
rect 24268 29996 24274 30048
rect 25314 29996 25320 30048
rect 25372 30036 25378 30048
rect 26252 30036 26280 30076
rect 25372 30008 26280 30036
rect 25372 29996 25378 30008
rect 26326 29996 26332 30048
rect 26384 29996 26390 30048
rect 27540 30036 27568 30076
rect 27614 30064 27620 30116
rect 27672 30104 27678 30116
rect 27890 30104 27896 30116
rect 27672 30076 27896 30104
rect 27672 30064 27678 30076
rect 27890 30064 27896 30076
rect 27948 30064 27954 30116
rect 27982 30064 27988 30116
rect 28040 30104 28046 30116
rect 28626 30104 28632 30116
rect 28040 30076 28632 30104
rect 28040 30064 28046 30076
rect 28626 30064 28632 30076
rect 28684 30104 28690 30116
rect 28902 30104 28908 30116
rect 28684 30076 28908 30104
rect 28684 30064 28690 30076
rect 28902 30064 28908 30076
rect 28960 30064 28966 30116
rect 31588 30104 31616 30144
rect 30208 30076 31616 30104
rect 28166 30036 28172 30048
rect 27540 30008 28172 30036
rect 28166 29996 28172 30008
rect 28224 29996 28230 30048
rect 28718 29996 28724 30048
rect 28776 30036 28782 30048
rect 30208 30036 30236 30076
rect 31938 30064 31944 30116
rect 31996 30104 32002 30116
rect 33321 30107 33379 30113
rect 33321 30104 33333 30107
rect 31996 30076 33333 30104
rect 31996 30064 32002 30076
rect 33321 30073 33333 30076
rect 33367 30073 33379 30107
rect 33321 30067 33379 30073
rect 28776 30008 30236 30036
rect 31849 30039 31907 30045
rect 28776 29996 28782 30008
rect 31849 30005 31861 30039
rect 31895 30036 31907 30039
rect 32582 30036 32588 30048
rect 31895 30008 32588 30036
rect 31895 30005 31907 30008
rect 31849 29999 31907 30005
rect 32582 29996 32588 30008
rect 32640 30036 32646 30048
rect 32858 30036 32864 30048
rect 32640 30008 32864 30036
rect 32640 29996 32646 30008
rect 32858 29996 32864 30008
rect 32916 30036 32922 30048
rect 33796 30036 33824 30212
rect 33873 30209 33885 30212
rect 33919 30209 33931 30243
rect 36078 30240 36084 30252
rect 35558 30226 36084 30240
rect 33873 30203 33931 30209
rect 35544 30212 36084 30226
rect 34146 30132 34152 30184
rect 34204 30132 34210 30184
rect 34425 30175 34483 30181
rect 34425 30172 34437 30175
rect 34256 30144 34437 30172
rect 34057 30107 34115 30113
rect 34057 30073 34069 30107
rect 34103 30104 34115 30107
rect 34256 30104 34284 30144
rect 34425 30141 34437 30144
rect 34471 30141 34483 30175
rect 34425 30135 34483 30141
rect 34103 30076 34284 30104
rect 34103 30073 34115 30076
rect 34057 30067 34115 30073
rect 32916 30008 33824 30036
rect 32916 29996 32922 30008
rect 34422 29996 34428 30048
rect 34480 30036 34486 30048
rect 35544 30036 35572 30212
rect 36078 30200 36084 30212
rect 36136 30200 36142 30252
rect 34480 30008 35572 30036
rect 34480 29996 34486 30008
rect 1104 29946 36524 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 36524 29946
rect 1104 29872 36524 29894
rect 6273 29835 6331 29841
rect 6273 29801 6285 29835
rect 6319 29832 6331 29835
rect 6638 29832 6644 29844
rect 6319 29804 6644 29832
rect 6319 29801 6331 29804
rect 6273 29795 6331 29801
rect 6638 29792 6644 29804
rect 6696 29792 6702 29844
rect 9674 29832 9680 29844
rect 6932 29804 9680 29832
rect 3068 29736 6868 29764
rect 3068 29708 3096 29736
rect 3050 29656 3056 29708
rect 3108 29656 3114 29708
rect 4893 29699 4951 29705
rect 4893 29665 4905 29699
rect 4939 29696 4951 29699
rect 6270 29696 6276 29708
rect 4939 29668 6276 29696
rect 4939 29665 4951 29668
rect 4893 29659 4951 29665
rect 6270 29656 6276 29668
rect 6328 29656 6334 29708
rect 6840 29705 6868 29736
rect 6825 29699 6883 29705
rect 6825 29665 6837 29699
rect 6871 29665 6883 29699
rect 6825 29659 6883 29665
rect 6932 29640 6960 29804
rect 9674 29792 9680 29804
rect 9732 29792 9738 29844
rect 9953 29835 10011 29841
rect 9953 29801 9965 29835
rect 9999 29832 10011 29835
rect 10686 29832 10692 29844
rect 9999 29804 10692 29832
rect 9999 29801 10011 29804
rect 9953 29795 10011 29801
rect 10686 29792 10692 29804
rect 10744 29792 10750 29844
rect 16669 29835 16727 29841
rect 16669 29801 16681 29835
rect 16715 29801 16727 29835
rect 16669 29795 16727 29801
rect 8018 29724 8024 29776
rect 8076 29764 8082 29776
rect 9309 29767 9367 29773
rect 8076 29736 9168 29764
rect 8076 29724 8082 29736
rect 8202 29656 8208 29708
rect 8260 29656 8266 29708
rect 2869 29631 2927 29637
rect 2869 29597 2881 29631
rect 2915 29628 2927 29631
rect 4338 29628 4344 29640
rect 2915 29600 4344 29628
rect 2915 29597 2927 29600
rect 2869 29591 2927 29597
rect 4338 29588 4344 29600
rect 4396 29588 4402 29640
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29628 5227 29631
rect 5258 29628 5264 29640
rect 5215 29600 5264 29628
rect 5215 29597 5227 29600
rect 5169 29591 5227 29597
rect 5258 29588 5264 29600
rect 5316 29588 5322 29640
rect 6641 29631 6699 29637
rect 6641 29597 6653 29631
rect 6687 29628 6699 29631
rect 6914 29628 6920 29640
rect 6687 29600 6920 29628
rect 6687 29597 6699 29600
rect 6641 29591 6699 29597
rect 6914 29588 6920 29600
rect 6972 29588 6978 29640
rect 7650 29588 7656 29640
rect 7708 29588 7714 29640
rect 7837 29631 7895 29637
rect 7837 29597 7849 29631
rect 7883 29628 7895 29631
rect 7926 29628 7932 29640
rect 7883 29600 7932 29628
rect 7883 29597 7895 29600
rect 7837 29591 7895 29597
rect 7926 29588 7932 29600
rect 7984 29628 7990 29640
rect 8294 29628 8300 29640
rect 7984 29600 8300 29628
rect 7984 29588 7990 29600
rect 8294 29588 8300 29600
rect 8352 29588 8358 29640
rect 8386 29588 8392 29640
rect 8444 29588 8450 29640
rect 8573 29631 8631 29637
rect 8573 29597 8585 29631
rect 8619 29628 8631 29631
rect 8662 29628 8668 29640
rect 8619 29600 8668 29628
rect 8619 29597 8631 29600
rect 8573 29591 8631 29597
rect 8662 29588 8668 29600
rect 8720 29588 8726 29640
rect 9140 29637 9168 29736
rect 9309 29733 9321 29767
rect 9355 29764 9367 29767
rect 10042 29764 10048 29776
rect 9355 29736 10048 29764
rect 9355 29733 9367 29736
rect 9309 29727 9367 29733
rect 10042 29724 10048 29736
rect 10100 29724 10106 29776
rect 10505 29767 10563 29773
rect 10505 29733 10517 29767
rect 10551 29733 10563 29767
rect 14921 29767 14979 29773
rect 14921 29764 14933 29767
rect 10505 29727 10563 29733
rect 11072 29736 14933 29764
rect 10520 29696 10548 29727
rect 11072 29708 11100 29736
rect 14921 29733 14933 29736
rect 14967 29733 14979 29767
rect 16684 29764 16712 29795
rect 17494 29792 17500 29844
rect 17552 29792 17558 29844
rect 18598 29832 18604 29844
rect 17788 29804 18604 29832
rect 17218 29764 17224 29776
rect 14921 29727 14979 29733
rect 15120 29736 16068 29764
rect 16684 29736 17224 29764
rect 10244 29668 10548 29696
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29597 9183 29631
rect 9125 29591 9183 29597
rect 9306 29588 9312 29640
rect 9364 29588 9370 29640
rect 10137 29631 10195 29637
rect 10137 29597 10149 29631
rect 10183 29622 10195 29631
rect 10244 29622 10272 29668
rect 11054 29656 11060 29708
rect 11112 29656 11118 29708
rect 12434 29656 12440 29708
rect 12492 29696 12498 29708
rect 13354 29696 13360 29708
rect 12492 29668 13360 29696
rect 12492 29656 12498 29668
rect 13354 29656 13360 29668
rect 13412 29656 13418 29708
rect 13446 29656 13452 29708
rect 13504 29696 13510 29708
rect 15120 29696 15148 29736
rect 13504 29668 15148 29696
rect 13504 29656 13510 29668
rect 10183 29597 10272 29622
rect 10137 29594 10272 29597
rect 10137 29591 10195 29594
rect 10318 29588 10324 29640
rect 10376 29588 10382 29640
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29597 10471 29631
rect 10413 29591 10471 29597
rect 4709 29563 4767 29569
rect 4709 29560 4721 29563
rect 2884 29532 4721 29560
rect 2884 29504 2912 29532
rect 4709 29529 4721 29532
rect 4755 29560 4767 29563
rect 5442 29560 5448 29572
rect 4755 29532 5448 29560
rect 4755 29529 4767 29532
rect 4709 29523 4767 29529
rect 5442 29520 5448 29532
rect 5500 29520 5506 29572
rect 6733 29563 6791 29569
rect 6733 29529 6745 29563
rect 6779 29560 6791 29563
rect 7558 29560 7564 29572
rect 6779 29532 7564 29560
rect 6779 29529 6791 29532
rect 6733 29523 6791 29529
rect 7558 29520 7564 29532
rect 7616 29560 7622 29572
rect 8110 29560 8116 29572
rect 7616 29532 8116 29560
rect 7616 29520 7622 29532
rect 8110 29520 8116 29532
rect 8168 29560 8174 29572
rect 10428 29560 10456 29591
rect 10502 29588 10508 29640
rect 10560 29628 10566 29640
rect 10689 29631 10747 29637
rect 10689 29628 10701 29631
rect 10560 29600 10701 29628
rect 10560 29588 10566 29600
rect 10689 29597 10701 29600
rect 10735 29597 10747 29631
rect 10689 29591 10747 29597
rect 10781 29631 10839 29637
rect 10781 29597 10793 29631
rect 10827 29628 10839 29631
rect 10870 29628 10876 29640
rect 10827 29600 10876 29628
rect 10827 29597 10839 29600
rect 10781 29591 10839 29597
rect 10870 29588 10876 29600
rect 10928 29588 10934 29640
rect 12710 29637 12716 29640
rect 12708 29628 12716 29637
rect 12671 29600 12716 29628
rect 12708 29591 12716 29600
rect 12710 29588 12716 29591
rect 12768 29588 12774 29640
rect 13078 29628 13084 29640
rect 13039 29600 13084 29628
rect 13078 29588 13084 29600
rect 13136 29588 13142 29640
rect 13173 29631 13231 29637
rect 13173 29597 13185 29631
rect 13219 29628 13231 29631
rect 13630 29628 13636 29640
rect 13219 29600 13636 29628
rect 13219 29597 13231 29600
rect 13173 29591 13231 29597
rect 13630 29588 13636 29600
rect 13688 29588 13694 29640
rect 15120 29637 15148 29668
rect 15194 29656 15200 29708
rect 15252 29696 15258 29708
rect 15930 29696 15936 29708
rect 15252 29668 15936 29696
rect 15252 29656 15258 29668
rect 15488 29637 15516 29668
rect 15930 29656 15936 29668
rect 15988 29656 15994 29708
rect 16040 29696 16068 29736
rect 17218 29724 17224 29736
rect 17276 29724 17282 29776
rect 17402 29696 17408 29708
rect 16040 29668 17408 29696
rect 17402 29656 17408 29668
rect 17460 29656 17466 29708
rect 15100 29631 15158 29637
rect 15100 29597 15112 29631
rect 15146 29597 15158 29631
rect 15472 29631 15530 29637
rect 15100 29591 15158 29597
rect 15212 29600 15424 29628
rect 10594 29560 10600 29572
rect 8168 29532 10364 29560
rect 10428 29532 10600 29560
rect 8168 29520 8174 29532
rect 1762 29452 1768 29504
rect 1820 29492 1826 29504
rect 2409 29495 2467 29501
rect 2409 29492 2421 29495
rect 1820 29464 2421 29492
rect 1820 29452 1826 29464
rect 2409 29461 2421 29464
rect 2455 29461 2467 29495
rect 2409 29455 2467 29461
rect 2777 29495 2835 29501
rect 2777 29461 2789 29495
rect 2823 29492 2835 29495
rect 2866 29492 2872 29504
rect 2823 29464 2872 29492
rect 2823 29461 2835 29464
rect 2777 29455 2835 29461
rect 2866 29452 2872 29464
rect 2924 29452 2930 29504
rect 4154 29452 4160 29504
rect 4212 29492 4218 29504
rect 4249 29495 4307 29501
rect 4249 29492 4261 29495
rect 4212 29464 4261 29492
rect 4212 29452 4218 29464
rect 4249 29461 4261 29464
rect 4295 29461 4307 29495
rect 4249 29455 4307 29461
rect 4614 29452 4620 29504
rect 4672 29452 4678 29504
rect 5718 29452 5724 29504
rect 5776 29452 5782 29504
rect 7098 29452 7104 29504
rect 7156 29452 7162 29504
rect 7282 29452 7288 29504
rect 7340 29492 7346 29504
rect 10134 29492 10140 29504
rect 7340 29464 10140 29492
rect 7340 29452 7346 29464
rect 10134 29452 10140 29464
rect 10192 29452 10198 29504
rect 10336 29492 10364 29532
rect 10594 29520 10600 29532
rect 10652 29520 10658 29572
rect 10962 29520 10968 29572
rect 11020 29560 11026 29572
rect 11149 29563 11207 29569
rect 11149 29560 11161 29563
rect 11020 29532 11161 29560
rect 11020 29520 11026 29532
rect 11149 29529 11161 29532
rect 11195 29529 11207 29563
rect 11149 29523 11207 29529
rect 11238 29520 11244 29572
rect 11296 29560 11302 29572
rect 12618 29560 12624 29572
rect 11296 29532 12624 29560
rect 11296 29520 11302 29532
rect 12618 29520 12624 29532
rect 12676 29560 12682 29572
rect 12805 29563 12863 29569
rect 12805 29560 12817 29563
rect 12676 29532 12817 29560
rect 12676 29520 12682 29532
rect 12805 29529 12817 29532
rect 12851 29529 12863 29563
rect 12805 29523 12863 29529
rect 12897 29563 12955 29569
rect 12897 29529 12909 29563
rect 12943 29560 12955 29563
rect 13722 29560 13728 29572
rect 12943 29532 13728 29560
rect 12943 29529 12955 29532
rect 12897 29523 12955 29529
rect 13722 29520 13728 29532
rect 13780 29560 13786 29572
rect 15212 29569 15240 29600
rect 15197 29563 15255 29569
rect 13780 29532 14596 29560
rect 13780 29520 13786 29532
rect 11330 29492 11336 29504
rect 10336 29464 11336 29492
rect 11330 29452 11336 29464
rect 11388 29452 11394 29504
rect 12526 29452 12532 29504
rect 12584 29452 12590 29504
rect 13814 29452 13820 29504
rect 13872 29492 13878 29504
rect 14458 29492 14464 29504
rect 13872 29464 14464 29492
rect 13872 29452 13878 29464
rect 14458 29452 14464 29464
rect 14516 29452 14522 29504
rect 14568 29492 14596 29532
rect 15197 29529 15209 29563
rect 15243 29529 15255 29563
rect 15197 29523 15255 29529
rect 15286 29520 15292 29572
rect 15344 29520 15350 29572
rect 15396 29560 15424 29600
rect 15472 29597 15484 29631
rect 15518 29597 15530 29631
rect 15472 29591 15530 29597
rect 15562 29588 15568 29640
rect 15620 29588 15626 29640
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 17494 29628 17500 29640
rect 15804 29600 17500 29628
rect 15804 29588 15810 29600
rect 17494 29588 17500 29600
rect 17552 29588 17558 29640
rect 17678 29588 17684 29640
rect 17736 29588 17742 29640
rect 17788 29637 17816 29804
rect 18598 29792 18604 29804
rect 18656 29832 18662 29844
rect 18656 29804 18736 29832
rect 18656 29792 18662 29804
rect 17954 29724 17960 29776
rect 18012 29764 18018 29776
rect 18708 29764 18736 29804
rect 18782 29792 18788 29844
rect 18840 29792 18846 29844
rect 19886 29792 19892 29844
rect 19944 29832 19950 29844
rect 22097 29835 22155 29841
rect 22097 29832 22109 29835
rect 19944 29804 22109 29832
rect 19944 29792 19950 29804
rect 22097 29801 22109 29804
rect 22143 29832 22155 29835
rect 22143 29804 24900 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 21818 29764 21824 29776
rect 18012 29736 18644 29764
rect 18708 29736 21824 29764
rect 18012 29724 18018 29736
rect 17972 29696 18000 29724
rect 17972 29668 18092 29696
rect 17773 29631 17831 29637
rect 17773 29597 17785 29631
rect 17819 29597 17831 29631
rect 17773 29591 17831 29597
rect 17954 29588 17960 29640
rect 18012 29588 18018 29640
rect 18064 29637 18092 29668
rect 18414 29656 18420 29708
rect 18472 29656 18478 29708
rect 18616 29696 18644 29736
rect 21818 29724 21824 29736
rect 21876 29724 21882 29776
rect 21910 29724 21916 29776
rect 21968 29764 21974 29776
rect 22554 29764 22560 29776
rect 21968 29736 22560 29764
rect 21968 29724 21974 29736
rect 22554 29724 22560 29736
rect 22612 29724 22618 29776
rect 24872 29764 24900 29804
rect 24946 29792 24952 29844
rect 25004 29792 25010 29844
rect 25869 29835 25927 29841
rect 25869 29801 25881 29835
rect 25915 29832 25927 29835
rect 27614 29832 27620 29844
rect 25915 29804 27620 29832
rect 25915 29801 25927 29804
rect 25869 29795 25927 29801
rect 27614 29792 27620 29804
rect 27672 29792 27678 29844
rect 28258 29792 28264 29844
rect 28316 29832 28322 29844
rect 29270 29832 29276 29844
rect 28316 29804 29276 29832
rect 28316 29792 28322 29804
rect 29270 29792 29276 29804
rect 29328 29792 29334 29844
rect 29362 29792 29368 29844
rect 29420 29792 29426 29844
rect 29822 29792 29828 29844
rect 29880 29832 29886 29844
rect 30285 29835 30343 29841
rect 30285 29832 30297 29835
rect 29880 29804 30297 29832
rect 29880 29792 29886 29804
rect 30285 29801 30297 29804
rect 30331 29801 30343 29835
rect 30285 29795 30343 29801
rect 31478 29792 31484 29844
rect 31536 29832 31542 29844
rect 32861 29835 32919 29841
rect 32861 29832 32873 29835
rect 31536 29804 32873 29832
rect 31536 29792 31542 29804
rect 32861 29801 32873 29804
rect 32907 29801 32919 29835
rect 32861 29795 32919 29801
rect 33686 29792 33692 29844
rect 33744 29832 33750 29844
rect 35069 29835 35127 29841
rect 35069 29832 35081 29835
rect 33744 29804 35081 29832
rect 33744 29792 33750 29804
rect 35069 29801 35081 29804
rect 35115 29801 35127 29835
rect 35069 29795 35127 29801
rect 26326 29764 26332 29776
rect 24872 29736 26332 29764
rect 26326 29724 26332 29736
rect 26384 29724 26390 29776
rect 28721 29767 28779 29773
rect 28721 29733 28733 29767
rect 28767 29764 28779 29767
rect 31570 29764 31576 29776
rect 28767 29736 30144 29764
rect 28767 29733 28779 29736
rect 28721 29727 28779 29733
rect 18690 29696 18696 29708
rect 18616 29668 18696 29696
rect 18690 29656 18696 29668
rect 18748 29656 18754 29708
rect 22094 29656 22100 29708
rect 22152 29696 22158 29708
rect 22152 29668 22416 29696
rect 22152 29656 22158 29668
rect 18049 29631 18107 29637
rect 18049 29597 18061 29631
rect 18095 29597 18107 29631
rect 18049 29591 18107 29597
rect 18138 29588 18144 29640
rect 18196 29588 18202 29640
rect 18230 29588 18236 29640
rect 18288 29588 18294 29640
rect 18432 29628 18460 29656
rect 18606 29631 18664 29637
rect 18606 29628 18618 29631
rect 18432 29600 18618 29628
rect 18606 29597 18618 29600
rect 18652 29597 18664 29631
rect 18606 29591 18664 29597
rect 20438 29588 20444 29640
rect 20496 29588 20502 29640
rect 20898 29588 20904 29640
rect 20956 29588 20962 29640
rect 21634 29588 21640 29640
rect 21692 29588 21698 29640
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 21959 29600 22094 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 15654 29560 15660 29572
rect 15396 29532 15660 29560
rect 15654 29520 15660 29532
rect 15712 29520 15718 29572
rect 16206 29520 16212 29572
rect 16264 29560 16270 29572
rect 16637 29563 16695 29569
rect 16637 29560 16649 29563
rect 16264 29532 16649 29560
rect 16264 29520 16270 29532
rect 16637 29529 16649 29532
rect 16683 29529 16695 29563
rect 16637 29523 16695 29529
rect 16850 29520 16856 29572
rect 16908 29520 16914 29572
rect 18417 29563 18475 29569
rect 18417 29529 18429 29563
rect 18463 29529 18475 29563
rect 18417 29523 18475 29529
rect 15304 29492 15332 29520
rect 14568 29464 15332 29492
rect 15378 29452 15384 29504
rect 15436 29492 15442 29504
rect 16485 29495 16543 29501
rect 16485 29492 16497 29495
rect 15436 29464 16497 29492
rect 15436 29452 15442 29464
rect 16485 29461 16497 29464
rect 16531 29461 16543 29495
rect 16868 29492 16896 29520
rect 18046 29492 18052 29504
rect 16868 29464 18052 29492
rect 16485 29455 16543 29461
rect 18046 29452 18052 29464
rect 18104 29452 18110 29504
rect 18322 29452 18328 29504
rect 18380 29492 18386 29504
rect 18432 29492 18460 29523
rect 18506 29520 18512 29572
rect 18564 29520 18570 29572
rect 21177 29563 21235 29569
rect 21177 29560 21189 29563
rect 18616 29532 21189 29560
rect 18616 29492 18644 29532
rect 21177 29529 21189 29532
rect 21223 29529 21235 29563
rect 22066 29560 22094 29600
rect 22186 29588 22192 29640
rect 22244 29588 22250 29640
rect 22278 29588 22284 29640
rect 22336 29588 22342 29640
rect 22388 29628 22416 29668
rect 22462 29656 22468 29708
rect 22520 29656 22526 29708
rect 22738 29656 22744 29708
rect 22796 29656 22802 29708
rect 24210 29656 24216 29708
rect 24268 29696 24274 29708
rect 24854 29696 24860 29708
rect 24268 29668 24440 29696
rect 24268 29656 24274 29668
rect 22388 29600 22784 29628
rect 22462 29560 22468 29572
rect 22066 29532 22468 29560
rect 21177 29523 21235 29529
rect 22462 29520 22468 29532
rect 22520 29520 22526 29572
rect 22756 29560 22784 29600
rect 22830 29588 22836 29640
rect 22888 29588 22894 29640
rect 24302 29628 24308 29640
rect 23584 29600 24308 29628
rect 23584 29560 23612 29600
rect 24302 29588 24308 29600
rect 24360 29588 24366 29640
rect 24412 29637 24440 29668
rect 24688 29668 24860 29696
rect 24688 29637 24716 29668
rect 24854 29656 24860 29668
rect 24912 29656 24918 29708
rect 26878 29696 26884 29708
rect 26160 29668 26884 29696
rect 24397 29631 24455 29637
rect 24397 29597 24409 29631
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 24669 29631 24727 29637
rect 24669 29597 24681 29631
rect 24715 29597 24727 29631
rect 24669 29591 24727 29597
rect 24762 29588 24768 29640
rect 24820 29628 24826 29640
rect 26160 29628 26188 29668
rect 26878 29656 26884 29668
rect 26936 29656 26942 29708
rect 26973 29699 27031 29705
rect 26973 29665 26985 29699
rect 27019 29696 27031 29699
rect 27982 29696 27988 29708
rect 27019 29668 27988 29696
rect 27019 29665 27031 29668
rect 26973 29659 27031 29665
rect 27982 29656 27988 29668
rect 28040 29656 28046 29708
rect 28736 29696 28764 29727
rect 28644 29668 28764 29696
rect 24820 29600 26188 29628
rect 26237 29631 26295 29637
rect 24820 29588 24826 29600
rect 26237 29597 26249 29631
rect 26283 29628 26295 29631
rect 26602 29628 26608 29640
rect 26283 29600 26608 29628
rect 26283 29597 26295 29600
rect 26237 29591 26295 29597
rect 26602 29588 26608 29600
rect 26660 29588 26666 29640
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29597 26755 29631
rect 26697 29591 26755 29597
rect 22756 29532 23612 29560
rect 23658 29520 23664 29572
rect 23716 29560 23722 29572
rect 24581 29563 24639 29569
rect 24581 29560 24593 29563
rect 23716 29532 24593 29560
rect 23716 29520 23722 29532
rect 24581 29529 24593 29532
rect 24627 29529 24639 29563
rect 24581 29523 24639 29529
rect 26050 29520 26056 29572
rect 26108 29520 26114 29572
rect 26329 29563 26387 29569
rect 26329 29529 26341 29563
rect 26375 29529 26387 29563
rect 26329 29523 26387 29529
rect 18380 29464 18644 29492
rect 18380 29452 18386 29464
rect 20622 29452 20628 29504
rect 20680 29492 20686 29504
rect 21729 29495 21787 29501
rect 21729 29492 21741 29495
rect 20680 29464 21741 29492
rect 20680 29452 20686 29464
rect 21729 29461 21741 29464
rect 21775 29461 21787 29495
rect 21729 29455 21787 29461
rect 21818 29452 21824 29504
rect 21876 29492 21882 29504
rect 22094 29492 22100 29504
rect 21876 29464 22100 29492
rect 21876 29452 21882 29464
rect 22094 29452 22100 29464
rect 22152 29452 22158 29504
rect 22186 29452 22192 29504
rect 22244 29492 22250 29504
rect 23934 29492 23940 29504
rect 22244 29464 23940 29492
rect 22244 29452 22250 29464
rect 23934 29452 23940 29464
rect 23992 29492 23998 29504
rect 26344 29492 26372 29523
rect 23992 29464 26372 29492
rect 26712 29492 26740 29591
rect 26878 29520 26884 29572
rect 26936 29520 26942 29572
rect 27246 29520 27252 29572
rect 27304 29520 27310 29572
rect 28534 29560 28540 29572
rect 28474 29532 28540 29560
rect 28534 29520 28540 29532
rect 28592 29520 28598 29572
rect 27154 29492 27160 29504
rect 26712 29464 27160 29492
rect 23992 29452 23998 29464
rect 27154 29452 27160 29464
rect 27212 29492 27218 29504
rect 28644 29492 28672 29668
rect 28994 29656 29000 29708
rect 29052 29696 29058 29708
rect 30006 29696 30012 29708
rect 29052 29668 30012 29696
rect 29052 29656 29058 29668
rect 30006 29656 30012 29668
rect 30064 29656 30070 29708
rect 30116 29705 30144 29736
rect 30944 29736 31576 29764
rect 30101 29699 30159 29705
rect 30101 29665 30113 29699
rect 30147 29665 30159 29699
rect 30101 29659 30159 29665
rect 30466 29656 30472 29708
rect 30524 29656 30530 29708
rect 30944 29705 30972 29736
rect 31570 29724 31576 29736
rect 31628 29764 31634 29776
rect 32306 29764 32312 29776
rect 31628 29736 32312 29764
rect 31628 29724 31634 29736
rect 32306 29724 32312 29736
rect 32364 29724 32370 29776
rect 34517 29767 34575 29773
rect 34517 29733 34529 29767
rect 34563 29764 34575 29767
rect 34698 29764 34704 29776
rect 34563 29736 34704 29764
rect 34563 29733 34575 29736
rect 34517 29727 34575 29733
rect 34698 29724 34704 29736
rect 34756 29724 34762 29776
rect 30929 29699 30987 29705
rect 30929 29665 30941 29699
rect 30975 29665 30987 29699
rect 30929 29659 30987 29665
rect 31662 29656 31668 29708
rect 31720 29656 31726 29708
rect 32416 29668 34376 29696
rect 32416 29640 32444 29668
rect 28718 29588 28724 29640
rect 28776 29628 28782 29640
rect 28813 29631 28871 29637
rect 28813 29628 28825 29631
rect 28776 29600 28825 29628
rect 28776 29588 28782 29600
rect 28813 29597 28825 29600
rect 28859 29597 28871 29631
rect 28813 29591 28871 29597
rect 28902 29588 28908 29640
rect 28960 29628 28966 29640
rect 29181 29631 29239 29637
rect 29181 29628 29193 29631
rect 28960 29600 29193 29628
rect 28960 29588 28966 29600
rect 29181 29597 29193 29600
rect 29227 29597 29239 29631
rect 29181 29591 29239 29597
rect 30190 29588 30196 29640
rect 30248 29628 30254 29640
rect 30561 29631 30619 29637
rect 30561 29628 30573 29631
rect 30248 29600 30573 29628
rect 30248 29588 30254 29600
rect 30561 29597 30573 29600
rect 30607 29597 30619 29631
rect 30561 29591 30619 29597
rect 30742 29588 30748 29640
rect 30800 29588 30806 29640
rect 30834 29588 30840 29640
rect 30892 29628 30898 29640
rect 30892 29600 31156 29628
rect 30892 29588 30898 29600
rect 28994 29520 29000 29572
rect 29052 29520 29058 29572
rect 29089 29563 29147 29569
rect 29089 29529 29101 29563
rect 29135 29560 29147 29563
rect 29270 29560 29276 29572
rect 29135 29532 29276 29560
rect 29135 29529 29147 29532
rect 29089 29523 29147 29529
rect 29270 29520 29276 29532
rect 29328 29520 29334 29572
rect 30760 29560 30788 29588
rect 31021 29563 31079 29569
rect 31021 29560 31033 29563
rect 30760 29532 31033 29560
rect 31021 29529 31033 29532
rect 31067 29529 31079 29563
rect 31128 29560 31156 29600
rect 31202 29588 31208 29640
rect 31260 29588 31266 29640
rect 31386 29588 31392 29640
rect 31444 29588 31450 29640
rect 32122 29588 32128 29640
rect 32180 29588 32186 29640
rect 32398 29588 32404 29640
rect 32456 29588 32462 29640
rect 32493 29631 32551 29637
rect 32493 29597 32505 29631
rect 32539 29628 32551 29631
rect 32674 29628 32680 29640
rect 32539 29600 32680 29628
rect 32539 29597 32551 29600
rect 32493 29591 32551 29597
rect 32674 29588 32680 29600
rect 32732 29628 32738 29640
rect 34348 29637 34376 29668
rect 34532 29668 35020 29696
rect 34532 29640 34560 29668
rect 32769 29631 32827 29637
rect 32769 29628 32781 29631
rect 32732 29600 32781 29628
rect 32732 29588 32738 29600
rect 32769 29597 32781 29600
rect 32815 29597 32827 29631
rect 32769 29591 32827 29597
rect 34333 29631 34391 29637
rect 34333 29597 34345 29631
rect 34379 29597 34391 29631
rect 34333 29591 34391 29597
rect 34514 29588 34520 29640
rect 34572 29588 34578 29640
rect 34606 29588 34612 29640
rect 34664 29628 34670 29640
rect 34992 29637 35020 29668
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34664 29600 34897 29628
rect 34664 29588 34670 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 34977 29631 35035 29637
rect 34977 29597 34989 29631
rect 35023 29597 35035 29631
rect 34977 29591 35035 29597
rect 35618 29588 35624 29640
rect 35676 29588 35682 29640
rect 31297 29563 31355 29569
rect 31297 29560 31309 29563
rect 31128 29532 31309 29560
rect 31021 29523 31079 29529
rect 31297 29529 31309 29532
rect 31343 29529 31355 29563
rect 31297 29523 31355 29529
rect 31527 29563 31585 29569
rect 31527 29529 31539 29563
rect 31573 29560 31585 29563
rect 32582 29560 32588 29572
rect 31573 29532 32588 29560
rect 31573 29529 31585 29532
rect 31527 29523 31585 29529
rect 32582 29520 32588 29532
rect 32640 29520 32646 29572
rect 33778 29520 33784 29572
rect 33836 29560 33842 29572
rect 34793 29563 34851 29569
rect 34793 29560 34805 29563
rect 33836 29532 34805 29560
rect 33836 29520 33842 29532
rect 34793 29529 34805 29532
rect 34839 29529 34851 29563
rect 34793 29523 34851 29529
rect 35805 29563 35863 29569
rect 35805 29529 35817 29563
rect 35851 29529 35863 29563
rect 35805 29523 35863 29529
rect 27212 29464 28672 29492
rect 27212 29452 27218 29464
rect 28810 29452 28816 29504
rect 28868 29492 28874 29504
rect 29549 29495 29607 29501
rect 29549 29492 29561 29495
rect 28868 29464 29561 29492
rect 28868 29452 28874 29464
rect 29549 29461 29561 29464
rect 29595 29461 29607 29495
rect 29549 29455 29607 29461
rect 30282 29452 30288 29504
rect 30340 29492 30346 29504
rect 30653 29495 30711 29501
rect 30653 29492 30665 29495
rect 30340 29464 30665 29492
rect 30340 29452 30346 29464
rect 30653 29461 30665 29464
rect 30699 29461 30711 29495
rect 30653 29455 30711 29461
rect 30742 29452 30748 29504
rect 30800 29492 30806 29504
rect 30837 29495 30895 29501
rect 30837 29492 30849 29495
rect 30800 29464 30849 29492
rect 30800 29452 30806 29464
rect 30837 29461 30849 29464
rect 30883 29461 30895 29495
rect 30837 29455 30895 29461
rect 31662 29452 31668 29504
rect 31720 29492 31726 29504
rect 32122 29492 32128 29504
rect 31720 29464 32128 29492
rect 31720 29452 31726 29464
rect 32122 29452 32128 29464
rect 32180 29452 32186 29504
rect 32214 29452 32220 29504
rect 32272 29452 32278 29504
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 33042 29492 33048 29504
rect 32456 29464 33048 29492
rect 32456 29452 32462 29464
rect 33042 29452 33048 29464
rect 33100 29492 33106 29504
rect 34054 29492 34060 29504
rect 33100 29464 34060 29492
rect 33100 29452 33106 29464
rect 34054 29452 34060 29464
rect 34112 29452 34118 29504
rect 34330 29452 34336 29504
rect 34388 29492 34394 29504
rect 35437 29495 35495 29501
rect 35437 29492 35449 29495
rect 34388 29464 35449 29492
rect 34388 29452 34394 29464
rect 35437 29461 35449 29464
rect 35483 29492 35495 29495
rect 35820 29492 35848 29523
rect 35483 29464 35848 29492
rect 35483 29461 35495 29464
rect 35437 29455 35495 29461
rect 36078 29452 36084 29504
rect 36136 29452 36142 29504
rect 1104 29402 36524 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 36524 29402
rect 1104 29328 36524 29350
rect 4062 29288 4068 29300
rect 3804 29260 4068 29288
rect 1762 29180 1768 29232
rect 1820 29180 1826 29232
rect 3804 29220 3832 29260
rect 4062 29248 4068 29260
rect 4120 29288 4126 29300
rect 4798 29288 4804 29300
rect 4120 29260 4804 29288
rect 4120 29248 4126 29260
rect 2990 29192 3832 29220
rect 3881 29223 3939 29229
rect 3881 29189 3893 29223
rect 3927 29220 3939 29223
rect 4154 29220 4160 29232
rect 3927 29192 4160 29220
rect 3927 29189 3939 29192
rect 3881 29183 3939 29189
rect 4154 29180 4160 29192
rect 4212 29180 4218 29232
rect 4264 29220 4292 29260
rect 4798 29248 4804 29260
rect 4856 29248 4862 29300
rect 5718 29248 5724 29300
rect 5776 29288 5782 29300
rect 5813 29291 5871 29297
rect 5813 29288 5825 29291
rect 5776 29260 5825 29288
rect 5776 29248 5782 29260
rect 5813 29257 5825 29260
rect 5859 29257 5871 29291
rect 5813 29251 5871 29257
rect 6733 29291 6791 29297
rect 6733 29257 6745 29291
rect 6779 29288 6791 29291
rect 7098 29288 7104 29300
rect 6779 29260 7104 29288
rect 6779 29257 6791 29260
rect 6733 29251 6791 29257
rect 7098 29248 7104 29260
rect 7156 29248 7162 29300
rect 7745 29291 7803 29297
rect 7745 29257 7757 29291
rect 7791 29257 7803 29291
rect 7745 29251 7803 29257
rect 7837 29291 7895 29297
rect 7837 29257 7849 29291
rect 7883 29288 7895 29291
rect 8018 29288 8024 29300
rect 7883 29260 8024 29288
rect 7883 29257 7895 29260
rect 7837 29251 7895 29257
rect 5905 29223 5963 29229
rect 4264 29192 4370 29220
rect 5905 29189 5917 29223
rect 5951 29220 5963 29223
rect 6638 29220 6644 29232
rect 5951 29192 6644 29220
rect 5951 29189 5963 29192
rect 5905 29183 5963 29189
rect 6638 29180 6644 29192
rect 6696 29180 6702 29232
rect 6825 29223 6883 29229
rect 6825 29189 6837 29223
rect 6871 29220 6883 29223
rect 6914 29220 6920 29232
rect 6871 29192 6920 29220
rect 6871 29189 6883 29192
rect 6825 29183 6883 29189
rect 6914 29180 6920 29192
rect 6972 29180 6978 29232
rect 7469 29223 7527 29229
rect 7469 29189 7481 29223
rect 7515 29220 7527 29223
rect 7650 29220 7656 29232
rect 7515 29192 7656 29220
rect 7515 29189 7527 29192
rect 7469 29183 7527 29189
rect 7650 29180 7656 29192
rect 7708 29180 7714 29232
rect 7760 29220 7788 29251
rect 8018 29248 8024 29260
rect 8076 29248 8082 29300
rect 8312 29260 8616 29288
rect 8312 29220 8340 29260
rect 7760 29192 8340 29220
rect 5258 29112 5264 29164
rect 5316 29152 5322 29164
rect 7193 29155 7251 29161
rect 5316 29124 7052 29152
rect 5316 29112 5322 29124
rect 1394 29044 1400 29096
rect 1452 29084 1458 29096
rect 1489 29087 1547 29093
rect 1489 29084 1501 29087
rect 1452 29056 1501 29084
rect 1452 29044 1458 29056
rect 1489 29053 1501 29056
rect 1535 29084 1547 29087
rect 3605 29087 3663 29093
rect 3605 29084 3617 29087
rect 1535 29056 3617 29084
rect 1535 29053 1547 29056
rect 1489 29047 1547 29053
rect 3605 29053 3617 29056
rect 3651 29053 3663 29087
rect 4338 29084 4344 29096
rect 3605 29047 3663 29053
rect 3712 29056 4344 29084
rect 3237 29019 3295 29025
rect 3237 28985 3249 29019
rect 3283 29016 3295 29019
rect 3712 29016 3740 29056
rect 4338 29044 4344 29056
rect 4396 29044 4402 29096
rect 6089 29087 6147 29093
rect 6089 29053 6101 29087
rect 6135 29084 6147 29087
rect 6270 29084 6276 29096
rect 6135 29056 6276 29084
rect 6135 29053 6147 29056
rect 6089 29047 6147 29053
rect 6270 29044 6276 29056
rect 6328 29084 6334 29096
rect 6917 29087 6975 29093
rect 6917 29084 6929 29087
rect 6328 29056 6929 29084
rect 6328 29044 6334 29056
rect 6917 29053 6929 29056
rect 6963 29053 6975 29087
rect 7024 29084 7052 29124
rect 7193 29121 7205 29155
rect 7239 29152 7251 29155
rect 7282 29152 7288 29164
rect 7239 29124 7288 29152
rect 7239 29121 7251 29124
rect 7193 29115 7251 29121
rect 7282 29112 7288 29124
rect 7340 29112 7346 29164
rect 7374 29112 7380 29164
rect 7432 29112 7438 29164
rect 7561 29155 7619 29161
rect 7561 29121 7573 29155
rect 7607 29152 7619 29155
rect 7742 29152 7748 29164
rect 7607 29124 7748 29152
rect 7607 29121 7619 29124
rect 7561 29115 7619 29121
rect 7742 29112 7748 29124
rect 7800 29152 7806 29164
rect 7975 29155 8033 29161
rect 7975 29152 7987 29155
rect 7800 29124 7987 29152
rect 7800 29112 7806 29124
rect 7975 29121 7987 29124
rect 8021 29121 8033 29155
rect 7975 29115 8033 29121
rect 8113 29155 8171 29161
rect 8113 29121 8125 29155
rect 8159 29121 8171 29155
rect 8113 29115 8171 29121
rect 8205 29155 8263 29161
rect 8205 29121 8217 29155
rect 8251 29121 8263 29155
rect 8205 29115 8263 29121
rect 8128 29084 8156 29115
rect 7024 29056 8156 29084
rect 6917 29047 6975 29053
rect 3283 28988 3740 29016
rect 3283 28985 3295 28988
rect 3237 28979 3295 28985
rect 5258 28976 5264 29028
rect 5316 29016 5322 29028
rect 5445 29019 5503 29025
rect 5445 29016 5457 29019
rect 5316 28988 5457 29016
rect 5316 28976 5322 28988
rect 5445 28985 5457 28988
rect 5491 28985 5503 29019
rect 5445 28979 5503 28985
rect 7374 28976 7380 29028
rect 7432 29016 7438 29028
rect 8018 29016 8024 29028
rect 7432 28988 8024 29016
rect 7432 28976 7438 28988
rect 8018 28976 8024 28988
rect 8076 29016 8082 29028
rect 8220 29016 8248 29115
rect 8294 29112 8300 29164
rect 8352 29161 8358 29164
rect 8588 29161 8616 29260
rect 8864 29260 8984 29288
rect 8864 29229 8892 29260
rect 8849 29223 8907 29229
rect 8849 29189 8861 29223
rect 8895 29189 8907 29223
rect 8956 29220 8984 29260
rect 9030 29248 9036 29300
rect 9088 29288 9094 29300
rect 9217 29291 9275 29297
rect 9217 29288 9229 29291
rect 9088 29260 9229 29288
rect 9088 29248 9094 29260
rect 9217 29257 9229 29260
rect 9263 29257 9275 29291
rect 9217 29251 9275 29257
rect 9306 29248 9312 29300
rect 9364 29248 9370 29300
rect 10045 29291 10103 29297
rect 10045 29257 10057 29291
rect 10091 29288 10103 29291
rect 10226 29288 10232 29300
rect 10091 29260 10232 29288
rect 10091 29257 10103 29260
rect 10045 29251 10103 29257
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 10318 29248 10324 29300
rect 10376 29288 10382 29300
rect 11606 29288 11612 29300
rect 10376 29260 11612 29288
rect 10376 29248 10382 29260
rect 11606 29248 11612 29260
rect 11664 29248 11670 29300
rect 13078 29288 13084 29300
rect 11900 29260 13084 29288
rect 9398 29220 9404 29232
rect 8956 29192 9404 29220
rect 8849 29183 8907 29189
rect 9398 29180 9404 29192
rect 9456 29220 9462 29232
rect 9677 29223 9735 29229
rect 9677 29220 9689 29223
rect 9456 29192 9689 29220
rect 9456 29180 9462 29192
rect 9677 29189 9689 29192
rect 9723 29189 9735 29223
rect 11238 29220 11244 29232
rect 9677 29183 9735 29189
rect 9876 29192 11244 29220
rect 8352 29155 8391 29161
rect 8379 29121 8391 29155
rect 8352 29115 8391 29121
rect 8456 29155 8514 29161
rect 8456 29121 8468 29155
rect 8502 29152 8514 29155
rect 8562 29155 8620 29161
rect 8502 29121 8524 29152
rect 8456 29115 8524 29121
rect 8562 29121 8574 29155
rect 8608 29121 8620 29155
rect 8562 29115 8620 29121
rect 8721 29155 8779 29161
rect 8721 29121 8733 29155
rect 8767 29121 8779 29155
rect 8721 29115 8779 29121
rect 8352 29112 8358 29115
rect 8496 29084 8524 29115
rect 8076 28988 8248 29016
rect 8404 29056 8524 29084
rect 8404 28994 8432 29056
rect 8736 29016 8764 29115
rect 8938 29112 8944 29164
rect 8996 29112 9002 29164
rect 9122 29161 9128 29164
rect 9079 29155 9128 29161
rect 9079 29121 9091 29155
rect 9125 29121 9128 29155
rect 9079 29115 9128 29121
rect 9122 29112 9128 29115
rect 9180 29152 9186 29164
rect 9493 29155 9551 29161
rect 9493 29152 9505 29155
rect 9180 29124 9505 29152
rect 9180 29112 9186 29124
rect 9493 29121 9505 29124
rect 9539 29121 9551 29155
rect 9493 29115 9551 29121
rect 9582 29112 9588 29164
rect 9640 29112 9646 29164
rect 9876 29161 9904 29192
rect 11238 29180 11244 29192
rect 11296 29180 11302 29232
rect 11330 29180 11336 29232
rect 11388 29220 11394 29232
rect 11900 29229 11928 29260
rect 13078 29248 13084 29260
rect 13136 29248 13142 29300
rect 13814 29288 13820 29300
rect 13188 29260 13820 29288
rect 11885 29223 11943 29229
rect 11388 29192 11652 29220
rect 11388 29180 11394 29192
rect 9861 29155 9919 29161
rect 9861 29121 9873 29155
rect 9907 29121 9919 29155
rect 9861 29115 9919 29121
rect 10042 29112 10048 29164
rect 10100 29152 10106 29164
rect 10229 29155 10287 29161
rect 10229 29152 10241 29155
rect 10100 29124 10241 29152
rect 10100 29112 10106 29124
rect 10229 29121 10241 29124
rect 10275 29121 10287 29155
rect 10229 29115 10287 29121
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29121 10471 29155
rect 10413 29115 10471 29121
rect 10505 29155 10563 29161
rect 10505 29121 10517 29155
rect 10551 29152 10563 29155
rect 10594 29152 10600 29164
rect 10551 29124 10600 29152
rect 10551 29121 10563 29124
rect 10505 29115 10563 29121
rect 10134 29084 10140 29096
rect 9140 29056 10140 29084
rect 9140 29016 9168 29056
rect 10134 29044 10140 29056
rect 10192 29044 10198 29096
rect 8076 28976 8082 28988
rect 8404 28966 8616 28994
rect 8736 28988 9168 29016
rect 9214 28976 9220 29028
rect 9272 29016 9278 29028
rect 10226 29016 10232 29028
rect 9272 28988 10232 29016
rect 9272 28976 9278 28988
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 5350 28908 5356 28960
rect 5408 28908 5414 28960
rect 6086 28908 6092 28960
rect 6144 28948 6150 28960
rect 6365 28951 6423 28957
rect 6365 28948 6377 28951
rect 6144 28920 6377 28948
rect 6144 28908 6150 28920
rect 6365 28917 6377 28920
rect 6411 28917 6423 28951
rect 8588 28948 8616 28966
rect 8662 28948 8668 28960
rect 8588 28920 8668 28948
rect 6365 28911 6423 28917
rect 8662 28908 8668 28920
rect 8720 28908 8726 28960
rect 10318 28908 10324 28960
rect 10376 28948 10382 28960
rect 10428 28948 10456 29115
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 10870 29112 10876 29164
rect 10928 29112 10934 29164
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29152 11207 29155
rect 11514 29152 11520 29164
rect 11195 29124 11520 29152
rect 11195 29121 11207 29124
rect 11149 29115 11207 29121
rect 11514 29112 11520 29124
rect 11572 29112 11578 29164
rect 11624 29161 11652 29192
rect 11885 29189 11897 29223
rect 11931 29189 11943 29223
rect 11885 29183 11943 29189
rect 12641 29223 12699 29229
rect 12641 29189 12653 29223
rect 12687 29220 12699 29223
rect 12986 29220 12992 29232
rect 12687 29192 12992 29220
rect 12687 29189 12699 29192
rect 12641 29183 12699 29189
rect 12986 29180 12992 29192
rect 13044 29180 13050 29232
rect 13188 29220 13216 29260
rect 13814 29248 13820 29260
rect 13872 29248 13878 29300
rect 15562 29288 15568 29300
rect 14016 29260 15568 29288
rect 13265 29223 13323 29229
rect 13265 29220 13277 29223
rect 13188 29192 13277 29220
rect 13265 29189 13277 29192
rect 13311 29189 13323 29223
rect 13265 29183 13323 29189
rect 13357 29223 13415 29229
rect 13357 29189 13369 29223
rect 13403 29220 13415 29223
rect 13722 29220 13728 29232
rect 13403 29192 13728 29220
rect 13403 29189 13415 29192
rect 13357 29183 13415 29189
rect 13722 29180 13728 29192
rect 13780 29180 13786 29232
rect 11609 29155 11667 29161
rect 11609 29121 11621 29155
rect 11655 29121 11667 29155
rect 11609 29115 11667 29121
rect 11793 29155 11851 29161
rect 11793 29121 11805 29155
rect 11839 29121 11851 29155
rect 11793 29115 11851 29121
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29152 12035 29155
rect 12066 29152 12072 29164
rect 12023 29124 12072 29152
rect 12023 29121 12035 29124
rect 11977 29115 12035 29121
rect 10778 29044 10784 29096
rect 10836 29044 10842 29096
rect 10962 29044 10968 29096
rect 11020 29084 11026 29096
rect 11241 29087 11299 29093
rect 11241 29084 11253 29087
rect 11020 29056 11253 29084
rect 11020 29044 11026 29056
rect 11241 29053 11253 29056
rect 11287 29053 11299 29087
rect 11241 29047 11299 29053
rect 10597 29019 10655 29025
rect 10597 28985 10609 29019
rect 10643 29016 10655 29019
rect 10686 29016 10692 29028
rect 10643 28988 10692 29016
rect 10643 28985 10655 28988
rect 10597 28979 10655 28985
rect 10686 28976 10692 28988
rect 10744 28976 10750 29028
rect 11808 29016 11836 29115
rect 12066 29112 12072 29124
rect 12124 29112 12130 29164
rect 12253 29155 12311 29161
rect 12253 29121 12265 29155
rect 12299 29121 12311 29155
rect 12253 29115 12311 29121
rect 11882 29044 11888 29096
rect 11940 29084 11946 29096
rect 12268 29084 12296 29115
rect 12342 29112 12348 29164
rect 12400 29112 12406 29164
rect 12529 29155 12587 29161
rect 12529 29153 12541 29155
rect 12452 29125 12541 29153
rect 11940 29056 12296 29084
rect 12452 29084 12480 29125
rect 12529 29121 12541 29125
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 12757 29155 12815 29161
rect 12757 29121 12769 29155
rect 12803 29152 12815 29155
rect 12894 29152 12900 29164
rect 12803 29124 12900 29152
rect 12803 29121 12815 29124
rect 12757 29115 12815 29121
rect 12894 29112 12900 29124
rect 12952 29112 12958 29164
rect 13170 29161 13176 29164
rect 13168 29152 13176 29161
rect 13131 29124 13176 29152
rect 13168 29115 13176 29124
rect 13170 29112 13176 29115
rect 13228 29112 13234 29164
rect 13446 29112 13452 29164
rect 13504 29112 13510 29164
rect 13540 29155 13598 29161
rect 13540 29121 13552 29155
rect 13586 29121 13598 29155
rect 13540 29115 13598 29121
rect 13464 29084 13492 29112
rect 12452 29056 13492 29084
rect 13556 29084 13584 29115
rect 13630 29112 13636 29164
rect 13688 29152 13694 29164
rect 14016 29152 14044 29260
rect 15562 29248 15568 29260
rect 15620 29288 15626 29300
rect 16669 29291 16727 29297
rect 16669 29288 16681 29291
rect 15620 29260 16681 29288
rect 15620 29248 15626 29260
rect 16669 29257 16681 29260
rect 16715 29257 16727 29291
rect 17586 29288 17592 29300
rect 16669 29251 16727 29257
rect 16960 29260 17592 29288
rect 14369 29223 14427 29229
rect 14369 29189 14381 29223
rect 14415 29220 14427 29223
rect 15194 29220 15200 29232
rect 14415 29192 15200 29220
rect 14415 29189 14427 29192
rect 14369 29183 14427 29189
rect 15194 29180 15200 29192
rect 15252 29180 15258 29232
rect 15378 29220 15384 29232
rect 15304 29192 15384 29220
rect 13688 29124 14044 29152
rect 13688 29112 13694 29124
rect 14090 29112 14096 29164
rect 14148 29112 14154 29164
rect 14277 29155 14335 29161
rect 14277 29121 14289 29155
rect 14323 29121 14335 29155
rect 14277 29115 14335 29121
rect 13814 29084 13820 29096
rect 13556 29056 13820 29084
rect 11940 29044 11946 29056
rect 12452 29016 12480 29056
rect 13814 29044 13820 29056
rect 13872 29084 13878 29096
rect 14182 29084 14188 29096
rect 13872 29056 14188 29084
rect 13872 29044 13878 29056
rect 14182 29044 14188 29056
rect 14240 29044 14246 29096
rect 11808 28988 12480 29016
rect 12897 29019 12955 29025
rect 12897 28985 12909 29019
rect 12943 29016 12955 29019
rect 13446 29016 13452 29028
rect 12943 28988 13452 29016
rect 12943 28985 12955 28988
rect 12897 28979 12955 28985
rect 13446 28976 13452 28988
rect 13504 28976 13510 29028
rect 13538 28976 13544 29028
rect 13596 29016 13602 29028
rect 14292 29016 14320 29115
rect 14458 29112 14464 29164
rect 14516 29112 14522 29164
rect 14734 29112 14740 29164
rect 14792 29112 14798 29164
rect 14826 29112 14832 29164
rect 14884 29152 14890 29164
rect 15304 29161 15332 29192
rect 15378 29180 15384 29192
rect 15436 29180 15442 29232
rect 16209 29223 16267 29229
rect 16209 29189 16221 29223
rect 16255 29220 16267 29223
rect 16850 29220 16856 29232
rect 16255 29192 16856 29220
rect 16255 29189 16267 29192
rect 16209 29183 16267 29189
rect 16850 29180 16856 29192
rect 16908 29180 16914 29232
rect 15013 29155 15071 29161
rect 15013 29152 15025 29155
rect 14884 29124 15025 29152
rect 14884 29112 14890 29124
rect 15013 29121 15025 29124
rect 15059 29121 15071 29155
rect 15013 29115 15071 29121
rect 15289 29155 15347 29161
rect 15289 29121 15301 29155
rect 15335 29121 15347 29155
rect 15289 29115 15347 29121
rect 15470 29112 15476 29164
rect 15528 29112 15534 29164
rect 16114 29112 16120 29164
rect 16172 29112 16178 29164
rect 16298 29112 16304 29164
rect 16356 29112 16362 29164
rect 16465 29155 16523 29161
rect 16465 29121 16477 29155
rect 16511 29152 16523 29155
rect 16511 29121 16528 29152
rect 16465 29115 16528 29121
rect 15105 29087 15163 29093
rect 15105 29053 15117 29087
rect 15151 29084 15163 29087
rect 15378 29084 15384 29096
rect 15151 29056 15384 29084
rect 15151 29053 15163 29056
rect 15105 29047 15163 29053
rect 15378 29044 15384 29056
rect 15436 29044 15442 29096
rect 15654 29044 15660 29096
rect 15712 29084 15718 29096
rect 16500 29084 16528 29115
rect 16574 29112 16580 29164
rect 16632 29152 16638 29164
rect 16960 29152 16988 29260
rect 17586 29248 17592 29260
rect 17644 29248 17650 29300
rect 17954 29248 17960 29300
rect 18012 29288 18018 29300
rect 18325 29291 18383 29297
rect 18325 29288 18337 29291
rect 18012 29260 18337 29288
rect 18012 29248 18018 29260
rect 18325 29257 18337 29260
rect 18371 29257 18383 29291
rect 22094 29288 22100 29300
rect 18325 29251 18383 29257
rect 20088 29260 22100 29288
rect 17405 29223 17463 29229
rect 17405 29189 17417 29223
rect 17451 29220 17463 29223
rect 17494 29220 17500 29232
rect 17451 29192 17500 29220
rect 17451 29189 17463 29192
rect 17405 29183 17463 29189
rect 17494 29180 17500 29192
rect 17552 29180 17558 29232
rect 18506 29220 18512 29232
rect 18064 29192 18512 29220
rect 18064 29152 18092 29192
rect 18506 29180 18512 29192
rect 18564 29180 18570 29232
rect 20088 29220 20116 29260
rect 22094 29248 22100 29260
rect 22152 29288 22158 29300
rect 22554 29288 22560 29300
rect 22152 29260 22232 29288
rect 22152 29248 22158 29260
rect 19996 29192 20116 29220
rect 19996 29164 20024 29192
rect 20438 29180 20444 29232
rect 20496 29220 20502 29232
rect 20809 29223 20867 29229
rect 20809 29220 20821 29223
rect 20496 29192 20821 29220
rect 20496 29180 20502 29192
rect 20809 29189 20821 29192
rect 20855 29189 20867 29223
rect 21818 29220 21824 29232
rect 20809 29183 20867 29189
rect 21284 29192 21824 29220
rect 18325 29155 18383 29161
rect 18325 29152 18337 29155
rect 16632 29124 16988 29152
rect 17328 29124 18092 29152
rect 18156 29124 18337 29152
rect 16632 29112 16638 29124
rect 15712 29056 16528 29084
rect 15712 29044 15718 29056
rect 13596 28988 14320 29016
rect 14645 29019 14703 29025
rect 13596 28976 13602 28988
rect 14645 28985 14657 29019
rect 14691 29016 14703 29019
rect 15197 29019 15255 29025
rect 15197 29016 15209 29019
rect 14691 28988 15209 29016
rect 14691 28985 14703 28988
rect 14645 28979 14703 28985
rect 15197 28985 15209 28988
rect 15243 28985 15255 29019
rect 15197 28979 15255 28985
rect 10376 28920 10456 28948
rect 10376 28908 10382 28920
rect 12158 28908 12164 28960
rect 12216 28908 12222 28960
rect 12802 28908 12808 28960
rect 12860 28948 12866 28960
rect 12989 28951 13047 28957
rect 12989 28948 13001 28951
rect 12860 28920 13001 28948
rect 12860 28908 12866 28920
rect 12989 28917 13001 28920
rect 13035 28917 13047 28951
rect 12989 28911 13047 28917
rect 15930 28908 15936 28960
rect 15988 28908 15994 28960
rect 16500 28948 16528 29056
rect 16853 29087 16911 29093
rect 16853 29053 16865 29087
rect 16899 29053 16911 29087
rect 16853 29047 16911 29053
rect 16945 29087 17003 29093
rect 16945 29053 16957 29087
rect 16991 29084 17003 29087
rect 17126 29084 17132 29096
rect 16991 29056 17132 29084
rect 16991 29053 17003 29056
rect 16945 29047 17003 29053
rect 16868 29016 16896 29047
rect 17126 29044 17132 29056
rect 17184 29044 17190 29096
rect 17328 29028 17356 29124
rect 18156 29028 18184 29124
rect 18325 29121 18337 29124
rect 18371 29121 18383 29155
rect 18325 29115 18383 29121
rect 19426 29112 19432 29164
rect 19484 29152 19490 29164
rect 19797 29155 19855 29161
rect 19797 29152 19809 29155
rect 19484 29124 19809 29152
rect 19484 29112 19490 29124
rect 19797 29121 19809 29124
rect 19843 29121 19855 29155
rect 19797 29115 19855 29121
rect 19886 29112 19892 29164
rect 19944 29112 19950 29164
rect 19978 29112 19984 29164
rect 20036 29112 20042 29164
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29152 20131 29155
rect 20346 29152 20352 29164
rect 20119 29124 20352 29152
rect 20119 29121 20131 29124
rect 20073 29115 20131 29121
rect 20346 29112 20352 29124
rect 20404 29112 20410 29164
rect 20533 29155 20591 29161
rect 20533 29121 20545 29155
rect 20579 29121 20591 29155
rect 20533 29115 20591 29121
rect 18230 29044 18236 29096
rect 18288 29084 18294 29096
rect 18601 29087 18659 29093
rect 18601 29084 18613 29087
rect 18288 29056 18613 29084
rect 18288 29044 18294 29056
rect 18601 29053 18613 29056
rect 18647 29053 18659 29087
rect 20548 29084 20576 29115
rect 20622 29112 20628 29164
rect 20680 29112 20686 29164
rect 20898 29112 20904 29164
rect 20956 29112 20962 29164
rect 21082 29112 21088 29164
rect 21140 29112 21146 29164
rect 21174 29112 21180 29164
rect 21232 29112 21238 29164
rect 21284 29084 21312 29192
rect 21818 29180 21824 29192
rect 21876 29180 21882 29232
rect 22204 29229 22232 29260
rect 22480 29260 22560 29288
rect 22189 29223 22247 29229
rect 22189 29189 22201 29223
rect 22235 29189 22247 29223
rect 22480 29220 22508 29260
rect 22554 29248 22560 29260
rect 22612 29248 22618 29300
rect 23106 29248 23112 29300
rect 23164 29288 23170 29300
rect 23753 29291 23811 29297
rect 23753 29288 23765 29291
rect 23164 29260 23765 29288
rect 23164 29248 23170 29260
rect 23753 29257 23765 29260
rect 23799 29257 23811 29291
rect 23753 29251 23811 29257
rect 22646 29220 22652 29232
rect 22189 29183 22247 29189
rect 22479 29192 22508 29220
rect 22572 29192 22652 29220
rect 21361 29155 21419 29161
rect 21361 29121 21373 29155
rect 21407 29121 21419 29155
rect 21361 29115 21419 29121
rect 21453 29155 21511 29161
rect 21453 29121 21465 29155
rect 21499 29121 21511 29155
rect 21453 29115 21511 29121
rect 20548 29056 21312 29084
rect 18601 29047 18659 29053
rect 17310 29016 17316 29028
rect 16868 28988 17316 29016
rect 17310 28976 17316 28988
rect 17368 28976 17374 29028
rect 17402 28976 17408 29028
rect 17460 29016 17466 29028
rect 17862 29016 17868 29028
rect 17460 28988 17868 29016
rect 17460 28976 17466 28988
rect 17862 28976 17868 28988
rect 17920 28976 17926 29028
rect 18138 28976 18144 29028
rect 18196 28976 18202 29028
rect 18414 28976 18420 29028
rect 18472 28976 18478 29028
rect 20254 28976 20260 29028
rect 20312 28976 20318 29028
rect 20349 29019 20407 29025
rect 20349 28985 20361 29019
rect 20395 29016 20407 29019
rect 21266 29016 21272 29028
rect 20395 28988 21272 29016
rect 20395 28985 20407 28988
rect 20349 28979 20407 28985
rect 21266 28976 21272 28988
rect 21324 28976 21330 29028
rect 19150 28948 19156 28960
rect 16500 28920 19156 28948
rect 19150 28908 19156 28920
rect 19208 28908 19214 28960
rect 20622 28908 20628 28960
rect 20680 28948 20686 28960
rect 20809 28951 20867 28957
rect 20809 28948 20821 28951
rect 20680 28920 20821 28948
rect 20680 28908 20686 28920
rect 20809 28917 20821 28920
rect 20855 28948 20867 28951
rect 21376 28948 21404 29115
rect 21468 29084 21496 29115
rect 22002 29112 22008 29164
rect 22060 29161 22066 29164
rect 22479 29161 22507 29192
rect 22572 29161 22600 29192
rect 22646 29180 22652 29192
rect 22704 29220 22710 29232
rect 23768 29220 23796 29251
rect 24302 29248 24308 29300
rect 24360 29288 24366 29300
rect 25130 29288 25136 29300
rect 24360 29260 25136 29288
rect 24360 29248 24366 29260
rect 25130 29248 25136 29260
rect 25188 29288 25194 29300
rect 25409 29291 25467 29297
rect 25409 29288 25421 29291
rect 25188 29260 25421 29288
rect 25188 29248 25194 29260
rect 25409 29257 25421 29260
rect 25455 29257 25467 29291
rect 25409 29251 25467 29257
rect 26510 29248 26516 29300
rect 26568 29288 26574 29300
rect 26973 29291 27031 29297
rect 26973 29288 26985 29291
rect 26568 29260 26985 29288
rect 26568 29248 26574 29260
rect 26973 29257 26985 29260
rect 27019 29257 27031 29291
rect 26973 29251 27031 29257
rect 27246 29248 27252 29300
rect 27304 29288 27310 29300
rect 27985 29291 28043 29297
rect 27985 29288 27997 29291
rect 27304 29260 27997 29288
rect 27304 29248 27310 29260
rect 27985 29257 27997 29260
rect 28031 29257 28043 29291
rect 27985 29251 28043 29257
rect 28166 29248 28172 29300
rect 28224 29288 28230 29300
rect 28350 29288 28356 29300
rect 28224 29260 28356 29288
rect 28224 29248 28230 29260
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 28442 29248 28448 29300
rect 28500 29288 28506 29300
rect 28902 29288 28908 29300
rect 28500 29260 28908 29288
rect 28500 29248 28506 29260
rect 28902 29248 28908 29260
rect 28960 29248 28966 29300
rect 30190 29288 30196 29300
rect 29472 29260 30196 29288
rect 22704 29192 23612 29220
rect 23768 29192 24072 29220
rect 22704 29180 22710 29192
rect 22060 29155 22109 29161
rect 22060 29121 22063 29155
rect 22097 29152 22109 29155
rect 22281 29155 22339 29161
rect 22097 29124 22153 29152
rect 22097 29121 22109 29124
rect 22060 29115 22109 29121
rect 22281 29121 22293 29155
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 22436 29155 22507 29161
rect 22436 29121 22448 29155
rect 22482 29124 22507 29155
rect 22557 29155 22615 29161
rect 22482 29121 22494 29124
rect 22436 29115 22494 29121
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22557 29115 22615 29121
rect 22833 29155 22891 29161
rect 22833 29121 22845 29155
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 23017 29155 23075 29161
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 23290 29152 23296 29164
rect 23063 29124 23296 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 22060 29112 22066 29115
rect 22186 29084 22192 29096
rect 21468 29056 22192 29084
rect 22186 29044 22192 29056
rect 22244 29044 22250 29096
rect 22296 29084 22324 29115
rect 22649 29087 22707 29093
rect 22649 29084 22661 29087
rect 22296 29056 22661 29084
rect 22572 29028 22600 29056
rect 22649 29053 22661 29056
rect 22695 29053 22707 29087
rect 22848 29084 22876 29115
rect 23290 29112 23296 29124
rect 23348 29112 23354 29164
rect 23385 29155 23443 29161
rect 23385 29121 23397 29155
rect 23431 29121 23443 29155
rect 23385 29115 23443 29121
rect 22848 29056 23060 29084
rect 22649 29047 22707 29053
rect 23032 29028 23060 29056
rect 23106 29044 23112 29096
rect 23164 29084 23170 29096
rect 23400 29084 23428 29115
rect 23164 29056 23428 29084
rect 23477 29087 23535 29093
rect 23164 29044 23170 29056
rect 23477 29053 23489 29087
rect 23523 29053 23535 29087
rect 23584 29084 23612 29192
rect 23934 29112 23940 29164
rect 23992 29112 23998 29164
rect 24044 29161 24072 29192
rect 24118 29180 24124 29232
rect 24176 29220 24182 29232
rect 26050 29220 26056 29232
rect 24176 29192 26056 29220
rect 24176 29180 24182 29192
rect 26050 29180 26056 29192
rect 26108 29180 26114 29232
rect 26789 29223 26847 29229
rect 26789 29189 26801 29223
rect 26835 29220 26847 29223
rect 26835 29192 27660 29220
rect 26835 29189 26847 29192
rect 26789 29183 26847 29189
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29121 24087 29155
rect 24029 29115 24087 29121
rect 24136 29124 24440 29152
rect 24136 29084 24164 29124
rect 23584 29056 24164 29084
rect 24213 29087 24271 29093
rect 23477 29047 23535 29053
rect 24213 29053 24225 29087
rect 24259 29084 24271 29087
rect 24305 29087 24363 29093
rect 24305 29084 24317 29087
rect 24259 29056 24317 29084
rect 24259 29053 24271 29056
rect 24213 29047 24271 29053
rect 24305 29053 24317 29056
rect 24351 29053 24363 29087
rect 24412 29084 24440 29124
rect 24486 29112 24492 29164
rect 24544 29112 24550 29164
rect 24578 29112 24584 29164
rect 24636 29112 24642 29164
rect 24762 29112 24768 29164
rect 24820 29112 24826 29164
rect 24857 29155 24915 29161
rect 24857 29121 24869 29155
rect 24903 29152 24915 29155
rect 25222 29152 25228 29164
rect 24903 29124 25228 29152
rect 24903 29121 24915 29124
rect 24857 29115 24915 29121
rect 25222 29112 25228 29124
rect 25280 29112 25286 29164
rect 25314 29112 25320 29164
rect 25372 29112 25378 29164
rect 26145 29155 26203 29161
rect 26145 29121 26157 29155
rect 26191 29152 26203 29155
rect 26234 29152 26240 29164
rect 26191 29124 26240 29152
rect 26191 29121 26203 29124
rect 26145 29115 26203 29121
rect 26234 29112 26240 29124
rect 26292 29112 26298 29164
rect 26326 29112 26332 29164
rect 26384 29112 26390 29164
rect 27154 29161 27160 29164
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29121 26479 29155
rect 26421 29115 26479 29121
rect 26513 29155 26571 29161
rect 26513 29121 26525 29155
rect 26559 29121 26571 29155
rect 27152 29152 27160 29161
rect 27115 29124 27160 29152
rect 26513 29115 26571 29121
rect 27152 29115 27160 29124
rect 25038 29084 25044 29096
rect 24412 29056 25044 29084
rect 24305 29047 24363 29053
rect 21913 29019 21971 29025
rect 21913 28985 21925 29019
rect 21959 29016 21971 29019
rect 22278 29016 22284 29028
rect 21959 28988 22284 29016
rect 21959 28985 21971 28988
rect 21913 28979 21971 28985
rect 22278 28976 22284 28988
rect 22336 28976 22342 29028
rect 22554 28976 22560 29028
rect 22612 28976 22618 29028
rect 23014 28976 23020 29028
rect 23072 28976 23078 29028
rect 23492 29016 23520 29047
rect 25038 29044 25044 29056
rect 25096 29044 25102 29096
rect 24026 29016 24032 29028
rect 23124 28988 24032 29016
rect 20855 28920 21404 28948
rect 20855 28917 20867 28920
rect 20809 28911 20867 28917
rect 22370 28908 22376 28960
rect 22428 28948 22434 28960
rect 23124 28948 23152 28988
rect 24026 28976 24032 28988
rect 24084 28976 24090 29028
rect 24121 29019 24179 29025
rect 24121 28985 24133 29019
rect 24167 29016 24179 29019
rect 26436 29016 26464 29115
rect 26528 29084 26556 29115
rect 27154 29112 27160 29115
rect 27212 29112 27218 29164
rect 27249 29155 27307 29161
rect 27249 29121 27261 29155
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 26970 29084 26976 29096
rect 26528 29056 26976 29084
rect 26970 29044 26976 29056
rect 27028 29084 27034 29096
rect 27264 29084 27292 29115
rect 27338 29112 27344 29164
rect 27396 29112 27402 29164
rect 27522 29112 27528 29164
rect 27580 29112 27586 29164
rect 27632 29161 27660 29192
rect 27798 29180 27804 29232
rect 27856 29180 27862 29232
rect 29472 29220 29500 29260
rect 30190 29248 30196 29260
rect 30248 29248 30254 29300
rect 30561 29291 30619 29297
rect 30561 29257 30573 29291
rect 30607 29288 30619 29291
rect 30650 29288 30656 29300
rect 30607 29260 30656 29288
rect 30607 29257 30619 29260
rect 30561 29251 30619 29257
rect 30650 29248 30656 29260
rect 30708 29248 30714 29300
rect 30926 29288 30932 29300
rect 30760 29260 30932 29288
rect 28092 29192 29500 29220
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29121 27675 29155
rect 27617 29115 27675 29121
rect 27706 29112 27712 29164
rect 27764 29152 27770 29164
rect 28092 29152 28120 29192
rect 27764 29124 28120 29152
rect 28169 29155 28227 29161
rect 27764 29112 27770 29124
rect 28169 29121 28181 29155
rect 28215 29121 28227 29155
rect 28169 29115 28227 29121
rect 28261 29155 28319 29161
rect 28261 29121 28273 29155
rect 28307 29121 28319 29155
rect 28261 29115 28319 29121
rect 27028 29056 27292 29084
rect 27028 29044 27034 29056
rect 26786 29016 26792 29028
rect 24167 28988 24992 29016
rect 26436 28988 26792 29016
rect 24167 28985 24179 28988
rect 24121 28979 24179 28985
rect 24964 28960 24992 28988
rect 26786 28976 26792 28988
rect 26844 28976 26850 29028
rect 26878 28976 26884 29028
rect 26936 29016 26942 29028
rect 28184 29016 28212 29115
rect 28276 29084 28304 29115
rect 28350 29112 28356 29164
rect 28408 29112 28414 29164
rect 28442 29112 28448 29164
rect 28500 29161 28506 29164
rect 28500 29155 28529 29161
rect 28517 29121 28529 29155
rect 28500 29115 28529 29121
rect 28629 29155 28687 29161
rect 28629 29121 28641 29155
rect 28675 29152 28687 29155
rect 28810 29152 28816 29164
rect 28675 29124 28816 29152
rect 28675 29121 28687 29124
rect 28629 29115 28687 29121
rect 28500 29112 28506 29115
rect 28810 29112 28816 29124
rect 28868 29112 28874 29164
rect 28902 29112 28908 29164
rect 28960 29112 28966 29164
rect 29472 29161 29500 29192
rect 29656 29192 30604 29220
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29121 29515 29155
rect 29457 29115 29515 29121
rect 29546 29112 29552 29164
rect 29604 29152 29610 29164
rect 29656 29161 29684 29192
rect 29641 29155 29699 29161
rect 29641 29152 29653 29155
rect 29604 29124 29653 29152
rect 29604 29112 29610 29124
rect 29641 29121 29653 29124
rect 29687 29121 29699 29155
rect 29641 29115 29699 29121
rect 29730 29112 29736 29164
rect 29788 29152 29794 29164
rect 30009 29155 30067 29161
rect 30009 29152 30021 29155
rect 29788 29124 30021 29152
rect 29788 29112 29794 29124
rect 30009 29121 30021 29124
rect 30055 29121 30067 29155
rect 30009 29115 30067 29121
rect 30101 29155 30159 29161
rect 30101 29121 30113 29155
rect 30147 29121 30159 29155
rect 30101 29115 30159 29121
rect 29178 29084 29184 29096
rect 28276 29056 29184 29084
rect 29178 29044 29184 29056
rect 29236 29044 29242 29096
rect 29362 29044 29368 29096
rect 29420 29084 29426 29096
rect 30116 29084 30144 29115
rect 30190 29112 30196 29164
rect 30248 29152 30254 29164
rect 30285 29155 30343 29161
rect 30285 29152 30297 29155
rect 30248 29124 30297 29152
rect 30248 29112 30254 29124
rect 30285 29121 30297 29124
rect 30331 29121 30343 29155
rect 30285 29115 30343 29121
rect 30374 29112 30380 29164
rect 30432 29112 30438 29164
rect 30469 29155 30527 29161
rect 30469 29121 30481 29155
rect 30515 29121 30527 29155
rect 30469 29115 30527 29121
rect 30484 29084 30512 29115
rect 29420 29056 30512 29084
rect 30576 29084 30604 29192
rect 30760 29161 30788 29260
rect 30926 29248 30932 29260
rect 30984 29248 30990 29300
rect 31662 29288 31668 29300
rect 31496 29260 31668 29288
rect 30837 29223 30895 29229
rect 30837 29189 30849 29223
rect 30883 29220 30895 29223
rect 31202 29220 31208 29232
rect 30883 29192 31208 29220
rect 30883 29189 30895 29192
rect 30837 29183 30895 29189
rect 31202 29180 31208 29192
rect 31260 29180 31266 29232
rect 30745 29155 30803 29161
rect 30745 29121 30757 29155
rect 30791 29121 30803 29155
rect 30745 29115 30803 29121
rect 30929 29155 30987 29161
rect 30929 29121 30941 29155
rect 30975 29152 30987 29155
rect 31018 29152 31024 29164
rect 30975 29124 31024 29152
rect 30975 29121 30987 29124
rect 30929 29115 30987 29121
rect 31018 29112 31024 29124
rect 31076 29112 31082 29164
rect 31496 29152 31524 29260
rect 31662 29248 31668 29260
rect 31720 29248 31726 29300
rect 31849 29291 31907 29297
rect 31849 29257 31861 29291
rect 31895 29257 31907 29291
rect 31849 29251 31907 29257
rect 31570 29180 31576 29232
rect 31628 29220 31634 29232
rect 31864 29220 31892 29251
rect 32030 29248 32036 29300
rect 32088 29288 32094 29300
rect 32306 29288 32312 29300
rect 32088 29260 32312 29288
rect 32088 29248 32094 29260
rect 32306 29248 32312 29260
rect 32364 29248 32370 29300
rect 32766 29248 32772 29300
rect 32824 29248 32830 29300
rect 33042 29288 33048 29300
rect 32968 29260 33048 29288
rect 31628 29192 31892 29220
rect 31628 29180 31634 29192
rect 32122 29180 32128 29232
rect 32180 29220 32186 29232
rect 32493 29223 32551 29229
rect 32493 29220 32505 29223
rect 32180 29192 32505 29220
rect 32180 29180 32186 29192
rect 32493 29189 32505 29192
rect 32539 29220 32551 29223
rect 32861 29223 32919 29229
rect 32861 29220 32873 29223
rect 32539 29192 32873 29220
rect 32539 29189 32551 29192
rect 32493 29183 32551 29189
rect 32861 29189 32873 29192
rect 32907 29189 32919 29223
rect 32861 29183 32919 29189
rect 31843 29158 31901 29161
rect 31938 29158 31944 29164
rect 31843 29155 31944 29158
rect 31496 29124 31708 29152
rect 31386 29084 31392 29096
rect 30576 29056 31392 29084
rect 29420 29044 29426 29056
rect 31386 29044 31392 29056
rect 31444 29044 31450 29096
rect 31570 29044 31576 29096
rect 31628 29044 31634 29096
rect 28534 29016 28540 29028
rect 26936 28988 28120 29016
rect 28184 28988 28540 29016
rect 26936 28976 26942 28988
rect 22428 28920 23152 28948
rect 22428 28908 22434 28920
rect 23474 28908 23480 28960
rect 23532 28948 23538 28960
rect 24578 28948 24584 28960
rect 23532 28920 24584 28948
rect 23532 28908 23538 28920
rect 24578 28908 24584 28920
rect 24636 28908 24642 28960
rect 24946 28908 24952 28960
rect 25004 28908 25010 28960
rect 26234 28908 26240 28960
rect 26292 28948 26298 28960
rect 27798 28948 27804 28960
rect 26292 28920 27804 28948
rect 26292 28908 26298 28920
rect 27798 28908 27804 28920
rect 27856 28908 27862 28960
rect 28092 28948 28120 28988
rect 28534 28976 28540 28988
rect 28592 28976 28598 29028
rect 29454 29016 29460 29028
rect 28644 28988 29460 29016
rect 28644 28948 28672 28988
rect 29454 28976 29460 28988
rect 29512 28976 29518 29028
rect 31680 29016 31708 29124
rect 31843 29121 31855 29155
rect 31889 29130 31944 29155
rect 31889 29121 31901 29130
rect 31843 29115 31901 29121
rect 31938 29112 31944 29130
rect 31996 29112 32002 29164
rect 32283 29155 32341 29161
rect 32283 29121 32295 29155
rect 32329 29152 32341 29155
rect 32329 29121 32352 29152
rect 32283 29115 32352 29121
rect 32125 29087 32183 29093
rect 32125 29053 32137 29087
rect 32171 29084 32183 29087
rect 32324 29084 32352 29115
rect 32398 29112 32404 29164
rect 32456 29112 32462 29164
rect 32582 29112 32588 29164
rect 32640 29112 32646 29164
rect 32968 29161 32996 29260
rect 33042 29248 33048 29260
rect 33100 29248 33106 29300
rect 34057 29291 34115 29297
rect 34057 29257 34069 29291
rect 34103 29288 34115 29291
rect 34514 29288 34520 29300
rect 34103 29260 34520 29288
rect 34103 29257 34115 29260
rect 34057 29251 34115 29257
rect 34514 29248 34520 29260
rect 34572 29248 34578 29300
rect 35342 29288 35348 29300
rect 34808 29260 35348 29288
rect 33410 29180 33416 29232
rect 33468 29180 33474 29232
rect 34808 29220 34836 29260
rect 35342 29248 35348 29260
rect 35400 29248 35406 29300
rect 36078 29220 36084 29232
rect 33704 29192 34836 29220
rect 35650 29192 36084 29220
rect 32953 29155 33011 29161
rect 32953 29121 32965 29155
rect 32999 29121 33011 29155
rect 32953 29115 33011 29121
rect 33137 29155 33195 29161
rect 33137 29121 33149 29155
rect 33183 29152 33195 29155
rect 33704 29152 33732 29192
rect 36078 29180 36084 29192
rect 36136 29180 36142 29232
rect 33183 29124 33732 29152
rect 33183 29121 33195 29124
rect 33137 29115 33195 29121
rect 32766 29084 32772 29096
rect 32171 29056 32260 29084
rect 32324 29056 32772 29084
rect 32171 29053 32183 29056
rect 32125 29047 32183 29053
rect 31757 29019 31815 29025
rect 31757 29016 31769 29019
rect 31680 28988 31769 29016
rect 31757 28985 31769 28988
rect 31803 28985 31815 29019
rect 31757 28979 31815 28985
rect 31938 28976 31944 29028
rect 31996 28994 32002 29028
rect 32232 29016 32260 29056
rect 32766 29044 32772 29056
rect 32824 29044 32830 29096
rect 32858 29044 32864 29096
rect 32916 29084 32922 29096
rect 33152 29084 33180 29115
rect 33778 29112 33784 29164
rect 33836 29112 33842 29164
rect 33873 29155 33931 29161
rect 33873 29121 33885 29155
rect 33919 29121 33931 29155
rect 33873 29115 33931 29121
rect 32916 29056 33180 29084
rect 32916 29044 32922 29056
rect 33318 29044 33324 29096
rect 33376 29084 33382 29096
rect 33888 29084 33916 29115
rect 33376 29056 33916 29084
rect 33376 29044 33382 29056
rect 33226 29016 33232 29028
rect 31996 28976 32076 28994
rect 32232 28988 33232 29016
rect 33226 28976 33232 28988
rect 33284 28976 33290 29028
rect 31956 28966 32076 28976
rect 28092 28920 28672 28948
rect 28810 28908 28816 28960
rect 28868 28948 28874 28960
rect 29181 28951 29239 28957
rect 29181 28948 29193 28951
rect 28868 28920 29193 28948
rect 28868 28908 28874 28920
rect 29181 28917 29193 28920
rect 29227 28948 29239 28951
rect 29270 28948 29276 28960
rect 29227 28920 29276 28948
rect 29227 28917 29239 28920
rect 29181 28911 29239 28917
rect 29270 28908 29276 28920
rect 29328 28948 29334 28960
rect 29546 28948 29552 28960
rect 29328 28920 29552 28948
rect 29328 28908 29334 28920
rect 29546 28908 29552 28920
rect 29604 28908 29610 28960
rect 29825 28951 29883 28957
rect 29825 28917 29837 28951
rect 29871 28948 29883 28951
rect 30466 28948 30472 28960
rect 29871 28920 30472 28948
rect 29871 28917 29883 28920
rect 29825 28911 29883 28917
rect 30466 28908 30472 28920
rect 30524 28908 30530 28960
rect 32048 28948 32076 28966
rect 32306 28948 32312 28960
rect 32048 28920 32312 28948
rect 32306 28908 32312 28920
rect 32364 28908 32370 28960
rect 33042 28908 33048 28960
rect 33100 28948 33106 28960
rect 33505 28951 33563 28957
rect 33505 28948 33517 28951
rect 33100 28920 33517 28948
rect 33100 28908 33106 28920
rect 33505 28917 33517 28920
rect 33551 28917 33563 28951
rect 33888 28948 33916 29056
rect 34146 29044 34152 29096
rect 34204 29044 34210 29096
rect 34422 29044 34428 29096
rect 34480 29044 34486 29096
rect 36170 29044 36176 29096
rect 36228 29044 36234 29096
rect 34790 28948 34796 28960
rect 33888 28920 34796 28948
rect 33505 28911 33563 28917
rect 34790 28908 34796 28920
rect 34848 28908 34854 28960
rect 1104 28858 36524 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 36524 28858
rect 1104 28784 36524 28806
rect 3789 28747 3847 28753
rect 3789 28713 3801 28747
rect 3835 28744 3847 28747
rect 4246 28744 4252 28756
rect 3835 28716 4252 28744
rect 3835 28713 3847 28716
rect 3789 28707 3847 28713
rect 4246 28704 4252 28716
rect 4304 28744 4310 28756
rect 5166 28744 5172 28756
rect 4304 28716 5172 28744
rect 4304 28704 4310 28716
rect 5166 28704 5172 28716
rect 5224 28704 5230 28756
rect 5442 28704 5448 28756
rect 5500 28744 5506 28756
rect 7561 28747 7619 28753
rect 5500 28716 7144 28744
rect 5500 28704 5506 28716
rect 7116 28676 7144 28716
rect 7561 28713 7573 28747
rect 7607 28744 7619 28747
rect 7650 28744 7656 28756
rect 7607 28716 7656 28744
rect 7607 28713 7619 28716
rect 7561 28707 7619 28713
rect 7650 28704 7656 28716
rect 7708 28704 7714 28756
rect 7742 28704 7748 28756
rect 7800 28744 7806 28756
rect 8110 28744 8116 28756
rect 7800 28716 8116 28744
rect 7800 28704 7806 28716
rect 8110 28704 8116 28716
rect 8168 28704 8174 28756
rect 8297 28747 8355 28753
rect 8297 28713 8309 28747
rect 8343 28744 8355 28747
rect 8386 28744 8392 28756
rect 8343 28716 8392 28744
rect 8343 28713 8355 28716
rect 8297 28707 8355 28713
rect 8386 28704 8392 28716
rect 8444 28704 8450 28756
rect 15930 28744 15936 28756
rect 10060 28716 15936 28744
rect 9401 28679 9459 28685
rect 9401 28676 9413 28679
rect 7116 28648 9413 28676
rect 9401 28645 9413 28648
rect 9447 28645 9459 28679
rect 9401 28639 9459 28645
rect 4522 28568 4528 28620
rect 4580 28608 4586 28620
rect 4706 28608 4712 28620
rect 4580 28580 4712 28608
rect 4580 28568 4586 28580
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 5258 28568 5264 28620
rect 5316 28568 5322 28620
rect 5537 28611 5595 28617
rect 5537 28577 5549 28611
rect 5583 28608 5595 28611
rect 5810 28608 5816 28620
rect 5583 28580 5816 28608
rect 5583 28577 5595 28580
rect 5537 28571 5595 28577
rect 5810 28568 5816 28580
rect 5868 28568 5874 28620
rect 6086 28568 6092 28620
rect 6144 28568 6150 28620
rect 6638 28568 6644 28620
rect 6696 28608 6702 28620
rect 10060 28608 10088 28716
rect 15930 28704 15936 28716
rect 15988 28704 15994 28756
rect 16574 28704 16580 28756
rect 16632 28744 16638 28756
rect 16761 28747 16819 28753
rect 16761 28744 16773 28747
rect 16632 28716 16773 28744
rect 16632 28704 16638 28716
rect 16761 28713 16773 28716
rect 16807 28744 16819 28747
rect 17218 28744 17224 28756
rect 16807 28716 17224 28744
rect 16807 28713 16819 28716
rect 16761 28707 16819 28713
rect 17218 28704 17224 28716
rect 17276 28704 17282 28756
rect 18233 28747 18291 28753
rect 18233 28713 18245 28747
rect 18279 28744 18291 28747
rect 18414 28744 18420 28756
rect 18279 28716 18420 28744
rect 18279 28713 18291 28716
rect 18233 28707 18291 28713
rect 18414 28704 18420 28716
rect 18472 28704 18478 28756
rect 20438 28704 20444 28756
rect 20496 28704 20502 28756
rect 21726 28744 21732 28756
rect 20548 28716 21732 28744
rect 10226 28636 10232 28688
rect 10284 28636 10290 28688
rect 10965 28679 11023 28685
rect 10965 28676 10977 28679
rect 10704 28648 10977 28676
rect 10704 28617 10732 28648
rect 10965 28645 10977 28648
rect 11011 28645 11023 28679
rect 10965 28639 11023 28645
rect 11238 28636 11244 28688
rect 11296 28676 11302 28688
rect 12250 28676 12256 28688
rect 11296 28648 12256 28676
rect 11296 28636 11302 28648
rect 12250 28636 12256 28648
rect 12308 28636 12314 28688
rect 12526 28636 12532 28688
rect 12584 28636 12590 28688
rect 14550 28636 14556 28688
rect 14608 28676 14614 28688
rect 20548 28676 20576 28716
rect 21726 28704 21732 28716
rect 21784 28704 21790 28756
rect 24949 28747 25007 28753
rect 24949 28713 24961 28747
rect 24995 28744 25007 28747
rect 25038 28744 25044 28756
rect 24995 28716 25044 28744
rect 24995 28713 25007 28716
rect 24949 28707 25007 28713
rect 25038 28704 25044 28716
rect 25096 28704 25102 28756
rect 26234 28744 26240 28756
rect 25240 28716 26240 28744
rect 20901 28679 20959 28685
rect 20901 28676 20913 28679
rect 14608 28648 17264 28676
rect 14608 28636 14614 28648
rect 6696 28580 7420 28608
rect 6696 28568 6702 28580
rect 1394 28500 1400 28552
rect 1452 28500 1458 28552
rect 1670 28432 1676 28484
rect 1728 28432 1734 28484
rect 2898 28444 4016 28472
rect 3142 28364 3148 28416
rect 3200 28364 3206 28416
rect 3988 28404 4016 28444
rect 4798 28432 4804 28484
rect 4856 28472 4862 28484
rect 7392 28472 7420 28580
rect 7668 28580 10088 28608
rect 10689 28611 10747 28617
rect 7668 28549 7696 28580
rect 10689 28577 10701 28611
rect 10735 28577 10747 28611
rect 10689 28571 10747 28577
rect 10778 28568 10784 28620
rect 10836 28568 10842 28620
rect 11146 28568 11152 28620
rect 11204 28568 11210 28620
rect 11514 28568 11520 28620
rect 11572 28608 11578 28620
rect 11609 28611 11667 28617
rect 11609 28608 11621 28611
rect 11572 28580 11621 28608
rect 11572 28568 11578 28580
rect 11609 28577 11621 28580
rect 11655 28577 11667 28611
rect 11609 28571 11667 28577
rect 12158 28568 12164 28620
rect 12216 28568 12222 28620
rect 13262 28608 13268 28620
rect 13096 28580 13268 28608
rect 7653 28543 7711 28549
rect 7653 28509 7665 28543
rect 7699 28509 7711 28543
rect 7653 28503 7711 28509
rect 7746 28543 7804 28549
rect 7746 28509 7758 28543
rect 7792 28509 7804 28543
rect 8021 28543 8079 28549
rect 8021 28540 8033 28543
rect 7746 28503 7804 28509
rect 7852 28512 8033 28540
rect 7760 28472 7788 28503
rect 4856 28444 6578 28472
rect 7392 28444 7788 28472
rect 4856 28432 4862 28444
rect 4908 28404 4936 28444
rect 3988 28376 4936 28404
rect 5442 28364 5448 28416
rect 5500 28404 5506 28416
rect 7852 28404 7880 28512
rect 8021 28509 8033 28512
rect 8067 28509 8079 28543
rect 8021 28503 8079 28509
rect 8110 28500 8116 28552
rect 8168 28549 8174 28552
rect 8168 28540 8176 28549
rect 8168 28512 8213 28540
rect 8168 28503 8176 28512
rect 8168 28500 8174 28503
rect 8294 28500 8300 28552
rect 8352 28500 8358 28552
rect 9582 28500 9588 28552
rect 9640 28540 9646 28552
rect 10796 28540 10824 28568
rect 11241 28543 11299 28549
rect 11241 28540 11253 28543
rect 9640 28512 11253 28540
rect 9640 28500 9646 28512
rect 11241 28509 11253 28512
rect 11287 28509 11299 28543
rect 11241 28503 11299 28509
rect 11882 28500 11888 28552
rect 11940 28540 11946 28552
rect 12069 28543 12127 28549
rect 12069 28540 12081 28543
rect 11940 28512 12081 28540
rect 11940 28500 11946 28512
rect 12069 28509 12081 28512
rect 12115 28509 12127 28543
rect 12069 28503 12127 28509
rect 12250 28500 12256 28552
rect 12308 28500 12314 28552
rect 12342 28500 12348 28552
rect 12400 28500 12406 28552
rect 12710 28549 12716 28552
rect 12708 28540 12716 28549
rect 12671 28512 12716 28540
rect 12708 28503 12716 28512
rect 12710 28500 12716 28503
rect 12768 28500 12774 28552
rect 13096 28549 13124 28580
rect 13262 28568 13268 28580
rect 13320 28568 13326 28620
rect 14182 28568 14188 28620
rect 14240 28608 14246 28620
rect 16850 28608 16856 28620
rect 14240 28580 16856 28608
rect 14240 28568 14246 28580
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 16942 28568 16948 28620
rect 17000 28608 17006 28620
rect 17000 28580 17080 28608
rect 17000 28568 17006 28580
rect 13080 28543 13138 28549
rect 13080 28509 13092 28543
rect 13126 28509 13138 28543
rect 13080 28503 13138 28509
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28540 13231 28543
rect 13630 28540 13636 28552
rect 13219 28512 13636 28540
rect 13219 28509 13231 28512
rect 13173 28503 13231 28509
rect 13630 28500 13636 28512
rect 13688 28500 13694 28552
rect 7929 28475 7987 28481
rect 7929 28441 7941 28475
rect 7975 28472 7987 28475
rect 8312 28472 8340 28500
rect 9030 28472 9036 28484
rect 7975 28444 9036 28472
rect 7975 28441 7987 28444
rect 7929 28435 7987 28441
rect 9030 28432 9036 28444
rect 9088 28432 9094 28484
rect 9674 28432 9680 28484
rect 9732 28432 9738 28484
rect 9953 28475 10011 28481
rect 9953 28441 9965 28475
rect 9999 28472 10011 28475
rect 10226 28472 10232 28484
rect 9999 28444 10232 28472
rect 9999 28441 10011 28444
rect 9953 28435 10011 28441
rect 10226 28432 10232 28444
rect 10284 28472 10290 28484
rect 10781 28475 10839 28481
rect 10781 28472 10793 28475
rect 10284 28444 10793 28472
rect 10284 28432 10290 28444
rect 10781 28441 10793 28444
rect 10827 28441 10839 28475
rect 10781 28435 10839 28441
rect 11514 28432 11520 28484
rect 11572 28432 11578 28484
rect 11606 28432 11612 28484
rect 11664 28472 11670 28484
rect 12805 28475 12863 28481
rect 12805 28472 12817 28475
rect 11664 28444 12817 28472
rect 11664 28432 11670 28444
rect 12805 28441 12817 28444
rect 12851 28441 12863 28475
rect 12805 28435 12863 28441
rect 12897 28475 12955 28481
rect 12897 28441 12909 28475
rect 12943 28472 12955 28475
rect 13722 28472 13728 28484
rect 12943 28444 13728 28472
rect 12943 28441 12955 28444
rect 12897 28435 12955 28441
rect 5500 28376 7880 28404
rect 5500 28364 5506 28376
rect 9766 28364 9772 28416
rect 9824 28404 9830 28416
rect 9861 28407 9919 28413
rect 9861 28404 9873 28407
rect 9824 28376 9873 28404
rect 9824 28364 9830 28376
rect 9861 28373 9873 28376
rect 9907 28373 9919 28407
rect 9861 28367 9919 28373
rect 10318 28364 10324 28416
rect 10376 28404 10382 28416
rect 10689 28407 10747 28413
rect 10689 28404 10701 28407
rect 10376 28376 10701 28404
rect 10376 28364 10382 28376
rect 10689 28373 10701 28376
rect 10735 28404 10747 28407
rect 11422 28404 11428 28416
rect 10735 28376 11428 28404
rect 10735 28373 10747 28376
rect 10689 28367 10747 28373
rect 11422 28364 11428 28376
rect 11480 28404 11486 28416
rect 11885 28407 11943 28413
rect 11885 28404 11897 28407
rect 11480 28376 11897 28404
rect 11480 28364 11486 28376
rect 11885 28373 11897 28376
rect 11931 28373 11943 28407
rect 11885 28367 11943 28373
rect 12158 28364 12164 28416
rect 12216 28404 12222 28416
rect 12912 28404 12940 28435
rect 13722 28432 13728 28444
rect 13780 28432 13786 28484
rect 16206 28432 16212 28484
rect 16264 28472 16270 28484
rect 16729 28475 16787 28481
rect 16729 28472 16741 28475
rect 16264 28444 16741 28472
rect 16264 28432 16270 28444
rect 16729 28441 16741 28444
rect 16775 28472 16787 28475
rect 16775 28441 16804 28472
rect 16729 28435 16804 28441
rect 12216 28376 12940 28404
rect 12216 28364 12222 28376
rect 15286 28364 15292 28416
rect 15344 28404 15350 28416
rect 16577 28407 16635 28413
rect 16577 28404 16589 28407
rect 15344 28376 16589 28404
rect 15344 28364 15350 28376
rect 16577 28373 16589 28376
rect 16623 28373 16635 28407
rect 16776 28404 16804 28435
rect 16942 28432 16948 28484
rect 17000 28432 17006 28484
rect 17052 28481 17080 28580
rect 17236 28552 17264 28648
rect 19306 28648 20576 28676
rect 20640 28648 20913 28676
rect 19306 28608 19334 28648
rect 20640 28608 20668 28648
rect 20901 28645 20913 28648
rect 20947 28645 20959 28679
rect 25240 28676 25268 28716
rect 26234 28704 26240 28716
rect 26292 28704 26298 28756
rect 26326 28704 26332 28756
rect 26384 28744 26390 28756
rect 27341 28747 27399 28753
rect 27341 28744 27353 28747
rect 26384 28716 27353 28744
rect 26384 28704 26390 28716
rect 27341 28713 27353 28716
rect 27387 28713 27399 28747
rect 27341 28707 27399 28713
rect 27522 28704 27528 28756
rect 27580 28744 27586 28756
rect 28169 28747 28227 28753
rect 28169 28744 28181 28747
rect 27580 28716 28181 28744
rect 27580 28704 27586 28716
rect 28169 28713 28181 28716
rect 28215 28713 28227 28747
rect 28169 28707 28227 28713
rect 28810 28704 28816 28756
rect 28868 28704 28874 28756
rect 28902 28704 28908 28756
rect 28960 28744 28966 28756
rect 33226 28744 33232 28756
rect 28960 28716 33232 28744
rect 28960 28704 28966 28716
rect 33226 28704 33232 28716
rect 33284 28704 33290 28756
rect 33962 28704 33968 28756
rect 34020 28744 34026 28756
rect 34793 28747 34851 28753
rect 34793 28744 34805 28747
rect 34020 28716 34805 28744
rect 34020 28704 34026 28716
rect 34793 28713 34805 28716
rect 34839 28713 34851 28747
rect 34793 28707 34851 28713
rect 20901 28639 20959 28645
rect 21928 28648 25268 28676
rect 25317 28679 25375 28685
rect 17972 28580 19334 28608
rect 19536 28580 20668 28608
rect 20732 28580 21036 28608
rect 17218 28500 17224 28552
rect 17276 28540 17282 28552
rect 17681 28543 17739 28549
rect 17681 28540 17693 28543
rect 17276 28512 17693 28540
rect 17276 28500 17282 28512
rect 17681 28509 17693 28512
rect 17727 28509 17739 28543
rect 17681 28503 17739 28509
rect 17770 28500 17776 28552
rect 17828 28540 17834 28552
rect 17972 28549 18000 28580
rect 17957 28543 18015 28549
rect 17957 28540 17969 28543
rect 17828 28512 17969 28540
rect 17828 28500 17834 28512
rect 17957 28509 17969 28512
rect 18003 28509 18015 28543
rect 17957 28503 18015 28509
rect 18046 28500 18052 28552
rect 18104 28500 18110 28552
rect 19536 28549 19564 28580
rect 19521 28543 19579 28549
rect 19521 28509 19533 28543
rect 19567 28509 19579 28543
rect 19521 28503 19579 28509
rect 19702 28500 19708 28552
rect 19760 28500 19766 28552
rect 20625 28543 20683 28549
rect 20625 28540 20637 28543
rect 19812 28512 20637 28540
rect 17037 28475 17095 28481
rect 17037 28441 17049 28475
rect 17083 28441 17095 28475
rect 17037 28435 17095 28441
rect 17586 28432 17592 28484
rect 17644 28472 17650 28484
rect 17865 28475 17923 28481
rect 17865 28472 17877 28475
rect 17644 28444 17877 28472
rect 17644 28432 17650 28444
rect 17865 28441 17877 28444
rect 17911 28441 17923 28475
rect 17865 28435 17923 28441
rect 18874 28432 18880 28484
rect 18932 28472 18938 28484
rect 19812 28472 19840 28512
rect 20625 28509 20637 28512
rect 20671 28540 20683 28543
rect 20732 28540 20760 28580
rect 20671 28512 20760 28540
rect 20809 28543 20867 28549
rect 20671 28509 20683 28512
rect 20625 28503 20683 28509
rect 20809 28509 20821 28543
rect 20855 28540 20867 28543
rect 20898 28540 20904 28552
rect 20855 28512 20904 28540
rect 20855 28509 20867 28512
rect 20809 28503 20867 28509
rect 20898 28500 20904 28512
rect 20956 28500 20962 28552
rect 21008 28540 21036 28580
rect 21174 28568 21180 28620
rect 21232 28568 21238 28620
rect 21266 28568 21272 28620
rect 21324 28608 21330 28620
rect 21324 28580 21588 28608
rect 21324 28568 21330 28580
rect 21080 28543 21138 28549
rect 21080 28540 21092 28543
rect 21008 28512 21092 28540
rect 21080 28509 21092 28512
rect 21126 28509 21138 28543
rect 21192 28540 21220 28568
rect 21450 28540 21456 28552
rect 21192 28512 21456 28540
rect 21080 28503 21138 28509
rect 21450 28500 21456 28512
rect 21508 28500 21514 28552
rect 21560 28549 21588 28580
rect 21726 28568 21732 28620
rect 21784 28608 21790 28620
rect 21928 28608 21956 28648
rect 25317 28645 25329 28679
rect 25363 28676 25375 28679
rect 25363 28648 26556 28676
rect 25363 28645 25375 28648
rect 25317 28639 25375 28645
rect 21784 28580 21956 28608
rect 21784 28568 21790 28580
rect 22002 28568 22008 28620
rect 22060 28608 22066 28620
rect 24486 28608 24492 28620
rect 22060 28580 24492 28608
rect 22060 28568 22066 28580
rect 21545 28543 21603 28549
rect 21545 28509 21557 28543
rect 21591 28509 21603 28543
rect 21545 28503 21603 28509
rect 18932 28444 19840 28472
rect 18932 28432 18938 28444
rect 20346 28432 20352 28484
rect 20404 28472 20410 28484
rect 21174 28472 21180 28484
rect 20404 28444 21180 28472
rect 20404 28432 20410 28444
rect 21174 28432 21180 28444
rect 21232 28432 21238 28484
rect 21269 28475 21327 28481
rect 21269 28441 21281 28475
rect 21315 28472 21327 28475
rect 22020 28472 22048 28568
rect 22186 28549 22192 28552
rect 22184 28540 22192 28549
rect 22147 28512 22192 28540
rect 22184 28503 22192 28512
rect 22186 28500 22192 28503
rect 22244 28500 22250 28552
rect 22388 28549 22416 28580
rect 24486 28568 24492 28580
rect 24544 28568 24550 28620
rect 25130 28568 25136 28620
rect 25188 28608 25194 28620
rect 25225 28611 25283 28617
rect 25225 28608 25237 28611
rect 25188 28580 25237 28608
rect 25188 28568 25194 28580
rect 25225 28577 25237 28580
rect 25271 28577 25283 28611
rect 25225 28571 25283 28577
rect 25409 28611 25467 28617
rect 25409 28577 25421 28611
rect 25455 28608 25467 28611
rect 26421 28611 26479 28617
rect 26421 28608 26433 28611
rect 25455 28580 26433 28608
rect 25455 28577 25467 28580
rect 25409 28571 25467 28577
rect 26421 28577 26433 28580
rect 26467 28577 26479 28611
rect 26528 28608 26556 28648
rect 26878 28636 26884 28688
rect 26936 28636 26942 28688
rect 27706 28636 27712 28688
rect 27764 28676 27770 28688
rect 28828 28676 28856 28704
rect 27764 28648 28856 28676
rect 27764 28636 27770 28648
rect 31938 28636 31944 28688
rect 31996 28636 32002 28688
rect 32674 28676 32680 28688
rect 32324 28648 32680 28676
rect 26602 28608 26608 28620
rect 26528 28580 26608 28608
rect 26421 28571 26479 28577
rect 26602 28568 26608 28580
rect 26660 28608 26666 28620
rect 26660 28580 28028 28608
rect 26660 28568 26666 28580
rect 22373 28543 22431 28549
rect 22373 28509 22385 28543
rect 22419 28509 22431 28543
rect 22554 28540 22560 28552
rect 22515 28512 22560 28540
rect 22373 28503 22431 28509
rect 22554 28500 22560 28512
rect 22612 28500 22618 28552
rect 22649 28543 22707 28549
rect 22649 28509 22661 28543
rect 22695 28540 22707 28543
rect 23293 28543 23351 28549
rect 22695 28512 23152 28540
rect 22695 28509 22707 28512
rect 22649 28503 22707 28509
rect 21315 28444 22048 28472
rect 22281 28475 22339 28481
rect 21315 28441 21327 28444
rect 21269 28435 21327 28441
rect 22281 28441 22293 28475
rect 22327 28441 22339 28475
rect 22281 28435 22339 28441
rect 17237 28407 17295 28413
rect 17237 28404 17249 28407
rect 16776 28376 17249 28404
rect 16577 28367 16635 28373
rect 17237 28373 17249 28376
rect 17283 28373 17295 28407
rect 17237 28367 17295 28373
rect 17402 28364 17408 28416
rect 17460 28364 17466 28416
rect 17770 28364 17776 28416
rect 17828 28404 17834 28416
rect 19337 28407 19395 28413
rect 19337 28404 19349 28407
rect 17828 28376 19349 28404
rect 17828 28364 17834 28376
rect 19337 28373 19349 28376
rect 19383 28373 19395 28407
rect 21284 28404 21312 28435
rect 21358 28404 21364 28416
rect 21284 28376 21364 28404
rect 19337 28367 19395 28373
rect 21358 28364 21364 28376
rect 21416 28364 21422 28416
rect 22005 28407 22063 28413
rect 22005 28373 22017 28407
rect 22051 28404 22063 28407
rect 22186 28404 22192 28416
rect 22051 28376 22192 28404
rect 22051 28373 22063 28376
rect 22005 28367 22063 28373
rect 22186 28364 22192 28376
rect 22244 28364 22250 28416
rect 22296 28404 22324 28435
rect 23124 28416 23152 28512
rect 23293 28509 23305 28543
rect 23339 28509 23351 28543
rect 23293 28503 23351 28509
rect 23308 28472 23336 28503
rect 23382 28500 23388 28552
rect 23440 28540 23446 28552
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 23440 28512 23581 28540
rect 23440 28500 23446 28512
rect 23569 28509 23581 28512
rect 23615 28540 23627 28543
rect 25685 28543 25743 28549
rect 23615 28512 25636 28540
rect 23615 28509 23627 28512
rect 23569 28503 23627 28509
rect 23308 28444 23428 28472
rect 23400 28416 23428 28444
rect 25608 28416 25636 28512
rect 25685 28509 25697 28543
rect 25731 28509 25743 28543
rect 25685 28503 25743 28509
rect 25700 28472 25728 28503
rect 25866 28500 25872 28552
rect 25924 28540 25930 28552
rect 26050 28540 26056 28552
rect 25924 28512 26056 28540
rect 25924 28500 25930 28512
rect 26050 28500 26056 28512
rect 26108 28540 26114 28552
rect 26145 28543 26203 28549
rect 26145 28540 26157 28543
rect 26108 28512 26157 28540
rect 26108 28500 26114 28512
rect 26145 28509 26157 28512
rect 26191 28509 26203 28543
rect 26145 28503 26203 28509
rect 26234 28500 26240 28552
rect 26292 28540 26298 28552
rect 26292 28512 26556 28540
rect 26292 28500 26298 28512
rect 26418 28472 26424 28484
rect 25700 28444 26424 28472
rect 26418 28432 26424 28444
rect 26476 28432 26482 28484
rect 26528 28472 26556 28512
rect 26694 28500 26700 28552
rect 26752 28500 26758 28552
rect 26786 28500 26792 28552
rect 26844 28500 26850 28552
rect 26970 28500 26976 28552
rect 27028 28500 27034 28552
rect 27614 28500 27620 28552
rect 27672 28540 27678 28552
rect 28000 28549 28028 28580
rect 31018 28568 31024 28620
rect 31076 28608 31082 28620
rect 31956 28608 31984 28636
rect 31076 28580 31984 28608
rect 31076 28568 31082 28580
rect 27709 28543 27767 28549
rect 27709 28540 27721 28543
rect 27672 28512 27721 28540
rect 27672 28500 27678 28512
rect 27709 28509 27721 28512
rect 27755 28509 27767 28543
rect 27709 28503 27767 28509
rect 27985 28543 28043 28549
rect 27985 28509 27997 28543
rect 28031 28509 28043 28543
rect 27985 28503 28043 28509
rect 29089 28543 29147 28549
rect 29089 28509 29101 28543
rect 29135 28540 29147 28543
rect 29178 28540 29184 28552
rect 29135 28512 29184 28540
rect 29135 28509 29147 28512
rect 29089 28503 29147 28509
rect 29178 28500 29184 28512
rect 29236 28500 29242 28552
rect 30466 28500 30472 28552
rect 30524 28540 30530 28552
rect 31110 28540 31116 28552
rect 30524 28512 31116 28540
rect 30524 28500 30530 28512
rect 31110 28500 31116 28512
rect 31168 28500 31174 28552
rect 31956 28549 31984 28580
rect 31941 28543 31999 28549
rect 31941 28509 31953 28543
rect 31987 28509 31999 28543
rect 31941 28503 31999 28509
rect 32030 28500 32036 28552
rect 32088 28500 32094 28552
rect 32122 28500 32128 28552
rect 32180 28500 32186 28552
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32324 28540 32352 28648
rect 32674 28636 32680 28648
rect 32732 28676 32738 28688
rect 32769 28679 32827 28685
rect 32769 28676 32781 28679
rect 32732 28648 32781 28676
rect 32732 28636 32738 28648
rect 32769 28645 32781 28648
rect 32815 28645 32827 28679
rect 32769 28639 32827 28645
rect 33134 28636 33140 28688
rect 33192 28676 33198 28688
rect 33594 28676 33600 28688
rect 33192 28648 33600 28676
rect 33192 28636 33198 28648
rect 33594 28636 33600 28648
rect 33652 28636 33658 28688
rect 32876 28580 33824 28608
rect 32493 28543 32551 28549
rect 32493 28540 32505 28543
rect 32324 28512 32505 28540
rect 32217 28503 32275 28509
rect 32493 28509 32505 28512
rect 32539 28509 32551 28543
rect 32493 28503 32551 28509
rect 27249 28475 27307 28481
rect 27249 28472 27261 28475
rect 26528 28444 27261 28472
rect 27249 28441 27261 28444
rect 27295 28441 27307 28475
rect 28258 28472 28264 28484
rect 27249 28435 27307 28441
rect 27724 28444 28264 28472
rect 22554 28404 22560 28416
rect 22296 28376 22560 28404
rect 22554 28364 22560 28376
rect 22612 28364 22618 28416
rect 23106 28364 23112 28416
rect 23164 28364 23170 28416
rect 23382 28364 23388 28416
rect 23440 28364 23446 28416
rect 23477 28407 23535 28413
rect 23477 28373 23489 28407
rect 23523 28404 23535 28407
rect 23842 28404 23848 28416
rect 23523 28376 23848 28404
rect 23523 28373 23535 28376
rect 23477 28367 23535 28373
rect 23842 28364 23848 28376
rect 23900 28364 23906 28416
rect 25590 28364 25596 28416
rect 25648 28364 25654 28416
rect 25774 28364 25780 28416
rect 25832 28364 25838 28416
rect 26510 28364 26516 28416
rect 26568 28364 26574 28416
rect 26786 28364 26792 28416
rect 26844 28404 26850 28416
rect 27724 28404 27752 28444
rect 28258 28432 28264 28444
rect 28316 28432 28322 28484
rect 28350 28432 28356 28484
rect 28408 28472 28414 28484
rect 28445 28475 28503 28481
rect 28445 28472 28457 28475
rect 28408 28444 28457 28472
rect 28408 28432 28414 28444
rect 28445 28441 28457 28444
rect 28491 28472 28503 28475
rect 31386 28472 31392 28484
rect 28491 28444 31392 28472
rect 28491 28441 28503 28444
rect 28445 28435 28503 28441
rect 31386 28432 31392 28444
rect 31444 28432 31450 28484
rect 32048 28472 32076 28500
rect 32232 28472 32260 28503
rect 32674 28500 32680 28552
rect 32732 28500 32738 28552
rect 32876 28549 32904 28580
rect 33796 28552 33824 28580
rect 34054 28568 34060 28620
rect 34112 28568 34118 28620
rect 34606 28568 34612 28620
rect 34664 28608 34670 28620
rect 35161 28611 35219 28617
rect 35161 28608 35173 28611
rect 34664 28580 35173 28608
rect 34664 28568 34670 28580
rect 35161 28577 35173 28580
rect 35207 28608 35219 28611
rect 35805 28611 35863 28617
rect 35805 28608 35817 28611
rect 35207 28580 35817 28608
rect 35207 28577 35219 28580
rect 35161 28571 35219 28577
rect 35805 28577 35817 28580
rect 35851 28577 35863 28611
rect 35805 28571 35863 28577
rect 32861 28543 32919 28549
rect 32861 28509 32873 28543
rect 32907 28509 32919 28543
rect 32861 28503 32919 28509
rect 33226 28500 33232 28552
rect 33284 28500 33290 28552
rect 33410 28500 33416 28552
rect 33468 28500 33474 28552
rect 33505 28543 33563 28549
rect 33505 28509 33517 28543
rect 33551 28509 33563 28543
rect 33505 28503 33563 28509
rect 33520 28472 33548 28503
rect 33778 28500 33784 28552
rect 33836 28500 33842 28552
rect 34241 28543 34299 28549
rect 34241 28509 34253 28543
rect 34287 28540 34299 28543
rect 34698 28540 34704 28552
rect 34287 28512 34704 28540
rect 34287 28509 34299 28512
rect 34241 28503 34299 28509
rect 34698 28500 34704 28512
rect 34756 28500 34762 28552
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 34974 28540 34980 28552
rect 34848 28512 34980 28540
rect 34848 28500 34854 28512
rect 34974 28500 34980 28512
rect 35032 28500 35038 28552
rect 35066 28500 35072 28552
rect 35124 28500 35130 28552
rect 35250 28500 35256 28552
rect 35308 28500 35314 28552
rect 32048 28444 32260 28472
rect 33428 28444 33548 28472
rect 33428 28416 33456 28444
rect 35434 28432 35440 28484
rect 35492 28472 35498 28484
rect 35529 28475 35587 28481
rect 35529 28472 35541 28475
rect 35492 28444 35541 28472
rect 35492 28432 35498 28444
rect 35529 28441 35541 28444
rect 35575 28441 35587 28475
rect 35529 28435 35587 28441
rect 26844 28376 27752 28404
rect 26844 28364 26850 28376
rect 27798 28364 27804 28416
rect 27856 28364 27862 28416
rect 28810 28364 28816 28416
rect 28868 28413 28874 28416
rect 28868 28404 28880 28413
rect 28868 28376 28913 28404
rect 28868 28367 28880 28376
rect 28868 28364 28874 28367
rect 29178 28364 29184 28416
rect 29236 28404 29242 28416
rect 29730 28404 29736 28416
rect 29236 28376 29736 28404
rect 29236 28364 29242 28376
rect 29730 28364 29736 28376
rect 29788 28404 29794 28416
rect 30834 28404 30840 28416
rect 29788 28376 30840 28404
rect 29788 28364 29794 28376
rect 30834 28364 30840 28376
rect 30892 28404 30898 28416
rect 31570 28404 31576 28416
rect 30892 28376 31576 28404
rect 30892 28364 30898 28376
rect 31570 28364 31576 28376
rect 31628 28364 31634 28416
rect 32030 28364 32036 28416
rect 32088 28364 32094 28416
rect 32493 28407 32551 28413
rect 32493 28373 32505 28407
rect 32539 28404 32551 28407
rect 32858 28404 32864 28416
rect 32539 28376 32864 28404
rect 32539 28373 32551 28376
rect 32493 28367 32551 28373
rect 32858 28364 32864 28376
rect 32916 28364 32922 28416
rect 33321 28407 33379 28413
rect 33321 28373 33333 28407
rect 33367 28404 33379 28407
rect 33410 28404 33416 28416
rect 33367 28376 33416 28404
rect 33367 28373 33379 28376
rect 33321 28367 33379 28373
rect 33410 28364 33416 28376
rect 33468 28364 33474 28416
rect 34330 28364 34336 28416
rect 34388 28404 34394 28416
rect 34425 28407 34483 28413
rect 34425 28404 34437 28407
rect 34388 28376 34437 28404
rect 34388 28364 34394 28376
rect 34425 28373 34437 28376
rect 34471 28373 34483 28407
rect 34425 28367 34483 28373
rect 1104 28314 36524 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 36524 28314
rect 1104 28240 36524 28262
rect 1670 28160 1676 28212
rect 1728 28200 1734 28212
rect 2409 28203 2467 28209
rect 2409 28200 2421 28203
rect 1728 28172 2421 28200
rect 1728 28160 1734 28172
rect 2409 28169 2421 28172
rect 2455 28169 2467 28203
rect 2409 28163 2467 28169
rect 3988 28172 4660 28200
rect 3988 28141 4016 28172
rect 3973 28135 4031 28141
rect 3973 28101 3985 28135
rect 4019 28101 4031 28135
rect 3973 28095 4031 28101
rect 4065 28135 4123 28141
rect 4065 28101 4077 28135
rect 4111 28132 4123 28135
rect 4246 28132 4252 28144
rect 4111 28104 4252 28132
rect 4111 28101 4123 28104
rect 4065 28095 4123 28101
rect 4246 28092 4252 28104
rect 4304 28092 4310 28144
rect 4632 28076 4660 28172
rect 4798 28160 4804 28212
rect 4856 28200 4862 28212
rect 5077 28203 5135 28209
rect 5077 28200 5089 28203
rect 4856 28172 5089 28200
rect 4856 28160 4862 28172
rect 5077 28169 5089 28172
rect 5123 28169 5135 28203
rect 5077 28163 5135 28169
rect 6840 28172 7788 28200
rect 4709 28135 4767 28141
rect 4709 28101 4721 28135
rect 4755 28132 4767 28135
rect 4755 28104 5488 28132
rect 4755 28101 4767 28104
rect 4709 28095 4767 28101
rect 5460 28076 5488 28104
rect 2774 28024 2780 28076
rect 2832 28024 2838 28076
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28064 2927 28067
rect 3142 28064 3148 28076
rect 2915 28036 3148 28064
rect 2915 28033 2927 28036
rect 2869 28027 2927 28033
rect 3142 28024 3148 28036
rect 3200 28064 3206 28076
rect 3789 28067 3847 28073
rect 3789 28064 3801 28067
rect 3200 28036 3801 28064
rect 3200 28024 3206 28036
rect 3789 28033 3801 28036
rect 3835 28033 3847 28067
rect 3789 28027 3847 28033
rect 3050 27956 3056 28008
rect 3108 27956 3114 28008
rect 3804 27996 3832 28027
rect 4154 28024 4160 28076
rect 4212 28024 4218 28076
rect 4430 28024 4436 28076
rect 4488 28024 4494 28076
rect 4614 28024 4620 28076
rect 4672 28024 4678 28076
rect 4801 28067 4859 28073
rect 4801 28033 4813 28067
rect 4847 28064 4859 28067
rect 4982 28064 4988 28076
rect 4847 28036 4988 28064
rect 4847 28033 4859 28036
rect 4801 28027 4859 28033
rect 4982 28024 4988 28036
rect 5040 28024 5046 28076
rect 5442 28024 5448 28076
rect 5500 28064 5506 28076
rect 5629 28067 5687 28073
rect 5629 28064 5641 28067
rect 5500 28036 5641 28064
rect 5500 28024 5506 28036
rect 5629 28033 5641 28036
rect 5675 28033 5687 28067
rect 5629 28027 5687 28033
rect 5718 28024 5724 28076
rect 5776 28064 5782 28076
rect 6733 28067 6791 28073
rect 6733 28064 6745 28067
rect 5776 28036 6745 28064
rect 5776 28024 5782 28036
rect 6733 28033 6745 28036
rect 6779 28033 6791 28067
rect 6733 28027 6791 28033
rect 6840 27996 6868 28172
rect 7650 28132 7656 28144
rect 7116 28104 7656 28132
rect 7116 28073 7144 28104
rect 7650 28092 7656 28104
rect 7708 28092 7714 28144
rect 7760 28132 7788 28172
rect 8478 28160 8484 28212
rect 8536 28160 8542 28212
rect 9674 28160 9680 28212
rect 9732 28200 9738 28212
rect 10229 28203 10287 28209
rect 10229 28200 10241 28203
rect 9732 28172 10241 28200
rect 9732 28160 9738 28172
rect 10229 28169 10241 28172
rect 10275 28169 10287 28203
rect 11514 28200 11520 28212
rect 10229 28163 10287 28169
rect 10796 28172 11520 28200
rect 7760 28104 10640 28132
rect 7101 28067 7159 28073
rect 7101 28033 7113 28067
rect 7147 28033 7159 28067
rect 7285 28067 7343 28073
rect 7285 28064 7297 28067
rect 7101 28027 7159 28033
rect 7208 28036 7297 28064
rect 3804 27968 6868 27996
rect 5810 27888 5816 27940
rect 5868 27928 5874 27940
rect 7208 27928 7236 28036
rect 7285 28033 7297 28036
rect 7331 28033 7343 28067
rect 7285 28027 7343 28033
rect 7558 28024 7564 28076
rect 7616 28024 7622 28076
rect 8386 28024 8392 28076
rect 8444 28024 8450 28076
rect 8573 28067 8631 28073
rect 8573 28033 8585 28067
rect 8619 28064 8631 28067
rect 8938 28064 8944 28076
rect 8619 28036 8944 28064
rect 8619 28033 8631 28036
rect 8573 28027 8631 28033
rect 8938 28024 8944 28036
rect 8996 28024 9002 28076
rect 10502 28024 10508 28076
rect 10560 28024 10566 28076
rect 10612 28064 10640 28104
rect 10686 28092 10692 28144
rect 10744 28132 10750 28144
rect 10796 28141 10824 28172
rect 11514 28160 11520 28172
rect 11572 28160 11578 28212
rect 12250 28160 12256 28212
rect 12308 28200 12314 28212
rect 16669 28203 16727 28209
rect 16669 28200 16681 28203
rect 12308 28172 16681 28200
rect 12308 28160 12314 28172
rect 16669 28169 16681 28172
rect 16715 28169 16727 28203
rect 16669 28163 16727 28169
rect 17678 28160 17684 28212
rect 17736 28200 17742 28212
rect 17773 28203 17831 28209
rect 17773 28200 17785 28203
rect 17736 28172 17785 28200
rect 17736 28160 17742 28172
rect 17773 28169 17785 28172
rect 17819 28169 17831 28203
rect 17773 28163 17831 28169
rect 18046 28160 18052 28212
rect 18104 28200 18110 28212
rect 19061 28203 19119 28209
rect 19061 28200 19073 28203
rect 18104 28172 19073 28200
rect 18104 28160 18110 28172
rect 19061 28169 19073 28172
rect 19107 28169 19119 28203
rect 19061 28163 19119 28169
rect 19150 28160 19156 28212
rect 19208 28200 19214 28212
rect 28810 28200 28816 28212
rect 19208 28172 28816 28200
rect 19208 28160 19214 28172
rect 28810 28160 28816 28172
rect 28868 28160 28874 28212
rect 29086 28160 29092 28212
rect 29144 28160 29150 28212
rect 29717 28203 29775 28209
rect 29717 28200 29729 28203
rect 29564 28172 29729 28200
rect 10781 28135 10839 28141
rect 10781 28132 10793 28135
rect 10744 28104 10793 28132
rect 10744 28092 10750 28104
rect 10781 28101 10793 28104
rect 10827 28101 10839 28135
rect 10781 28095 10839 28101
rect 10873 28135 10931 28141
rect 10873 28101 10885 28135
rect 10919 28132 10931 28135
rect 11054 28132 11060 28144
rect 10919 28104 11060 28132
rect 10919 28101 10931 28104
rect 10873 28095 10931 28101
rect 11054 28092 11060 28104
rect 11112 28092 11118 28144
rect 14826 28132 14832 28144
rect 12636 28104 14832 28132
rect 11238 28064 11244 28076
rect 10612 28036 11244 28064
rect 11238 28024 11244 28036
rect 11296 28024 11302 28076
rect 12342 28024 12348 28076
rect 12400 28064 12406 28076
rect 12636 28073 12664 28104
rect 14826 28092 14832 28104
rect 14884 28092 14890 28144
rect 16945 28135 17003 28141
rect 16945 28101 16957 28135
rect 16991 28132 17003 28135
rect 28350 28132 28356 28144
rect 16991 28104 21440 28132
rect 16991 28101 17003 28104
rect 16945 28095 17003 28101
rect 12621 28067 12679 28073
rect 12621 28064 12633 28067
rect 12400 28036 12633 28064
rect 12400 28024 12406 28036
rect 12621 28033 12633 28036
rect 12667 28033 12679 28067
rect 12621 28027 12679 28033
rect 16666 28024 16672 28076
rect 16724 28064 16730 28076
rect 16807 28067 16865 28073
rect 16807 28064 16819 28067
rect 16724 28036 16819 28064
rect 16724 28024 16730 28036
rect 16807 28033 16819 28036
rect 16853 28033 16865 28067
rect 16807 28027 16865 28033
rect 10134 27956 10140 28008
rect 10192 27996 10198 28008
rect 10413 27999 10471 28005
rect 10413 27996 10425 27999
rect 10192 27968 10425 27996
rect 10192 27956 10198 27968
rect 10413 27965 10425 27968
rect 10459 27996 10471 27999
rect 11146 27996 11152 28008
rect 10459 27968 11152 27996
rect 10459 27965 10471 27968
rect 10413 27959 10471 27965
rect 11146 27956 11152 27968
rect 11204 27956 11210 28008
rect 11698 27956 11704 28008
rect 11756 27996 11762 28008
rect 12802 27996 12808 28008
rect 11756 27968 12808 27996
rect 11756 27956 11762 27968
rect 12802 27956 12808 27968
rect 12860 27956 12866 28008
rect 12894 27956 12900 28008
rect 12952 27956 12958 28008
rect 5868 27900 7236 27928
rect 5868 27888 5874 27900
rect 7374 27888 7380 27940
rect 7432 27888 7438 27940
rect 11606 27888 11612 27940
rect 11664 27928 11670 27940
rect 16960 27928 16988 28095
rect 17037 28067 17095 28073
rect 17037 28033 17049 28067
rect 17083 28033 17095 28067
rect 17218 28064 17224 28076
rect 17179 28036 17224 28064
rect 17037 28027 17095 28033
rect 11664 27900 16988 27928
rect 11664 27888 11670 27900
rect 2498 27820 2504 27872
rect 2556 27860 2562 27872
rect 4341 27863 4399 27869
rect 4341 27860 4353 27863
rect 2556 27832 4353 27860
rect 2556 27820 2562 27832
rect 4341 27829 4353 27832
rect 4387 27829 4399 27863
rect 4341 27823 4399 27829
rect 4706 27820 4712 27872
rect 4764 27860 4770 27872
rect 4985 27863 5043 27869
rect 4985 27860 4997 27863
rect 4764 27832 4997 27860
rect 4764 27820 4770 27832
rect 4985 27829 4997 27832
rect 5031 27829 5043 27863
rect 4985 27823 5043 27829
rect 11238 27820 11244 27872
rect 11296 27860 11302 27872
rect 12437 27863 12495 27869
rect 12437 27860 12449 27863
rect 11296 27832 12449 27860
rect 11296 27820 11302 27832
rect 12437 27829 12449 27832
rect 12483 27829 12495 27863
rect 12437 27823 12495 27829
rect 12805 27863 12863 27869
rect 12805 27829 12817 27863
rect 12851 27860 12863 27863
rect 16390 27860 16396 27872
rect 12851 27832 16396 27860
rect 12851 27829 12863 27832
rect 12805 27823 12863 27829
rect 16390 27820 16396 27832
rect 16448 27820 16454 27872
rect 16850 27820 16856 27872
rect 16908 27860 16914 27872
rect 17052 27860 17080 28027
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 17313 28067 17371 28073
rect 17313 28033 17325 28067
rect 17359 28064 17371 28067
rect 17402 28064 17408 28076
rect 17359 28036 17408 28064
rect 17359 28033 17371 28036
rect 17313 28027 17371 28033
rect 17402 28024 17408 28036
rect 17460 28024 17466 28076
rect 17681 28067 17739 28073
rect 17681 28033 17693 28067
rect 17727 28033 17739 28067
rect 17681 28027 17739 28033
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28033 17923 28067
rect 17865 28027 17923 28033
rect 17696 27928 17724 28027
rect 17880 27996 17908 28027
rect 18046 28024 18052 28076
rect 18104 28064 18110 28076
rect 18141 28067 18199 28073
rect 18141 28064 18153 28067
rect 18104 28036 18153 28064
rect 18104 28024 18110 28036
rect 18141 28033 18153 28036
rect 18187 28033 18199 28067
rect 18141 28027 18199 28033
rect 18322 28024 18328 28076
rect 18380 28024 18386 28076
rect 18414 28024 18420 28076
rect 18472 28024 18478 28076
rect 18601 28067 18659 28073
rect 18601 28033 18613 28067
rect 18647 28033 18659 28067
rect 18601 28027 18659 28033
rect 18877 28067 18935 28073
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 19521 28067 19579 28073
rect 19521 28033 19533 28067
rect 19567 28064 19579 28067
rect 19567 28036 19748 28064
rect 19567 28033 19579 28036
rect 19521 28027 19579 28033
rect 17957 27999 18015 28005
rect 17957 27996 17969 27999
rect 17880 27968 17969 27996
rect 17957 27965 17969 27968
rect 18003 27996 18015 27999
rect 18616 27996 18644 28027
rect 18003 27968 18644 27996
rect 18003 27965 18015 27968
rect 17957 27959 18015 27965
rect 18690 27956 18696 28008
rect 18748 27956 18754 28008
rect 18138 27928 18144 27940
rect 17696 27900 18144 27928
rect 18138 27888 18144 27900
rect 18196 27888 18202 27940
rect 16908 27832 17080 27860
rect 16908 27820 16914 27832
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 18892 27860 18920 28027
rect 18966 27956 18972 28008
rect 19024 27996 19030 28008
rect 19613 27999 19671 28005
rect 19613 27996 19625 27999
rect 19024 27968 19625 27996
rect 19024 27956 19030 27968
rect 19613 27965 19625 27968
rect 19659 27965 19671 27999
rect 19613 27959 19671 27965
rect 18012 27832 18920 27860
rect 18012 27820 18018 27832
rect 19518 27820 19524 27872
rect 19576 27820 19582 27872
rect 19610 27820 19616 27872
rect 19668 27860 19674 27872
rect 19720 27860 19748 28036
rect 19886 28024 19892 28076
rect 19944 28064 19950 28076
rect 20993 28067 21051 28073
rect 19944 28062 20760 28064
rect 20993 28062 21005 28067
rect 19944 28036 21005 28062
rect 19944 28024 19950 28036
rect 20732 28034 21005 28036
rect 20993 28033 21005 28034
rect 21039 28033 21051 28067
rect 20993 28027 21051 28033
rect 21082 28024 21088 28076
rect 21140 28024 21146 28076
rect 20622 27956 20628 28008
rect 20680 27996 20686 28008
rect 20809 27999 20867 28005
rect 20809 27996 20821 27999
rect 20680 27968 20821 27996
rect 20680 27956 20686 27968
rect 20809 27965 20821 27968
rect 20855 27965 20867 27999
rect 21412 27996 21440 28104
rect 23308 28104 28356 28132
rect 21542 28024 21548 28076
rect 21600 28064 21606 28076
rect 22738 28064 22744 28076
rect 21600 28036 22744 28064
rect 21600 28024 21606 28036
rect 22738 28024 22744 28036
rect 22796 28024 22802 28076
rect 23308 27996 23336 28104
rect 28350 28092 28356 28104
rect 28408 28092 28414 28144
rect 28994 28092 29000 28144
rect 29052 28132 29058 28144
rect 29564 28132 29592 28172
rect 29717 28169 29729 28172
rect 29763 28200 29775 28203
rect 29763 28172 30420 28200
rect 29763 28169 29775 28172
rect 29717 28163 29775 28169
rect 29052 28104 29592 28132
rect 29052 28092 29058 28104
rect 29914 28092 29920 28144
rect 29972 28092 29978 28144
rect 30006 28092 30012 28144
rect 30064 28132 30070 28144
rect 30064 28104 30328 28132
rect 30064 28092 30070 28104
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28064 23719 28067
rect 23934 28064 23940 28076
rect 23707 28036 23940 28064
rect 23707 28033 23719 28036
rect 23661 28027 23719 28033
rect 23934 28024 23940 28036
rect 23992 28024 23998 28076
rect 24213 28067 24271 28073
rect 24213 28033 24225 28067
rect 24259 28064 24271 28067
rect 24302 28064 24308 28076
rect 24259 28036 24308 28064
rect 24259 28033 24271 28036
rect 24213 28027 24271 28033
rect 24302 28024 24308 28036
rect 24360 28024 24366 28076
rect 24397 28067 24455 28073
rect 24397 28033 24409 28067
rect 24443 28033 24455 28067
rect 24397 28027 24455 28033
rect 21412 27968 23336 27996
rect 20809 27959 20867 27965
rect 23382 27956 23388 28008
rect 23440 27996 23446 28008
rect 23477 27999 23535 28005
rect 23477 27996 23489 27999
rect 23440 27968 23489 27996
rect 23440 27956 23446 27968
rect 23477 27965 23489 27968
rect 23523 27996 23535 27999
rect 24412 27996 24440 28027
rect 25590 28024 25596 28076
rect 25648 28064 25654 28076
rect 25958 28064 25964 28076
rect 25648 28036 25964 28064
rect 25648 28024 25654 28036
rect 25958 28024 25964 28036
rect 26016 28064 26022 28076
rect 26053 28067 26111 28073
rect 26053 28064 26065 28067
rect 26016 28036 26065 28064
rect 26016 28024 26022 28036
rect 26053 28033 26065 28036
rect 26099 28064 26111 28067
rect 27798 28064 27804 28076
rect 26099 28036 27804 28064
rect 26099 28033 26111 28036
rect 26053 28027 26111 28033
rect 27798 28024 27804 28036
rect 27856 28024 27862 28076
rect 28077 28067 28135 28073
rect 28077 28033 28089 28067
rect 28123 28064 28135 28067
rect 28445 28067 28503 28073
rect 28445 28064 28457 28067
rect 28123 28036 28457 28064
rect 28123 28033 28135 28036
rect 28077 28027 28135 28033
rect 28445 28033 28457 28036
rect 28491 28033 28503 28067
rect 28445 28027 28503 28033
rect 28902 28024 28908 28076
rect 28960 28024 28966 28076
rect 29089 28067 29147 28073
rect 29089 28033 29101 28067
rect 29135 28064 29147 28067
rect 29178 28064 29184 28076
rect 29135 28036 29184 28064
rect 29135 28033 29147 28036
rect 29089 28027 29147 28033
rect 29178 28024 29184 28036
rect 29236 28024 29242 28076
rect 29270 28024 29276 28076
rect 29328 28064 29334 28076
rect 30300 28073 30328 28104
rect 30193 28067 30251 28073
rect 30193 28064 30205 28067
rect 29328 28036 30205 28064
rect 29328 28024 29334 28036
rect 30193 28033 30205 28036
rect 30239 28033 30251 28067
rect 30193 28027 30251 28033
rect 30285 28067 30343 28073
rect 30285 28033 30297 28067
rect 30331 28033 30343 28067
rect 30392 28064 30420 28172
rect 30466 28160 30472 28212
rect 30524 28200 30530 28212
rect 30745 28203 30803 28209
rect 30745 28200 30757 28203
rect 30524 28172 30757 28200
rect 30524 28160 30530 28172
rect 30745 28169 30757 28172
rect 30791 28169 30803 28203
rect 30745 28163 30803 28169
rect 31570 28160 31576 28212
rect 31628 28160 31634 28212
rect 32122 28160 32128 28212
rect 32180 28200 32186 28212
rect 32180 28172 32450 28200
rect 32180 28160 32186 28172
rect 30653 28135 30711 28141
rect 30653 28101 30665 28135
rect 30699 28132 30711 28135
rect 31294 28132 31300 28144
rect 30699 28104 31300 28132
rect 30699 28101 30711 28104
rect 30653 28095 30711 28101
rect 31294 28092 31300 28104
rect 31352 28092 31358 28144
rect 31588 28132 31616 28160
rect 32422 28132 32450 28172
rect 32490 28160 32496 28212
rect 32548 28160 32554 28212
rect 33511 28203 33569 28209
rect 32600 28172 33364 28200
rect 32600 28132 32628 28172
rect 33336 28141 33364 28172
rect 33511 28169 33523 28203
rect 33557 28200 33569 28203
rect 33870 28200 33876 28212
rect 33557 28172 33876 28200
rect 33557 28169 33569 28172
rect 33511 28163 33569 28169
rect 33870 28160 33876 28172
rect 33928 28160 33934 28212
rect 31588 28104 31984 28132
rect 32422 28104 32628 28132
rect 33295 28135 33364 28141
rect 30392 28036 30696 28064
rect 30285 28027 30343 28033
rect 23523 27968 24440 27996
rect 23523 27965 23535 27968
rect 23477 27959 23535 27965
rect 24578 27956 24584 28008
rect 24636 27996 24642 28008
rect 24673 27999 24731 28005
rect 24673 27996 24685 27999
rect 24636 27968 24685 27996
rect 24636 27956 24642 27968
rect 24673 27965 24685 27968
rect 24719 27965 24731 27999
rect 24673 27959 24731 27965
rect 25314 27956 25320 28008
rect 25372 27996 25378 28008
rect 25866 27996 25872 28008
rect 25372 27968 25872 27996
rect 25372 27956 25378 27968
rect 25866 27956 25872 27968
rect 25924 27996 25930 28008
rect 26329 27999 26387 28005
rect 26329 27996 26341 27999
rect 25924 27968 26341 27996
rect 25924 27956 25930 27968
rect 26329 27965 26341 27968
rect 26375 27965 26387 27999
rect 26329 27959 26387 27965
rect 19889 27931 19947 27937
rect 19889 27897 19901 27931
rect 19935 27928 19947 27931
rect 23658 27928 23664 27940
rect 19935 27900 23664 27928
rect 19935 27897 19947 27900
rect 19889 27891 19947 27897
rect 23658 27888 23664 27900
rect 23716 27888 23722 27940
rect 24489 27931 24547 27937
rect 24489 27928 24501 27931
rect 23768 27900 24501 27928
rect 21542 27860 21548 27872
rect 19668 27832 21548 27860
rect 19668 27820 19674 27832
rect 21542 27820 21548 27832
rect 21600 27820 21606 27872
rect 22278 27820 22284 27872
rect 22336 27860 22342 27872
rect 23768 27860 23796 27900
rect 24489 27897 24501 27900
rect 24535 27928 24547 27931
rect 25406 27928 25412 27940
rect 24535 27900 25412 27928
rect 24535 27897 24547 27900
rect 24489 27891 24547 27897
rect 25406 27888 25412 27900
rect 25464 27888 25470 27940
rect 26344 27928 26372 27959
rect 26878 27956 26884 28008
rect 26936 27996 26942 28008
rect 27433 27999 27491 28005
rect 27433 27996 27445 27999
rect 26936 27968 27445 27996
rect 26936 27956 26942 27968
rect 27433 27965 27445 27968
rect 27479 27965 27491 27999
rect 27433 27959 27491 27965
rect 28350 27956 28356 28008
rect 28408 27956 28414 28008
rect 28813 27999 28871 28005
rect 28813 27965 28825 27999
rect 28859 27996 28871 27999
rect 30098 27996 30104 28008
rect 28859 27968 30104 27996
rect 28859 27965 28871 27968
rect 28813 27959 28871 27965
rect 30098 27956 30104 27968
rect 30156 27956 30162 28008
rect 30466 27956 30472 28008
rect 30524 27996 30530 28008
rect 30561 27999 30619 28005
rect 30561 27996 30573 27999
rect 30524 27968 30573 27996
rect 30524 27956 30530 27968
rect 30561 27965 30573 27968
rect 30607 27965 30619 27999
rect 30561 27959 30619 27965
rect 29454 27928 29460 27940
rect 26344 27900 29460 27928
rect 29454 27888 29460 27900
rect 29512 27888 29518 27940
rect 30668 27928 30696 28036
rect 31478 28024 31484 28076
rect 31536 28024 31542 28076
rect 31570 28024 31576 28076
rect 31628 28064 31634 28076
rect 31956 28073 31984 28104
rect 33091 28101 33149 28107
rect 33091 28098 33103 28101
rect 31757 28067 31815 28073
rect 31757 28064 31769 28067
rect 31628 28036 31769 28064
rect 31628 28024 31634 28036
rect 31757 28033 31769 28036
rect 31803 28033 31815 28067
rect 31757 28027 31815 28033
rect 31941 28067 31999 28073
rect 31941 28033 31953 28067
rect 31987 28033 31999 28067
rect 31941 28027 31999 28033
rect 32401 28067 32459 28073
rect 32401 28033 32413 28067
rect 32447 28033 32459 28067
rect 32401 28027 32459 28033
rect 30926 27956 30932 28008
rect 30984 27956 30990 28008
rect 31021 27999 31079 28005
rect 31021 27965 31033 27999
rect 31067 27996 31079 27999
rect 31067 27968 31892 27996
rect 31067 27965 31079 27968
rect 31021 27959 31079 27965
rect 29564 27900 30604 27928
rect 30668 27900 31340 27928
rect 22336 27832 23796 27860
rect 24029 27863 24087 27869
rect 22336 27820 22342 27832
rect 24029 27829 24041 27863
rect 24075 27860 24087 27863
rect 24302 27860 24308 27872
rect 24075 27832 24308 27860
rect 24075 27829 24087 27832
rect 24029 27823 24087 27829
rect 24302 27820 24308 27832
rect 24360 27820 24366 27872
rect 24581 27863 24639 27869
rect 24581 27829 24593 27863
rect 24627 27860 24639 27863
rect 24854 27860 24860 27872
rect 24627 27832 24860 27860
rect 24627 27829 24639 27832
rect 24581 27823 24639 27829
rect 24854 27820 24860 27832
rect 24912 27820 24918 27872
rect 25866 27820 25872 27872
rect 25924 27820 25930 27872
rect 26237 27863 26295 27869
rect 26237 27829 26249 27863
rect 26283 27860 26295 27863
rect 26418 27860 26424 27872
rect 26283 27832 26424 27860
rect 26283 27829 26295 27832
rect 26237 27823 26295 27829
rect 26418 27820 26424 27832
rect 26476 27820 26482 27872
rect 28166 27820 28172 27872
rect 28224 27820 28230 27872
rect 29086 27820 29092 27872
rect 29144 27860 29150 27872
rect 29564 27869 29592 27900
rect 30576 27872 30604 27900
rect 31312 27872 31340 27900
rect 31662 27888 31668 27940
rect 31720 27928 31726 27940
rect 31754 27928 31760 27940
rect 31720 27900 31760 27928
rect 31720 27888 31726 27900
rect 31754 27888 31760 27900
rect 31812 27888 31818 27940
rect 29549 27863 29607 27869
rect 29549 27860 29561 27863
rect 29144 27832 29561 27860
rect 29144 27820 29150 27832
rect 29549 27829 29561 27832
rect 29595 27829 29607 27863
rect 29549 27823 29607 27829
rect 29733 27863 29791 27869
rect 29733 27829 29745 27863
rect 29779 27860 29791 27863
rect 30009 27863 30067 27869
rect 30009 27860 30021 27863
rect 29779 27832 30021 27860
rect 29779 27829 29791 27832
rect 29733 27823 29791 27829
rect 30009 27829 30021 27832
rect 30055 27860 30067 27863
rect 30282 27860 30288 27872
rect 30055 27832 30288 27860
rect 30055 27829 30067 27832
rect 30009 27823 30067 27829
rect 30282 27820 30288 27832
rect 30340 27820 30346 27872
rect 30558 27820 30564 27872
rect 30616 27820 30622 27872
rect 30834 27820 30840 27872
rect 30892 27860 30898 27872
rect 31205 27863 31263 27869
rect 31205 27860 31217 27863
rect 30892 27832 31217 27860
rect 30892 27820 30898 27832
rect 31205 27829 31217 27832
rect 31251 27829 31263 27863
rect 31205 27823 31263 27829
rect 31294 27820 31300 27872
rect 31352 27860 31358 27872
rect 31389 27863 31447 27869
rect 31389 27860 31401 27863
rect 31352 27832 31401 27860
rect 31352 27820 31358 27832
rect 31389 27829 31401 27832
rect 31435 27829 31447 27863
rect 31864 27860 31892 27968
rect 32122 27956 32128 28008
rect 32180 27956 32186 28008
rect 31941 27931 31999 27937
rect 31941 27897 31953 27931
rect 31987 27928 31999 27931
rect 32140 27928 32168 27956
rect 32416 27928 32444 28027
rect 32490 28024 32496 28076
rect 32548 28064 32554 28076
rect 32585 28067 32643 28073
rect 33086 28070 33103 28098
rect 32585 28064 32597 28067
rect 32548 28036 32597 28064
rect 32548 28024 32554 28036
rect 32585 28033 32597 28036
rect 32631 28033 32643 28067
rect 32968 28067 33103 28070
rect 33137 28067 33149 28101
rect 33295 28101 33307 28135
rect 33341 28104 33364 28135
rect 33341 28101 33353 28104
rect 33295 28095 33353 28101
rect 33410 28092 33416 28144
rect 33468 28132 33474 28144
rect 33468 28104 33510 28132
rect 33468 28092 33474 28104
rect 32968 28064 33149 28067
rect 32585 28027 32643 28033
rect 32784 28061 33149 28064
rect 33597 28067 33655 28073
rect 32784 28042 33114 28061
rect 32784 28036 32996 28042
rect 32784 27928 32812 28036
rect 33597 28033 33609 28067
rect 33643 28033 33655 28067
rect 33597 28027 33655 28033
rect 32861 27999 32919 28005
rect 32861 27965 32873 27999
rect 32907 27996 32919 27999
rect 33226 27996 33232 28008
rect 32907 27968 33232 27996
rect 32907 27965 32919 27968
rect 32861 27959 32919 27965
rect 33226 27956 33232 27968
rect 33284 27996 33290 28008
rect 33612 27996 33640 28027
rect 33686 28024 33692 28076
rect 33744 28064 33750 28076
rect 34606 28064 34612 28076
rect 33744 28036 34612 28064
rect 33744 28024 33750 28036
rect 34606 28024 34612 28036
rect 34664 28024 34670 28076
rect 34974 28024 34980 28076
rect 35032 28024 35038 28076
rect 35066 28024 35072 28076
rect 35124 28024 35130 28076
rect 35250 28024 35256 28076
rect 35308 28064 35314 28076
rect 35526 28064 35532 28076
rect 35308 28036 35532 28064
rect 35308 28024 35314 28036
rect 35526 28024 35532 28036
rect 35584 28024 35590 28076
rect 36170 28024 36176 28076
rect 36228 28024 36234 28076
rect 33284 27968 33640 27996
rect 35866 27968 36032 27996
rect 33284 27956 33290 27968
rect 31987 27900 32812 27928
rect 31987 27897 31999 27900
rect 31941 27891 31999 27897
rect 33502 27888 33508 27940
rect 33560 27928 33566 27940
rect 33560 27900 34928 27928
rect 33560 27888 33566 27900
rect 32125 27863 32183 27869
rect 32125 27860 32137 27863
rect 31864 27832 32137 27860
rect 31389 27823 31447 27829
rect 32125 27829 32137 27832
rect 32171 27860 32183 27863
rect 32582 27860 32588 27872
rect 32171 27832 32588 27860
rect 32171 27829 32183 27832
rect 32125 27823 32183 27829
rect 32582 27820 32588 27832
rect 32640 27820 32646 27872
rect 32674 27820 32680 27872
rect 32732 27860 32738 27872
rect 32769 27863 32827 27869
rect 32769 27860 32781 27863
rect 32732 27832 32781 27860
rect 32732 27820 32738 27832
rect 32769 27829 32781 27832
rect 32815 27829 32827 27863
rect 32769 27823 32827 27829
rect 32950 27820 32956 27872
rect 33008 27820 33014 27872
rect 33134 27820 33140 27872
rect 33192 27860 33198 27872
rect 33962 27860 33968 27872
rect 33192 27832 33968 27860
rect 33192 27820 33198 27832
rect 33962 27820 33968 27832
rect 34020 27820 34026 27872
rect 34330 27820 34336 27872
rect 34388 27860 34394 27872
rect 34900 27869 34928 27900
rect 34974 27888 34980 27940
rect 35032 27928 35038 27940
rect 35866 27928 35894 27968
rect 36004 27937 36032 27968
rect 35032 27900 35894 27928
rect 35989 27931 36047 27937
rect 35032 27888 35038 27900
rect 35989 27897 36001 27931
rect 36035 27897 36047 27931
rect 35989 27891 36047 27897
rect 34425 27863 34483 27869
rect 34425 27860 34437 27863
rect 34388 27832 34437 27860
rect 34388 27820 34394 27832
rect 34425 27829 34437 27832
rect 34471 27829 34483 27863
rect 34425 27823 34483 27829
rect 34885 27863 34943 27869
rect 34885 27829 34897 27863
rect 34931 27860 34943 27863
rect 35161 27863 35219 27869
rect 35161 27860 35173 27863
rect 34931 27832 35173 27860
rect 34931 27829 34943 27832
rect 34885 27823 34943 27829
rect 35161 27829 35173 27832
rect 35207 27829 35219 27863
rect 35161 27823 35219 27829
rect 1104 27770 36524 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 36524 27770
rect 1104 27696 36524 27718
rect 2774 27616 2780 27668
rect 2832 27656 2838 27668
rect 6914 27656 6920 27668
rect 2832 27628 6920 27656
rect 2832 27616 2838 27628
rect 6914 27616 6920 27628
rect 6972 27616 6978 27668
rect 8018 27616 8024 27668
rect 8076 27656 8082 27668
rect 8846 27656 8852 27668
rect 8076 27628 8852 27656
rect 8076 27616 8082 27628
rect 8846 27616 8852 27628
rect 8904 27616 8910 27668
rect 8938 27616 8944 27668
rect 8996 27616 9002 27668
rect 9646 27628 12848 27656
rect 9646 27588 9674 27628
rect 6932 27560 9674 27588
rect 9953 27591 10011 27597
rect 2682 27480 2688 27532
rect 2740 27520 2746 27532
rect 3145 27523 3203 27529
rect 3145 27520 3157 27523
rect 2740 27492 3157 27520
rect 2740 27480 2746 27492
rect 3145 27489 3157 27492
rect 3191 27520 3203 27523
rect 6932 27520 6960 27560
rect 9953 27557 9965 27591
rect 9999 27588 10011 27591
rect 10410 27588 10416 27600
rect 9999 27560 10416 27588
rect 9999 27557 10011 27560
rect 9953 27551 10011 27557
rect 10410 27548 10416 27560
rect 10468 27548 10474 27600
rect 10505 27591 10563 27597
rect 10505 27557 10517 27591
rect 10551 27557 10563 27591
rect 10505 27551 10563 27557
rect 3191 27492 6960 27520
rect 7009 27523 7067 27529
rect 3191 27489 3203 27492
rect 3145 27483 3203 27489
rect 1394 27412 1400 27464
rect 1452 27412 1458 27464
rect 4632 27461 4660 27492
rect 7009 27489 7021 27523
rect 7055 27520 7067 27523
rect 7190 27520 7196 27532
rect 7055 27492 7196 27520
rect 7055 27489 7067 27492
rect 7009 27483 7067 27489
rect 7190 27480 7196 27492
rect 7248 27480 7254 27532
rect 7466 27480 7472 27532
rect 7524 27520 7530 27532
rect 7926 27520 7932 27532
rect 7524 27492 7932 27520
rect 7524 27480 7530 27492
rect 7926 27480 7932 27492
rect 7984 27520 7990 27532
rect 8665 27523 8723 27529
rect 7984 27492 8524 27520
rect 7984 27480 7990 27492
rect 4617 27455 4675 27461
rect 4617 27421 4629 27455
rect 4663 27421 4675 27455
rect 4617 27415 4675 27421
rect 4982 27412 4988 27464
rect 5040 27452 5046 27464
rect 5442 27452 5448 27464
rect 5040 27424 5448 27452
rect 5040 27412 5046 27424
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 7745 27455 7803 27461
rect 7745 27421 7757 27455
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 8021 27455 8079 27461
rect 8021 27421 8033 27455
rect 8067 27452 8079 27455
rect 8110 27452 8116 27464
rect 8067 27424 8116 27452
rect 8067 27421 8079 27424
rect 8021 27415 8079 27421
rect 1670 27344 1676 27396
rect 1728 27344 1734 27396
rect 2898 27356 3740 27384
rect 3712 27316 3740 27356
rect 3786 27344 3792 27396
rect 3844 27344 3850 27396
rect 4798 27344 4804 27396
rect 4856 27344 4862 27396
rect 4893 27387 4951 27393
rect 4893 27353 4905 27387
rect 4939 27384 4951 27387
rect 4939 27356 5304 27384
rect 4939 27353 4951 27356
rect 4893 27347 4951 27353
rect 4062 27316 4068 27328
rect 3712 27288 4068 27316
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 5166 27276 5172 27328
rect 5224 27276 5230 27328
rect 5276 27325 5304 27356
rect 6178 27344 6184 27396
rect 6236 27344 6242 27396
rect 6454 27344 6460 27396
rect 6512 27384 6518 27396
rect 6733 27387 6791 27393
rect 6733 27384 6745 27387
rect 6512 27356 6745 27384
rect 6512 27344 6518 27356
rect 6733 27353 6745 27356
rect 6779 27353 6791 27387
rect 7760 27384 7788 27415
rect 8110 27412 8116 27424
rect 8168 27412 8174 27464
rect 8202 27412 8208 27464
rect 8260 27412 8266 27464
rect 8496 27461 8524 27492
rect 8665 27489 8677 27523
rect 8711 27520 8723 27523
rect 8754 27520 8760 27532
rect 8711 27492 8760 27520
rect 8711 27489 8723 27492
rect 8665 27483 8723 27489
rect 8754 27480 8760 27492
rect 8812 27480 8818 27532
rect 10042 27520 10048 27532
rect 9094 27492 10048 27520
rect 8481 27455 8539 27461
rect 8481 27421 8493 27455
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 8570 27412 8576 27464
rect 8628 27452 8634 27464
rect 9094 27461 9122 27492
rect 10042 27480 10048 27492
rect 10100 27480 10106 27532
rect 10520 27520 10548 27551
rect 10152 27492 10548 27520
rect 9079 27455 9137 27461
rect 9079 27452 9091 27455
rect 8628 27424 9091 27452
rect 8628 27412 8634 27424
rect 9079 27421 9091 27424
rect 9125 27421 9137 27455
rect 9079 27415 9137 27421
rect 9492 27455 9550 27461
rect 9492 27421 9504 27455
rect 9538 27421 9550 27455
rect 9492 27415 9550 27421
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27452 9643 27455
rect 9950 27452 9956 27464
rect 9631 27424 9956 27452
rect 9631 27421 9643 27424
rect 9585 27415 9643 27421
rect 9217 27387 9275 27393
rect 9217 27384 9229 27387
rect 6733 27347 6791 27353
rect 6840 27356 9229 27384
rect 5261 27319 5319 27325
rect 5261 27285 5273 27319
rect 5307 27316 5319 27319
rect 6840 27316 6868 27356
rect 9217 27353 9229 27356
rect 9263 27353 9275 27387
rect 9217 27347 9275 27353
rect 9309 27387 9367 27393
rect 9309 27353 9321 27387
rect 9355 27353 9367 27387
rect 9508 27384 9536 27415
rect 9950 27412 9956 27424
rect 10008 27412 10014 27464
rect 10152 27461 10180 27492
rect 10962 27480 10968 27532
rect 11020 27520 11026 27532
rect 11149 27523 11207 27529
rect 11149 27520 11161 27523
rect 11020 27492 11161 27520
rect 11020 27480 11026 27492
rect 11149 27489 11161 27492
rect 11195 27489 11207 27523
rect 12820 27520 12848 27628
rect 12894 27616 12900 27668
rect 12952 27656 12958 27668
rect 13173 27659 13231 27665
rect 13173 27656 13185 27659
rect 12952 27628 13185 27656
rect 12952 27616 12958 27628
rect 13173 27625 13185 27628
rect 13219 27625 13231 27659
rect 13173 27619 13231 27625
rect 15930 27616 15936 27668
rect 15988 27656 15994 27668
rect 16209 27659 16267 27665
rect 16209 27656 16221 27659
rect 15988 27628 16221 27656
rect 15988 27616 15994 27628
rect 16209 27625 16221 27628
rect 16255 27656 16267 27659
rect 16574 27656 16580 27668
rect 16255 27628 16580 27656
rect 16255 27625 16267 27628
rect 16209 27619 16267 27625
rect 16574 27616 16580 27628
rect 16632 27616 16638 27668
rect 17402 27616 17408 27668
rect 17460 27656 17466 27668
rect 18414 27656 18420 27668
rect 17460 27628 18420 27656
rect 17460 27616 17466 27628
rect 18414 27616 18420 27628
rect 18472 27616 18478 27668
rect 24854 27616 24860 27668
rect 24912 27616 24918 27668
rect 25225 27659 25283 27665
rect 25225 27625 25237 27659
rect 25271 27656 25283 27659
rect 25774 27656 25780 27668
rect 25271 27628 25780 27656
rect 25271 27625 25283 27628
rect 25225 27619 25283 27625
rect 15378 27548 15384 27600
rect 15436 27548 15442 27600
rect 16485 27591 16543 27597
rect 16485 27557 16497 27591
rect 16531 27557 16543 27591
rect 16485 27551 16543 27557
rect 15562 27520 15568 27532
rect 12820 27492 13712 27520
rect 11149 27483 11207 27489
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27421 10195 27455
rect 10137 27415 10195 27421
rect 10318 27412 10324 27464
rect 10376 27412 10382 27464
rect 10410 27412 10416 27464
rect 10468 27452 10474 27464
rect 10594 27452 10600 27464
rect 10468 27424 10600 27452
rect 10468 27412 10474 27424
rect 10594 27412 10600 27424
rect 10652 27412 10658 27464
rect 10689 27455 10747 27461
rect 10689 27421 10701 27455
rect 10735 27421 10747 27455
rect 10689 27415 10747 27421
rect 10336 27384 10364 27412
rect 9508 27356 10364 27384
rect 10704 27384 10732 27415
rect 10778 27412 10784 27464
rect 10836 27412 10842 27464
rect 11057 27455 11115 27461
rect 11057 27421 11069 27455
rect 11103 27452 11115 27455
rect 11330 27452 11336 27464
rect 11103 27424 11336 27452
rect 11103 27421 11115 27424
rect 11057 27415 11115 27421
rect 11330 27412 11336 27424
rect 11388 27452 11394 27464
rect 12345 27455 12403 27461
rect 12345 27452 12357 27455
rect 11388 27424 12357 27452
rect 11388 27412 11394 27424
rect 12345 27421 12357 27424
rect 12391 27421 12403 27455
rect 12345 27415 12403 27421
rect 12526 27412 12532 27464
rect 12584 27412 12590 27464
rect 12713 27455 12771 27461
rect 12713 27421 12725 27455
rect 12759 27421 12771 27455
rect 12713 27415 12771 27421
rect 12805 27455 12863 27461
rect 12805 27421 12817 27455
rect 12851 27421 12863 27455
rect 12805 27415 12863 27421
rect 11146 27384 11152 27396
rect 10704 27356 11152 27384
rect 9309 27347 9367 27353
rect 5307 27288 6868 27316
rect 5307 27285 5319 27288
rect 5261 27279 5319 27285
rect 7098 27276 7104 27328
rect 7156 27276 7162 27328
rect 7558 27276 7564 27328
rect 7616 27316 7622 27328
rect 8478 27316 8484 27328
rect 7616 27288 8484 27316
rect 7616 27276 7622 27288
rect 8478 27276 8484 27288
rect 8536 27276 8542 27328
rect 8846 27276 8852 27328
rect 8904 27316 8910 27328
rect 9324 27316 9352 27347
rect 11146 27344 11152 27356
rect 11204 27344 11210 27396
rect 12728 27328 12756 27415
rect 12820 27384 12848 27415
rect 12894 27412 12900 27464
rect 12952 27412 12958 27464
rect 13081 27455 13139 27461
rect 13081 27421 13093 27455
rect 13127 27452 13139 27455
rect 13170 27452 13176 27464
rect 13127 27424 13176 27452
rect 13127 27421 13139 27424
rect 13081 27415 13139 27421
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 13262 27412 13268 27464
rect 13320 27461 13326 27464
rect 13684 27461 13712 27492
rect 13832 27492 15568 27520
rect 13832 27461 13860 27492
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 16390 27480 16396 27532
rect 16448 27520 16454 27532
rect 16500 27520 16528 27551
rect 17494 27548 17500 27600
rect 17552 27548 17558 27600
rect 18322 27588 18328 27600
rect 18202 27560 18328 27588
rect 16448 27492 16528 27520
rect 16448 27480 16454 27492
rect 16574 27480 16580 27532
rect 16632 27520 16638 27532
rect 17512 27520 17540 27548
rect 18202 27520 18230 27560
rect 18322 27548 18328 27560
rect 18380 27588 18386 27600
rect 18690 27588 18696 27600
rect 18380 27560 18696 27588
rect 18380 27548 18386 27560
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 20898 27588 20904 27600
rect 19996 27560 20904 27588
rect 19702 27520 19708 27532
rect 16632 27492 17816 27520
rect 16632 27480 16638 27492
rect 13320 27455 13369 27461
rect 13320 27421 13323 27455
rect 13357 27421 13369 27455
rect 13320 27415 13369 27421
rect 13669 27455 13727 27461
rect 13669 27421 13681 27455
rect 13715 27421 13727 27455
rect 13669 27415 13727 27421
rect 13817 27455 13875 27461
rect 13817 27421 13829 27455
rect 13863 27421 13875 27455
rect 13817 27415 13875 27421
rect 13320 27412 13326 27415
rect 14734 27412 14740 27464
rect 14792 27452 14798 27464
rect 14829 27455 14887 27461
rect 14829 27452 14841 27455
rect 14792 27424 14841 27452
rect 14792 27412 14798 27424
rect 14829 27421 14841 27424
rect 14875 27421 14887 27455
rect 14829 27415 14887 27421
rect 14918 27412 14924 27464
rect 14976 27452 14982 27464
rect 16666 27461 16672 27464
rect 15197 27455 15255 27461
rect 15197 27452 15209 27455
rect 14976 27424 15209 27452
rect 14976 27412 14982 27424
rect 15197 27421 15209 27424
rect 15243 27452 15255 27455
rect 16664 27452 16672 27461
rect 15243 27424 16672 27452
rect 15243 27421 15255 27424
rect 15197 27415 15255 27421
rect 16664 27415 16672 27424
rect 16666 27412 16672 27415
rect 16724 27412 16730 27464
rect 16758 27412 16764 27464
rect 16816 27412 16822 27464
rect 16850 27412 16856 27464
rect 16908 27412 16914 27464
rect 16942 27412 16948 27464
rect 17000 27461 17006 27464
rect 17000 27455 17039 27461
rect 17027 27421 17039 27455
rect 17000 27415 17039 27421
rect 17129 27455 17187 27461
rect 17129 27421 17141 27455
rect 17175 27452 17187 27455
rect 17310 27452 17316 27464
rect 17175 27424 17316 27452
rect 17175 27421 17187 27424
rect 17129 27415 17187 27421
rect 17000 27412 17006 27415
rect 17310 27412 17316 27424
rect 17368 27412 17374 27464
rect 17402 27412 17408 27464
rect 17460 27412 17466 27464
rect 17788 27461 17816 27492
rect 18156 27492 18230 27520
rect 18524 27492 19708 27520
rect 17497 27455 17555 27461
rect 17497 27421 17509 27455
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 17681 27455 17739 27461
rect 17681 27421 17693 27455
rect 17727 27421 17739 27455
rect 17681 27415 17739 27421
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27421 17831 27455
rect 17773 27415 17831 27421
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 18046 27452 18052 27464
rect 17911 27424 18052 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 13449 27387 13507 27393
rect 13449 27384 13461 27387
rect 12820 27356 13461 27384
rect 13449 27353 13461 27356
rect 13495 27353 13507 27387
rect 13449 27347 13507 27353
rect 9398 27316 9404 27328
rect 8904 27288 9404 27316
rect 8904 27276 8910 27288
rect 9398 27276 9404 27288
rect 9456 27276 9462 27328
rect 10318 27276 10324 27328
rect 10376 27276 10382 27328
rect 12710 27276 12716 27328
rect 12768 27276 12774 27328
rect 13464 27316 13492 27347
rect 13538 27344 13544 27396
rect 13596 27344 13602 27396
rect 15010 27344 15016 27396
rect 15068 27344 15074 27396
rect 15105 27387 15163 27393
rect 15105 27353 15117 27387
rect 15151 27384 15163 27387
rect 15654 27384 15660 27396
rect 15151 27356 15660 27384
rect 15151 27353 15163 27356
rect 15105 27347 15163 27353
rect 15654 27344 15660 27356
rect 15712 27344 15718 27396
rect 15838 27344 15844 27396
rect 15896 27384 15902 27396
rect 16025 27387 16083 27393
rect 16025 27384 16037 27387
rect 15896 27356 16037 27384
rect 15896 27344 15902 27356
rect 16025 27353 16037 27356
rect 16071 27353 16083 27387
rect 17512 27384 17540 27415
rect 16025 27347 16083 27353
rect 17144 27356 17540 27384
rect 17696 27384 17724 27415
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 18156 27461 18184 27492
rect 18141 27455 18199 27461
rect 18141 27421 18153 27455
rect 18187 27421 18199 27455
rect 18141 27415 18199 27421
rect 17696 27356 17908 27384
rect 17144 27328 17172 27356
rect 17880 27328 17908 27356
rect 18230 27344 18236 27396
rect 18288 27344 18294 27396
rect 18524 27393 18552 27492
rect 19702 27480 19708 27492
rect 19760 27480 19766 27532
rect 19337 27455 19395 27461
rect 19337 27421 19349 27455
rect 19383 27421 19395 27455
rect 19337 27415 19395 27421
rect 18509 27387 18567 27393
rect 18509 27353 18521 27387
rect 18555 27353 18567 27387
rect 18509 27347 18567 27353
rect 18693 27387 18751 27393
rect 18693 27353 18705 27387
rect 18739 27384 18751 27387
rect 19242 27384 19248 27396
rect 18739 27356 19248 27384
rect 18739 27353 18751 27356
rect 18693 27347 18751 27353
rect 13630 27316 13636 27328
rect 13464 27288 13636 27316
rect 13630 27276 13636 27288
rect 13688 27276 13694 27328
rect 16206 27276 16212 27328
rect 16264 27325 16270 27328
rect 16264 27319 16283 27325
rect 16271 27285 16283 27319
rect 16264 27279 16283 27285
rect 16264 27276 16270 27279
rect 16390 27276 16396 27328
rect 16448 27276 16454 27328
rect 17126 27276 17132 27328
rect 17184 27276 17190 27328
rect 17218 27276 17224 27328
rect 17276 27276 17282 27328
rect 17862 27276 17868 27328
rect 17920 27276 17926 27328
rect 18414 27276 18420 27328
rect 18472 27316 18478 27328
rect 18708 27316 18736 27347
rect 19242 27344 19248 27356
rect 19300 27384 19306 27396
rect 19352 27384 19380 27415
rect 19426 27412 19432 27464
rect 19484 27412 19490 27464
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27421 19579 27455
rect 19797 27455 19855 27461
rect 19797 27452 19809 27455
rect 19521 27415 19579 27421
rect 19720 27424 19809 27452
rect 19300 27356 19380 27384
rect 19300 27344 19306 27356
rect 18472 27288 18736 27316
rect 18472 27276 18478 27288
rect 18874 27276 18880 27328
rect 18932 27276 18938 27328
rect 19536 27316 19564 27415
rect 19720 27396 19748 27424
rect 19797 27421 19809 27424
rect 19843 27421 19855 27455
rect 19797 27415 19855 27421
rect 19889 27455 19947 27461
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 19996 27452 20024 27560
rect 20898 27548 20904 27560
rect 20956 27548 20962 27600
rect 21174 27548 21180 27600
rect 21232 27588 21238 27600
rect 21726 27588 21732 27600
rect 21232 27560 21732 27588
rect 21232 27548 21238 27560
rect 21726 27548 21732 27560
rect 21784 27548 21790 27600
rect 23106 27588 23112 27600
rect 22066 27560 23112 27588
rect 22066 27520 22094 27560
rect 23106 27548 23112 27560
rect 23164 27588 23170 27600
rect 24121 27591 24179 27597
rect 24121 27588 24133 27591
rect 23164 27560 24133 27588
rect 23164 27548 23170 27560
rect 24121 27557 24133 27560
rect 24167 27557 24179 27591
rect 24121 27551 24179 27557
rect 24302 27548 24308 27600
rect 24360 27588 24366 27600
rect 24360 27560 24624 27588
rect 24360 27548 24366 27560
rect 23293 27523 23351 27529
rect 23293 27520 23305 27523
rect 20088 27492 22094 27520
rect 22946 27492 23305 27520
rect 20088 27461 20116 27492
rect 19935 27424 20024 27452
rect 20073 27455 20131 27461
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 20073 27421 20085 27455
rect 20119 27421 20131 27455
rect 20073 27415 20131 27421
rect 21085 27455 21143 27461
rect 21085 27421 21097 27455
rect 21131 27452 21143 27455
rect 21266 27452 21272 27464
rect 21131 27424 21272 27452
rect 21131 27421 21143 27424
rect 21085 27415 21143 27421
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21358 27412 21364 27464
rect 21416 27412 21422 27464
rect 21450 27412 21456 27464
rect 21508 27452 21514 27464
rect 21821 27455 21879 27461
rect 21821 27452 21833 27455
rect 21508 27424 21833 27452
rect 21508 27412 21514 27424
rect 21821 27421 21833 27424
rect 21867 27452 21879 27455
rect 22946 27452 22974 27492
rect 23293 27489 23305 27492
rect 23339 27520 23351 27523
rect 23474 27520 23480 27532
rect 23339 27492 23480 27520
rect 23339 27489 23351 27492
rect 23293 27483 23351 27489
rect 23474 27480 23480 27492
rect 23532 27520 23538 27532
rect 23532 27492 23796 27520
rect 23532 27480 23538 27492
rect 21867 27424 22974 27452
rect 21867 27421 21879 27424
rect 21821 27415 21879 27421
rect 23014 27412 23020 27464
rect 23072 27412 23078 27464
rect 23109 27455 23167 27461
rect 23109 27421 23121 27455
rect 23155 27452 23167 27455
rect 23382 27452 23388 27464
rect 23155 27424 23388 27452
rect 23155 27421 23167 27424
rect 23109 27415 23167 27421
rect 19702 27344 19708 27396
rect 19760 27344 19766 27396
rect 21637 27387 21695 27393
rect 19812 27356 21588 27384
rect 19812 27316 19840 27356
rect 19536 27288 19840 27316
rect 19978 27276 19984 27328
rect 20036 27316 20042 27328
rect 20257 27319 20315 27325
rect 20257 27316 20269 27319
rect 20036 27288 20269 27316
rect 20036 27276 20042 27288
rect 20257 27285 20269 27288
rect 20303 27285 20315 27319
rect 20257 27279 20315 27285
rect 20530 27276 20536 27328
rect 20588 27316 20594 27328
rect 20901 27319 20959 27325
rect 20901 27316 20913 27319
rect 20588 27288 20913 27316
rect 20588 27276 20594 27288
rect 20901 27285 20913 27288
rect 20947 27285 20959 27319
rect 20901 27279 20959 27285
rect 21269 27319 21327 27325
rect 21269 27285 21281 27319
rect 21315 27316 21327 27319
rect 21450 27316 21456 27328
rect 21315 27288 21456 27316
rect 21315 27285 21327 27288
rect 21269 27279 21327 27285
rect 21450 27276 21456 27288
rect 21508 27276 21514 27328
rect 21560 27316 21588 27356
rect 21637 27353 21649 27387
rect 21683 27384 21695 27387
rect 21726 27384 21732 27396
rect 21683 27356 21732 27384
rect 21683 27353 21695 27356
rect 21637 27347 21695 27353
rect 21726 27344 21732 27356
rect 21784 27344 21790 27396
rect 22462 27344 22468 27396
rect 22520 27384 22526 27396
rect 23124 27384 23152 27415
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 23768 27396 23796 27492
rect 24210 27480 24216 27532
rect 24268 27520 24274 27532
rect 24489 27523 24547 27529
rect 24489 27520 24501 27523
rect 24268 27492 24501 27520
rect 24268 27480 24274 27492
rect 24489 27489 24501 27492
rect 24535 27489 24547 27523
rect 24489 27483 24547 27489
rect 24596 27520 24624 27560
rect 24872 27520 24900 27616
rect 24596 27492 24801 27520
rect 24872 27492 25360 27520
rect 24026 27412 24032 27464
rect 24084 27452 24090 27464
rect 24596 27461 24624 27492
rect 24397 27455 24455 27461
rect 24397 27452 24409 27455
rect 24084 27424 24409 27452
rect 24084 27412 24090 27424
rect 24397 27421 24409 27424
rect 24443 27421 24455 27455
rect 24397 27415 24455 27421
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 24670 27412 24676 27464
rect 24728 27412 24734 27464
rect 24773 27452 24801 27492
rect 24854 27452 24860 27464
rect 24773 27424 24860 27452
rect 24854 27412 24860 27424
rect 24912 27412 24918 27464
rect 25041 27455 25099 27461
rect 25041 27421 25053 27455
rect 25087 27452 25099 27455
rect 25130 27452 25136 27464
rect 25087 27424 25136 27452
rect 25087 27421 25099 27424
rect 25041 27415 25099 27421
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25332 27461 25360 27492
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27421 25375 27455
rect 25317 27415 25375 27421
rect 22520 27356 23152 27384
rect 22520 27344 22526 27356
rect 23750 27344 23756 27396
rect 23808 27344 23814 27396
rect 24118 27344 24124 27396
rect 24176 27344 24182 27396
rect 25424 27384 25452 27628
rect 25774 27616 25780 27628
rect 25832 27616 25838 27668
rect 26878 27616 26884 27668
rect 26936 27616 26942 27668
rect 28166 27616 28172 27668
rect 28224 27656 28230 27668
rect 28365 27659 28423 27665
rect 28365 27656 28377 27659
rect 28224 27628 28377 27656
rect 28224 27616 28230 27628
rect 28365 27625 28377 27628
rect 28411 27625 28423 27659
rect 28365 27619 28423 27625
rect 29181 27659 29239 27665
rect 29181 27625 29193 27659
rect 29227 27656 29239 27659
rect 29546 27656 29552 27668
rect 29227 27628 29552 27656
rect 29227 27625 29239 27628
rect 29181 27619 29239 27625
rect 29546 27616 29552 27628
rect 29604 27656 29610 27668
rect 29822 27656 29828 27668
rect 29604 27628 29828 27656
rect 29604 27616 29610 27628
rect 29822 27616 29828 27628
rect 29880 27616 29886 27668
rect 30098 27616 30104 27668
rect 30156 27656 30162 27668
rect 30193 27659 30251 27665
rect 30193 27656 30205 27659
rect 30156 27628 30205 27656
rect 30156 27616 30162 27628
rect 30193 27625 30205 27628
rect 30239 27625 30251 27659
rect 30742 27656 30748 27668
rect 30193 27619 30251 27625
rect 30484 27628 30748 27656
rect 30374 27588 30380 27600
rect 28552 27560 28764 27588
rect 28258 27480 28264 27532
rect 28316 27520 28322 27532
rect 28552 27520 28580 27560
rect 28316 27492 28580 27520
rect 28316 27480 28322 27492
rect 28626 27480 28632 27532
rect 28684 27480 28690 27532
rect 28736 27520 28764 27560
rect 29656 27560 30380 27588
rect 29656 27520 29684 27560
rect 30116 27529 30144 27560
rect 30374 27548 30380 27560
rect 30432 27548 30438 27600
rect 28736 27492 29684 27520
rect 30101 27523 30159 27529
rect 30101 27489 30113 27523
rect 30147 27489 30159 27523
rect 30484 27520 30512 27628
rect 30742 27616 30748 27628
rect 30800 27616 30806 27668
rect 31846 27616 31852 27668
rect 31904 27656 31910 27668
rect 32122 27656 32128 27668
rect 31904 27628 32128 27656
rect 31904 27616 31910 27628
rect 32122 27616 32128 27628
rect 32180 27616 32186 27668
rect 33962 27616 33968 27668
rect 34020 27656 34026 27668
rect 34020 27628 34284 27656
rect 34020 27616 34026 27628
rect 32306 27588 32312 27600
rect 30101 27483 30159 27489
rect 30392 27492 30512 27520
rect 30668 27560 32312 27588
rect 30392 27464 30420 27492
rect 25498 27412 25504 27464
rect 25556 27412 25562 27464
rect 26786 27452 26792 27464
rect 25608 27424 26792 27452
rect 24412 27356 25452 27384
rect 22278 27316 22284 27328
rect 21560 27288 22284 27316
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 22738 27276 22744 27328
rect 22796 27316 22802 27328
rect 23293 27319 23351 27325
rect 23293 27316 23305 27319
rect 22796 27288 23305 27316
rect 22796 27276 22802 27288
rect 23293 27285 23305 27288
rect 23339 27285 23351 27319
rect 23293 27279 23351 27285
rect 23382 27276 23388 27328
rect 23440 27276 23446 27328
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 23569 27319 23627 27325
rect 23569 27316 23581 27319
rect 23532 27288 23581 27316
rect 23532 27276 23538 27288
rect 23569 27285 23581 27288
rect 23615 27285 23627 27319
rect 23569 27279 23627 27285
rect 23661 27319 23719 27325
rect 23661 27285 23673 27319
rect 23707 27316 23719 27319
rect 24412 27316 24440 27356
rect 23707 27288 24440 27316
rect 23707 27285 23719 27288
rect 23661 27279 23719 27285
rect 24762 27276 24768 27328
rect 24820 27316 24826 27328
rect 25608 27316 25636 27424
rect 26786 27412 26792 27424
rect 26844 27412 26850 27464
rect 29825 27455 29883 27461
rect 29217 27424 29684 27452
rect 29217 27421 29285 27424
rect 25774 27344 25780 27396
rect 25832 27384 25838 27396
rect 25869 27387 25927 27393
rect 25869 27384 25881 27387
rect 25832 27356 25881 27384
rect 25832 27344 25838 27356
rect 25869 27353 25881 27356
rect 25915 27353 25927 27387
rect 25869 27347 25927 27353
rect 26050 27344 26056 27396
rect 26108 27344 26114 27396
rect 27062 27344 27068 27396
rect 27120 27384 27126 27396
rect 27120 27356 27186 27384
rect 27120 27344 27126 27356
rect 28994 27344 29000 27396
rect 29052 27344 29058 27396
rect 29217 27390 29239 27421
rect 29227 27387 29239 27390
rect 29273 27387 29285 27421
rect 29227 27381 29285 27387
rect 24820 27288 25636 27316
rect 24820 27276 24826 27288
rect 25682 27276 25688 27328
rect 25740 27276 25746 27328
rect 26234 27276 26240 27328
rect 26292 27276 26298 27328
rect 27430 27276 27436 27328
rect 27488 27316 27494 27328
rect 29012 27316 29040 27344
rect 27488 27288 29040 27316
rect 27488 27276 27494 27288
rect 29270 27276 29276 27328
rect 29328 27316 29334 27328
rect 29365 27319 29423 27325
rect 29365 27316 29377 27319
rect 29328 27288 29377 27316
rect 29328 27276 29334 27288
rect 29365 27285 29377 27288
rect 29411 27285 29423 27319
rect 29365 27279 29423 27285
rect 29454 27276 29460 27328
rect 29512 27316 29518 27328
rect 29549 27319 29607 27325
rect 29549 27316 29561 27319
rect 29512 27288 29561 27316
rect 29512 27276 29518 27288
rect 29549 27285 29561 27288
rect 29595 27285 29607 27319
rect 29656 27316 29684 27424
rect 29825 27421 29837 27455
rect 29871 27452 29883 27455
rect 29871 27424 30328 27452
rect 29871 27421 29883 27424
rect 29825 27415 29883 27421
rect 30300 27396 30328 27424
rect 30374 27412 30380 27464
rect 30432 27412 30438 27464
rect 30668 27461 30696 27560
rect 32306 27548 32312 27560
rect 32364 27548 32370 27600
rect 31478 27520 31484 27532
rect 31036 27492 31484 27520
rect 30469 27455 30527 27461
rect 30469 27421 30481 27455
rect 30515 27421 30527 27455
rect 30469 27415 30527 27421
rect 30653 27455 30711 27461
rect 30653 27421 30665 27455
rect 30699 27421 30711 27455
rect 30653 27415 30711 27421
rect 30745 27455 30803 27461
rect 30745 27421 30757 27455
rect 30791 27452 30803 27455
rect 30926 27452 30932 27464
rect 30791 27424 30932 27452
rect 30791 27421 30803 27424
rect 30745 27415 30803 27421
rect 29730 27344 29736 27396
rect 29788 27344 29794 27396
rect 29914 27344 29920 27396
rect 29972 27344 29978 27396
rect 30282 27344 30288 27396
rect 30340 27384 30346 27396
rect 30484 27384 30512 27415
rect 30926 27412 30932 27424
rect 30984 27412 30990 27464
rect 31036 27461 31064 27492
rect 31478 27480 31484 27492
rect 31536 27520 31542 27532
rect 33134 27520 33140 27532
rect 31536 27492 33140 27520
rect 31536 27480 31542 27492
rect 31021 27455 31079 27461
rect 31021 27421 31033 27455
rect 31067 27421 31079 27455
rect 31021 27415 31079 27421
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27452 31263 27455
rect 31754 27452 31760 27464
rect 31251 27424 31760 27452
rect 31251 27421 31263 27424
rect 31205 27415 31263 27421
rect 31754 27412 31760 27424
rect 31812 27412 31818 27464
rect 31846 27412 31852 27464
rect 31904 27412 31910 27464
rect 31956 27461 31984 27492
rect 33134 27480 33140 27492
rect 33192 27480 33198 27532
rect 34256 27529 34284 27628
rect 34330 27616 34336 27668
rect 34388 27616 34394 27668
rect 34422 27616 34428 27668
rect 34480 27656 34486 27668
rect 34977 27659 35035 27665
rect 34977 27656 34989 27659
rect 34480 27628 34989 27656
rect 34480 27616 34486 27628
rect 34977 27625 34989 27628
rect 35023 27625 35035 27659
rect 34977 27619 35035 27625
rect 35342 27616 35348 27668
rect 35400 27656 35406 27668
rect 35989 27659 36047 27665
rect 35989 27656 36001 27659
rect 35400 27628 36001 27656
rect 35400 27616 35406 27628
rect 35989 27625 36001 27628
rect 36035 27625 36047 27659
rect 35989 27619 36047 27625
rect 34348 27588 34376 27616
rect 34348 27560 34468 27588
rect 34241 27523 34299 27529
rect 34241 27489 34253 27523
rect 34287 27489 34299 27523
rect 34241 27483 34299 27489
rect 34330 27480 34336 27532
rect 34388 27480 34394 27532
rect 31956 27455 32019 27461
rect 31956 27424 31973 27455
rect 31961 27421 31973 27424
rect 32007 27421 32019 27455
rect 31961 27415 32019 27421
rect 34054 27412 34060 27464
rect 34112 27412 34118 27464
rect 34149 27455 34207 27461
rect 34149 27421 34161 27455
rect 34195 27452 34207 27455
rect 34440 27452 34468 27560
rect 34517 27523 34575 27529
rect 34517 27489 34529 27523
rect 34563 27489 34575 27523
rect 34517 27483 34575 27489
rect 34195 27424 34468 27452
rect 34532 27452 34560 27483
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 34532 27424 34713 27452
rect 34195 27421 34207 27424
rect 34149 27415 34207 27421
rect 34701 27421 34713 27424
rect 34747 27421 34759 27455
rect 34701 27415 34759 27421
rect 35161 27455 35219 27461
rect 35161 27421 35173 27455
rect 35207 27421 35219 27455
rect 35161 27415 35219 27421
rect 30340 27356 30512 27384
rect 30340 27344 30346 27356
rect 31662 27344 31668 27396
rect 31720 27344 31726 27396
rect 32217 27387 32275 27393
rect 32217 27384 32229 27387
rect 31864 27356 32229 27384
rect 30558 27316 30564 27328
rect 29656 27288 30564 27316
rect 29549 27279 29607 27285
rect 30558 27276 30564 27288
rect 30616 27316 30622 27328
rect 30929 27319 30987 27325
rect 30929 27316 30941 27319
rect 30616 27288 30941 27316
rect 30616 27276 30622 27288
rect 30929 27285 30941 27288
rect 30975 27285 30987 27319
rect 30929 27279 30987 27285
rect 31478 27276 31484 27328
rect 31536 27316 31542 27328
rect 31864 27316 31892 27356
rect 32217 27353 32229 27356
rect 32263 27353 32275 27387
rect 32217 27347 32275 27353
rect 32766 27344 32772 27396
rect 32824 27384 32830 27396
rect 35176 27384 35204 27415
rect 35250 27412 35256 27464
rect 35308 27412 35314 27464
rect 35342 27412 35348 27464
rect 35400 27452 35406 27464
rect 35437 27455 35495 27461
rect 35437 27452 35449 27455
rect 35400 27424 35449 27452
rect 35400 27412 35406 27424
rect 35437 27421 35449 27424
rect 35483 27421 35495 27455
rect 35437 27415 35495 27421
rect 35529 27455 35587 27461
rect 35529 27421 35541 27455
rect 35575 27452 35587 27455
rect 35986 27452 35992 27464
rect 35575 27424 35992 27452
rect 35575 27421 35587 27424
rect 35529 27415 35587 27421
rect 35986 27412 35992 27424
rect 36044 27412 36050 27464
rect 36173 27455 36231 27461
rect 36173 27421 36185 27455
rect 36219 27452 36231 27455
rect 36262 27452 36268 27464
rect 36219 27424 36268 27452
rect 36219 27421 36231 27424
rect 36173 27415 36231 27421
rect 36262 27412 36268 27424
rect 36320 27412 36326 27464
rect 36078 27384 36084 27396
rect 32824 27356 36084 27384
rect 32824 27344 32830 27356
rect 36078 27344 36084 27356
rect 36136 27344 36142 27396
rect 31536 27288 31892 27316
rect 31536 27276 31542 27288
rect 32030 27276 32036 27328
rect 32088 27276 32094 27328
rect 33594 27276 33600 27328
rect 33652 27316 33658 27328
rect 34330 27316 34336 27328
rect 33652 27288 34336 27316
rect 33652 27276 33658 27288
rect 34330 27276 34336 27288
rect 34388 27276 34394 27328
rect 34793 27319 34851 27325
rect 34793 27285 34805 27319
rect 34839 27316 34851 27319
rect 35250 27316 35256 27328
rect 34839 27288 35256 27316
rect 34839 27285 34851 27288
rect 34793 27279 34851 27285
rect 35250 27276 35256 27288
rect 35308 27276 35314 27328
rect 1104 27226 36524 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 36524 27226
rect 1104 27152 36524 27174
rect 1670 27072 1676 27124
rect 1728 27112 1734 27124
rect 2225 27115 2283 27121
rect 2225 27112 2237 27115
rect 1728 27084 2237 27112
rect 1728 27072 1734 27084
rect 2225 27081 2237 27084
rect 2271 27081 2283 27115
rect 2225 27075 2283 27081
rect 2682 27072 2688 27124
rect 2740 27072 2746 27124
rect 3694 27112 3700 27124
rect 3160 27084 3700 27112
rect 2593 27047 2651 27053
rect 2593 27013 2605 27047
rect 2639 27044 2651 27047
rect 3160 27044 3188 27084
rect 3694 27072 3700 27084
rect 3752 27072 3758 27124
rect 4798 27072 4804 27124
rect 4856 27112 4862 27124
rect 5810 27112 5816 27124
rect 4856 27084 5816 27112
rect 4856 27072 4862 27084
rect 5810 27072 5816 27084
rect 5868 27072 5874 27124
rect 6365 27115 6423 27121
rect 6365 27081 6377 27115
rect 6411 27112 6423 27115
rect 6454 27112 6460 27124
rect 6411 27084 6460 27112
rect 6411 27081 6423 27084
rect 6365 27075 6423 27081
rect 6454 27072 6460 27084
rect 6512 27072 6518 27124
rect 6733 27115 6791 27121
rect 6733 27081 6745 27115
rect 6779 27112 6791 27115
rect 7098 27112 7104 27124
rect 6779 27084 7104 27112
rect 6779 27081 6791 27084
rect 6733 27075 6791 27081
rect 7098 27072 7104 27084
rect 7156 27072 7162 27124
rect 7558 27072 7564 27124
rect 7616 27072 7622 27124
rect 8018 27072 8024 27124
rect 8076 27112 8082 27124
rect 8076 27084 8524 27112
rect 8076 27072 8082 27084
rect 3786 27044 3792 27056
rect 2639 27016 3188 27044
rect 3252 27016 3792 27044
rect 2639 27013 2651 27016
rect 2593 27007 2651 27013
rect 3252 26985 3280 27016
rect 3786 27004 3792 27016
rect 3844 27004 3850 27056
rect 4062 27004 4068 27056
rect 4120 27004 4126 27056
rect 8496 27053 8524 27084
rect 8679 27084 10088 27112
rect 8389 27047 8447 27053
rect 8389 27044 8401 27047
rect 5828 27016 8401 27044
rect 5828 26985 5856 27016
rect 8389 27013 8401 27016
rect 8435 27013 8447 27047
rect 8389 27007 8447 27013
rect 8481 27047 8539 27053
rect 8481 27013 8493 27047
rect 8527 27013 8539 27047
rect 8481 27007 8539 27013
rect 3237 26979 3295 26985
rect 3237 26945 3249 26979
rect 3283 26945 3295 26979
rect 3237 26939 3295 26945
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26976 5871 26979
rect 5902 26976 5908 26988
rect 5859 26948 5908 26976
rect 5859 26945 5871 26948
rect 5813 26939 5871 26945
rect 2869 26911 2927 26917
rect 2869 26877 2881 26911
rect 2915 26908 2927 26911
rect 3050 26908 3056 26920
rect 2915 26880 3056 26908
rect 2915 26877 2927 26880
rect 2869 26871 2927 26877
rect 3050 26868 3056 26880
rect 3108 26868 3114 26920
rect 1394 26800 1400 26852
rect 1452 26840 1458 26852
rect 3252 26840 3280 26939
rect 3513 26911 3571 26917
rect 3513 26877 3525 26911
rect 3559 26908 3571 26911
rect 4798 26908 4804 26920
rect 3559 26880 4804 26908
rect 3559 26877 3571 26880
rect 3513 26871 3571 26877
rect 4798 26868 4804 26880
rect 4856 26868 4862 26920
rect 4985 26911 5043 26917
rect 4985 26877 4997 26911
rect 5031 26908 5043 26911
rect 5828 26908 5856 26939
rect 5902 26936 5908 26948
rect 5960 26936 5966 26988
rect 6178 26936 6184 26988
rect 6236 26976 6242 26988
rect 7098 26976 7104 26988
rect 6236 26948 7104 26976
rect 6236 26936 6242 26948
rect 7098 26936 7104 26948
rect 7156 26936 7162 26988
rect 7466 26936 7472 26988
rect 7524 26936 7530 26988
rect 7742 26936 7748 26988
rect 7800 26976 7806 26988
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 7800 26948 7849 26976
rect 7800 26936 7806 26948
rect 7837 26945 7849 26948
rect 7883 26945 7895 26979
rect 8251 26979 8309 26985
rect 8251 26976 8263 26979
rect 7837 26939 7895 26945
rect 7944 26948 8263 26976
rect 6822 26908 6828 26920
rect 5031 26880 5856 26908
rect 5920 26880 6828 26908
rect 5031 26877 5043 26880
rect 4985 26871 5043 26877
rect 5920 26840 5948 26880
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7009 26911 7067 26917
rect 7009 26877 7021 26911
rect 7055 26877 7067 26911
rect 7009 26871 7067 26877
rect 1452 26812 3280 26840
rect 5092 26812 5948 26840
rect 1452 26800 1458 26812
rect 3694 26732 3700 26784
rect 3752 26772 3758 26784
rect 5092 26772 5120 26812
rect 6270 26800 6276 26852
rect 6328 26840 6334 26852
rect 7024 26840 7052 26871
rect 7650 26868 7656 26920
rect 7708 26908 7714 26920
rect 7944 26908 7972 26948
rect 8251 26945 8263 26948
rect 8297 26976 8309 26979
rect 8570 26976 8576 26988
rect 8297 26948 8576 26976
rect 8297 26945 8309 26948
rect 8251 26939 8309 26945
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 8679 26985 8707 27084
rect 8664 26979 8722 26985
rect 8664 26945 8676 26979
rect 8710 26945 8722 26979
rect 8664 26939 8722 26945
rect 8754 26936 8760 26988
rect 8812 26976 8818 26988
rect 9950 26976 9956 26988
rect 8812 26948 9956 26976
rect 8812 26936 8818 26948
rect 9950 26936 9956 26948
rect 10008 26936 10014 26988
rect 7708 26880 7972 26908
rect 8021 26911 8079 26917
rect 7708 26868 7714 26880
rect 8021 26877 8033 26911
rect 8067 26908 8079 26911
rect 8772 26908 8800 26936
rect 8067 26880 8800 26908
rect 8067 26877 8079 26880
rect 8021 26871 8079 26877
rect 6328 26812 7052 26840
rect 6328 26800 6334 26812
rect 3752 26744 5120 26772
rect 3752 26732 3758 26744
rect 5166 26732 5172 26784
rect 5224 26732 5230 26784
rect 8018 26732 8024 26784
rect 8076 26772 8082 26784
rect 8113 26775 8171 26781
rect 8113 26772 8125 26775
rect 8076 26744 8125 26772
rect 8076 26732 8082 26744
rect 8113 26741 8125 26744
rect 8159 26741 8171 26775
rect 8113 26735 8171 26741
rect 8846 26732 8852 26784
rect 8904 26772 8910 26784
rect 9953 26775 10011 26781
rect 9953 26772 9965 26775
rect 8904 26744 9965 26772
rect 8904 26732 8910 26744
rect 9953 26741 9965 26744
rect 9999 26741 10011 26775
rect 10060 26772 10088 27084
rect 10686 27072 10692 27124
rect 10744 27112 10750 27124
rect 10870 27112 10876 27124
rect 10744 27084 10876 27112
rect 10744 27072 10750 27084
rect 10870 27072 10876 27084
rect 10928 27112 10934 27124
rect 12437 27115 12495 27121
rect 10928 27084 11284 27112
rect 10928 27072 10934 27084
rect 10318 27004 10324 27056
rect 10376 27044 10382 27056
rect 11256 27053 11284 27084
rect 12437 27081 12449 27115
rect 12483 27112 12495 27115
rect 12710 27112 12716 27124
rect 12483 27084 12716 27112
rect 12483 27081 12495 27084
rect 12437 27075 12495 27081
rect 12710 27072 12716 27084
rect 12768 27072 12774 27124
rect 13906 27112 13912 27124
rect 13096 27084 13912 27112
rect 10413 27047 10471 27053
rect 10413 27044 10425 27047
rect 10376 27016 10425 27044
rect 10376 27004 10382 27016
rect 10413 27013 10425 27016
rect 10459 27044 10471 27047
rect 11241 27047 11299 27053
rect 10459 27016 10640 27044
rect 10459 27013 10471 27016
rect 10413 27007 10471 27013
rect 10226 26936 10232 26988
rect 10284 26976 10290 26988
rect 10505 26979 10563 26985
rect 10505 26976 10517 26979
rect 10284 26948 10517 26976
rect 10284 26936 10290 26948
rect 10505 26945 10517 26948
rect 10551 26945 10563 26979
rect 10505 26939 10563 26945
rect 10413 26911 10471 26917
rect 10413 26877 10425 26911
rect 10459 26877 10471 26911
rect 10612 26908 10640 27016
rect 11241 27013 11253 27047
rect 11287 27013 11299 27047
rect 11241 27007 11299 27013
rect 11330 27004 11336 27056
rect 11388 27004 11394 27056
rect 12728 27044 12756 27072
rect 12728 27016 13032 27044
rect 10686 26936 10692 26988
rect 10744 26976 10750 26988
rect 10873 26979 10931 26985
rect 10873 26976 10885 26979
rect 10744 26948 10885 26976
rect 10744 26936 10750 26948
rect 10873 26945 10885 26948
rect 10919 26945 10931 26979
rect 10873 26939 10931 26945
rect 10965 26979 11023 26985
rect 10965 26945 10977 26979
rect 11011 26976 11023 26979
rect 11146 26976 11152 26988
rect 11011 26948 11152 26976
rect 11011 26945 11023 26948
rect 10965 26939 11023 26945
rect 11146 26936 11152 26948
rect 11204 26936 11210 26988
rect 12158 26936 12164 26988
rect 12216 26976 12222 26988
rect 12253 26979 12311 26985
rect 12253 26976 12265 26979
rect 12216 26948 12265 26976
rect 12216 26936 12222 26948
rect 12253 26945 12265 26948
rect 12299 26945 12311 26979
rect 12253 26939 12311 26945
rect 12526 26936 12532 26988
rect 12584 26936 12590 26988
rect 12802 26936 12808 26988
rect 12860 26936 12866 26988
rect 13004 26985 13032 27016
rect 12989 26979 13047 26985
rect 12989 26945 13001 26979
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 13096 26917 13124 27084
rect 13906 27072 13912 27084
rect 13964 27072 13970 27124
rect 14090 27072 14096 27124
rect 14148 27112 14154 27124
rect 18046 27112 18052 27124
rect 14148 27084 18052 27112
rect 14148 27072 14154 27084
rect 18046 27072 18052 27084
rect 18104 27072 18110 27124
rect 21450 27072 21456 27124
rect 21508 27112 21514 27124
rect 21979 27115 22037 27121
rect 21979 27112 21991 27115
rect 21508 27084 21991 27112
rect 21508 27072 21514 27084
rect 21979 27081 21991 27084
rect 22025 27081 22037 27115
rect 22462 27112 22468 27124
rect 21979 27075 22037 27081
rect 22204 27084 22468 27112
rect 13817 27047 13875 27053
rect 13817 27013 13829 27047
rect 13863 27044 13875 27047
rect 13924 27044 13952 27072
rect 13863 27016 13952 27044
rect 17957 27047 18015 27053
rect 13863 27013 13875 27016
rect 13817 27007 13875 27013
rect 17957 27013 17969 27047
rect 18003 27044 18015 27047
rect 18506 27044 18512 27056
rect 18003 27016 18512 27044
rect 18003 27013 18015 27016
rect 17957 27007 18015 27013
rect 18506 27004 18512 27016
rect 18564 27004 18570 27056
rect 19242 27004 19248 27056
rect 19300 27044 19306 27056
rect 19300 27016 21496 27044
rect 19300 27004 19306 27016
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13081 26911 13139 26917
rect 10612 26880 10824 26908
rect 10413 26871 10471 26877
rect 10428 26840 10456 26871
rect 10689 26843 10747 26849
rect 10689 26840 10701 26843
rect 10428 26812 10701 26840
rect 10689 26809 10701 26812
rect 10735 26809 10747 26843
rect 10796 26840 10824 26880
rect 13081 26877 13093 26911
rect 13127 26877 13139 26911
rect 13081 26871 13139 26877
rect 11330 26840 11336 26852
rect 10796 26812 11336 26840
rect 10689 26803 10747 26809
rect 11330 26800 11336 26812
rect 11388 26800 11394 26852
rect 12161 26843 12219 26849
rect 12161 26809 12173 26843
rect 12207 26840 12219 26843
rect 12894 26840 12900 26852
rect 12207 26812 12900 26840
rect 12207 26809 12219 26812
rect 12161 26803 12219 26809
rect 12894 26800 12900 26812
rect 12952 26840 12958 26852
rect 13188 26840 13216 26939
rect 13262 26936 13268 26988
rect 13320 26976 13326 26988
rect 13357 26979 13415 26985
rect 13357 26976 13369 26979
rect 13320 26948 13369 26976
rect 13320 26936 13326 26948
rect 13357 26945 13369 26948
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 13449 26939 13507 26945
rect 12952 26812 13216 26840
rect 13372 26840 13400 26939
rect 13464 26908 13492 26939
rect 13538 26936 13544 26988
rect 13596 26936 13602 26988
rect 13630 26936 13636 26988
rect 13688 26976 13694 26988
rect 13725 26979 13783 26985
rect 13725 26976 13737 26979
rect 13688 26948 13737 26976
rect 13688 26936 13694 26948
rect 13725 26945 13737 26948
rect 13771 26945 13783 26979
rect 13725 26939 13783 26945
rect 13906 26936 13912 26988
rect 13964 26985 13970 26988
rect 13964 26976 13972 26985
rect 13964 26948 14009 26976
rect 13964 26939 13972 26948
rect 13964 26936 13970 26939
rect 15746 26936 15752 26988
rect 15804 26976 15810 26988
rect 16206 26976 16212 26988
rect 15804 26948 16212 26976
rect 15804 26936 15810 26948
rect 16206 26936 16212 26948
rect 16264 26936 16270 26988
rect 16666 26936 16672 26988
rect 16724 26976 16730 26988
rect 17402 26976 17408 26988
rect 16724 26948 17408 26976
rect 16724 26936 16730 26948
rect 17402 26936 17408 26948
rect 17460 26936 17466 26988
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26976 18291 26979
rect 18322 26976 18328 26988
rect 18279 26948 18328 26976
rect 18279 26945 18291 26948
rect 18233 26939 18291 26945
rect 18322 26936 18328 26948
rect 18380 26976 18386 26988
rect 19518 26976 19524 26988
rect 18380 26948 19524 26976
rect 18380 26936 18386 26948
rect 19518 26936 19524 26948
rect 19576 26936 19582 26988
rect 19702 26936 19708 26988
rect 19760 26936 19766 26988
rect 19886 26936 19892 26988
rect 19944 26976 19950 26988
rect 20257 26979 20315 26985
rect 20257 26976 20269 26979
rect 19944 26948 20269 26976
rect 19944 26936 19950 26948
rect 20257 26945 20269 26948
rect 20303 26945 20315 26979
rect 20257 26939 20315 26945
rect 20438 26936 20444 26988
rect 20496 26936 20502 26988
rect 20898 26936 20904 26988
rect 20956 26936 20962 26988
rect 21082 26936 21088 26988
rect 21140 26976 21146 26988
rect 21361 26979 21419 26985
rect 21361 26976 21373 26979
rect 21140 26948 21373 26976
rect 21140 26936 21146 26948
rect 21361 26945 21373 26948
rect 21407 26945 21419 26979
rect 21361 26939 21419 26945
rect 14458 26908 14464 26920
rect 13464 26880 14464 26908
rect 14458 26868 14464 26880
rect 14516 26908 14522 26920
rect 15010 26908 15016 26920
rect 14516 26880 15016 26908
rect 14516 26868 14522 26880
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 16482 26868 16488 26920
rect 16540 26908 16546 26920
rect 17770 26908 17776 26920
rect 16540 26880 17776 26908
rect 16540 26868 16546 26880
rect 17770 26868 17776 26880
rect 17828 26868 17834 26920
rect 17972 26880 18276 26908
rect 13372 26812 14228 26840
rect 12952 26800 12958 26812
rect 11054 26772 11060 26784
rect 10060 26744 11060 26772
rect 9953 26735 10011 26741
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 12621 26775 12679 26781
rect 12621 26772 12633 26775
rect 11296 26744 12633 26772
rect 11296 26732 11302 26744
rect 12621 26741 12633 26744
rect 12667 26741 12679 26775
rect 12621 26735 12679 26741
rect 12802 26732 12808 26784
rect 12860 26772 12866 26784
rect 13906 26772 13912 26784
rect 12860 26744 13912 26772
rect 12860 26732 12866 26744
rect 13906 26732 13912 26744
rect 13964 26732 13970 26784
rect 14090 26732 14096 26784
rect 14148 26732 14154 26784
rect 14200 26772 14228 26812
rect 14366 26800 14372 26852
rect 14424 26840 14430 26852
rect 17972 26840 18000 26880
rect 18248 26852 18276 26880
rect 14424 26812 18000 26840
rect 14424 26800 14430 26812
rect 18138 26800 18144 26852
rect 18196 26800 18202 26852
rect 18230 26800 18236 26852
rect 18288 26800 18294 26852
rect 20070 26800 20076 26852
rect 20128 26800 20134 26852
rect 21376 26840 21404 26939
rect 21468 26908 21496 27016
rect 21542 27004 21548 27056
rect 21600 27044 21606 27056
rect 22204 27053 22232 27084
rect 22462 27072 22468 27084
rect 22520 27072 22526 27124
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 24026 27112 24032 27124
rect 23532 27084 24032 27112
rect 23532 27072 23538 27084
rect 24026 27072 24032 27084
rect 24084 27072 24090 27124
rect 24210 27072 24216 27124
rect 24268 27112 24274 27124
rect 24486 27112 24492 27124
rect 24268 27084 24492 27112
rect 24268 27072 24274 27084
rect 24486 27072 24492 27084
rect 24544 27072 24550 27124
rect 25958 27072 25964 27124
rect 26016 27072 26022 27124
rect 28350 27072 28356 27124
rect 28408 27112 28414 27124
rect 28445 27115 28503 27121
rect 28445 27112 28457 27115
rect 28408 27084 28457 27112
rect 28408 27072 28414 27084
rect 28445 27081 28457 27084
rect 28491 27112 28503 27115
rect 28902 27112 28908 27124
rect 28491 27084 28908 27112
rect 28491 27081 28503 27084
rect 28445 27075 28503 27081
rect 28902 27072 28908 27084
rect 28960 27072 28966 27124
rect 28994 27072 29000 27124
rect 29052 27112 29058 27124
rect 29362 27112 29368 27124
rect 29052 27084 29368 27112
rect 29052 27072 29058 27084
rect 29362 27072 29368 27084
rect 29420 27112 29426 27124
rect 29420 27084 31248 27112
rect 29420 27072 29426 27084
rect 22189 27047 22247 27053
rect 22189 27044 22201 27047
rect 21600 27016 22201 27044
rect 21600 27004 21606 27016
rect 22189 27013 22201 27016
rect 22235 27013 22247 27047
rect 22189 27007 22247 27013
rect 22738 27004 22744 27056
rect 22796 27044 22802 27056
rect 23661 27047 23719 27053
rect 23661 27044 23673 27047
rect 22796 27016 23673 27044
rect 22796 27004 22802 27016
rect 23661 27013 23673 27016
rect 23707 27013 23719 27047
rect 24578 27044 24584 27056
rect 23661 27007 23719 27013
rect 23768 27016 24584 27044
rect 22278 26936 22284 26988
rect 22336 26936 22342 26988
rect 23768 26976 23796 27016
rect 24578 27004 24584 27016
rect 24636 27044 24642 27056
rect 24636 27016 25084 27044
rect 24636 27004 24642 27016
rect 22388 26948 23796 26976
rect 23845 26979 23903 26985
rect 22388 26917 22416 26948
rect 23845 26945 23857 26979
rect 23891 26976 23903 26979
rect 24210 26976 24216 26988
rect 23891 26948 24216 26976
rect 23891 26945 23903 26948
rect 23845 26939 23903 26945
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24302 26936 24308 26988
rect 24360 26976 24366 26988
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24360 26948 24409 26976
rect 24360 26936 24366 26948
rect 24397 26945 24409 26948
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 24670 26936 24676 26988
rect 24728 26936 24734 26988
rect 25056 26985 25084 27016
rect 25130 27004 25136 27056
rect 25188 27044 25194 27056
rect 26326 27044 26332 27056
rect 25188 27016 26332 27044
rect 25188 27004 25194 27016
rect 26326 27004 26332 27016
rect 26384 27044 26390 27056
rect 26421 27047 26479 27053
rect 26421 27044 26433 27047
rect 26384 27016 26433 27044
rect 26384 27004 26390 27016
rect 26421 27013 26433 27016
rect 26467 27044 26479 27047
rect 26970 27044 26976 27056
rect 26467 27016 26976 27044
rect 26467 27013 26479 27016
rect 26421 27007 26479 27013
rect 26970 27004 26976 27016
rect 27028 27004 27034 27056
rect 30098 27044 30104 27056
rect 28368 27016 30104 27044
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 26786 26936 26792 26988
rect 26844 26936 26850 26988
rect 28258 26936 28264 26988
rect 28316 26976 28322 26988
rect 28368 26985 28396 27016
rect 30098 27004 30104 27016
rect 30156 27044 30162 27056
rect 30576 27053 30604 27084
rect 30377 27047 30435 27053
rect 30377 27044 30389 27047
rect 30156 27016 30389 27044
rect 30156 27004 30162 27016
rect 30377 27013 30389 27016
rect 30423 27013 30435 27047
rect 30377 27007 30435 27013
rect 30561 27047 30619 27053
rect 30561 27013 30573 27047
rect 30607 27013 30619 27047
rect 30561 27007 30619 27013
rect 30650 27004 30656 27056
rect 30708 27044 30714 27056
rect 31113 27047 31171 27053
rect 31113 27044 31125 27047
rect 30708 27016 31125 27044
rect 30708 27004 30714 27016
rect 31113 27013 31125 27016
rect 31159 27013 31171 27047
rect 31113 27007 31171 27013
rect 28353 26979 28411 26985
rect 28353 26976 28365 26979
rect 28316 26948 28365 26976
rect 28316 26936 28322 26948
rect 28353 26945 28365 26948
rect 28399 26945 28411 26979
rect 28353 26939 28411 26945
rect 28537 26979 28595 26985
rect 28537 26945 28549 26979
rect 28583 26976 28595 26979
rect 28994 26976 29000 26988
rect 28583 26948 29000 26976
rect 28583 26945 28595 26948
rect 28537 26939 28595 26945
rect 28994 26936 29000 26948
rect 29052 26936 29058 26988
rect 29454 26936 29460 26988
rect 29512 26976 29518 26988
rect 29917 26979 29975 26985
rect 29917 26976 29929 26979
rect 29512 26948 29929 26976
rect 29512 26936 29518 26948
rect 29917 26945 29929 26948
rect 29963 26945 29975 26979
rect 29917 26939 29975 26945
rect 30750 26936 30756 26988
rect 30808 26985 30814 26988
rect 30808 26979 30849 26985
rect 30837 26945 30849 26979
rect 30808 26939 30849 26945
rect 30808 26936 30814 26939
rect 31018 26936 31024 26988
rect 31076 26936 31082 26988
rect 22373 26911 22431 26917
rect 22373 26908 22385 26911
rect 21468 26880 22385 26908
rect 22373 26877 22385 26880
rect 22419 26877 22431 26911
rect 22373 26871 22431 26877
rect 22554 26868 22560 26920
rect 22612 26868 22618 26920
rect 24026 26868 24032 26920
rect 24084 26908 24090 26920
rect 24765 26911 24823 26917
rect 24765 26908 24777 26911
rect 24084 26880 24777 26908
rect 24084 26868 24090 26880
rect 24765 26877 24777 26880
rect 24811 26877 24823 26911
rect 24765 26871 24823 26877
rect 25590 26868 25596 26920
rect 25648 26908 25654 26920
rect 26973 26911 27031 26917
rect 26973 26908 26985 26911
rect 25648 26880 26985 26908
rect 25648 26868 25654 26880
rect 21376 26812 22048 26840
rect 17218 26772 17224 26784
rect 14200 26744 17224 26772
rect 17218 26732 17224 26744
rect 17276 26732 17282 26784
rect 17494 26732 17500 26784
rect 17552 26772 17558 26784
rect 17770 26772 17776 26784
rect 17552 26744 17776 26772
rect 17552 26732 17558 26744
rect 17770 26732 17776 26744
rect 17828 26732 17834 26784
rect 18046 26732 18052 26784
rect 18104 26732 18110 26784
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 21542 26772 21548 26784
rect 20496 26744 21548 26772
rect 20496 26732 20502 26744
rect 21542 26732 21548 26744
rect 21600 26732 21606 26784
rect 21726 26732 21732 26784
rect 21784 26772 21790 26784
rect 22020 26781 22048 26812
rect 23842 26800 23848 26852
rect 23900 26840 23906 26852
rect 24210 26840 24216 26852
rect 23900 26812 24216 26840
rect 23900 26800 23906 26812
rect 24210 26800 24216 26812
rect 24268 26800 24274 26852
rect 25498 26800 25504 26852
rect 25556 26840 25562 26852
rect 26620 26849 26648 26880
rect 26973 26877 26985 26880
rect 27019 26877 27031 26911
rect 26973 26871 27031 26877
rect 27249 26911 27307 26917
rect 27249 26877 27261 26911
rect 27295 26908 27307 26911
rect 27430 26908 27436 26920
rect 27295 26880 27436 26908
rect 27295 26877 27307 26880
rect 27249 26871 27307 26877
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 29546 26868 29552 26920
rect 29604 26908 29610 26920
rect 29733 26911 29791 26917
rect 29733 26908 29745 26911
rect 29604 26880 29745 26908
rect 29604 26868 29610 26880
rect 29733 26877 29745 26880
rect 29779 26877 29791 26911
rect 29733 26871 29791 26877
rect 26053 26843 26111 26849
rect 26053 26840 26065 26843
rect 25556 26812 26065 26840
rect 25556 26800 25562 26812
rect 26053 26809 26065 26812
rect 26099 26809 26111 26843
rect 26053 26803 26111 26809
rect 26605 26843 26663 26849
rect 26605 26809 26617 26843
rect 26651 26809 26663 26843
rect 26605 26803 26663 26809
rect 28994 26800 29000 26852
rect 29052 26840 29058 26852
rect 29564 26840 29592 26868
rect 29052 26812 29592 26840
rect 30193 26843 30251 26849
rect 29052 26800 29058 26812
rect 30193 26809 30205 26843
rect 30239 26840 30251 26843
rect 30374 26840 30380 26852
rect 30239 26812 30380 26840
rect 30239 26809 30251 26812
rect 30193 26803 30251 26809
rect 30374 26800 30380 26812
rect 30432 26800 30438 26852
rect 30650 26800 30656 26852
rect 30708 26840 30714 26852
rect 30745 26843 30803 26849
rect 30745 26840 30757 26843
rect 30708 26812 30757 26840
rect 30708 26800 30714 26812
rect 30745 26809 30757 26812
rect 30791 26809 30803 26843
rect 31220 26840 31248 27084
rect 31478 27072 31484 27124
rect 31536 27072 31542 27124
rect 32214 27072 32220 27124
rect 32272 27112 32278 27124
rect 32766 27112 32772 27124
rect 32272 27084 32772 27112
rect 32272 27072 32278 27084
rect 32766 27072 32772 27084
rect 32824 27072 32830 27124
rect 33428 27084 35020 27112
rect 31329 27047 31387 27053
rect 31329 27013 31341 27047
rect 31375 27044 31387 27047
rect 31570 27044 31576 27056
rect 31375 27016 31576 27044
rect 31375 27013 31387 27016
rect 31329 27007 31387 27013
rect 31570 27004 31576 27016
rect 31628 27004 31634 27056
rect 31846 27004 31852 27056
rect 31904 27044 31910 27056
rect 32398 27044 32404 27056
rect 31904 27016 32404 27044
rect 31904 27004 31910 27016
rect 32398 27004 32404 27016
rect 32456 27004 32462 27056
rect 32582 27004 32588 27056
rect 32640 27044 32646 27056
rect 32921 27047 32979 27053
rect 32921 27044 32933 27047
rect 32640 27016 32933 27044
rect 32640 27004 32646 27016
rect 32921 27013 32933 27016
rect 32967 27013 32979 27047
rect 32921 27007 32979 27013
rect 33134 27004 33140 27056
rect 33192 27004 33198 27056
rect 33428 27053 33456 27084
rect 33413 27047 33471 27053
rect 33413 27013 33425 27047
rect 33459 27013 33471 27047
rect 33413 27007 33471 27013
rect 34238 27004 34244 27056
rect 34296 27044 34302 27056
rect 34609 27047 34667 27053
rect 34609 27044 34621 27047
rect 34296 27016 34621 27044
rect 34296 27004 34302 27016
rect 34609 27013 34621 27016
rect 34655 27044 34667 27047
rect 34655 27016 34928 27044
rect 34655 27013 34667 27016
rect 34609 27007 34667 27013
rect 33226 26936 33232 26988
rect 33284 26936 33290 26988
rect 33594 26936 33600 26988
rect 33652 26976 33658 26988
rect 33689 26979 33747 26985
rect 33689 26976 33701 26979
rect 33652 26948 33701 26976
rect 33652 26936 33658 26948
rect 33689 26945 33701 26948
rect 33735 26945 33747 26979
rect 33689 26939 33747 26945
rect 33873 26979 33931 26985
rect 33873 26945 33885 26979
rect 33919 26976 33931 26979
rect 34330 26976 34336 26988
rect 33919 26948 34336 26976
rect 33919 26945 33931 26948
rect 33873 26939 33931 26945
rect 34330 26936 34336 26948
rect 34388 26936 34394 26988
rect 34422 26936 34428 26988
rect 34480 26976 34486 26988
rect 34480 26948 34652 26976
rect 34480 26936 34486 26948
rect 34624 26908 34652 26948
rect 34790 26936 34796 26988
rect 34848 26936 34854 26988
rect 34900 26985 34928 27016
rect 34885 26979 34943 26985
rect 34885 26945 34897 26979
rect 34931 26945 34943 26979
rect 34992 26976 35020 27084
rect 35066 27004 35072 27056
rect 35124 27044 35130 27056
rect 35253 27047 35311 27053
rect 35253 27044 35265 27047
rect 35124 27016 35265 27044
rect 35124 27004 35130 27016
rect 35253 27013 35265 27016
rect 35299 27013 35311 27047
rect 35253 27007 35311 27013
rect 35342 27004 35348 27056
rect 35400 27044 35406 27056
rect 35989 27047 36047 27053
rect 35989 27044 36001 27047
rect 35400 27016 36001 27044
rect 35400 27004 35406 27016
rect 35989 27013 36001 27016
rect 36035 27013 36047 27047
rect 35989 27007 36047 27013
rect 35526 26976 35532 26988
rect 34992 26948 35532 26976
rect 34885 26939 34943 26945
rect 35526 26936 35532 26948
rect 35584 26936 35590 26988
rect 35710 26936 35716 26988
rect 35768 26936 35774 26988
rect 35897 26979 35955 26985
rect 35897 26945 35909 26979
rect 35943 26976 35955 26979
rect 36078 26976 36084 26988
rect 35943 26948 36084 26976
rect 35943 26945 35955 26948
rect 35897 26939 35955 26945
rect 36078 26936 36084 26948
rect 36136 26936 36142 26988
rect 34624 26880 34928 26908
rect 33597 26843 33655 26849
rect 31220 26812 32996 26840
rect 30745 26803 30803 26809
rect 21821 26775 21879 26781
rect 21821 26772 21833 26775
rect 21784 26744 21833 26772
rect 21784 26732 21790 26744
rect 21821 26741 21833 26744
rect 21867 26741 21879 26775
rect 21821 26735 21879 26741
rect 22005 26775 22063 26781
rect 22005 26741 22017 26775
rect 22051 26772 22063 26775
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 22051 26744 22293 26772
rect 22051 26741 22063 26744
rect 22005 26735 22063 26741
rect 22281 26741 22293 26744
rect 22327 26741 22339 26775
rect 22281 26735 22339 26741
rect 22646 26732 22652 26784
rect 22704 26772 22710 26784
rect 26234 26772 26240 26784
rect 22704 26744 26240 26772
rect 22704 26732 22710 26744
rect 26234 26732 26240 26744
rect 26292 26732 26298 26784
rect 30098 26732 30104 26784
rect 30156 26732 30162 26784
rect 30282 26732 30288 26784
rect 30340 26772 30346 26784
rect 31297 26775 31355 26781
rect 31297 26772 31309 26775
rect 30340 26744 31309 26772
rect 30340 26732 30346 26744
rect 31297 26741 31309 26744
rect 31343 26741 31355 26775
rect 31297 26735 31355 26741
rect 32398 26732 32404 26784
rect 32456 26772 32462 26784
rect 32769 26775 32827 26781
rect 32769 26772 32781 26775
rect 32456 26744 32781 26772
rect 32456 26732 32462 26744
rect 32769 26741 32781 26744
rect 32815 26741 32827 26775
rect 32769 26735 32827 26741
rect 32858 26732 32864 26784
rect 32916 26772 32922 26784
rect 32968 26781 32996 26812
rect 33597 26809 33609 26843
rect 33643 26840 33655 26843
rect 33962 26840 33968 26852
rect 33643 26812 33968 26840
rect 33643 26809 33655 26812
rect 33597 26803 33655 26809
rect 33962 26800 33968 26812
rect 34020 26800 34026 26852
rect 34054 26800 34060 26852
rect 34112 26840 34118 26852
rect 34149 26843 34207 26849
rect 34149 26840 34161 26843
rect 34112 26812 34161 26840
rect 34112 26800 34118 26812
rect 34149 26809 34161 26812
rect 34195 26840 34207 26843
rect 34790 26840 34796 26852
rect 34195 26812 34796 26840
rect 34195 26809 34207 26812
rect 34149 26803 34207 26809
rect 34790 26800 34796 26812
rect 34848 26800 34854 26852
rect 34900 26840 34928 26880
rect 35805 26843 35863 26849
rect 35805 26840 35817 26843
rect 34900 26812 35817 26840
rect 35805 26809 35817 26812
rect 35851 26809 35863 26843
rect 35805 26803 35863 26809
rect 32953 26775 33011 26781
rect 32953 26772 32965 26775
rect 32916 26744 32965 26772
rect 32916 26732 32922 26744
rect 32953 26741 32965 26744
rect 32999 26741 33011 26775
rect 32953 26735 33011 26741
rect 33042 26732 33048 26784
rect 33100 26772 33106 26784
rect 33689 26775 33747 26781
rect 33689 26772 33701 26775
rect 33100 26744 33701 26772
rect 33100 26732 33106 26744
rect 33689 26741 33701 26744
rect 33735 26741 33747 26775
rect 34808 26772 34836 26800
rect 35253 26775 35311 26781
rect 35253 26772 35265 26775
rect 34808 26744 35265 26772
rect 33689 26735 33747 26741
rect 35253 26741 35265 26744
rect 35299 26741 35311 26775
rect 35253 26735 35311 26741
rect 35437 26775 35495 26781
rect 35437 26741 35449 26775
rect 35483 26772 35495 26775
rect 35986 26772 35992 26784
rect 35483 26744 35992 26772
rect 35483 26741 35495 26744
rect 35437 26735 35495 26741
rect 35986 26732 35992 26744
rect 36044 26732 36050 26784
rect 1104 26682 36524 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 36524 26682
rect 1104 26608 36524 26630
rect 4798 26528 4804 26580
rect 4856 26528 4862 26580
rect 6270 26568 6276 26580
rect 5368 26540 6276 26568
rect 3786 26392 3792 26444
rect 3844 26432 3850 26444
rect 5368 26441 5396 26540
rect 6270 26528 6276 26540
rect 6328 26528 6334 26580
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 8021 26571 8079 26577
rect 8021 26568 8033 26571
rect 7800 26540 8033 26568
rect 7800 26528 7806 26540
rect 8021 26537 8033 26540
rect 8067 26537 8079 26571
rect 8021 26531 8079 26537
rect 8386 26528 8392 26580
rect 8444 26568 8450 26580
rect 8941 26571 8999 26577
rect 8941 26568 8953 26571
rect 8444 26540 8953 26568
rect 8444 26528 8450 26540
rect 8941 26537 8953 26540
rect 8987 26537 8999 26571
rect 8941 26531 8999 26537
rect 9677 26571 9735 26577
rect 9677 26537 9689 26571
rect 9723 26568 9735 26571
rect 9858 26568 9864 26580
rect 9723 26540 9864 26568
rect 9723 26537 9735 26540
rect 9677 26531 9735 26537
rect 9858 26528 9864 26540
rect 9916 26528 9922 26580
rect 9950 26528 9956 26580
rect 10008 26568 10014 26580
rect 14366 26568 14372 26580
rect 10008 26540 14372 26568
rect 10008 26528 10014 26540
rect 14366 26528 14372 26540
rect 14424 26528 14430 26580
rect 14918 26568 14924 26580
rect 14568 26540 14924 26568
rect 5442 26460 5448 26512
rect 5500 26500 5506 26512
rect 5629 26503 5687 26509
rect 5629 26500 5641 26503
rect 5500 26472 5641 26500
rect 5500 26460 5506 26472
rect 5629 26469 5641 26472
rect 5675 26469 5687 26503
rect 9214 26500 9220 26512
rect 5629 26463 5687 26469
rect 6932 26472 9220 26500
rect 3881 26435 3939 26441
rect 3881 26432 3893 26435
rect 3844 26404 3893 26432
rect 3844 26392 3850 26404
rect 3881 26401 3893 26404
rect 3927 26401 3939 26435
rect 3881 26395 3939 26401
rect 5353 26435 5411 26441
rect 5353 26401 5365 26435
rect 5399 26401 5411 26435
rect 5994 26432 6000 26444
rect 5353 26395 5411 26401
rect 5736 26404 6000 26432
rect 4709 26367 4767 26373
rect 4709 26333 4721 26367
rect 4755 26364 4767 26367
rect 5736 26364 5764 26404
rect 5994 26392 6000 26404
rect 6052 26392 6058 26444
rect 4755 26336 5764 26364
rect 5813 26367 5871 26373
rect 4755 26333 4767 26336
rect 4709 26327 4767 26333
rect 5813 26333 5825 26367
rect 5859 26333 5871 26367
rect 5813 26327 5871 26333
rect 5166 26256 5172 26308
rect 5224 26256 5230 26308
rect 5718 26256 5724 26308
rect 5776 26296 5782 26308
rect 5828 26296 5856 26327
rect 5902 26324 5908 26376
rect 5960 26324 5966 26376
rect 6178 26324 6184 26376
rect 6236 26324 6242 26376
rect 6932 26373 6960 26472
rect 9214 26460 9220 26472
rect 9272 26460 9278 26512
rect 9398 26460 9404 26512
rect 9456 26500 9462 26512
rect 13262 26500 13268 26512
rect 9456 26472 13268 26500
rect 9456 26460 9462 26472
rect 13262 26460 13268 26472
rect 13320 26460 13326 26512
rect 13357 26503 13415 26509
rect 13357 26469 13369 26503
rect 13403 26469 13415 26503
rect 13357 26463 13415 26469
rect 7650 26392 7656 26444
rect 7708 26432 7714 26444
rect 8018 26432 8024 26444
rect 7708 26404 8024 26432
rect 7708 26392 7714 26404
rect 8018 26392 8024 26404
rect 8076 26432 8082 26444
rect 8076 26404 8202 26432
rect 8076 26392 8082 26404
rect 6917 26367 6975 26373
rect 6917 26333 6929 26367
rect 6963 26333 6975 26367
rect 6917 26327 6975 26333
rect 7926 26324 7932 26376
rect 7984 26324 7990 26376
rect 8174 26373 8202 26404
rect 8294 26392 8300 26444
rect 8352 26432 8358 26444
rect 13372 26432 13400 26463
rect 14274 26460 14280 26512
rect 14332 26500 14338 26512
rect 14568 26500 14596 26540
rect 14918 26528 14924 26540
rect 14976 26528 14982 26580
rect 17770 26528 17776 26580
rect 17828 26528 17834 26580
rect 20990 26528 20996 26580
rect 21048 26568 21054 26580
rect 21085 26571 21143 26577
rect 21085 26568 21097 26571
rect 21048 26540 21097 26568
rect 21048 26528 21054 26540
rect 21085 26537 21097 26540
rect 21131 26537 21143 26571
rect 21085 26531 21143 26537
rect 21910 26528 21916 26580
rect 21968 26568 21974 26580
rect 26142 26568 26148 26580
rect 21968 26540 26148 26568
rect 21968 26528 21974 26540
rect 26142 26528 26148 26540
rect 26200 26568 26206 26580
rect 26237 26571 26295 26577
rect 26237 26568 26249 26571
rect 26200 26540 26249 26568
rect 26200 26528 26206 26540
rect 26237 26537 26249 26540
rect 26283 26537 26295 26571
rect 26237 26531 26295 26537
rect 26602 26528 26608 26580
rect 26660 26568 26666 26580
rect 26697 26571 26755 26577
rect 26697 26568 26709 26571
rect 26660 26540 26709 26568
rect 26660 26528 26666 26540
rect 26697 26537 26709 26540
rect 26743 26537 26755 26571
rect 26697 26531 26755 26537
rect 26970 26528 26976 26580
rect 27028 26528 27034 26580
rect 27890 26528 27896 26580
rect 27948 26568 27954 26580
rect 29454 26568 29460 26580
rect 27948 26540 29460 26568
rect 27948 26528 27954 26540
rect 29454 26528 29460 26540
rect 29512 26528 29518 26580
rect 29730 26528 29736 26580
rect 29788 26568 29794 26580
rect 30193 26571 30251 26577
rect 30193 26568 30205 26571
rect 29788 26540 30205 26568
rect 29788 26528 29794 26540
rect 30193 26537 30205 26540
rect 30239 26568 30251 26571
rect 30466 26568 30472 26580
rect 30239 26540 30472 26568
rect 30239 26537 30251 26540
rect 30193 26531 30251 26537
rect 30466 26528 30472 26540
rect 30524 26528 30530 26580
rect 32585 26571 32643 26577
rect 32585 26537 32597 26571
rect 32631 26568 32643 26571
rect 32766 26568 32772 26580
rect 32631 26540 32772 26568
rect 32631 26537 32643 26540
rect 32585 26531 32643 26537
rect 32766 26528 32772 26540
rect 32824 26528 32830 26580
rect 33594 26528 33600 26580
rect 33652 26568 33658 26580
rect 33689 26571 33747 26577
rect 33689 26568 33701 26571
rect 33652 26540 33701 26568
rect 33652 26528 33658 26540
rect 33689 26537 33701 26540
rect 33735 26537 33747 26571
rect 33689 26531 33747 26537
rect 33870 26528 33876 26580
rect 33928 26568 33934 26580
rect 33928 26540 34192 26568
rect 33928 26528 33934 26540
rect 14332 26472 14596 26500
rect 14332 26460 14338 26472
rect 8352 26404 8432 26432
rect 8352 26392 8358 26404
rect 8404 26373 8432 26404
rect 8680 26404 13400 26432
rect 8159 26367 8217 26373
rect 8159 26333 8171 26367
rect 8205 26333 8217 26367
rect 8159 26327 8217 26333
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26333 8447 26367
rect 8570 26364 8576 26376
rect 8531 26336 8576 26364
rect 8389 26327 8447 26333
rect 5776 26268 5856 26296
rect 5997 26299 6055 26305
rect 5776 26256 5782 26268
rect 5997 26265 6009 26299
rect 6043 26265 6055 26299
rect 5997 26259 6055 26265
rect 4154 26188 4160 26240
rect 4212 26228 4218 26240
rect 5261 26231 5319 26237
rect 5261 26228 5273 26231
rect 4212 26200 5273 26228
rect 4212 26188 4218 26200
rect 5261 26197 5273 26200
rect 5307 26197 5319 26231
rect 5261 26191 5319 26197
rect 5810 26188 5816 26240
rect 5868 26228 5874 26240
rect 6012 26228 6040 26259
rect 6730 26256 6736 26308
rect 6788 26256 6794 26308
rect 7944 26296 7972 26324
rect 8297 26299 8355 26305
rect 8297 26296 8309 26299
rect 7944 26268 8309 26296
rect 8297 26265 8309 26268
rect 8343 26265 8355 26299
rect 8404 26296 8432 26327
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 8680 26373 8708 26404
rect 8665 26367 8723 26373
rect 8665 26333 8677 26367
rect 8711 26333 8723 26367
rect 8665 26327 8723 26333
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9493 26367 9551 26373
rect 9493 26333 9505 26367
rect 9539 26364 9551 26367
rect 9766 26364 9772 26376
rect 9539 26336 9772 26364
rect 9539 26333 9551 26336
rect 9493 26327 9551 26333
rect 8938 26296 8944 26308
rect 8404 26268 8944 26296
rect 8297 26259 8355 26265
rect 8938 26256 8944 26268
rect 8996 26296 9002 26308
rect 9140 26296 9168 26327
rect 9766 26324 9772 26336
rect 9824 26324 9830 26376
rect 9858 26324 9864 26376
rect 9916 26324 9922 26376
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26364 10195 26367
rect 10410 26364 10416 26376
rect 10183 26336 10416 26364
rect 10183 26333 10195 26336
rect 10137 26327 10195 26333
rect 10410 26324 10416 26336
rect 10468 26364 10474 26376
rect 10778 26364 10784 26376
rect 10468 26336 10784 26364
rect 10468 26324 10474 26336
rect 10778 26324 10784 26336
rect 10836 26324 10842 26376
rect 12526 26324 12532 26376
rect 12584 26324 12590 26376
rect 12710 26324 12716 26376
rect 12768 26324 12774 26376
rect 12805 26367 12863 26373
rect 12805 26333 12817 26367
rect 12851 26333 12863 26367
rect 12805 26327 12863 26333
rect 9217 26299 9275 26305
rect 9217 26296 9229 26299
rect 8996 26268 9168 26296
rect 8996 26256 9002 26268
rect 9198 26265 9229 26296
rect 9263 26265 9275 26299
rect 9198 26259 9275 26265
rect 5868 26200 6040 26228
rect 5868 26188 5874 26200
rect 7006 26188 7012 26240
rect 7064 26228 7070 26240
rect 7285 26231 7343 26237
rect 7285 26228 7297 26231
rect 7064 26200 7297 26228
rect 7064 26188 7070 26200
rect 7285 26197 7297 26200
rect 7331 26197 7343 26231
rect 7285 26191 7343 26197
rect 8846 26188 8852 26240
rect 8904 26228 8910 26240
rect 9198 26228 9226 26259
rect 9306 26256 9312 26308
rect 9364 26296 9370 26308
rect 9950 26296 9956 26308
rect 9364 26268 9956 26296
rect 9364 26256 9370 26268
rect 9950 26256 9956 26268
rect 10008 26256 10014 26308
rect 11054 26256 11060 26308
rect 11112 26296 11118 26308
rect 12345 26299 12403 26305
rect 12345 26296 12357 26299
rect 11112 26268 12357 26296
rect 11112 26256 11118 26268
rect 12345 26265 12357 26268
rect 12391 26265 12403 26299
rect 12345 26259 12403 26265
rect 12618 26256 12624 26308
rect 12676 26296 12682 26308
rect 12820 26296 12848 26327
rect 12894 26324 12900 26376
rect 12952 26324 12958 26376
rect 13078 26324 13084 26376
rect 13136 26324 13142 26376
rect 13262 26324 13268 26376
rect 13320 26364 13326 26376
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 13320 26336 13553 26364
rect 13320 26324 13326 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13633 26367 13691 26373
rect 13633 26333 13645 26367
rect 13679 26364 13691 26367
rect 13679 26336 13860 26364
rect 13679 26333 13691 26336
rect 13633 26327 13691 26333
rect 12676 26268 12848 26296
rect 13725 26299 13783 26305
rect 12676 26256 12682 26268
rect 13725 26265 13737 26299
rect 13771 26265 13783 26299
rect 13832 26296 13860 26336
rect 13906 26324 13912 26376
rect 13964 26324 13970 26376
rect 14090 26324 14096 26376
rect 14148 26364 14154 26376
rect 14366 26373 14372 26376
rect 14185 26367 14243 26373
rect 14185 26364 14197 26367
rect 14148 26336 14197 26364
rect 14148 26324 14154 26336
rect 14185 26333 14197 26336
rect 14231 26333 14243 26367
rect 14185 26327 14243 26333
rect 14333 26367 14372 26373
rect 14333 26333 14345 26367
rect 14333 26327 14372 26333
rect 14366 26324 14372 26327
rect 14424 26324 14430 26376
rect 14461 26367 14519 26373
rect 14461 26333 14473 26367
rect 14507 26364 14519 26367
rect 14568 26364 14596 26472
rect 14829 26503 14887 26509
rect 14829 26469 14841 26503
rect 14875 26500 14887 26503
rect 15289 26503 15347 26509
rect 15289 26500 15301 26503
rect 14875 26472 15301 26500
rect 14875 26469 14887 26472
rect 14829 26463 14887 26469
rect 15289 26469 15301 26472
rect 15335 26469 15347 26503
rect 15289 26463 15347 26469
rect 17512 26472 19334 26500
rect 14918 26392 14924 26444
rect 14976 26392 14982 26444
rect 15838 26392 15844 26444
rect 15896 26432 15902 26444
rect 17512 26432 17540 26472
rect 15896 26404 17540 26432
rect 15896 26392 15902 26404
rect 14507 26336 14596 26364
rect 14507 26333 14519 26336
rect 14461 26327 14519 26333
rect 14642 26324 14648 26376
rect 14700 26373 14706 26376
rect 14700 26364 14708 26373
rect 15105 26367 15163 26373
rect 14700 26336 14745 26364
rect 14700 26327 14708 26336
rect 15105 26333 15117 26367
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26364 15439 26367
rect 15562 26364 15568 26376
rect 15427 26336 15568 26364
rect 15427 26333 15439 26336
rect 15381 26327 15439 26333
rect 14700 26324 14706 26327
rect 13998 26296 14004 26308
rect 13832 26268 14004 26296
rect 13725 26259 13783 26265
rect 8904 26200 9226 26228
rect 8904 26188 8910 26200
rect 9766 26188 9772 26240
rect 9824 26228 9830 26240
rect 10045 26231 10103 26237
rect 10045 26228 10057 26231
rect 9824 26200 10057 26228
rect 9824 26188 9830 26200
rect 10045 26197 10057 26200
rect 10091 26228 10103 26231
rect 10594 26228 10600 26240
rect 10091 26200 10600 26228
rect 10091 26197 10103 26200
rect 10045 26191 10103 26197
rect 10594 26188 10600 26200
rect 10652 26228 10658 26240
rect 11146 26228 11152 26240
rect 10652 26200 11152 26228
rect 10652 26188 10658 26200
rect 11146 26188 11152 26200
rect 11204 26188 11210 26240
rect 13262 26188 13268 26240
rect 13320 26228 13326 26240
rect 13740 26228 13768 26259
rect 13998 26256 14004 26268
rect 14056 26296 14062 26308
rect 14553 26299 14611 26305
rect 14553 26296 14565 26299
rect 14056 26268 14565 26296
rect 14056 26256 14062 26268
rect 14553 26265 14565 26268
rect 14599 26265 14611 26299
rect 14553 26259 14611 26265
rect 14918 26256 14924 26308
rect 14976 26296 14982 26308
rect 15120 26296 15148 26327
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 16761 26367 16819 26373
rect 16761 26364 16773 26367
rect 16724 26336 16773 26364
rect 16724 26324 16730 26336
rect 16761 26333 16773 26336
rect 16807 26333 16819 26367
rect 16761 26327 16819 26333
rect 17037 26367 17095 26373
rect 17037 26333 17049 26367
rect 17083 26364 17095 26367
rect 17126 26364 17132 26376
rect 17083 26336 17132 26364
rect 17083 26333 17095 26336
rect 17037 26327 17095 26333
rect 17126 26324 17132 26336
rect 17184 26324 17190 26376
rect 17218 26324 17224 26376
rect 17276 26324 17282 26376
rect 17402 26373 17408 26376
rect 17400 26364 17408 26373
rect 17363 26336 17408 26364
rect 17400 26327 17408 26336
rect 17402 26324 17408 26327
rect 17460 26324 17466 26376
rect 17512 26373 17540 26404
rect 17586 26392 17592 26444
rect 17644 26392 17650 26444
rect 17497 26367 17555 26373
rect 17497 26333 17509 26367
rect 17543 26333 17555 26367
rect 17497 26327 17555 26333
rect 17604 26305 17632 26392
rect 19306 26364 19334 26472
rect 21174 26460 21180 26512
rect 21232 26500 21238 26512
rect 21269 26503 21327 26509
rect 21269 26500 21281 26503
rect 21232 26472 21281 26500
rect 21232 26460 21238 26472
rect 21269 26469 21281 26472
rect 21315 26500 21327 26503
rect 21315 26472 22692 26500
rect 21315 26469 21327 26472
rect 21269 26463 21327 26469
rect 20070 26392 20076 26444
rect 20128 26432 20134 26444
rect 21361 26435 21419 26441
rect 21361 26432 21373 26435
rect 20128 26404 21373 26432
rect 20128 26392 20134 26404
rect 21361 26401 21373 26404
rect 21407 26401 21419 26435
rect 21361 26395 21419 26401
rect 21726 26392 21732 26444
rect 21784 26392 21790 26444
rect 21818 26392 21824 26444
rect 21876 26432 21882 26444
rect 21876 26404 22600 26432
rect 21876 26392 21882 26404
rect 20162 26364 20168 26376
rect 19306 26336 20168 26364
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 22373 26367 22431 26373
rect 22373 26364 22385 26367
rect 22152 26336 22385 26364
rect 22152 26324 22158 26336
rect 22373 26333 22385 26336
rect 22419 26333 22431 26367
rect 22373 26327 22431 26333
rect 22462 26324 22468 26376
rect 22520 26324 22526 26376
rect 17589 26299 17647 26305
rect 17589 26296 17601 26299
rect 14976 26268 15148 26296
rect 15672 26268 17601 26296
rect 14976 26256 14982 26268
rect 15672 26228 15700 26268
rect 16776 26240 16804 26268
rect 17589 26265 17601 26268
rect 17635 26265 17647 26299
rect 17589 26259 17647 26265
rect 17678 26256 17684 26308
rect 17736 26296 17742 26308
rect 17773 26299 17831 26305
rect 17773 26296 17785 26299
rect 17736 26268 17785 26296
rect 17736 26256 17742 26268
rect 17773 26265 17785 26268
rect 17819 26265 17831 26299
rect 17773 26259 17831 26265
rect 18138 26256 18144 26308
rect 18196 26296 18202 26308
rect 20438 26296 20444 26308
rect 18196 26268 20444 26296
rect 18196 26256 18202 26268
rect 20438 26256 20444 26268
rect 20496 26296 20502 26308
rect 20901 26299 20959 26305
rect 20901 26296 20913 26299
rect 20496 26268 20913 26296
rect 20496 26256 20502 26268
rect 20901 26265 20913 26268
rect 20947 26265 20959 26299
rect 20901 26259 20959 26265
rect 21082 26256 21088 26308
rect 21140 26305 21146 26308
rect 21140 26299 21159 26305
rect 21147 26265 21159 26299
rect 21140 26259 21159 26265
rect 21140 26256 21146 26259
rect 21450 26256 21456 26308
rect 21508 26296 21514 26308
rect 22189 26299 22247 26305
rect 22189 26296 22201 26299
rect 21508 26268 22201 26296
rect 21508 26256 21514 26268
rect 22189 26265 22201 26268
rect 22235 26265 22247 26299
rect 22572 26296 22600 26404
rect 22664 26373 22692 26472
rect 24302 26460 24308 26512
rect 24360 26500 24366 26512
rect 24360 26472 28212 26500
rect 24360 26460 24366 26472
rect 26326 26392 26332 26444
rect 26384 26392 26390 26444
rect 26878 26432 26884 26444
rect 26528 26404 26884 26432
rect 22649 26367 22707 26373
rect 22649 26333 22661 26367
rect 22695 26333 22707 26367
rect 22649 26327 22707 26333
rect 22741 26367 22799 26373
rect 22741 26333 22753 26367
rect 22787 26364 22799 26367
rect 22922 26364 22928 26376
rect 22787 26336 22928 26364
rect 22787 26333 22799 26336
rect 22741 26327 22799 26333
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 25866 26324 25872 26376
rect 25924 26324 25930 26376
rect 26418 26324 26424 26376
rect 26476 26364 26482 26376
rect 26528 26373 26556 26404
rect 26878 26392 26884 26404
rect 26936 26392 26942 26444
rect 28184 26432 28212 26472
rect 29822 26460 29828 26512
rect 29880 26500 29886 26512
rect 32122 26500 32128 26512
rect 29880 26472 32128 26500
rect 29880 26460 29886 26472
rect 32122 26460 32128 26472
rect 32180 26460 32186 26512
rect 33781 26503 33839 26509
rect 33781 26500 33793 26503
rect 32692 26472 33793 26500
rect 28184 26404 28994 26432
rect 26513 26367 26571 26373
rect 26513 26364 26525 26367
rect 26476 26336 26525 26364
rect 26476 26324 26482 26336
rect 26513 26333 26525 26336
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 27430 26324 27436 26376
rect 27488 26324 27494 26376
rect 27801 26367 27859 26373
rect 27801 26333 27813 26367
rect 27847 26333 27859 26367
rect 27801 26327 27859 26333
rect 24762 26296 24768 26308
rect 22572 26268 24768 26296
rect 22189 26259 22247 26265
rect 24762 26256 24768 26268
rect 24820 26256 24826 26308
rect 26053 26299 26111 26305
rect 26053 26265 26065 26299
rect 26099 26296 26111 26299
rect 26602 26296 26608 26308
rect 26099 26268 26608 26296
rect 26099 26265 26111 26268
rect 26053 26259 26111 26265
rect 26602 26256 26608 26268
rect 26660 26256 26666 26308
rect 26694 26256 26700 26308
rect 26752 26296 26758 26308
rect 26881 26299 26939 26305
rect 26881 26296 26893 26299
rect 26752 26268 26893 26296
rect 26752 26256 26758 26268
rect 26881 26265 26893 26268
rect 26927 26296 26939 26299
rect 27816 26296 27844 26327
rect 27890 26324 27896 26376
rect 27948 26324 27954 26376
rect 28184 26373 28212 26404
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26333 28227 26367
rect 28169 26327 28227 26333
rect 28350 26324 28356 26376
rect 28408 26324 28414 26376
rect 28074 26296 28080 26308
rect 26927 26268 27292 26296
rect 27816 26268 28080 26296
rect 26927 26265 26939 26268
rect 26881 26259 26939 26265
rect 13320 26200 15700 26228
rect 13320 26188 13326 26200
rect 16298 26188 16304 26240
rect 16356 26228 16362 26240
rect 16577 26231 16635 26237
rect 16577 26228 16589 26231
rect 16356 26200 16589 26228
rect 16356 26188 16362 26200
rect 16577 26197 16589 26200
rect 16623 26197 16635 26231
rect 16577 26191 16635 26197
rect 16758 26188 16764 26240
rect 16816 26188 16822 26240
rect 17310 26188 17316 26240
rect 17368 26228 17374 26240
rect 18874 26228 18880 26240
rect 17368 26200 18880 26228
rect 17368 26188 17374 26200
rect 18874 26188 18880 26200
rect 18932 26188 18938 26240
rect 21545 26231 21603 26237
rect 21545 26197 21557 26231
rect 21591 26228 21603 26231
rect 24670 26228 24676 26240
rect 21591 26200 24676 26228
rect 21591 26197 21603 26200
rect 21545 26191 21603 26197
rect 24670 26188 24676 26200
rect 24728 26188 24734 26240
rect 27264 26237 27292 26268
rect 28074 26256 28080 26268
rect 28132 26256 28138 26308
rect 28258 26256 28264 26308
rect 28316 26256 28322 26308
rect 28966 26296 28994 26404
rect 29914 26392 29920 26444
rect 29972 26432 29978 26444
rect 30190 26432 30196 26444
rect 29972 26404 30196 26432
rect 29972 26392 29978 26404
rect 30190 26392 30196 26404
rect 30248 26392 30254 26444
rect 30374 26392 30380 26444
rect 30432 26432 30438 26444
rect 32692 26432 32720 26472
rect 33781 26469 33793 26472
rect 33827 26500 33839 26503
rect 34054 26500 34060 26512
rect 33827 26472 34060 26500
rect 33827 26469 33839 26472
rect 33781 26463 33839 26469
rect 34054 26460 34060 26472
rect 34112 26460 34118 26512
rect 33042 26432 33048 26444
rect 30432 26404 30604 26432
rect 30432 26392 30438 26404
rect 30576 26373 30604 26404
rect 31772 26404 32720 26432
rect 32784 26404 33048 26432
rect 31772 26376 31800 26404
rect 30561 26367 30619 26373
rect 30561 26333 30573 26367
rect 30607 26333 30619 26367
rect 30561 26327 30619 26333
rect 30837 26367 30895 26373
rect 30837 26333 30849 26367
rect 30883 26364 30895 26367
rect 31754 26364 31760 26376
rect 30883 26336 31760 26364
rect 30883 26333 30895 26336
rect 30837 26327 30895 26333
rect 31754 26324 31760 26336
rect 31812 26324 31818 26376
rect 32784 26373 32812 26404
rect 33042 26392 33048 26404
rect 33100 26392 33106 26444
rect 33134 26392 33140 26444
rect 33192 26432 33198 26444
rect 34164 26432 34192 26540
rect 34330 26528 34336 26580
rect 34388 26568 34394 26580
rect 35069 26571 35127 26577
rect 35069 26568 35081 26571
rect 34388 26540 35081 26568
rect 34388 26528 34394 26540
rect 35069 26537 35081 26540
rect 35115 26537 35127 26571
rect 35069 26531 35127 26537
rect 34514 26460 34520 26512
rect 34572 26500 34578 26512
rect 35989 26503 36047 26509
rect 35989 26500 36001 26503
rect 34572 26472 36001 26500
rect 34572 26460 34578 26472
rect 35989 26469 36001 26472
rect 36035 26469 36047 26503
rect 35989 26463 36047 26469
rect 33192 26404 33916 26432
rect 33192 26392 33198 26404
rect 32769 26367 32827 26373
rect 32769 26333 32781 26367
rect 32815 26333 32827 26367
rect 32769 26327 32827 26333
rect 32858 26324 32864 26376
rect 32916 26324 32922 26376
rect 32953 26367 33011 26373
rect 32953 26333 32965 26367
rect 32999 26364 33011 26367
rect 33152 26364 33180 26392
rect 33888 26376 33916 26404
rect 34072 26404 34192 26432
rect 34072 26376 34100 26404
rect 34790 26392 34796 26444
rect 34848 26392 34854 26444
rect 35158 26392 35164 26444
rect 35216 26432 35222 26444
rect 35529 26435 35587 26441
rect 35529 26432 35541 26435
rect 35216 26404 35541 26432
rect 35216 26392 35222 26404
rect 35529 26401 35541 26404
rect 35575 26401 35587 26435
rect 35529 26395 35587 26401
rect 32999 26336 33180 26364
rect 33229 26367 33287 26373
rect 32999 26333 33011 26336
rect 32953 26327 33011 26333
rect 33229 26333 33241 26367
rect 33275 26333 33287 26367
rect 33229 26327 33287 26333
rect 30377 26299 30435 26305
rect 30377 26296 30389 26299
rect 28966 26268 30389 26296
rect 30377 26265 30389 26268
rect 30423 26296 30435 26299
rect 31018 26296 31024 26308
rect 30423 26268 31024 26296
rect 30423 26265 30435 26268
rect 30377 26259 30435 26265
rect 31018 26256 31024 26268
rect 31076 26256 31082 26308
rect 32122 26256 32128 26308
rect 32180 26296 32186 26308
rect 33071 26299 33129 26305
rect 33071 26296 33083 26299
rect 32180 26268 33083 26296
rect 32180 26256 32186 26268
rect 33071 26265 33083 26268
rect 33117 26265 33129 26299
rect 33244 26296 33272 26327
rect 33318 26324 33324 26376
rect 33376 26324 33382 26376
rect 33594 26324 33600 26376
rect 33652 26324 33658 26376
rect 33870 26324 33876 26376
rect 33928 26324 33934 26376
rect 34054 26324 34060 26376
rect 34112 26324 34118 26376
rect 34238 26324 34244 26376
rect 34296 26364 34302 26376
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 34296 26336 34713 26364
rect 34296 26324 34302 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34808 26364 34836 26392
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34808 26336 34897 26364
rect 34701 26327 34759 26333
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 35250 26324 35256 26376
rect 35308 26324 35314 26376
rect 35437 26367 35495 26373
rect 35437 26333 35449 26367
rect 35483 26364 35495 26367
rect 35483 26336 35756 26364
rect 35483 26333 35495 26336
rect 35437 26327 35495 26333
rect 34606 26296 34612 26308
rect 33244 26268 34612 26296
rect 33071 26259 33129 26265
rect 34606 26256 34612 26268
rect 34664 26296 34670 26308
rect 34793 26299 34851 26305
rect 34793 26296 34805 26299
rect 34664 26268 34805 26296
rect 34664 26256 34670 26268
rect 34793 26265 34805 26268
rect 34839 26265 34851 26299
rect 35268 26296 35296 26324
rect 35618 26296 35624 26308
rect 35268 26268 35624 26296
rect 34793 26259 34851 26265
rect 35618 26256 35624 26268
rect 35676 26256 35682 26308
rect 35728 26296 35756 26336
rect 36170 26324 36176 26376
rect 36228 26324 36234 26376
rect 36354 26296 36360 26308
rect 35728 26268 36360 26296
rect 36354 26256 36360 26268
rect 36412 26256 36418 26308
rect 27249 26231 27307 26237
rect 27249 26197 27261 26231
rect 27295 26197 27307 26231
rect 27249 26191 27307 26197
rect 27982 26188 27988 26240
rect 28040 26228 28046 26240
rect 28902 26228 28908 26240
rect 28040 26200 28908 26228
rect 28040 26188 28046 26200
rect 28902 26188 28908 26200
rect 28960 26188 28966 26240
rect 30742 26188 30748 26240
rect 30800 26188 30806 26240
rect 31938 26188 31944 26240
rect 31996 26228 32002 26240
rect 32398 26228 32404 26240
rect 31996 26200 32404 26228
rect 31996 26188 32002 26200
rect 32398 26188 32404 26200
rect 32456 26188 32462 26240
rect 32490 26188 32496 26240
rect 32548 26228 32554 26240
rect 35066 26228 35072 26240
rect 32548 26200 35072 26228
rect 32548 26188 32554 26200
rect 35066 26188 35072 26200
rect 35124 26188 35130 26240
rect 35342 26188 35348 26240
rect 35400 26228 35406 26240
rect 35526 26228 35532 26240
rect 35400 26200 35532 26228
rect 35400 26188 35406 26200
rect 35526 26188 35532 26200
rect 35584 26188 35590 26240
rect 1104 26138 36524 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 36524 26138
rect 1104 26064 36524 26086
rect 3142 25984 3148 26036
rect 3200 25984 3206 26036
rect 4985 26027 5043 26033
rect 4985 25993 4997 26027
rect 5031 26024 5043 26027
rect 6178 26024 6184 26036
rect 5031 25996 6184 26024
rect 5031 25993 5043 25996
rect 4985 25987 5043 25993
rect 6178 25984 6184 25996
rect 6236 26024 6242 26036
rect 6236 25996 7972 26024
rect 6236 25984 6242 25996
rect 2958 25956 2964 25968
rect 2898 25928 2964 25956
rect 2958 25916 2964 25928
rect 3016 25956 3022 25968
rect 3970 25956 3976 25968
rect 3016 25928 3976 25956
rect 3016 25916 3022 25928
rect 3970 25916 3976 25928
rect 4028 25916 4034 25968
rect 5994 25916 6000 25968
rect 6052 25916 6058 25968
rect 6730 25956 6736 25968
rect 6104 25928 6736 25956
rect 6104 25888 6132 25928
rect 6730 25916 6736 25928
rect 6788 25956 6794 25968
rect 7944 25956 7972 25996
rect 8202 25984 8208 26036
rect 8260 25984 8266 26036
rect 9766 25984 9772 26036
rect 9824 25984 9830 26036
rect 10318 25984 10324 26036
rect 10376 26024 10382 26036
rect 11238 26024 11244 26036
rect 10376 25996 11244 26024
rect 10376 25984 10382 25996
rect 9861 25959 9919 25965
rect 6788 25928 7130 25956
rect 7944 25928 9444 25956
rect 6788 25916 6794 25928
rect 4646 25874 6132 25888
rect 4632 25860 6132 25874
rect 1394 25780 1400 25832
rect 1452 25780 1458 25832
rect 1673 25823 1731 25829
rect 1673 25789 1685 25823
rect 1719 25820 1731 25823
rect 2222 25820 2228 25832
rect 1719 25792 2228 25820
rect 1719 25789 1731 25792
rect 1673 25783 1731 25789
rect 2222 25780 2228 25792
rect 2280 25780 2286 25832
rect 2406 25780 2412 25832
rect 2464 25820 2470 25832
rect 3237 25823 3295 25829
rect 3237 25820 3249 25823
rect 2464 25792 3249 25820
rect 2464 25780 2470 25792
rect 3237 25789 3249 25792
rect 3283 25789 3295 25823
rect 3237 25783 3295 25789
rect 3513 25823 3571 25829
rect 3513 25789 3525 25823
rect 3559 25820 3571 25823
rect 3878 25820 3884 25832
rect 3559 25792 3884 25820
rect 3559 25789 3571 25792
rect 3513 25783 3571 25789
rect 3878 25780 3884 25792
rect 3936 25780 3942 25832
rect 4062 25780 4068 25832
rect 4120 25820 4126 25832
rect 4632 25820 4660 25860
rect 8294 25848 8300 25900
rect 8352 25888 8358 25900
rect 8389 25891 8447 25897
rect 8389 25888 8401 25891
rect 8352 25860 8401 25888
rect 8352 25848 8358 25860
rect 8389 25857 8401 25860
rect 8435 25857 8447 25891
rect 8389 25851 8447 25857
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25857 8539 25891
rect 8481 25851 8539 25857
rect 8573 25891 8631 25897
rect 8573 25857 8585 25891
rect 8619 25857 8631 25891
rect 8573 25851 8631 25857
rect 4120 25792 4660 25820
rect 4120 25780 4126 25792
rect 4706 25780 4712 25832
rect 4764 25820 4770 25832
rect 5169 25823 5227 25829
rect 5169 25820 5181 25823
rect 4764 25792 5181 25820
rect 4764 25780 4770 25792
rect 5169 25789 5181 25792
rect 5215 25820 5227 25823
rect 6365 25823 6423 25829
rect 6365 25820 6377 25823
rect 5215 25792 6377 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 6365 25789 6377 25792
rect 6411 25789 6423 25823
rect 6365 25783 6423 25789
rect 6638 25780 6644 25832
rect 6696 25780 6702 25832
rect 8496 25752 8524 25851
rect 8588 25820 8616 25851
rect 8754 25848 8760 25900
rect 8812 25848 8818 25900
rect 9306 25820 9312 25832
rect 8588 25792 9312 25820
rect 9306 25780 9312 25792
rect 9364 25780 9370 25832
rect 8662 25752 8668 25764
rect 8496 25724 8668 25752
rect 8662 25712 8668 25724
rect 8720 25712 8726 25764
rect 1394 25644 1400 25696
rect 1452 25684 1458 25696
rect 2406 25684 2412 25696
rect 1452 25656 2412 25684
rect 1452 25644 1458 25656
rect 2406 25644 2412 25656
rect 2464 25644 2470 25696
rect 7190 25644 7196 25696
rect 7248 25684 7254 25696
rect 7926 25684 7932 25696
rect 7248 25656 7932 25684
rect 7248 25644 7254 25656
rect 7926 25644 7932 25656
rect 7984 25684 7990 25696
rect 8113 25687 8171 25693
rect 8113 25684 8125 25687
rect 7984 25656 8125 25684
rect 7984 25644 7990 25656
rect 8113 25653 8125 25656
rect 8159 25653 8171 25687
rect 8113 25647 8171 25653
rect 9306 25644 9312 25696
rect 9364 25644 9370 25696
rect 9416 25684 9444 25928
rect 9861 25925 9873 25959
rect 9907 25956 9919 25959
rect 10226 25956 10232 25968
rect 9907 25928 10232 25956
rect 9907 25925 9919 25928
rect 9861 25919 9919 25925
rect 10226 25916 10232 25928
rect 10284 25956 10290 25968
rect 10704 25965 10732 25996
rect 11238 25984 11244 25996
rect 11296 25984 11302 26036
rect 11882 25984 11888 26036
rect 11940 26024 11946 26036
rect 16574 26024 16580 26036
rect 11940 25996 12480 26024
rect 11940 25984 11946 25996
rect 10689 25959 10747 25965
rect 10284 25928 10548 25956
rect 10284 25916 10290 25928
rect 9950 25848 9956 25900
rect 10008 25888 10014 25900
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 10008 25860 10333 25888
rect 10008 25848 10014 25860
rect 10321 25857 10333 25860
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 9769 25823 9827 25829
rect 9769 25789 9781 25823
rect 9815 25789 9827 25823
rect 9769 25783 9827 25789
rect 10229 25823 10287 25829
rect 10229 25789 10241 25823
rect 10275 25820 10287 25823
rect 10410 25820 10416 25832
rect 10275 25792 10416 25820
rect 10275 25789 10287 25792
rect 10229 25783 10287 25789
rect 9784 25752 9812 25783
rect 10410 25780 10416 25792
rect 10468 25780 10474 25832
rect 10520 25820 10548 25928
rect 10689 25925 10701 25959
rect 10735 25925 10747 25959
rect 10689 25919 10747 25925
rect 10778 25916 10784 25968
rect 10836 25916 10842 25968
rect 10980 25928 11928 25956
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25888 10655 25891
rect 10870 25888 10876 25900
rect 10643 25860 10876 25888
rect 10643 25857 10655 25860
rect 10597 25851 10655 25857
rect 10870 25848 10876 25860
rect 10928 25848 10934 25900
rect 10980 25897 11008 25928
rect 10965 25891 11023 25897
rect 10965 25857 10977 25891
rect 11011 25857 11023 25891
rect 10965 25851 11023 25857
rect 11514 25848 11520 25900
rect 11572 25848 11578 25900
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11146 25820 11152 25832
rect 10520 25792 11152 25820
rect 11146 25780 11152 25792
rect 11204 25780 11210 25832
rect 10045 25755 10103 25761
rect 10045 25752 10057 25755
rect 9784 25724 10057 25752
rect 10045 25721 10057 25724
rect 10091 25721 10103 25755
rect 10045 25715 10103 25721
rect 10134 25712 10140 25764
rect 10192 25752 10198 25764
rect 10686 25752 10692 25764
rect 10192 25724 10692 25752
rect 10192 25712 10198 25724
rect 10686 25712 10692 25724
rect 10744 25752 10750 25764
rect 11716 25752 11744 25851
rect 11900 25832 11928 25928
rect 12066 25848 12072 25900
rect 12124 25848 12130 25900
rect 12158 25848 12164 25900
rect 12216 25888 12222 25900
rect 12452 25897 12480 25996
rect 16240 25996 16580 26024
rect 12618 25916 12624 25968
rect 12676 25956 12682 25968
rect 12805 25959 12863 25965
rect 12805 25956 12817 25959
rect 12676 25928 12817 25956
rect 12676 25916 12682 25928
rect 12805 25925 12817 25928
rect 12851 25925 12863 25959
rect 12805 25919 12863 25925
rect 12253 25891 12311 25897
rect 12253 25888 12265 25891
rect 12216 25860 12265 25888
rect 12216 25848 12222 25860
rect 12253 25857 12265 25860
rect 12299 25857 12311 25891
rect 12253 25851 12311 25857
rect 12437 25891 12495 25897
rect 12437 25857 12449 25891
rect 12483 25857 12495 25891
rect 12437 25851 12495 25857
rect 11793 25823 11851 25829
rect 11793 25789 11805 25823
rect 11839 25789 11851 25823
rect 11793 25783 11851 25789
rect 10744 25724 11744 25752
rect 11808 25752 11836 25783
rect 11882 25780 11888 25832
rect 11940 25780 11946 25832
rect 12452 25820 12480 25851
rect 12526 25848 12532 25900
rect 12584 25848 12590 25900
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 12986 25897 12992 25900
rect 12943 25891 12992 25897
rect 12943 25857 12955 25891
rect 12989 25857 12992 25891
rect 12943 25851 12992 25857
rect 12986 25848 12992 25851
rect 13044 25888 13050 25900
rect 13630 25888 13636 25900
rect 13044 25860 13636 25888
rect 13044 25848 13050 25860
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 15746 25848 15752 25900
rect 15804 25848 15810 25900
rect 15930 25848 15936 25900
rect 15988 25888 15994 25900
rect 16114 25888 16120 25900
rect 15988 25860 16120 25888
rect 15988 25848 15994 25860
rect 16114 25848 16120 25860
rect 16172 25848 16178 25900
rect 16240 25897 16268 25996
rect 16574 25984 16580 25996
rect 16632 26024 16638 26036
rect 18877 26027 18935 26033
rect 16632 25996 17172 26024
rect 16632 25984 16638 25996
rect 16209 25891 16268 25897
rect 16209 25857 16221 25891
rect 16255 25860 16268 25891
rect 16255 25857 16267 25860
rect 16209 25851 16267 25857
rect 16298 25848 16304 25900
rect 16356 25848 16362 25900
rect 17144 25897 17172 25996
rect 18877 25993 18889 26027
rect 18923 26024 18935 26027
rect 19518 26024 19524 26036
rect 18923 25996 19524 26024
rect 18923 25993 18935 25996
rect 18877 25987 18935 25993
rect 17770 25916 17776 25968
rect 17828 25956 17834 25968
rect 18230 25965 18236 25968
rect 18224 25956 18236 25965
rect 17828 25928 18000 25956
rect 18191 25928 18236 25956
rect 17828 25916 17834 25928
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25888 17187 25891
rect 17402 25888 17408 25900
rect 17175 25860 17408 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17402 25848 17408 25860
rect 17460 25848 17466 25900
rect 17497 25891 17555 25897
rect 17497 25857 17509 25891
rect 17543 25888 17555 25891
rect 17586 25888 17592 25900
rect 17543 25860 17592 25888
rect 17543 25857 17555 25860
rect 17497 25851 17555 25857
rect 17586 25848 17592 25860
rect 17644 25848 17650 25900
rect 17681 25891 17739 25897
rect 17681 25857 17693 25891
rect 17727 25888 17739 25891
rect 17862 25888 17868 25900
rect 17727 25860 17868 25888
rect 17727 25857 17739 25860
rect 17681 25851 17739 25857
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 17972 25897 18000 25928
rect 18224 25919 18236 25928
rect 18230 25916 18236 25919
rect 18288 25916 18294 25968
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25857 18015 25891
rect 17957 25851 18015 25857
rect 18601 25891 18659 25897
rect 18601 25857 18613 25891
rect 18647 25888 18659 25891
rect 18693 25891 18751 25897
rect 18693 25888 18705 25891
rect 18647 25860 18705 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 18693 25857 18705 25860
rect 18739 25888 18751 25891
rect 18782 25888 18788 25900
rect 18739 25860 18788 25888
rect 18739 25857 18751 25860
rect 18693 25851 18751 25857
rect 18782 25848 18788 25860
rect 18840 25848 18846 25900
rect 12618 25820 12624 25832
rect 12452 25792 12624 25820
rect 12618 25780 12624 25792
rect 12676 25780 12682 25832
rect 16025 25823 16083 25829
rect 16025 25789 16037 25823
rect 16071 25789 16083 25823
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16025 25783 16083 25789
rect 16316 25792 16681 25820
rect 12158 25752 12164 25764
rect 11808 25724 12164 25752
rect 10744 25712 10750 25724
rect 12158 25712 12164 25724
rect 12216 25712 12222 25764
rect 12710 25712 12716 25764
rect 12768 25752 12774 25764
rect 13538 25752 13544 25764
rect 12768 25724 13544 25752
rect 12768 25712 12774 25724
rect 13538 25712 13544 25724
rect 13596 25712 13602 25764
rect 12526 25684 12532 25696
rect 9416 25656 12532 25684
rect 12526 25644 12532 25656
rect 12584 25644 12590 25696
rect 13081 25687 13139 25693
rect 13081 25653 13093 25687
rect 13127 25684 13139 25687
rect 13354 25684 13360 25696
rect 13127 25656 13360 25684
rect 13127 25653 13139 25656
rect 13081 25647 13139 25653
rect 13354 25644 13360 25656
rect 13412 25644 13418 25696
rect 14642 25644 14648 25696
rect 14700 25684 14706 25696
rect 15102 25684 15108 25696
rect 14700 25656 15108 25684
rect 14700 25644 14706 25656
rect 15102 25644 15108 25656
rect 15160 25684 15166 25696
rect 15565 25687 15623 25693
rect 15565 25684 15577 25687
rect 15160 25656 15577 25684
rect 15160 25644 15166 25656
rect 15565 25653 15577 25656
rect 15611 25653 15623 25687
rect 16040 25684 16068 25783
rect 16316 25761 16344 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 16669 25783 16727 25789
rect 17034 25780 17040 25832
rect 17092 25780 17098 25832
rect 17770 25780 17776 25832
rect 17828 25820 17834 25832
rect 18138 25820 18144 25832
rect 17828 25792 18144 25820
rect 17828 25780 17834 25792
rect 18138 25780 18144 25792
rect 18196 25780 18202 25832
rect 16301 25755 16359 25761
rect 16301 25721 16313 25755
rect 16347 25721 16359 25755
rect 16301 25715 16359 25721
rect 16390 25712 16396 25764
rect 16448 25752 16454 25764
rect 16761 25755 16819 25761
rect 16761 25752 16773 25755
rect 16448 25724 16773 25752
rect 16448 25712 16454 25724
rect 16761 25721 16773 25724
rect 16807 25721 16819 25755
rect 18892 25752 18920 25987
rect 19518 25984 19524 25996
rect 19576 26024 19582 26036
rect 19613 26027 19671 26033
rect 19613 26024 19625 26027
rect 19576 25996 19625 26024
rect 19576 25984 19582 25996
rect 19613 25993 19625 25996
rect 19659 25993 19671 26027
rect 19613 25987 19671 25993
rect 20346 25984 20352 26036
rect 20404 26024 20410 26036
rect 22094 26024 22100 26036
rect 20404 25996 22100 26024
rect 20404 25984 20410 25996
rect 22094 25984 22100 25996
rect 22152 26024 22158 26036
rect 23290 26024 23296 26036
rect 22152 25996 23296 26024
rect 22152 25984 22158 25996
rect 23290 25984 23296 25996
rect 23348 26024 23354 26036
rect 23401 26027 23459 26033
rect 23401 26024 23413 26027
rect 23348 25996 23413 26024
rect 23348 25984 23354 25996
rect 23401 25993 23413 25996
rect 23447 25993 23459 26027
rect 23401 25987 23459 25993
rect 23566 25984 23572 26036
rect 23624 25984 23630 26036
rect 23842 25984 23848 26036
rect 23900 26024 23906 26036
rect 24949 26027 25007 26033
rect 24949 26024 24961 26027
rect 23900 25996 24164 26024
rect 23900 25984 23906 25996
rect 24136 25965 24164 25996
rect 24780 25996 24961 26024
rect 23201 25959 23259 25965
rect 23201 25934 23213 25959
rect 23247 25934 23259 25959
rect 24121 25959 24179 25965
rect 18969 25891 19027 25897
rect 18969 25857 18981 25891
rect 19015 25888 19027 25891
rect 19058 25888 19064 25900
rect 19015 25860 19064 25888
rect 19015 25857 19027 25860
rect 18969 25851 19027 25857
rect 19058 25848 19064 25860
rect 19116 25848 19122 25900
rect 19613 25891 19671 25897
rect 19613 25857 19625 25891
rect 19659 25888 19671 25891
rect 19702 25888 19708 25900
rect 19659 25860 19708 25888
rect 19659 25857 19671 25860
rect 19613 25851 19671 25857
rect 19702 25848 19708 25860
rect 19760 25848 19766 25900
rect 23198 25882 23204 25934
rect 23256 25882 23262 25934
rect 24121 25925 24133 25959
rect 24167 25925 24179 25959
rect 24121 25919 24179 25925
rect 24213 25959 24271 25965
rect 24213 25925 24225 25959
rect 24259 25956 24271 25959
rect 24780 25956 24808 25996
rect 24949 25993 24961 25996
rect 24995 26024 25007 26027
rect 25130 26024 25136 26036
rect 24995 25996 25136 26024
rect 24995 25993 25007 25996
rect 24949 25987 25007 25993
rect 25130 25984 25136 25996
rect 25188 25984 25194 26036
rect 25774 25984 25780 26036
rect 25832 26024 25838 26036
rect 32030 26024 32036 26036
rect 25832 25996 32036 26024
rect 25832 25984 25838 25996
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 32122 25984 32128 26036
rect 32180 26024 32186 26036
rect 32490 26024 32496 26036
rect 32180 25996 32496 26024
rect 32180 25984 32186 25996
rect 32490 25984 32496 25996
rect 32548 26024 32554 26036
rect 32677 26027 32735 26033
rect 32677 26024 32689 26027
rect 32548 25996 32689 26024
rect 32548 25984 32554 25996
rect 32677 25993 32689 25996
rect 32723 25993 32735 26027
rect 33226 26024 33232 26036
rect 32677 25987 32735 25993
rect 33060 25996 33232 26024
rect 26418 25956 26424 25968
rect 24259 25928 24808 25956
rect 26160 25928 26424 25956
rect 24259 25925 24271 25928
rect 24213 25919 24271 25925
rect 23842 25848 23848 25900
rect 23900 25848 23906 25900
rect 23993 25891 24051 25897
rect 23993 25857 24005 25891
rect 24039 25888 24051 25891
rect 24039 25857 24072 25888
rect 23993 25851 24072 25857
rect 19426 25780 19432 25832
rect 19484 25780 19490 25832
rect 19978 25780 19984 25832
rect 20036 25780 20042 25832
rect 24044 25820 24072 25851
rect 24302 25848 24308 25900
rect 24360 25897 24366 25900
rect 24360 25851 24368 25897
rect 24360 25848 24366 25851
rect 24486 25848 24492 25900
rect 24544 25888 24550 25900
rect 24765 25891 24823 25897
rect 24765 25888 24777 25891
rect 24544 25860 24777 25888
rect 24544 25848 24550 25860
rect 24765 25857 24777 25860
rect 24811 25857 24823 25891
rect 24765 25851 24823 25857
rect 25041 25891 25099 25897
rect 25041 25857 25053 25891
rect 25087 25888 25099 25891
rect 25314 25888 25320 25900
rect 25087 25860 25320 25888
rect 25087 25857 25099 25860
rect 25041 25851 25099 25857
rect 24578 25820 24584 25832
rect 24044 25792 24584 25820
rect 16761 25715 16819 25721
rect 18248 25724 18920 25752
rect 17862 25684 17868 25696
rect 16040 25656 17868 25684
rect 15565 25647 15623 25653
rect 17862 25644 17868 25656
rect 17920 25644 17926 25696
rect 18248 25693 18276 25724
rect 19150 25712 19156 25764
rect 19208 25752 19214 25764
rect 21542 25752 21548 25764
rect 19208 25724 21548 25752
rect 19208 25712 19214 25724
rect 21542 25712 21548 25724
rect 21600 25712 21606 25764
rect 23750 25712 23756 25764
rect 23808 25752 23814 25764
rect 24044 25752 24072 25792
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 23808 25724 24072 25752
rect 23808 25712 23814 25724
rect 24486 25712 24492 25764
rect 24544 25712 24550 25764
rect 24762 25712 24768 25764
rect 24820 25752 24826 25764
rect 25056 25752 25084 25851
rect 25314 25848 25320 25860
rect 25372 25848 25378 25900
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25888 25651 25891
rect 25682 25888 25688 25900
rect 25639 25860 25688 25888
rect 25639 25857 25651 25860
rect 25593 25851 25651 25857
rect 25682 25848 25688 25860
rect 25740 25848 25746 25900
rect 25777 25891 25835 25897
rect 25777 25857 25789 25891
rect 25823 25888 25835 25891
rect 25958 25888 25964 25900
rect 25823 25860 25964 25888
rect 25823 25857 25835 25860
rect 25777 25851 25835 25857
rect 25958 25848 25964 25860
rect 26016 25848 26022 25900
rect 26160 25897 26188 25928
rect 26418 25916 26424 25928
rect 26476 25916 26482 25968
rect 26878 25916 26884 25968
rect 26936 25956 26942 25968
rect 27614 25956 27620 25968
rect 26936 25928 27384 25956
rect 26936 25916 26942 25928
rect 26145 25891 26203 25897
rect 26145 25857 26157 25891
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26234 25848 26240 25900
rect 26292 25848 26298 25900
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 26513 25891 26571 25897
rect 26513 25857 26525 25891
rect 26559 25888 26571 25891
rect 26970 25888 26976 25900
rect 26559 25860 26976 25888
rect 26559 25857 26571 25860
rect 26513 25851 26571 25857
rect 25406 25780 25412 25832
rect 25464 25820 25470 25832
rect 26344 25820 26372 25851
rect 26970 25848 26976 25860
rect 27028 25848 27034 25900
rect 27157 25891 27215 25897
rect 27157 25857 27169 25891
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 27249 25891 27307 25897
rect 27249 25857 27261 25891
rect 27295 25857 27307 25891
rect 27249 25851 27307 25857
rect 27172 25820 27200 25851
rect 25464 25792 27200 25820
rect 25464 25780 25470 25792
rect 24820 25724 25084 25752
rect 24820 25712 24826 25724
rect 25130 25712 25136 25764
rect 25188 25752 25194 25764
rect 25869 25755 25927 25761
rect 25869 25752 25881 25755
rect 25188 25724 25881 25752
rect 25188 25712 25194 25724
rect 25869 25721 25881 25724
rect 25915 25721 25927 25755
rect 27264 25752 27292 25851
rect 27356 25820 27384 25928
rect 27448 25928 27620 25956
rect 27448 25897 27476 25928
rect 27614 25916 27620 25928
rect 27672 25956 27678 25968
rect 27982 25956 27988 25968
rect 27672 25928 27988 25956
rect 27672 25916 27678 25928
rect 27982 25916 27988 25928
rect 28040 25916 28046 25968
rect 28997 25959 29055 25965
rect 28997 25925 29009 25959
rect 29043 25956 29055 25959
rect 29270 25956 29276 25968
rect 29043 25928 29276 25956
rect 29043 25925 29055 25928
rect 28997 25919 29055 25925
rect 29270 25916 29276 25928
rect 29328 25916 29334 25968
rect 29454 25916 29460 25968
rect 29512 25956 29518 25968
rect 30101 25959 30159 25965
rect 29512 25928 29776 25956
rect 29512 25916 29518 25928
rect 27433 25891 27491 25897
rect 27433 25857 27445 25891
rect 27479 25857 27491 25891
rect 27433 25851 27491 25857
rect 27522 25848 27528 25900
rect 27580 25848 27586 25900
rect 28718 25848 28724 25900
rect 28776 25897 28782 25900
rect 29748 25897 29776 25928
rect 30101 25925 30113 25959
rect 30147 25956 30159 25959
rect 30190 25956 30196 25968
rect 30147 25928 30196 25956
rect 30147 25925 30159 25928
rect 30101 25919 30159 25925
rect 30190 25916 30196 25928
rect 30248 25916 30254 25968
rect 30285 25959 30343 25965
rect 30285 25925 30297 25959
rect 30331 25925 30343 25959
rect 30285 25919 30343 25925
rect 31573 25959 31631 25965
rect 31573 25925 31585 25959
rect 31619 25956 31631 25959
rect 32217 25959 32275 25965
rect 32217 25956 32229 25959
rect 31619 25928 32229 25956
rect 31619 25925 31631 25928
rect 31573 25919 31631 25925
rect 32217 25925 32229 25928
rect 32263 25956 32275 25959
rect 32306 25956 32312 25968
rect 32263 25928 32312 25956
rect 32263 25925 32275 25928
rect 32217 25919 32275 25925
rect 28776 25891 28825 25897
rect 28776 25857 28779 25891
rect 28813 25857 28825 25891
rect 28776 25851 28825 25857
rect 28905 25891 28963 25897
rect 28905 25857 28917 25891
rect 28951 25857 28963 25891
rect 28905 25851 28963 25857
rect 29089 25891 29147 25897
rect 29089 25857 29101 25891
rect 29135 25857 29147 25891
rect 29089 25851 29147 25857
rect 29549 25891 29607 25897
rect 29549 25857 29561 25891
rect 29595 25857 29607 25891
rect 29549 25851 29607 25857
rect 29733 25891 29791 25897
rect 29733 25857 29745 25891
rect 29779 25888 29791 25891
rect 29914 25888 29920 25900
rect 29779 25860 29920 25888
rect 29779 25857 29791 25860
rect 29733 25851 29791 25857
rect 28776 25848 28782 25851
rect 28629 25823 28687 25829
rect 28629 25820 28641 25823
rect 27356 25792 28641 25820
rect 28629 25789 28641 25792
rect 28675 25789 28687 25823
rect 28920 25820 28948 25851
rect 28994 25820 29000 25832
rect 28920 25792 29000 25820
rect 28629 25783 28687 25789
rect 28994 25780 29000 25792
rect 29052 25780 29058 25832
rect 28166 25752 28172 25764
rect 27264 25724 28172 25752
rect 25869 25715 25927 25721
rect 28166 25712 28172 25724
rect 28224 25712 28230 25764
rect 29104 25752 29132 25851
rect 29564 25820 29592 25851
rect 29914 25848 29920 25860
rect 29972 25848 29978 25900
rect 30006 25848 30012 25900
rect 30064 25888 30070 25900
rect 30300 25888 30328 25919
rect 32306 25916 32312 25928
rect 32364 25916 32370 25968
rect 30064 25860 30328 25888
rect 30064 25848 30070 25860
rect 31754 25848 31760 25900
rect 31812 25848 31818 25900
rect 31938 25848 31944 25900
rect 31996 25848 32002 25900
rect 32122 25848 32128 25900
rect 32180 25888 32186 25900
rect 32401 25891 32459 25897
rect 32401 25888 32413 25891
rect 32180 25860 32413 25888
rect 32180 25848 32186 25860
rect 32401 25857 32413 25860
rect 32447 25857 32459 25891
rect 32401 25851 32459 25857
rect 32861 25891 32919 25897
rect 32861 25857 32873 25891
rect 32907 25888 32919 25891
rect 33060 25888 33088 25996
rect 33226 25984 33232 25996
rect 33284 25984 33290 26036
rect 33505 26027 33563 26033
rect 33505 25993 33517 26027
rect 33551 26024 33563 26027
rect 33594 26024 33600 26036
rect 33551 25996 33600 26024
rect 33551 25993 33563 25996
rect 33505 25987 33563 25993
rect 33594 25984 33600 25996
rect 33652 25984 33658 26036
rect 34514 25984 34520 26036
rect 34572 25984 34578 26036
rect 33962 25916 33968 25968
rect 34020 25916 34026 25968
rect 34532 25956 34560 25984
rect 34532 25928 34744 25956
rect 32907 25860 33088 25888
rect 32907 25857 32919 25860
rect 32861 25851 32919 25857
rect 33134 25848 33140 25900
rect 33192 25848 33198 25900
rect 33318 25848 33324 25900
rect 33376 25848 33382 25900
rect 33689 25891 33747 25897
rect 33689 25857 33701 25891
rect 33735 25888 33747 25891
rect 34054 25888 34060 25900
rect 33735 25860 34060 25888
rect 33735 25857 33747 25860
rect 33689 25851 33747 25857
rect 34054 25848 34060 25860
rect 34112 25848 34118 25900
rect 34238 25848 34244 25900
rect 34296 25888 34302 25900
rect 34425 25891 34483 25897
rect 34425 25888 34437 25891
rect 34296 25860 34437 25888
rect 34296 25848 34302 25860
rect 34425 25857 34437 25860
rect 34471 25857 34483 25891
rect 34425 25851 34483 25857
rect 34514 25848 34520 25900
rect 34572 25848 34578 25900
rect 34716 25897 34744 25928
rect 35066 25916 35072 25968
rect 35124 25956 35130 25968
rect 35618 25956 35624 25968
rect 35124 25928 35624 25956
rect 35124 25916 35130 25928
rect 35618 25916 35624 25928
rect 35676 25916 35682 25968
rect 34701 25891 34759 25897
rect 34701 25857 34713 25891
rect 34747 25888 34759 25891
rect 35161 25891 35219 25897
rect 35161 25888 35173 25891
rect 34747 25860 35173 25888
rect 34747 25857 34759 25860
rect 34701 25851 34759 25857
rect 35161 25857 35173 25860
rect 35207 25857 35219 25891
rect 35161 25851 35219 25857
rect 35250 25848 35256 25900
rect 35308 25888 35314 25900
rect 35437 25891 35495 25897
rect 35437 25888 35449 25891
rect 35308 25860 35449 25888
rect 35308 25848 35314 25860
rect 35437 25857 35449 25860
rect 35483 25888 35495 25891
rect 35710 25888 35716 25900
rect 35483 25860 35716 25888
rect 35483 25857 35495 25860
rect 35437 25851 35495 25857
rect 35710 25848 35716 25860
rect 35768 25848 35774 25900
rect 31018 25820 31024 25832
rect 29564 25792 31024 25820
rect 31018 25780 31024 25792
rect 31076 25820 31082 25832
rect 31849 25823 31907 25829
rect 31849 25820 31861 25823
rect 31076 25792 31861 25820
rect 31076 25780 31082 25792
rect 31849 25789 31861 25792
rect 31895 25789 31907 25823
rect 31849 25783 31907 25789
rect 33042 25780 33048 25832
rect 33100 25820 33106 25832
rect 33594 25820 33600 25832
rect 33100 25792 33600 25820
rect 33100 25780 33106 25792
rect 33594 25780 33600 25792
rect 33652 25780 33658 25832
rect 33781 25823 33839 25829
rect 33781 25789 33793 25823
rect 33827 25789 33839 25823
rect 33781 25783 33839 25789
rect 29104 25724 29408 25752
rect 18233 25687 18291 25693
rect 18233 25653 18245 25687
rect 18279 25653 18291 25687
rect 18233 25647 18291 25653
rect 18690 25644 18696 25696
rect 18748 25644 18754 25696
rect 19794 25644 19800 25696
rect 19852 25684 19858 25696
rect 23290 25684 23296 25696
rect 19852 25656 23296 25684
rect 19852 25644 19858 25656
rect 23290 25644 23296 25656
rect 23348 25644 23354 25696
rect 23382 25644 23388 25696
rect 23440 25644 23446 25696
rect 23658 25644 23664 25696
rect 23716 25684 23722 25696
rect 24581 25687 24639 25693
rect 24581 25684 24593 25687
rect 23716 25656 24593 25684
rect 23716 25644 23722 25656
rect 24581 25653 24593 25656
rect 24627 25653 24639 25687
rect 24581 25647 24639 25653
rect 26973 25687 27031 25693
rect 26973 25653 26985 25687
rect 27019 25684 27031 25687
rect 27338 25684 27344 25696
rect 27019 25656 27344 25684
rect 27019 25653 27031 25656
rect 26973 25647 27031 25653
rect 27338 25644 27344 25656
rect 27396 25644 27402 25696
rect 29270 25644 29276 25696
rect 29328 25644 29334 25696
rect 29380 25684 29408 25724
rect 29454 25712 29460 25764
rect 29512 25712 29518 25764
rect 29546 25712 29552 25764
rect 29604 25752 29610 25764
rect 32490 25752 32496 25764
rect 29604 25724 32496 25752
rect 29604 25712 29610 25724
rect 32490 25712 32496 25724
rect 32548 25712 32554 25764
rect 32674 25712 32680 25764
rect 32732 25752 32738 25764
rect 32858 25752 32864 25764
rect 32732 25724 32864 25752
rect 32732 25712 32738 25724
rect 32858 25712 32864 25724
rect 32916 25712 32922 25764
rect 33410 25712 33416 25764
rect 33468 25752 33474 25764
rect 33796 25752 33824 25783
rect 33962 25780 33968 25832
rect 34020 25820 34026 25832
rect 34333 25823 34391 25829
rect 34333 25820 34345 25823
rect 34020 25792 34345 25820
rect 34020 25780 34026 25792
rect 34333 25789 34345 25792
rect 34379 25820 34391 25823
rect 35342 25820 35348 25832
rect 34379 25792 35348 25820
rect 34379 25789 34391 25792
rect 34333 25783 34391 25789
rect 35342 25780 35348 25792
rect 35400 25780 35406 25832
rect 34422 25752 34428 25764
rect 33468 25724 33824 25752
rect 33980 25724 34428 25752
rect 33468 25712 33474 25724
rect 29730 25684 29736 25696
rect 29380 25656 29736 25684
rect 29730 25644 29736 25656
rect 29788 25644 29794 25696
rect 29914 25644 29920 25696
rect 29972 25644 29978 25696
rect 30101 25687 30159 25693
rect 30101 25653 30113 25687
rect 30147 25684 30159 25687
rect 30742 25684 30748 25696
rect 30147 25656 30748 25684
rect 30147 25653 30159 25656
rect 30101 25647 30159 25653
rect 30742 25644 30748 25656
rect 30800 25644 30806 25696
rect 31481 25687 31539 25693
rect 31481 25653 31493 25687
rect 31527 25684 31539 25687
rect 31846 25684 31852 25696
rect 31527 25656 31852 25684
rect 31527 25653 31539 25656
rect 31481 25647 31539 25653
rect 31846 25644 31852 25656
rect 31904 25644 31910 25696
rect 32214 25644 32220 25696
rect 32272 25684 32278 25696
rect 33980 25693 34008 25724
rect 34422 25712 34428 25724
rect 34480 25712 34486 25764
rect 35158 25712 35164 25764
rect 35216 25752 35222 25764
rect 35526 25752 35532 25764
rect 35216 25724 35532 25752
rect 35216 25712 35222 25724
rect 35526 25712 35532 25724
rect 35584 25712 35590 25764
rect 33321 25687 33379 25693
rect 33321 25684 33333 25687
rect 32272 25656 33333 25684
rect 32272 25644 32278 25656
rect 33321 25653 33333 25656
rect 33367 25653 33379 25687
rect 33321 25647 33379 25653
rect 33965 25687 34023 25693
rect 33965 25653 33977 25687
rect 34011 25653 34023 25687
rect 33965 25647 34023 25653
rect 34054 25644 34060 25696
rect 34112 25644 34118 25696
rect 34238 25644 34244 25696
rect 34296 25684 34302 25696
rect 34517 25687 34575 25693
rect 34517 25684 34529 25687
rect 34296 25656 34529 25684
rect 34296 25644 34302 25656
rect 34517 25653 34529 25656
rect 34563 25653 34575 25687
rect 34517 25647 34575 25653
rect 34790 25644 34796 25696
rect 34848 25684 34854 25696
rect 35345 25687 35403 25693
rect 35345 25684 35357 25687
rect 34848 25656 35357 25684
rect 34848 25644 34854 25656
rect 35345 25653 35357 25656
rect 35391 25653 35403 25687
rect 35345 25647 35403 25653
rect 1104 25594 36524 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 36524 25594
rect 1104 25520 36524 25542
rect 2222 25440 2228 25492
rect 2280 25440 2286 25492
rect 3878 25440 3884 25492
rect 3936 25440 3942 25492
rect 6638 25440 6644 25492
rect 6696 25480 6702 25492
rect 6825 25483 6883 25489
rect 6825 25480 6837 25483
rect 6696 25452 6837 25480
rect 6696 25440 6702 25452
rect 6825 25449 6837 25452
rect 6871 25449 6883 25483
rect 9306 25480 9312 25492
rect 6825 25443 6883 25449
rect 6932 25452 9312 25480
rect 2608 25384 6408 25412
rect 2406 25100 2412 25152
rect 2464 25140 2470 25152
rect 2608 25149 2636 25384
rect 2869 25347 2927 25353
rect 2869 25313 2881 25347
rect 2915 25344 2927 25347
rect 3050 25344 3056 25356
rect 2915 25316 3056 25344
rect 2915 25313 2927 25316
rect 2869 25307 2927 25313
rect 3050 25304 3056 25316
rect 3108 25344 3114 25356
rect 3786 25344 3792 25356
rect 3108 25316 3792 25344
rect 3108 25304 3114 25316
rect 3786 25304 3792 25316
rect 3844 25344 3850 25356
rect 4433 25347 4491 25353
rect 4433 25344 4445 25347
rect 3844 25316 4445 25344
rect 3844 25304 3850 25316
rect 4433 25313 4445 25316
rect 4479 25313 4491 25347
rect 4433 25307 4491 25313
rect 5353 25347 5411 25353
rect 5353 25313 5365 25347
rect 5399 25344 5411 25347
rect 6178 25344 6184 25356
rect 5399 25316 6184 25344
rect 5399 25313 5411 25316
rect 5353 25307 5411 25313
rect 6178 25304 6184 25316
rect 6236 25304 6242 25356
rect 6270 25304 6276 25356
rect 6328 25304 6334 25356
rect 6380 25353 6408 25384
rect 6365 25347 6423 25353
rect 6365 25313 6377 25347
rect 6411 25344 6423 25347
rect 6932 25344 6960 25452
rect 9306 25440 9312 25452
rect 9364 25440 9370 25492
rect 9769 25483 9827 25489
rect 9769 25449 9781 25483
rect 9815 25480 9827 25483
rect 9858 25480 9864 25492
rect 9815 25452 9864 25480
rect 9815 25449 9827 25452
rect 9769 25443 9827 25449
rect 9858 25440 9864 25452
rect 9916 25440 9922 25492
rect 10594 25440 10600 25492
rect 10652 25480 10658 25492
rect 11241 25483 11299 25489
rect 11241 25480 11253 25483
rect 10652 25452 11253 25480
rect 10652 25440 10658 25452
rect 11241 25449 11253 25452
rect 11287 25449 11299 25483
rect 11241 25443 11299 25449
rect 13630 25440 13636 25492
rect 13688 25480 13694 25492
rect 15194 25480 15200 25492
rect 13688 25452 15200 25480
rect 13688 25440 13694 25452
rect 15194 25440 15200 25452
rect 15252 25480 15258 25492
rect 15470 25480 15476 25492
rect 15252 25452 15476 25480
rect 15252 25440 15258 25452
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 17221 25483 17279 25489
rect 17221 25449 17233 25483
rect 17267 25480 17279 25483
rect 17494 25480 17500 25492
rect 17267 25452 17500 25480
rect 17267 25449 17279 25452
rect 17221 25443 17279 25449
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 17862 25440 17868 25492
rect 17920 25480 17926 25492
rect 17920 25452 19104 25480
rect 17920 25440 17926 25452
rect 7760 25384 8340 25412
rect 7650 25344 7656 25356
rect 6411 25316 6960 25344
rect 7274 25316 7656 25344
rect 6411 25313 6423 25316
rect 6365 25307 6423 25313
rect 2685 25279 2743 25285
rect 2685 25245 2697 25279
rect 2731 25276 2743 25279
rect 3142 25276 3148 25288
rect 2731 25248 3148 25276
rect 2731 25245 2743 25248
rect 2685 25239 2743 25245
rect 3142 25236 3148 25248
rect 3200 25236 3206 25288
rect 5626 25236 5632 25288
rect 5684 25236 5690 25288
rect 5721 25279 5779 25285
rect 5721 25245 5733 25279
rect 5767 25276 5779 25279
rect 5767 25248 5948 25276
rect 5767 25245 5779 25248
rect 5721 25239 5779 25245
rect 5920 25220 5948 25248
rect 5994 25236 6000 25288
rect 6052 25236 6058 25288
rect 6457 25279 6515 25285
rect 6457 25245 6469 25279
rect 6503 25276 6515 25279
rect 7006 25276 7012 25288
rect 6503 25248 7012 25276
rect 6503 25245 6515 25248
rect 6457 25239 6515 25245
rect 7006 25236 7012 25248
rect 7064 25236 7070 25288
rect 7274 25285 7302 25316
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 7101 25279 7159 25285
rect 7101 25245 7113 25279
rect 7147 25245 7159 25279
rect 7101 25239 7159 25245
rect 7259 25279 7317 25285
rect 7259 25245 7271 25279
rect 7305 25245 7317 25279
rect 7259 25239 7317 25245
rect 7561 25279 7619 25285
rect 7561 25245 7573 25279
rect 7607 25276 7619 25279
rect 7760 25276 7788 25384
rect 7837 25347 7895 25353
rect 7837 25313 7849 25347
rect 7883 25344 7895 25347
rect 8202 25344 8208 25356
rect 7883 25316 8208 25344
rect 7883 25313 7895 25316
rect 7837 25307 7895 25313
rect 8202 25304 8208 25316
rect 8260 25304 8266 25356
rect 8312 25285 8340 25384
rect 8478 25372 8484 25424
rect 8536 25372 8542 25424
rect 8938 25372 8944 25424
rect 8996 25372 9002 25424
rect 11606 25412 11612 25424
rect 9324 25384 11612 25412
rect 9324 25353 9352 25384
rect 11606 25372 11612 25384
rect 11664 25372 11670 25424
rect 14093 25415 14151 25421
rect 14093 25381 14105 25415
rect 14139 25381 14151 25415
rect 15378 25412 15384 25424
rect 14093 25375 14151 25381
rect 15304 25384 15384 25412
rect 9309 25347 9367 25353
rect 9309 25313 9321 25347
rect 9355 25313 9367 25347
rect 9309 25307 9367 25313
rect 8297 25279 8355 25285
rect 7607 25248 7788 25276
rect 7852 25248 8248 25276
rect 7607 25245 7619 25248
rect 7561 25239 7619 25245
rect 5810 25168 5816 25220
rect 5868 25168 5874 25220
rect 5902 25168 5908 25220
rect 5960 25208 5966 25220
rect 7116 25208 7144 25239
rect 5960 25180 7144 25208
rect 7377 25211 7435 25217
rect 5960 25168 5966 25180
rect 7377 25177 7389 25211
rect 7423 25177 7435 25211
rect 7377 25171 7435 25177
rect 7469 25211 7527 25217
rect 7469 25177 7481 25211
rect 7515 25208 7527 25211
rect 7852 25208 7880 25248
rect 8018 25217 8024 25220
rect 7515 25180 7880 25208
rect 7995 25211 8024 25217
rect 7515 25177 7527 25180
rect 7469 25171 7527 25177
rect 7995 25177 8007 25211
rect 7995 25171 8024 25177
rect 2593 25143 2651 25149
rect 2593 25140 2605 25143
rect 2464 25112 2605 25140
rect 2464 25100 2470 25112
rect 2593 25109 2605 25112
rect 2639 25109 2651 25143
rect 2593 25103 2651 25109
rect 3970 25100 3976 25152
rect 4028 25140 4034 25152
rect 4249 25143 4307 25149
rect 4249 25140 4261 25143
rect 4028 25112 4261 25140
rect 4028 25100 4034 25112
rect 4249 25109 4261 25112
rect 4295 25109 4307 25143
rect 4249 25103 4307 25109
rect 4341 25143 4399 25149
rect 4341 25109 4353 25143
rect 4387 25140 4399 25143
rect 4709 25143 4767 25149
rect 4709 25140 4721 25143
rect 4387 25112 4721 25140
rect 4387 25109 4399 25112
rect 4341 25103 4399 25109
rect 4709 25109 4721 25112
rect 4755 25109 4767 25143
rect 4709 25103 4767 25109
rect 5445 25143 5503 25149
rect 5445 25109 5457 25143
rect 5491 25140 5503 25143
rect 5626 25140 5632 25152
rect 5491 25112 5632 25140
rect 5491 25109 5503 25112
rect 5445 25103 5503 25109
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 6454 25100 6460 25152
rect 6512 25140 6518 25152
rect 7392 25140 7420 25171
rect 8018 25168 8024 25171
rect 8076 25168 8082 25220
rect 8110 25168 8116 25220
rect 8168 25168 8174 25220
rect 8220 25217 8248 25248
rect 8297 25245 8309 25279
rect 8343 25276 8355 25279
rect 9122 25276 9128 25288
rect 8343 25248 9128 25276
rect 8343 25245 8355 25248
rect 8297 25239 8355 25245
rect 9122 25236 9128 25248
rect 9180 25236 9186 25288
rect 8205 25211 8263 25217
rect 8205 25177 8217 25211
rect 8251 25208 8263 25211
rect 9324 25208 9352 25307
rect 10318 25304 10324 25356
rect 10376 25304 10382 25356
rect 10413 25347 10471 25353
rect 10413 25313 10425 25347
rect 10459 25344 10471 25347
rect 12526 25344 12532 25356
rect 10459 25316 12532 25344
rect 10459 25313 10471 25316
rect 10413 25307 10471 25313
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 9950 25236 9956 25288
rect 10008 25236 10014 25288
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25276 10103 25279
rect 10226 25276 10232 25288
rect 10091 25248 10232 25276
rect 10091 25245 10103 25248
rect 10045 25239 10103 25245
rect 10226 25236 10232 25248
rect 10284 25236 10290 25288
rect 10505 25279 10563 25285
rect 10505 25245 10517 25279
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25276 10655 25279
rect 10781 25279 10839 25285
rect 10781 25276 10793 25279
rect 10643 25248 10793 25276
rect 10643 25245 10655 25248
rect 10597 25239 10655 25245
rect 10781 25245 10793 25248
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25276 11023 25279
rect 11057 25279 11115 25285
rect 11057 25276 11069 25279
rect 11011 25248 11069 25276
rect 11011 25245 11023 25248
rect 10965 25239 11023 25245
rect 11057 25245 11069 25248
rect 11103 25276 11115 25279
rect 11606 25276 11612 25288
rect 11103 25248 11612 25276
rect 11103 25245 11115 25248
rect 11057 25239 11115 25245
rect 8251 25180 9352 25208
rect 8251 25177 8263 25180
rect 8205 25171 8263 25177
rect 10134 25168 10140 25220
rect 10192 25208 10198 25220
rect 10520 25208 10548 25239
rect 10192 25180 10548 25208
rect 10796 25208 10824 25239
rect 11606 25236 11612 25248
rect 11664 25236 11670 25288
rect 11882 25236 11888 25288
rect 11940 25236 11946 25288
rect 12066 25236 12072 25288
rect 12124 25236 12130 25288
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25276 12679 25279
rect 12986 25276 12992 25288
rect 12667 25248 12992 25276
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 12986 25236 12992 25248
rect 13044 25236 13050 25288
rect 13078 25236 13084 25288
rect 13136 25236 13142 25288
rect 13173 25279 13231 25285
rect 13173 25245 13185 25279
rect 13219 25245 13231 25279
rect 13173 25239 13231 25245
rect 10796 25180 11008 25208
rect 10192 25168 10198 25180
rect 6512 25112 7420 25140
rect 6512 25100 6518 25112
rect 7742 25100 7748 25152
rect 7800 25100 7806 25152
rect 7834 25100 7840 25152
rect 7892 25140 7898 25152
rect 10594 25140 10600 25152
rect 7892 25112 10600 25140
rect 7892 25100 7898 25112
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 10778 25100 10784 25152
rect 10836 25140 10842 25152
rect 10873 25143 10931 25149
rect 10873 25140 10885 25143
rect 10836 25112 10885 25140
rect 10836 25100 10842 25112
rect 10873 25109 10885 25112
rect 10919 25109 10931 25143
rect 10980 25140 11008 25180
rect 11146 25168 11152 25220
rect 11204 25208 11210 25220
rect 12084 25208 12112 25236
rect 11204 25180 12112 25208
rect 11204 25168 11210 25180
rect 12710 25168 12716 25220
rect 12768 25208 12774 25220
rect 13188 25208 13216 25239
rect 13354 25236 13360 25288
rect 13412 25236 13418 25288
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25276 13507 25279
rect 14108 25276 14136 25375
rect 13495 25248 14136 25276
rect 13495 25245 13507 25248
rect 13449 25239 13507 25245
rect 14274 25236 14280 25288
rect 14332 25236 14338 25288
rect 14458 25236 14464 25288
rect 14516 25236 14522 25288
rect 14642 25236 14648 25288
rect 14700 25236 14706 25288
rect 15304 25285 15332 25384
rect 15378 25372 15384 25384
rect 15436 25372 15442 25424
rect 16574 25372 16580 25424
rect 16632 25412 16638 25424
rect 17405 25415 17463 25421
rect 17405 25412 17417 25415
rect 16632 25384 17417 25412
rect 16632 25372 16638 25384
rect 17405 25381 17417 25384
rect 17451 25381 17463 25415
rect 18230 25412 18236 25424
rect 17405 25375 17463 25381
rect 17880 25384 18236 25412
rect 17034 25344 17040 25356
rect 15396 25316 17040 25344
rect 15396 25285 15424 25316
rect 17034 25304 17040 25316
rect 17092 25304 17098 25356
rect 15105 25279 15163 25285
rect 15105 25245 15117 25279
rect 15151 25245 15163 25279
rect 15105 25239 15163 25245
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25245 15347 25279
rect 15289 25239 15347 25245
rect 15381 25279 15439 25285
rect 15381 25245 15393 25279
rect 15427 25245 15439 25279
rect 15381 25239 15439 25245
rect 12768 25180 13216 25208
rect 12768 25168 12774 25180
rect 13722 25168 13728 25220
rect 13780 25208 13786 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 13780 25180 14381 25208
rect 13780 25168 13786 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 11790 25140 11796 25152
rect 10980 25112 11796 25140
rect 10873 25103 10931 25109
rect 11790 25100 11796 25112
rect 11848 25100 11854 25152
rect 12434 25100 12440 25152
rect 12492 25140 12498 25152
rect 12529 25143 12587 25149
rect 12529 25140 12541 25143
rect 12492 25112 12541 25140
rect 12492 25100 12498 25112
rect 12529 25109 12541 25112
rect 12575 25109 12587 25143
rect 12529 25103 12587 25109
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 12897 25143 12955 25149
rect 12897 25140 12909 25143
rect 12860 25112 12909 25140
rect 12860 25100 12866 25112
rect 12897 25109 12909 25112
rect 12943 25109 12955 25143
rect 12897 25103 12955 25109
rect 13354 25100 13360 25152
rect 13412 25140 13418 25152
rect 15120 25140 15148 25239
rect 15470 25236 15476 25288
rect 15528 25236 15534 25288
rect 16758 25236 16764 25288
rect 16816 25276 16822 25288
rect 17880 25285 17908 25384
rect 18230 25372 18236 25384
rect 18288 25412 18294 25424
rect 18966 25412 18972 25424
rect 18288 25384 18972 25412
rect 18288 25372 18294 25384
rect 18966 25372 18972 25384
rect 19024 25372 19030 25424
rect 19076 25412 19104 25452
rect 19426 25440 19432 25492
rect 19484 25480 19490 25492
rect 19613 25483 19671 25489
rect 19613 25480 19625 25483
rect 19484 25452 19625 25480
rect 19484 25440 19490 25452
rect 19613 25449 19625 25452
rect 19659 25449 19671 25483
rect 19613 25443 19671 25449
rect 23477 25483 23535 25489
rect 23477 25449 23489 25483
rect 23523 25480 23535 25483
rect 23842 25480 23848 25492
rect 23523 25452 23848 25480
rect 23523 25449 23535 25452
rect 23477 25443 23535 25449
rect 23842 25440 23848 25452
rect 23900 25440 23906 25492
rect 24213 25483 24271 25489
rect 24213 25449 24225 25483
rect 24259 25480 24271 25483
rect 24394 25480 24400 25492
rect 24259 25452 24400 25480
rect 24259 25449 24271 25452
rect 24213 25443 24271 25449
rect 24394 25440 24400 25452
rect 24452 25440 24458 25492
rect 24670 25440 24676 25492
rect 24728 25480 24734 25492
rect 28166 25480 28172 25492
rect 24728 25452 28172 25480
rect 24728 25440 24734 25452
rect 20809 25415 20867 25421
rect 20809 25412 20821 25415
rect 19076 25384 20821 25412
rect 20809 25381 20821 25384
rect 20855 25381 20867 25415
rect 21358 25412 21364 25424
rect 20809 25375 20867 25381
rect 21008 25384 21364 25412
rect 21008 25353 21036 25384
rect 21358 25372 21364 25384
rect 21416 25372 21422 25424
rect 22186 25372 22192 25424
rect 22244 25412 22250 25424
rect 22738 25412 22744 25424
rect 22244 25384 22744 25412
rect 22244 25372 22250 25384
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 24762 25412 24768 25424
rect 23124 25384 24768 25412
rect 20993 25347 21051 25353
rect 18248 25316 19472 25344
rect 18248 25285 18276 25316
rect 17589 25279 17647 25285
rect 17589 25276 17601 25279
rect 16816 25248 17601 25276
rect 16816 25236 16822 25248
rect 17589 25245 17601 25248
rect 17635 25245 17647 25279
rect 17589 25239 17647 25245
rect 17865 25279 17923 25285
rect 17865 25245 17877 25279
rect 17911 25245 17923 25279
rect 17865 25239 17923 25245
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25245 18291 25279
rect 18233 25239 18291 25245
rect 18506 25236 18512 25288
rect 18564 25236 18570 25288
rect 18874 25236 18880 25288
rect 18932 25276 18938 25288
rect 19444 25285 19472 25316
rect 20993 25313 21005 25347
rect 21039 25313 21051 25347
rect 20993 25307 21051 25313
rect 21177 25347 21235 25353
rect 21177 25313 21189 25347
rect 21223 25344 21235 25347
rect 23014 25344 23020 25356
rect 21223 25316 23020 25344
rect 21223 25313 21235 25316
rect 21177 25307 21235 25313
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 18932 25248 19257 25276
rect 18932 25236 18938 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19429 25279 19487 25285
rect 19429 25245 19441 25279
rect 19475 25276 19487 25279
rect 19518 25276 19524 25288
rect 19475 25248 19524 25276
rect 19475 25245 19487 25248
rect 19429 25239 19487 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 19794 25236 19800 25288
rect 19852 25236 19858 25288
rect 19978 25236 19984 25288
rect 20036 25276 20042 25288
rect 20073 25279 20131 25285
rect 20073 25276 20085 25279
rect 20036 25248 20085 25276
rect 20036 25236 20042 25248
rect 20073 25245 20085 25248
rect 20119 25245 20131 25279
rect 20073 25239 20131 25245
rect 20257 25279 20315 25285
rect 20257 25245 20269 25279
rect 20303 25276 20315 25279
rect 20438 25276 20444 25288
rect 20303 25248 20444 25276
rect 20303 25245 20315 25248
rect 20257 25239 20315 25245
rect 20438 25236 20444 25248
rect 20496 25236 20502 25288
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 16850 25168 16856 25220
rect 16908 25168 16914 25220
rect 18138 25168 18144 25220
rect 18196 25208 18202 25220
rect 19337 25211 19395 25217
rect 19337 25208 19349 25211
rect 18196 25180 19349 25208
rect 18196 25168 18202 25180
rect 19337 25177 19349 25180
rect 19383 25177 19395 25211
rect 21284 25208 21312 25239
rect 21358 25236 21364 25288
rect 21416 25276 21422 25288
rect 22020 25285 22048 25316
rect 23014 25304 23020 25316
rect 23072 25304 23078 25356
rect 21637 25279 21695 25285
rect 21637 25276 21649 25279
rect 21416 25248 21649 25276
rect 21416 25236 21422 25248
rect 21637 25245 21649 25248
rect 21683 25245 21695 25279
rect 21637 25239 21695 25245
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25245 22063 25279
rect 22005 25239 22063 25245
rect 22462 25236 22468 25288
rect 22520 25236 22526 25288
rect 23124 25285 23152 25384
rect 24762 25372 24768 25384
rect 24820 25372 24826 25424
rect 23658 25304 23664 25356
rect 23716 25304 23722 25356
rect 25056 25353 25084 25452
rect 28166 25440 28172 25452
rect 28224 25440 28230 25492
rect 29730 25440 29736 25492
rect 29788 25440 29794 25492
rect 30929 25483 30987 25489
rect 30929 25449 30941 25483
rect 30975 25480 30987 25483
rect 33042 25480 33048 25492
rect 30975 25452 33048 25480
rect 30975 25449 30987 25452
rect 30929 25443 30987 25449
rect 33042 25440 33048 25452
rect 33100 25440 33106 25492
rect 33226 25440 33232 25492
rect 33284 25480 33290 25492
rect 34238 25480 34244 25492
rect 33284 25452 34244 25480
rect 33284 25440 33290 25452
rect 34238 25440 34244 25452
rect 34296 25440 34302 25492
rect 34330 25440 34336 25492
rect 34388 25480 34394 25492
rect 35069 25483 35127 25489
rect 34388 25452 34652 25480
rect 34388 25440 34394 25452
rect 25774 25372 25780 25424
rect 25832 25372 25838 25424
rect 28902 25372 28908 25424
rect 28960 25412 28966 25424
rect 29914 25412 29920 25424
rect 28960 25384 29920 25412
rect 28960 25372 28966 25384
rect 29914 25372 29920 25384
rect 29972 25372 29978 25424
rect 32214 25412 32220 25424
rect 32140 25384 32220 25412
rect 25041 25347 25099 25353
rect 25041 25313 25053 25347
rect 25087 25313 25099 25347
rect 25714 25316 27292 25344
rect 25041 25307 25099 25313
rect 23109 25279 23167 25285
rect 23109 25245 23121 25279
rect 23155 25245 23167 25279
rect 23109 25239 23167 25245
rect 23474 25236 23480 25288
rect 23532 25276 23538 25288
rect 23937 25279 23995 25285
rect 23937 25276 23949 25279
rect 23532 25248 23949 25276
rect 23532 25236 23538 25248
rect 23937 25245 23949 25248
rect 23983 25245 23995 25279
rect 23937 25239 23995 25245
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25276 24087 25279
rect 24486 25276 24492 25288
rect 24075 25248 24492 25276
rect 24075 25245 24087 25248
rect 24029 25239 24087 25245
rect 24486 25236 24492 25248
rect 24544 25236 24550 25288
rect 24854 25236 24860 25288
rect 24912 25276 24918 25288
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 24912 25248 24961 25276
rect 24912 25236 24918 25248
rect 24949 25245 24961 25248
rect 24995 25276 25007 25279
rect 25314 25276 25320 25288
rect 24995 25248 25320 25276
rect 24995 25245 25007 25248
rect 24949 25239 25007 25245
rect 25314 25236 25320 25248
rect 25372 25236 25378 25288
rect 25593 25279 25651 25285
rect 25593 25245 25605 25279
rect 25639 25276 25651 25279
rect 25958 25276 25964 25288
rect 25639 25248 25964 25276
rect 25639 25245 25651 25248
rect 25593 25239 25651 25245
rect 25958 25236 25964 25248
rect 26016 25236 26022 25288
rect 26418 25276 26424 25288
rect 26252 25248 26424 25276
rect 22480 25208 22508 25236
rect 21284 25180 22508 25208
rect 19337 25171 19395 25177
rect 22922 25168 22928 25220
rect 22980 25168 22986 25220
rect 23569 25211 23627 25217
rect 23569 25177 23581 25211
rect 23615 25208 23627 25211
rect 25406 25208 25412 25220
rect 23615 25180 25412 25208
rect 23615 25177 23627 25180
rect 23569 25171 23627 25177
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 26252 25208 26280 25248
rect 26418 25236 26424 25248
rect 26476 25236 26482 25288
rect 27264 25276 27292 25316
rect 27338 25304 27344 25356
rect 27396 25304 27402 25356
rect 27709 25347 27767 25353
rect 27709 25313 27721 25347
rect 27755 25344 27767 25347
rect 28626 25344 28632 25356
rect 27755 25316 28632 25344
rect 27755 25313 27767 25316
rect 27709 25307 27767 25313
rect 28626 25304 28632 25316
rect 28684 25304 28690 25356
rect 28994 25304 29000 25356
rect 29052 25344 29058 25356
rect 31665 25347 31723 25353
rect 31665 25344 31677 25347
rect 29052 25316 29960 25344
rect 29052 25304 29058 25316
rect 27798 25276 27804 25288
rect 27264 25248 27804 25276
rect 27798 25236 27804 25248
rect 27856 25276 27862 25288
rect 29012 25276 29040 25304
rect 27856 25248 29040 25276
rect 27856 25236 27862 25248
rect 27985 25211 28043 25217
rect 25792 25180 26280 25208
rect 27002 25180 27108 25208
rect 13412 25112 15148 25140
rect 13412 25100 13418 25112
rect 15654 25100 15660 25152
rect 15712 25100 15718 25152
rect 17230 25143 17288 25149
rect 17230 25109 17242 25143
rect 17276 25140 17288 25143
rect 17402 25140 17408 25152
rect 17276 25112 17408 25140
rect 17276 25109 17288 25112
rect 17230 25103 17288 25109
rect 17402 25100 17408 25112
rect 17460 25100 17466 25152
rect 17494 25100 17500 25152
rect 17552 25140 17558 25152
rect 21361 25143 21419 25149
rect 21361 25140 21373 25143
rect 17552 25112 21373 25140
rect 17552 25100 17558 25112
rect 21361 25109 21373 25112
rect 21407 25109 21419 25143
rect 21361 25103 21419 25109
rect 23198 25100 23204 25152
rect 23256 25100 23262 25152
rect 23293 25143 23351 25149
rect 23293 25109 23305 25143
rect 23339 25140 23351 25143
rect 23382 25140 23388 25152
rect 23339 25112 23388 25140
rect 23339 25109 23351 25112
rect 23293 25103 23351 25109
rect 23382 25100 23388 25112
rect 23440 25140 23446 25152
rect 25792 25140 25820 25180
rect 27080 25152 27108 25180
rect 27985 25177 27997 25211
rect 28031 25208 28043 25211
rect 28994 25208 29000 25220
rect 28031 25180 29000 25208
rect 28031 25177 28043 25180
rect 27985 25171 28043 25177
rect 28994 25168 29000 25180
rect 29052 25168 29058 25220
rect 29932 25217 29960 25316
rect 31496 25316 31677 25344
rect 30837 25279 30895 25285
rect 30837 25245 30849 25279
rect 30883 25276 30895 25279
rect 31018 25276 31024 25288
rect 30883 25248 31024 25276
rect 30883 25245 30895 25248
rect 30837 25239 30895 25245
rect 31018 25236 31024 25248
rect 31076 25236 31082 25288
rect 31113 25279 31171 25285
rect 31113 25245 31125 25279
rect 31159 25245 31171 25279
rect 31113 25239 31171 25245
rect 29917 25211 29975 25217
rect 29917 25177 29929 25211
rect 29963 25177 29975 25211
rect 31128 25208 31156 25239
rect 31202 25236 31208 25288
rect 31260 25236 31266 25288
rect 31294 25236 31300 25288
rect 31352 25236 31358 25288
rect 31496 25285 31524 25316
rect 31665 25313 31677 25316
rect 31711 25313 31723 25347
rect 31665 25307 31723 25313
rect 32030 25304 32036 25356
rect 32088 25304 32094 25356
rect 32140 25353 32168 25384
rect 32214 25372 32220 25384
rect 32272 25372 32278 25424
rect 32309 25415 32367 25421
rect 32309 25381 32321 25415
rect 32355 25412 32367 25415
rect 33410 25412 33416 25424
rect 32355 25384 33416 25412
rect 32355 25381 32367 25384
rect 32309 25375 32367 25381
rect 33410 25372 33416 25384
rect 33468 25372 33474 25424
rect 33686 25372 33692 25424
rect 33744 25412 33750 25424
rect 33873 25415 33931 25421
rect 33873 25412 33885 25415
rect 33744 25384 33885 25412
rect 33744 25372 33750 25384
rect 33873 25381 33885 25384
rect 33919 25412 33931 25415
rect 34514 25412 34520 25424
rect 33919 25384 34520 25412
rect 33919 25381 33931 25384
rect 33873 25375 33931 25381
rect 34514 25372 34520 25384
rect 34572 25372 34578 25424
rect 34624 25412 34652 25452
rect 35069 25449 35081 25483
rect 35115 25480 35127 25483
rect 35342 25480 35348 25492
rect 35115 25452 35348 25480
rect 35115 25449 35127 25452
rect 35069 25443 35127 25449
rect 35342 25440 35348 25452
rect 35400 25440 35406 25492
rect 35526 25440 35532 25492
rect 35584 25440 35590 25492
rect 36538 25480 36544 25492
rect 35636 25452 36544 25480
rect 35636 25412 35664 25452
rect 36538 25440 36544 25452
rect 36596 25440 36602 25492
rect 34624 25384 35664 25412
rect 35710 25372 35716 25424
rect 35768 25372 35774 25424
rect 35802 25372 35808 25424
rect 35860 25412 35866 25424
rect 35897 25415 35955 25421
rect 35897 25412 35909 25415
rect 35860 25384 35909 25412
rect 35860 25372 35866 25384
rect 35897 25381 35909 25384
rect 35943 25381 35955 25415
rect 35897 25375 35955 25381
rect 32125 25347 32183 25353
rect 32125 25313 32137 25347
rect 32171 25313 32183 25347
rect 32125 25307 32183 25313
rect 32398 25304 32404 25356
rect 32456 25344 32462 25356
rect 34054 25344 34060 25356
rect 32456 25316 32904 25344
rect 32456 25304 32462 25316
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25245 31539 25279
rect 31481 25239 31539 25245
rect 31573 25279 31631 25285
rect 31573 25245 31585 25279
rect 31619 25276 31631 25279
rect 31754 25276 31760 25288
rect 31619 25248 31760 25276
rect 31619 25245 31631 25248
rect 31573 25239 31631 25245
rect 31754 25236 31760 25248
rect 31812 25236 31818 25288
rect 31846 25236 31852 25288
rect 31904 25236 31910 25288
rect 31941 25279 31999 25285
rect 31941 25245 31953 25279
rect 31987 25276 31999 25279
rect 31987 25270 32004 25276
rect 31987 25245 32260 25270
rect 31941 25242 32260 25245
rect 31941 25239 31999 25242
rect 29917 25171 29975 25177
rect 30668 25180 31156 25208
rect 32232 25208 32260 25242
rect 32490 25236 32496 25288
rect 32548 25236 32554 25288
rect 32876 25285 32904 25316
rect 33428 25316 34060 25344
rect 32769 25279 32827 25285
rect 32769 25278 32781 25279
rect 32692 25276 32781 25278
rect 32600 25250 32781 25276
rect 32600 25248 32720 25250
rect 32398 25208 32404 25220
rect 32232 25180 32404 25208
rect 23440 25112 25820 25140
rect 25915 25143 25973 25149
rect 23440 25100 23446 25112
rect 25915 25109 25927 25143
rect 25961 25140 25973 25143
rect 26050 25140 26056 25152
rect 25961 25112 26056 25140
rect 25961 25109 25973 25112
rect 25915 25103 25973 25109
rect 26050 25100 26056 25112
rect 26108 25140 26114 25152
rect 26786 25140 26792 25152
rect 26108 25112 26792 25140
rect 26108 25100 26114 25112
rect 26786 25100 26792 25112
rect 26844 25100 26850 25152
rect 27062 25100 27068 25152
rect 27120 25100 27126 25152
rect 27893 25143 27951 25149
rect 27893 25109 27905 25143
rect 27939 25140 27951 25143
rect 28350 25140 28356 25152
rect 27939 25112 28356 25140
rect 27939 25109 27951 25112
rect 27893 25103 27951 25109
rect 28350 25100 28356 25112
rect 28408 25100 28414 25152
rect 28626 25100 28632 25152
rect 28684 25140 28690 25152
rect 29549 25143 29607 25149
rect 29549 25140 29561 25143
rect 28684 25112 29561 25140
rect 28684 25100 28690 25112
rect 29549 25109 29561 25112
rect 29595 25109 29607 25143
rect 29549 25103 29607 25109
rect 29717 25143 29775 25149
rect 29717 25109 29729 25143
rect 29763 25140 29775 25143
rect 30668 25140 30696 25180
rect 29763 25112 30696 25140
rect 29763 25109 29775 25112
rect 29717 25103 29775 25109
rect 30742 25100 30748 25152
rect 30800 25100 30806 25152
rect 31128 25140 31156 25180
rect 32398 25168 32404 25180
rect 32456 25168 32462 25220
rect 32600 25208 32628 25248
rect 32769 25245 32781 25250
rect 32815 25245 32827 25279
rect 32769 25239 32827 25245
rect 32861 25279 32919 25285
rect 32861 25245 32873 25279
rect 32907 25245 32919 25279
rect 32861 25239 32919 25245
rect 32953 25279 33011 25285
rect 32953 25245 32965 25279
rect 32999 25245 33011 25279
rect 32953 25239 33011 25245
rect 33045 25279 33103 25285
rect 33045 25245 33057 25279
rect 33091 25276 33103 25279
rect 33137 25279 33195 25285
rect 33137 25276 33149 25279
rect 33091 25248 33149 25276
rect 33091 25245 33103 25248
rect 33045 25239 33103 25245
rect 33137 25245 33149 25248
rect 33183 25276 33195 25279
rect 33336 25276 33385 25278
rect 33428 25276 33456 25316
rect 34054 25304 34060 25316
rect 34112 25304 34118 25356
rect 35728 25344 35756 25372
rect 34256 25316 35756 25344
rect 33183 25248 33456 25276
rect 33505 25279 33563 25285
rect 33183 25245 33195 25248
rect 33137 25239 33195 25245
rect 33505 25245 33517 25279
rect 33551 25245 33563 25279
rect 33505 25239 33563 25245
rect 32968 25208 32996 25239
rect 32600 25180 32996 25208
rect 33520 25208 33548 25239
rect 33686 25236 33692 25288
rect 33744 25236 33750 25288
rect 33778 25236 33784 25288
rect 33836 25236 33842 25288
rect 33965 25279 34023 25285
rect 33965 25245 33977 25279
rect 34011 25276 34023 25279
rect 34256 25276 34284 25316
rect 34011 25248 34284 25276
rect 34011 25245 34023 25248
rect 33965 25239 34023 25245
rect 34790 25236 34796 25288
rect 34848 25276 34854 25288
rect 35069 25279 35127 25285
rect 35069 25276 35081 25279
rect 34848 25248 35081 25276
rect 34848 25236 34854 25248
rect 35069 25245 35081 25248
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 33870 25208 33876 25220
rect 33520 25180 33876 25208
rect 32600 25140 32628 25180
rect 33870 25168 33876 25180
rect 33928 25208 33934 25220
rect 34808 25208 34836 25236
rect 33928 25180 34836 25208
rect 35084 25208 35112 25239
rect 35250 25236 35256 25288
rect 35308 25276 35314 25288
rect 35618 25276 35624 25288
rect 35308 25248 35624 25276
rect 35308 25236 35314 25248
rect 35618 25236 35624 25248
rect 35676 25236 35682 25288
rect 35710 25236 35716 25288
rect 35768 25236 35774 25288
rect 35986 25236 35992 25288
rect 36044 25276 36050 25288
rect 36081 25279 36139 25285
rect 36081 25276 36093 25279
rect 36044 25248 36093 25276
rect 36044 25236 36050 25248
rect 36081 25245 36093 25248
rect 36127 25245 36139 25279
rect 36081 25239 36139 25245
rect 35342 25208 35348 25220
rect 35084 25180 35348 25208
rect 33928 25168 33934 25180
rect 35342 25168 35348 25180
rect 35400 25168 35406 25220
rect 31128 25112 32628 25140
rect 32677 25143 32735 25149
rect 32677 25109 32689 25143
rect 32723 25140 32735 25143
rect 32950 25140 32956 25152
rect 32723 25112 32956 25140
rect 32723 25109 32735 25112
rect 32677 25103 32735 25109
rect 32950 25100 32956 25112
rect 33008 25100 33014 25152
rect 33226 25100 33232 25152
rect 33284 25100 33290 25152
rect 1104 25050 36524 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 36524 25050
rect 1104 24976 36524 24998
rect 3237 24939 3295 24945
rect 3237 24905 3249 24939
rect 3283 24905 3295 24939
rect 3237 24899 3295 24905
rect 4080 24908 4844 24936
rect 2958 24868 2964 24880
rect 2898 24840 2964 24868
rect 2958 24828 2964 24840
rect 3016 24828 3022 24880
rect 1394 24692 1400 24744
rect 1452 24692 1458 24744
rect 1673 24735 1731 24741
rect 1673 24701 1685 24735
rect 1719 24732 1731 24735
rect 3252 24732 3280 24899
rect 3602 24828 3608 24880
rect 3660 24828 3666 24880
rect 4080 24812 4108 24908
rect 4706 24868 4712 24880
rect 4172 24840 4712 24868
rect 1719 24704 3280 24732
rect 3620 24772 4016 24800
rect 1719 24701 1731 24704
rect 1673 24695 1731 24701
rect 2774 24624 2780 24676
rect 2832 24664 2838 24676
rect 3620 24664 3648 24772
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24701 3755 24735
rect 3697 24695 3755 24701
rect 2832 24636 3648 24664
rect 2832 24624 2838 24636
rect 3145 24599 3203 24605
rect 3145 24565 3157 24599
rect 3191 24596 3203 24599
rect 3712 24596 3740 24695
rect 3786 24692 3792 24744
rect 3844 24692 3850 24744
rect 3988 24732 4016 24772
rect 4062 24760 4068 24812
rect 4120 24760 4126 24812
rect 4172 24741 4200 24840
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 4816 24868 4844 24908
rect 5902 24896 5908 24948
rect 5960 24896 5966 24948
rect 5994 24896 6000 24948
rect 6052 24936 6058 24948
rect 6052 24908 8064 24936
rect 6052 24896 6058 24908
rect 4816 24840 4922 24868
rect 5718 24828 5724 24880
rect 5776 24868 5782 24880
rect 6454 24868 6460 24880
rect 5776 24840 6460 24868
rect 5776 24828 5782 24840
rect 6454 24828 6460 24840
rect 6512 24828 6518 24880
rect 7006 24828 7012 24880
rect 7064 24868 7070 24880
rect 8036 24868 8064 24908
rect 9030 24896 9036 24948
rect 9088 24936 9094 24948
rect 9582 24936 9588 24948
rect 9088 24908 9588 24936
rect 9088 24896 9094 24908
rect 9582 24896 9588 24908
rect 9640 24896 9646 24948
rect 9677 24939 9735 24945
rect 9677 24905 9689 24939
rect 9723 24936 9735 24939
rect 10042 24936 10048 24948
rect 9723 24908 10048 24936
rect 9723 24905 9735 24908
rect 9677 24899 9735 24905
rect 10042 24896 10048 24908
rect 10100 24896 10106 24948
rect 11882 24896 11888 24948
rect 11940 24936 11946 24948
rect 12161 24939 12219 24945
rect 12161 24936 12173 24939
rect 11940 24908 12173 24936
rect 11940 24896 11946 24908
rect 12161 24905 12173 24908
rect 12207 24905 12219 24939
rect 13354 24936 13360 24948
rect 12161 24899 12219 24905
rect 12361 24908 13360 24936
rect 12361 24868 12389 24908
rect 13354 24896 13360 24908
rect 13412 24896 13418 24948
rect 13538 24896 13544 24948
rect 13596 24936 13602 24948
rect 15378 24936 15384 24948
rect 13596 24908 15384 24936
rect 13596 24896 13602 24908
rect 15378 24896 15384 24908
rect 15436 24896 15442 24948
rect 15838 24896 15844 24948
rect 15896 24896 15902 24948
rect 17402 24896 17408 24948
rect 17460 24896 17466 24948
rect 18141 24939 18199 24945
rect 18141 24905 18153 24939
rect 18187 24936 18199 24939
rect 18874 24936 18880 24948
rect 18187 24908 18880 24936
rect 18187 24905 18199 24908
rect 18141 24899 18199 24905
rect 18874 24896 18880 24908
rect 18932 24896 18938 24948
rect 19260 24908 22692 24936
rect 7064 24840 7222 24868
rect 8036 24840 12389 24868
rect 7064 24828 7070 24840
rect 13078 24828 13084 24880
rect 13136 24868 13142 24880
rect 15102 24868 15108 24880
rect 13136 24840 15108 24868
rect 13136 24828 13142 24840
rect 9674 24800 9680 24812
rect 9635 24772 9680 24800
rect 9674 24760 9680 24772
rect 9732 24760 9738 24812
rect 9766 24760 9772 24812
rect 9824 24800 9830 24812
rect 11146 24800 11152 24812
rect 9824 24772 11152 24800
rect 9824 24760 9830 24772
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 11348 24772 12296 24800
rect 4157 24735 4215 24741
rect 4157 24732 4169 24735
rect 3988 24704 4169 24732
rect 4157 24701 4169 24704
rect 4203 24701 4215 24735
rect 4157 24695 4215 24701
rect 4433 24735 4491 24741
rect 4433 24701 4445 24735
rect 4479 24732 4491 24735
rect 4522 24732 4528 24744
rect 4479 24704 4528 24732
rect 4479 24701 4491 24704
rect 4433 24695 4491 24701
rect 4522 24692 4528 24704
rect 4580 24692 4586 24744
rect 4798 24692 4804 24744
rect 4856 24732 4862 24744
rect 6457 24735 6515 24741
rect 6457 24732 6469 24735
rect 4856 24704 6469 24732
rect 4856 24692 4862 24704
rect 6457 24701 6469 24704
rect 6503 24701 6515 24735
rect 6457 24695 6515 24701
rect 6733 24735 6791 24741
rect 6733 24701 6745 24735
rect 6779 24732 6791 24735
rect 7282 24732 7288 24744
rect 6779 24704 7288 24732
rect 6779 24701 6791 24704
rect 6733 24695 6791 24701
rect 7282 24692 7288 24704
rect 7340 24692 7346 24744
rect 8202 24692 8208 24744
rect 8260 24732 8266 24744
rect 8941 24735 8999 24741
rect 8941 24732 8953 24735
rect 8260 24704 8953 24732
rect 8260 24692 8266 24704
rect 8941 24701 8953 24704
rect 8987 24732 8999 24735
rect 9214 24732 9220 24744
rect 8987 24704 9220 24732
rect 8987 24701 8999 24704
rect 8941 24695 8999 24701
rect 9214 24692 9220 24704
rect 9272 24692 9278 24744
rect 10137 24735 10195 24741
rect 10137 24701 10149 24735
rect 10183 24732 10195 24735
rect 10226 24732 10232 24744
rect 10183 24704 10232 24732
rect 10183 24701 10195 24704
rect 10137 24695 10195 24701
rect 10226 24692 10232 24704
rect 10284 24692 10290 24744
rect 9122 24624 9128 24676
rect 9180 24664 9186 24676
rect 11348 24664 11376 24772
rect 11422 24692 11428 24744
rect 11480 24732 11486 24744
rect 11609 24735 11667 24741
rect 11609 24732 11621 24735
rect 11480 24704 11621 24732
rect 11480 24692 11486 24704
rect 11609 24701 11621 24704
rect 11655 24701 11667 24735
rect 11609 24695 11667 24701
rect 11701 24735 11759 24741
rect 11701 24701 11713 24735
rect 11747 24701 11759 24735
rect 11701 24695 11759 24701
rect 9180 24636 11376 24664
rect 11716 24664 11744 24695
rect 11790 24692 11796 24744
rect 11848 24692 11854 24744
rect 11882 24692 11888 24744
rect 11940 24692 11946 24744
rect 11974 24692 11980 24744
rect 12032 24732 12038 24744
rect 12069 24735 12127 24741
rect 12069 24732 12081 24735
rect 12032 24704 12081 24732
rect 12032 24692 12038 24704
rect 12069 24701 12081 24704
rect 12115 24701 12127 24735
rect 12069 24695 12127 24701
rect 12158 24664 12164 24676
rect 11716 24636 12164 24664
rect 9180 24624 9186 24636
rect 12158 24624 12164 24636
rect 12216 24624 12222 24676
rect 12268 24664 12296 24772
rect 12342 24760 12348 24812
rect 12400 24760 12406 24812
rect 12434 24760 12440 24812
rect 12492 24760 12498 24812
rect 12710 24760 12716 24812
rect 12768 24760 12774 24812
rect 13280 24809 13308 24840
rect 15102 24828 15108 24840
rect 15160 24868 15166 24880
rect 19061 24871 19119 24877
rect 19061 24868 19073 24871
rect 15160 24840 15976 24868
rect 15160 24828 15166 24840
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24769 13323 24803
rect 13265 24763 13323 24769
rect 13354 24760 13360 24812
rect 13412 24760 13418 24812
rect 13446 24760 13452 24812
rect 13504 24800 13510 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 13504 24772 13553 24800
rect 13504 24760 13510 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 14090 24800 14096 24812
rect 13679 24772 14096 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14090 24760 14096 24772
rect 14148 24760 14154 24812
rect 15565 24803 15623 24809
rect 15565 24769 15577 24803
rect 15611 24800 15623 24803
rect 15654 24800 15660 24812
rect 15611 24772 15660 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 15948 24809 15976 24840
rect 18800 24840 19073 24868
rect 15933 24803 15991 24809
rect 15933 24769 15945 24803
rect 15979 24769 15991 24803
rect 15933 24763 15991 24769
rect 17589 24803 17647 24809
rect 17589 24769 17601 24803
rect 17635 24800 17647 24803
rect 17678 24800 17684 24812
rect 17635 24772 17684 24800
rect 17635 24769 17647 24772
rect 17589 24763 17647 24769
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 17862 24760 17868 24812
rect 17920 24760 17926 24812
rect 18506 24760 18512 24812
rect 18564 24800 18570 24812
rect 18800 24809 18828 24840
rect 19061 24837 19073 24840
rect 19107 24837 19119 24871
rect 19260 24868 19288 24908
rect 19061 24831 19119 24837
rect 19168 24840 19288 24868
rect 18785 24803 18843 24809
rect 18785 24800 18797 24803
rect 18564 24772 18797 24800
rect 18564 24760 18570 24772
rect 18785 24769 18797 24772
rect 18831 24769 18843 24803
rect 18785 24763 18843 24769
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19168 24800 19196 24840
rect 19426 24828 19432 24880
rect 19484 24828 19490 24880
rect 19981 24871 20039 24877
rect 19981 24837 19993 24871
rect 20027 24868 20039 24871
rect 20806 24868 20812 24880
rect 20027 24840 20812 24868
rect 20027 24837 20039 24840
rect 19981 24831 20039 24837
rect 19024 24772 19196 24800
rect 19245 24803 19303 24809
rect 19024 24760 19030 24772
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19444 24800 19472 24828
rect 19291 24772 19472 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 19886 24760 19892 24812
rect 19944 24760 19950 24812
rect 12894 24692 12900 24744
rect 12952 24732 12958 24744
rect 15197 24735 15255 24741
rect 15197 24732 15209 24735
rect 12952 24704 15209 24732
rect 12952 24692 12958 24704
rect 15197 24701 15209 24704
rect 15243 24701 15255 24735
rect 15197 24695 15255 24701
rect 17773 24735 17831 24741
rect 17773 24701 17785 24735
rect 17819 24732 17831 24735
rect 18690 24732 18696 24744
rect 17819 24704 18696 24732
rect 17819 24701 17831 24704
rect 17773 24695 17831 24701
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 19429 24735 19487 24741
rect 19429 24701 19441 24735
rect 19475 24732 19487 24735
rect 19518 24732 19524 24744
rect 19475 24704 19524 24732
rect 19475 24701 19487 24704
rect 19429 24695 19487 24701
rect 19518 24692 19524 24704
rect 19576 24692 19582 24744
rect 18601 24667 18659 24673
rect 18601 24664 18613 24667
rect 12268 24636 18613 24664
rect 18601 24633 18613 24636
rect 18647 24633 18659 24667
rect 18601 24627 18659 24633
rect 19242 24624 19248 24676
rect 19300 24664 19306 24676
rect 19996 24664 20024 24831
rect 20806 24828 20812 24840
rect 20864 24828 20870 24880
rect 21637 24871 21695 24877
rect 21407 24837 21465 24843
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 20088 24732 20116 24763
rect 20162 24760 20168 24812
rect 20220 24800 20226 24812
rect 20257 24803 20315 24809
rect 20257 24800 20269 24803
rect 20220 24772 20269 24800
rect 20220 24760 20226 24772
rect 20257 24769 20269 24772
rect 20303 24800 20315 24803
rect 20622 24800 20628 24812
rect 20303 24772 20628 24800
rect 20303 24769 20315 24772
rect 20257 24763 20315 24769
rect 20622 24760 20628 24772
rect 20680 24760 20686 24812
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 21407 24803 21419 24837
rect 21453 24803 21465 24837
rect 21637 24837 21649 24871
rect 21683 24868 21695 24871
rect 21726 24868 21732 24880
rect 21683 24840 21732 24868
rect 21683 24837 21695 24840
rect 21637 24831 21695 24837
rect 21726 24828 21732 24840
rect 21784 24828 21790 24880
rect 21818 24828 21824 24880
rect 21876 24868 21882 24880
rect 22664 24877 22692 24908
rect 26970 24896 26976 24948
rect 27028 24936 27034 24948
rect 27341 24939 27399 24945
rect 27341 24936 27353 24939
rect 27028 24908 27353 24936
rect 27028 24896 27034 24908
rect 27341 24905 27353 24908
rect 27387 24905 27399 24939
rect 27341 24899 27399 24905
rect 28810 24896 28816 24948
rect 28868 24896 28874 24948
rect 28920 24908 29776 24936
rect 22649 24871 22707 24877
rect 21876 24840 22140 24868
rect 21876 24828 21882 24840
rect 22112 24809 22140 24840
rect 22649 24837 22661 24871
rect 22695 24837 22707 24871
rect 22649 24831 22707 24837
rect 24762 24828 24768 24880
rect 24820 24868 24826 24880
rect 26234 24868 26240 24880
rect 24820 24840 26240 24868
rect 24820 24828 24826 24840
rect 26234 24828 26240 24840
rect 26292 24828 26298 24880
rect 26344 24840 26740 24868
rect 21407 24800 21465 24803
rect 20772 24797 21465 24800
rect 22097 24803 22155 24809
rect 20772 24772 21450 24797
rect 20772 24760 20778 24772
rect 22097 24769 22109 24803
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 23290 24760 23296 24812
rect 23348 24760 23354 24812
rect 23382 24760 23388 24812
rect 23440 24760 23446 24812
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 23753 24803 23811 24809
rect 23753 24800 23765 24803
rect 23624 24772 23765 24800
rect 23624 24760 23630 24772
rect 23753 24769 23765 24772
rect 23799 24769 23811 24803
rect 23753 24763 23811 24769
rect 20346 24732 20352 24744
rect 20088 24704 20352 24732
rect 20346 24692 20352 24704
rect 20404 24692 20410 24744
rect 21358 24732 21364 24744
rect 21284 24704 21364 24732
rect 21284 24673 21312 24704
rect 21358 24692 21364 24704
rect 21416 24692 21422 24744
rect 21726 24692 21732 24744
rect 21784 24732 21790 24744
rect 22005 24735 22063 24741
rect 22005 24732 22017 24735
rect 21784 24704 22017 24732
rect 21784 24692 21790 24704
rect 22005 24701 22017 24704
rect 22051 24701 22063 24735
rect 22005 24695 22063 24701
rect 22189 24735 22247 24741
rect 22189 24701 22201 24735
rect 22235 24701 22247 24735
rect 22189 24695 22247 24701
rect 22281 24735 22339 24741
rect 22281 24701 22293 24735
rect 22327 24732 22339 24735
rect 22738 24732 22744 24744
rect 22327 24704 22744 24732
rect 22327 24701 22339 24704
rect 22281 24695 22339 24701
rect 19300 24636 20024 24664
rect 21269 24667 21327 24673
rect 19300 24624 19306 24636
rect 21269 24633 21281 24667
rect 21315 24633 21327 24667
rect 22204 24664 22232 24695
rect 22738 24692 22744 24704
rect 22796 24692 22802 24744
rect 22925 24735 22983 24741
rect 22925 24701 22937 24735
rect 22971 24732 22983 24735
rect 23014 24732 23020 24744
rect 22971 24704 23020 24732
rect 22971 24701 22983 24704
rect 22925 24695 22983 24701
rect 23014 24692 23020 24704
rect 23072 24692 23078 24744
rect 24118 24692 24124 24744
rect 24176 24732 24182 24744
rect 24673 24735 24731 24741
rect 24673 24732 24685 24735
rect 24176 24704 24685 24732
rect 24176 24692 24182 24704
rect 24673 24701 24685 24704
rect 24719 24701 24731 24735
rect 24780 24732 24808 24828
rect 24857 24803 24915 24809
rect 24857 24769 24869 24803
rect 24903 24800 24915 24803
rect 25222 24800 25228 24812
rect 24903 24772 25228 24800
rect 24903 24769 24915 24772
rect 24857 24763 24915 24769
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 26344 24800 26372 24840
rect 26712 24812 26740 24840
rect 28718 24828 28724 24880
rect 28776 24868 28782 24880
rect 28920 24868 28948 24908
rect 29748 24880 29776 24908
rect 30190 24896 30196 24948
rect 30248 24936 30254 24948
rect 30926 24936 30932 24948
rect 30248 24908 30932 24936
rect 30248 24896 30254 24908
rect 30926 24896 30932 24908
rect 30984 24896 30990 24948
rect 31497 24939 31555 24945
rect 31497 24936 31509 24939
rect 31036 24908 31509 24936
rect 28776 24840 28948 24868
rect 29380 24840 29592 24868
rect 28776 24828 28782 24840
rect 26191 24772 26372 24800
rect 26421 24803 26479 24809
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 26421 24769 26433 24803
rect 26467 24800 26479 24803
rect 26602 24800 26608 24812
rect 26467 24772 26608 24800
rect 26467 24769 26479 24772
rect 26421 24763 26479 24769
rect 26602 24760 26608 24772
rect 26660 24760 26666 24812
rect 26694 24760 26700 24812
rect 26752 24800 26758 24812
rect 26752 24772 27844 24800
rect 26752 24760 26758 24772
rect 24949 24735 25007 24741
rect 24949 24732 24961 24735
rect 24780 24704 24961 24732
rect 24673 24695 24731 24701
rect 24949 24701 24961 24704
rect 24995 24701 25007 24735
rect 24949 24695 25007 24701
rect 25041 24735 25099 24741
rect 25041 24701 25053 24735
rect 25087 24701 25099 24735
rect 25041 24695 25099 24701
rect 25133 24735 25191 24741
rect 25133 24701 25145 24735
rect 25179 24732 25191 24735
rect 25866 24732 25872 24744
rect 25179 24704 25872 24732
rect 25179 24701 25191 24704
rect 25133 24695 25191 24701
rect 22370 24664 22376 24676
rect 22204 24636 22376 24664
rect 21269 24627 21327 24633
rect 22370 24624 22376 24636
rect 22428 24664 22434 24676
rect 25056 24664 25084 24695
rect 25866 24692 25872 24704
rect 25924 24732 25930 24744
rect 26329 24735 26387 24741
rect 26329 24732 26341 24735
rect 25924 24704 26341 24732
rect 25924 24692 25930 24704
rect 26329 24701 26341 24704
rect 26375 24701 26387 24735
rect 26329 24695 26387 24701
rect 27154 24692 27160 24744
rect 27212 24692 27218 24744
rect 27249 24735 27307 24741
rect 27249 24701 27261 24735
rect 27295 24701 27307 24735
rect 27249 24695 27307 24701
rect 22428 24636 25084 24664
rect 22428 24624 22434 24636
rect 26234 24624 26240 24676
rect 26292 24664 26298 24676
rect 27264 24664 27292 24695
rect 26292 24636 27292 24664
rect 26292 24624 26298 24636
rect 27522 24624 27528 24676
rect 27580 24664 27586 24676
rect 27709 24667 27767 24673
rect 27709 24664 27721 24667
rect 27580 24636 27721 24664
rect 27580 24624 27586 24636
rect 27709 24633 27721 24636
rect 27755 24633 27767 24667
rect 27816 24664 27844 24772
rect 28074 24760 28080 24812
rect 28132 24760 28138 24812
rect 28258 24760 28264 24812
rect 28316 24760 28322 24812
rect 28534 24760 28540 24812
rect 28592 24760 28598 24812
rect 29086 24760 29092 24812
rect 29144 24760 29150 24812
rect 29178 24760 29184 24812
rect 29236 24760 29242 24812
rect 29380 24809 29408 24840
rect 29365 24803 29423 24809
rect 29365 24769 29377 24803
rect 29411 24769 29423 24803
rect 29365 24763 29423 24769
rect 29457 24803 29515 24809
rect 29457 24769 29469 24803
rect 29503 24769 29515 24803
rect 29564 24800 29592 24840
rect 29730 24828 29736 24880
rect 29788 24868 29794 24880
rect 30719 24871 30777 24877
rect 30719 24868 30731 24871
rect 29788 24840 30731 24868
rect 29788 24828 29794 24840
rect 30719 24837 30731 24840
rect 30765 24868 30777 24871
rect 31036 24868 31064 24908
rect 31497 24905 31509 24908
rect 31543 24936 31555 24939
rect 31846 24936 31852 24948
rect 31543 24908 31852 24936
rect 31543 24905 31555 24908
rect 31497 24899 31555 24905
rect 31846 24896 31852 24908
rect 31904 24896 31910 24948
rect 32125 24939 32183 24945
rect 32125 24905 32137 24939
rect 32171 24936 32183 24939
rect 32490 24936 32496 24948
rect 32171 24908 32496 24936
rect 32171 24905 32183 24908
rect 32125 24899 32183 24905
rect 32490 24896 32496 24908
rect 32548 24896 32554 24948
rect 33045 24939 33103 24945
rect 33045 24905 33057 24939
rect 33091 24936 33103 24939
rect 33134 24936 33140 24948
rect 33091 24908 33140 24936
rect 33091 24905 33103 24908
rect 33045 24899 33103 24905
rect 33134 24896 33140 24908
rect 33192 24896 33198 24948
rect 35250 24896 35256 24948
rect 35308 24936 35314 24948
rect 35802 24936 35808 24948
rect 35308 24908 35808 24936
rect 35308 24896 35314 24908
rect 35802 24896 35808 24908
rect 35860 24896 35866 24948
rect 30765 24840 31064 24868
rect 30765 24837 30777 24840
rect 30719 24831 30777 24837
rect 31294 24828 31300 24880
rect 31352 24868 31358 24880
rect 31352 24840 31892 24868
rect 31352 24828 31358 24840
rect 30374 24800 30380 24812
rect 29564 24772 30380 24800
rect 29457 24763 29515 24769
rect 28166 24692 28172 24744
rect 28224 24732 28230 24744
rect 29472 24732 29500 24763
rect 30374 24760 30380 24772
rect 30432 24760 30438 24812
rect 30837 24803 30895 24809
rect 30837 24769 30849 24803
rect 30883 24800 30895 24803
rect 30883 24769 30896 24800
rect 30837 24763 30896 24769
rect 28224 24704 29500 24732
rect 30561 24735 30619 24741
rect 28224 24692 28230 24704
rect 30561 24701 30573 24735
rect 30607 24701 30619 24735
rect 30561 24695 30619 24701
rect 30576 24664 30604 24695
rect 27816 24636 30604 24664
rect 30868 24664 30896 24763
rect 30926 24760 30932 24812
rect 30984 24760 30990 24812
rect 31021 24803 31079 24809
rect 31021 24769 31033 24803
rect 31067 24800 31079 24803
rect 31864 24800 31892 24840
rect 31938 24828 31944 24880
rect 31996 24868 32002 24880
rect 31996 24840 33088 24868
rect 31996 24828 32002 24840
rect 32122 24800 32128 24812
rect 31067 24772 31524 24800
rect 31864 24772 32128 24800
rect 31067 24769 31079 24772
rect 31021 24763 31079 24769
rect 31496 24744 31524 24772
rect 32122 24760 32128 24772
rect 32180 24760 32186 24812
rect 32306 24760 32312 24812
rect 32364 24760 32370 24812
rect 32398 24760 32404 24812
rect 32456 24760 32462 24812
rect 32493 24803 32551 24809
rect 32493 24769 32505 24803
rect 32539 24769 32551 24803
rect 32493 24763 32551 24769
rect 31478 24692 31484 24744
rect 31536 24732 31542 24744
rect 32508 24732 32536 24763
rect 32582 24760 32588 24812
rect 32640 24800 32646 24812
rect 32677 24803 32735 24809
rect 32677 24800 32689 24803
rect 32640 24772 32689 24800
rect 32640 24760 32646 24772
rect 32677 24769 32689 24772
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 32858 24760 32864 24812
rect 32916 24760 32922 24812
rect 33060 24809 33088 24840
rect 35158 24828 35164 24880
rect 35216 24828 35222 24880
rect 33045 24803 33103 24809
rect 33045 24769 33057 24803
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33318 24760 33324 24812
rect 33376 24800 33382 24812
rect 33686 24800 33692 24812
rect 33376 24772 33692 24800
rect 33376 24760 33382 24772
rect 33686 24760 33692 24772
rect 33744 24760 33750 24812
rect 33781 24803 33839 24809
rect 33781 24769 33793 24803
rect 33827 24800 33839 24803
rect 33962 24800 33968 24812
rect 33827 24772 33968 24800
rect 33827 24769 33839 24772
rect 33781 24763 33839 24769
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 34146 24760 34152 24812
rect 34204 24760 34210 24812
rect 31536 24704 32536 24732
rect 33597 24735 33655 24741
rect 31536 24692 31542 24704
rect 33597 24701 33609 24735
rect 33643 24701 33655 24735
rect 33597 24695 33655 24701
rect 33873 24735 33931 24741
rect 33873 24701 33885 24735
rect 33919 24732 33931 24735
rect 33919 24704 34284 24732
rect 33919 24701 33931 24704
rect 33873 24695 33931 24701
rect 31665 24667 31723 24673
rect 30868 24636 31616 24664
rect 27709 24627 27767 24633
rect 5994 24596 6000 24608
rect 3191 24568 6000 24596
rect 3191 24565 3203 24568
rect 3145 24559 3203 24565
rect 5994 24556 6000 24568
rect 6052 24556 6058 24608
rect 6178 24556 6184 24608
rect 6236 24596 6242 24608
rect 7834 24596 7840 24608
rect 6236 24568 7840 24596
rect 6236 24556 6242 24568
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 8018 24556 8024 24608
rect 8076 24596 8082 24608
rect 8297 24599 8355 24605
rect 8297 24596 8309 24599
rect 8076 24568 8309 24596
rect 8076 24556 8082 24568
rect 8297 24565 8309 24568
rect 8343 24565 8355 24599
rect 8297 24559 8355 24565
rect 8478 24556 8484 24608
rect 8536 24596 8542 24608
rect 9493 24599 9551 24605
rect 9493 24596 9505 24599
rect 8536 24568 9505 24596
rect 8536 24556 8542 24568
rect 9493 24565 9505 24568
rect 9539 24565 9551 24599
rect 9493 24559 9551 24565
rect 10045 24599 10103 24605
rect 10045 24565 10057 24599
rect 10091 24596 10103 24599
rect 10410 24596 10416 24608
rect 10091 24568 10416 24596
rect 10091 24565 10103 24568
rect 10045 24559 10103 24565
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 11698 24556 11704 24608
rect 11756 24596 11762 24608
rect 11974 24596 11980 24608
rect 11756 24568 11980 24596
rect 11756 24556 11762 24568
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 12250 24556 12256 24608
rect 12308 24596 12314 24608
rect 12621 24599 12679 24605
rect 12621 24596 12633 24599
rect 12308 24568 12633 24596
rect 12308 24556 12314 24568
rect 12621 24565 12633 24568
rect 12667 24565 12679 24599
rect 12621 24559 12679 24565
rect 12986 24556 12992 24608
rect 13044 24596 13050 24608
rect 13081 24599 13139 24605
rect 13081 24596 13093 24599
rect 13044 24568 13093 24596
rect 13044 24556 13050 24568
rect 13081 24565 13093 24568
rect 13127 24565 13139 24599
rect 13081 24559 13139 24565
rect 15470 24556 15476 24608
rect 15528 24556 15534 24608
rect 15654 24556 15660 24608
rect 15712 24556 15718 24608
rect 17865 24599 17923 24605
rect 17865 24565 17877 24599
rect 17911 24596 17923 24599
rect 17954 24596 17960 24608
rect 17911 24568 17960 24596
rect 17911 24565 17923 24568
rect 17865 24559 17923 24565
rect 17954 24556 17960 24568
rect 18012 24556 18018 24608
rect 18138 24556 18144 24608
rect 18196 24556 18202 24608
rect 18690 24556 18696 24608
rect 18748 24596 18754 24608
rect 19610 24596 19616 24608
rect 18748 24568 19616 24596
rect 18748 24556 18754 24568
rect 19610 24556 19616 24568
rect 19668 24556 19674 24608
rect 19702 24556 19708 24608
rect 19760 24556 19766 24608
rect 19794 24556 19800 24608
rect 19852 24596 19858 24608
rect 21358 24596 21364 24608
rect 19852 24568 21364 24596
rect 19852 24556 19858 24568
rect 21358 24556 21364 24568
rect 21416 24556 21422 24608
rect 21450 24556 21456 24608
rect 21508 24556 21514 24608
rect 21542 24556 21548 24608
rect 21600 24596 21606 24608
rect 21821 24599 21879 24605
rect 21821 24596 21833 24599
rect 21600 24568 21833 24596
rect 21600 24556 21606 24568
rect 21821 24565 21833 24568
rect 21867 24565 21879 24599
rect 21821 24559 21879 24565
rect 24118 24556 24124 24608
rect 24176 24596 24182 24608
rect 25038 24596 25044 24608
rect 24176 24568 25044 24596
rect 24176 24556 24182 24568
rect 25038 24556 25044 24568
rect 25096 24596 25102 24608
rect 25866 24596 25872 24608
rect 25096 24568 25872 24596
rect 25096 24556 25102 24568
rect 25866 24556 25872 24568
rect 25924 24556 25930 24608
rect 25958 24556 25964 24608
rect 26016 24556 26022 24608
rect 27154 24556 27160 24608
rect 27212 24596 27218 24608
rect 28350 24596 28356 24608
rect 27212 24568 28356 24596
rect 27212 24556 27218 24568
rect 28350 24556 28356 24568
rect 28408 24596 28414 24608
rect 29270 24596 29276 24608
rect 28408 24568 29276 24596
rect 28408 24556 28414 24568
rect 29270 24556 29276 24568
rect 29328 24556 29334 24608
rect 29641 24599 29699 24605
rect 29641 24565 29653 24599
rect 29687 24596 29699 24599
rect 30926 24596 30932 24608
rect 29687 24568 30932 24596
rect 29687 24565 29699 24568
rect 29641 24559 29699 24565
rect 30926 24556 30932 24568
rect 30984 24556 30990 24608
rect 31018 24556 31024 24608
rect 31076 24596 31082 24608
rect 31205 24599 31263 24605
rect 31205 24596 31217 24599
rect 31076 24568 31217 24596
rect 31076 24556 31082 24568
rect 31205 24565 31217 24568
rect 31251 24565 31263 24599
rect 31205 24559 31263 24565
rect 31294 24556 31300 24608
rect 31352 24596 31358 24608
rect 31481 24599 31539 24605
rect 31481 24596 31493 24599
rect 31352 24568 31493 24596
rect 31352 24556 31358 24568
rect 31481 24565 31493 24568
rect 31527 24565 31539 24599
rect 31588 24596 31616 24636
rect 31665 24633 31677 24667
rect 31711 24664 31723 24667
rect 33612 24664 33640 24695
rect 31711 24636 33640 24664
rect 31711 24633 31723 24636
rect 31665 24627 31723 24633
rect 31754 24596 31760 24608
rect 31588 24568 31760 24596
rect 31481 24559 31539 24565
rect 31754 24556 31760 24568
rect 31812 24596 31818 24608
rect 31938 24596 31944 24608
rect 31812 24568 31944 24596
rect 31812 24556 31818 24568
rect 31938 24556 31944 24568
rect 31996 24556 32002 24608
rect 32122 24556 32128 24608
rect 32180 24596 32186 24608
rect 32398 24596 32404 24608
rect 32180 24568 32404 24596
rect 32180 24556 32186 24568
rect 32398 24556 32404 24568
rect 32456 24556 32462 24608
rect 32582 24556 32588 24608
rect 32640 24596 32646 24608
rect 33226 24596 33232 24608
rect 32640 24568 33232 24596
rect 32640 24556 32646 24568
rect 33226 24556 33232 24568
rect 33284 24556 33290 24608
rect 34054 24556 34060 24608
rect 34112 24556 34118 24608
rect 34256 24596 34284 24704
rect 34422 24692 34428 24744
rect 34480 24692 34486 24744
rect 36170 24692 36176 24744
rect 36228 24692 36234 24744
rect 34606 24596 34612 24608
rect 34256 24568 34612 24596
rect 34606 24556 34612 24568
rect 34664 24556 34670 24608
rect 1104 24506 36524 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 36524 24506
rect 1104 24432 36524 24454
rect 4614 24352 4620 24404
rect 4672 24392 4678 24404
rect 4709 24395 4767 24401
rect 4709 24392 4721 24395
rect 4672 24364 4721 24392
rect 4672 24352 4678 24364
rect 4709 24361 4721 24364
rect 4755 24361 4767 24395
rect 7098 24392 7104 24404
rect 4709 24355 4767 24361
rect 5276 24364 7104 24392
rect 4062 24284 4068 24336
rect 4120 24324 4126 24336
rect 5276 24324 5304 24364
rect 7098 24352 7104 24364
rect 7156 24352 7162 24404
rect 7282 24352 7288 24404
rect 7340 24352 7346 24404
rect 11422 24352 11428 24404
rect 11480 24352 11486 24404
rect 11606 24352 11612 24404
rect 11664 24392 11670 24404
rect 12161 24395 12219 24401
rect 12161 24392 12173 24395
rect 11664 24364 12173 24392
rect 11664 24352 11670 24364
rect 12161 24361 12173 24364
rect 12207 24361 12219 24395
rect 12161 24355 12219 24361
rect 12345 24395 12403 24401
rect 12345 24361 12357 24395
rect 12391 24392 12403 24395
rect 12526 24392 12532 24404
rect 12391 24364 12532 24392
rect 12391 24361 12403 24364
rect 12345 24355 12403 24361
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 14090 24352 14096 24404
rect 14148 24352 14154 24404
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 15749 24395 15807 24401
rect 15749 24392 15761 24395
rect 14516 24364 15761 24392
rect 14516 24352 14522 24364
rect 6270 24324 6276 24336
rect 4120 24296 5304 24324
rect 5368 24296 6276 24324
rect 4120 24284 4126 24296
rect 3602 24216 3608 24268
rect 3660 24256 3666 24268
rect 5368 24265 5396 24296
rect 6270 24284 6276 24296
rect 6328 24324 6334 24336
rect 6328 24296 7880 24324
rect 6328 24284 6334 24296
rect 7852 24268 7880 24296
rect 8386 24284 8392 24336
rect 8444 24284 8450 24336
rect 10134 24284 10140 24336
rect 10192 24324 10198 24336
rect 10229 24327 10287 24333
rect 10229 24324 10241 24327
rect 10192 24296 10241 24324
rect 10192 24284 10198 24296
rect 10229 24293 10241 24296
rect 10275 24293 10287 24327
rect 10229 24287 10287 24293
rect 10318 24284 10324 24336
rect 10376 24324 10382 24336
rect 12710 24324 12716 24336
rect 10376 24296 12716 24324
rect 10376 24284 10382 24296
rect 5353 24259 5411 24265
rect 3660 24228 5212 24256
rect 3660 24216 3666 24228
rect 3418 24148 3424 24200
rect 3476 24148 3482 24200
rect 4522 24148 4528 24200
rect 4580 24148 4586 24200
rect 5184 24197 5212 24228
rect 5353 24225 5365 24259
rect 5399 24225 5411 24259
rect 5353 24219 5411 24225
rect 5902 24216 5908 24268
rect 5960 24256 5966 24268
rect 6089 24259 6147 24265
rect 6089 24256 6101 24259
rect 5960 24228 6101 24256
rect 5960 24216 5966 24228
rect 6089 24225 6101 24228
rect 6135 24225 6147 24259
rect 7190 24256 7196 24268
rect 6089 24219 6147 24225
rect 6564 24228 7196 24256
rect 5169 24191 5227 24197
rect 5169 24157 5181 24191
rect 5215 24188 5227 24191
rect 6178 24188 6184 24200
rect 5215 24160 6184 24188
rect 5215 24157 5227 24160
rect 5169 24151 5227 24157
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 6454 24148 6460 24200
rect 6512 24148 6518 24200
rect 6564 24197 6592 24228
rect 7190 24216 7196 24228
rect 7248 24216 7254 24268
rect 7834 24216 7840 24268
rect 7892 24216 7898 24268
rect 8757 24259 8815 24265
rect 8757 24225 8769 24259
rect 8803 24256 8815 24259
rect 8803 24228 10364 24256
rect 8803 24225 8815 24228
rect 8757 24219 8815 24225
rect 10336 24200 10364 24228
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24157 6607 24191
rect 6549 24151 6607 24157
rect 6822 24148 6828 24200
rect 6880 24148 6886 24200
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24188 7711 24191
rect 8018 24188 8024 24200
rect 7699 24160 8024 24188
rect 7699 24157 7711 24160
rect 7653 24151 7711 24157
rect 8018 24148 8024 24160
rect 8076 24148 8082 24200
rect 8573 24191 8631 24197
rect 8573 24157 8585 24191
rect 8619 24157 8631 24191
rect 8573 24151 8631 24157
rect 9585 24191 9643 24197
rect 9585 24157 9597 24191
rect 9631 24188 9643 24191
rect 9766 24188 9772 24200
rect 9631 24160 9772 24188
rect 9631 24157 9643 24160
rect 9585 24151 9643 24157
rect 5077 24123 5135 24129
rect 5077 24089 5089 24123
rect 5123 24120 5135 24123
rect 5537 24123 5595 24129
rect 5537 24120 5549 24123
rect 5123 24092 5549 24120
rect 5123 24089 5135 24092
rect 5077 24083 5135 24089
rect 5537 24089 5549 24092
rect 5583 24089 5595 24123
rect 5537 24083 5595 24089
rect 6638 24080 6644 24132
rect 6696 24080 6702 24132
rect 8205 24123 8263 24129
rect 8205 24089 8217 24123
rect 8251 24120 8263 24123
rect 8478 24120 8484 24132
rect 8251 24092 8484 24120
rect 8251 24089 8263 24092
rect 8205 24083 8263 24089
rect 8478 24080 8484 24092
rect 8536 24080 8542 24132
rect 2314 24012 2320 24064
rect 2372 24052 2378 24064
rect 2777 24055 2835 24061
rect 2777 24052 2789 24055
rect 2372 24024 2789 24052
rect 2372 24012 2378 24024
rect 2777 24021 2789 24024
rect 2823 24021 2835 24055
rect 2777 24015 2835 24021
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 4614 24052 4620 24064
rect 4019 24024 4620 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 6270 24012 6276 24064
rect 6328 24012 6334 24064
rect 7745 24055 7803 24061
rect 7745 24021 7757 24055
rect 7791 24052 7803 24055
rect 8386 24052 8392 24064
rect 7791 24024 8392 24052
rect 7791 24021 7803 24024
rect 7745 24015 7803 24021
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 8588 24052 8616 24151
rect 9766 24148 9772 24160
rect 9824 24148 9830 24200
rect 9953 24191 10011 24197
rect 9953 24157 9965 24191
rect 9999 24188 10011 24191
rect 10134 24188 10140 24200
rect 9999 24160 10140 24188
rect 9999 24157 10011 24160
rect 9953 24151 10011 24157
rect 10134 24148 10140 24160
rect 10192 24148 10198 24200
rect 10318 24148 10324 24200
rect 10376 24148 10382 24200
rect 10612 24188 10640 24296
rect 12710 24284 12716 24296
rect 12768 24284 12774 24336
rect 10689 24259 10747 24265
rect 10689 24225 10701 24259
rect 10735 24256 10747 24259
rect 10870 24256 10876 24268
rect 10735 24228 10876 24256
rect 10735 24225 10747 24228
rect 10689 24219 10747 24225
rect 10870 24216 10876 24228
rect 10928 24256 10934 24268
rect 11609 24259 11667 24265
rect 11609 24256 11621 24259
rect 10928 24228 11621 24256
rect 10928 24216 10934 24228
rect 11609 24225 11621 24228
rect 11655 24225 11667 24259
rect 11609 24219 11667 24225
rect 11974 24216 11980 24268
rect 12032 24216 12038 24268
rect 13538 24256 13544 24268
rect 13096 24228 13544 24256
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 10612 24160 10793 24188
rect 9858 24080 9864 24132
rect 9916 24120 9922 24132
rect 10704 24120 10732 24160
rect 10781 24157 10793 24160
rect 10827 24157 10839 24191
rect 11152 24191 11210 24197
rect 11152 24188 11164 24191
rect 10781 24151 10839 24157
rect 11072 24160 11164 24188
rect 9916 24092 10732 24120
rect 9916 24080 9922 24092
rect 10042 24052 10048 24064
rect 8588 24024 10048 24052
rect 10042 24012 10048 24024
rect 10100 24012 10106 24064
rect 10594 24012 10600 24064
rect 10652 24052 10658 24064
rect 10778 24052 10784 24064
rect 10652 24024 10784 24052
rect 10652 24012 10658 24024
rect 10778 24012 10784 24024
rect 10836 24052 10842 24064
rect 11072 24052 11100 24160
rect 11152 24157 11164 24160
rect 11198 24157 11210 24191
rect 11152 24151 11210 24157
rect 11698 24148 11704 24200
rect 11756 24148 11762 24200
rect 11992 24120 12020 24216
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12400 24160 12664 24188
rect 12400 24148 12406 24160
rect 11164 24092 12020 24120
rect 12069 24123 12127 24129
rect 11164 24061 11192 24092
rect 12069 24089 12081 24123
rect 12115 24089 12127 24123
rect 12069 24083 12127 24089
rect 10836 24024 11100 24052
rect 11149 24055 11207 24061
rect 10836 24012 10842 24024
rect 11149 24021 11161 24055
rect 11195 24021 11207 24055
rect 11149 24015 11207 24021
rect 11333 24055 11391 24061
rect 11333 24021 11345 24055
rect 11379 24052 11391 24055
rect 11882 24052 11888 24064
rect 11379 24024 11888 24052
rect 11379 24021 11391 24024
rect 11333 24015 11391 24021
rect 11882 24012 11888 24024
rect 11940 24012 11946 24064
rect 11974 24012 11980 24064
rect 12032 24052 12038 24064
rect 12084 24052 12112 24083
rect 12158 24080 12164 24132
rect 12216 24120 12222 24132
rect 12529 24123 12587 24129
rect 12529 24120 12541 24123
rect 12216 24092 12541 24120
rect 12216 24080 12222 24092
rect 12529 24089 12541 24092
rect 12575 24089 12587 24123
rect 12636 24120 12664 24160
rect 12710 24148 12716 24200
rect 12768 24148 12774 24200
rect 12806 24191 12864 24197
rect 12806 24157 12818 24191
rect 12852 24157 12864 24191
rect 12806 24151 12864 24157
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24188 13047 24191
rect 13096 24188 13124 24228
rect 13538 24216 13544 24228
rect 13596 24216 13602 24268
rect 15396 24256 15424 24364
rect 15749 24361 15761 24364
rect 15795 24361 15807 24395
rect 15749 24355 15807 24361
rect 15933 24395 15991 24401
rect 15933 24361 15945 24395
rect 15979 24392 15991 24395
rect 16390 24392 16396 24404
rect 15979 24364 16396 24392
rect 15979 24361 15991 24364
rect 15933 24355 15991 24361
rect 16390 24352 16396 24364
rect 16448 24352 16454 24404
rect 17034 24352 17040 24404
rect 17092 24392 17098 24404
rect 19702 24392 19708 24404
rect 17092 24364 19708 24392
rect 17092 24352 17098 24364
rect 19702 24352 19708 24364
rect 19760 24352 19766 24404
rect 19812 24364 22324 24392
rect 15470 24284 15476 24336
rect 15528 24324 15534 24336
rect 16209 24327 16267 24333
rect 16209 24324 16221 24327
rect 15528 24296 16221 24324
rect 15528 24284 15534 24296
rect 16209 24293 16221 24296
rect 16255 24293 16267 24327
rect 16209 24287 16267 24293
rect 19426 24284 19432 24336
rect 19484 24324 19490 24336
rect 19812 24324 19840 24364
rect 19484 24296 19840 24324
rect 19484 24284 19490 24296
rect 19886 24284 19892 24336
rect 19944 24324 19950 24336
rect 20073 24327 20131 24333
rect 20073 24324 20085 24327
rect 19944 24296 20085 24324
rect 19944 24284 19950 24296
rect 20073 24293 20085 24296
rect 20119 24293 20131 24327
rect 22296 24324 22324 24364
rect 22370 24352 22376 24404
rect 22428 24352 22434 24404
rect 22922 24352 22928 24404
rect 22980 24392 22986 24404
rect 23382 24392 23388 24404
rect 22980 24364 23388 24392
rect 22980 24352 22986 24364
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 25958 24352 25964 24404
rect 26016 24401 26022 24404
rect 26016 24395 26065 24401
rect 26016 24361 26019 24395
rect 26053 24361 26065 24395
rect 26016 24355 26065 24361
rect 26145 24395 26203 24401
rect 26145 24361 26157 24395
rect 26191 24392 26203 24395
rect 26510 24392 26516 24404
rect 26191 24364 26516 24392
rect 26191 24361 26203 24364
rect 26145 24355 26203 24361
rect 26016 24352 26022 24355
rect 26510 24352 26516 24364
rect 26568 24352 26574 24404
rect 27617 24395 27675 24401
rect 27617 24361 27629 24395
rect 27663 24361 27675 24395
rect 27617 24355 27675 24361
rect 27632 24324 27660 24355
rect 28350 24352 28356 24404
rect 28408 24392 28414 24404
rect 28721 24395 28779 24401
rect 28721 24392 28733 24395
rect 28408 24364 28733 24392
rect 28408 24352 28414 24364
rect 28721 24361 28733 24364
rect 28767 24361 28779 24395
rect 28721 24355 28779 24361
rect 28994 24352 29000 24404
rect 29052 24352 29058 24404
rect 29178 24352 29184 24404
rect 29236 24352 29242 24404
rect 30374 24352 30380 24404
rect 30432 24392 30438 24404
rect 31662 24392 31668 24404
rect 30432 24364 31668 24392
rect 30432 24352 30438 24364
rect 31662 24352 31668 24364
rect 31720 24352 31726 24404
rect 32600 24364 33272 24392
rect 32600 24324 32628 24364
rect 22296 24296 32628 24324
rect 32677 24327 32735 24333
rect 20073 24287 20131 24293
rect 32677 24293 32689 24327
rect 32723 24324 32735 24327
rect 33042 24324 33048 24336
rect 32723 24296 33048 24324
rect 32723 24293 32735 24296
rect 32677 24287 32735 24293
rect 33042 24284 33048 24296
rect 33100 24284 33106 24336
rect 33244 24324 33272 24364
rect 33318 24352 33324 24404
rect 33376 24352 33382 24404
rect 33428 24364 33732 24392
rect 33428 24324 33456 24364
rect 33244 24296 33456 24324
rect 33597 24327 33655 24333
rect 33597 24293 33609 24327
rect 33643 24293 33655 24327
rect 33704 24324 33732 24364
rect 33778 24352 33784 24404
rect 33836 24352 33842 24404
rect 34422 24352 34428 24404
rect 34480 24392 34486 24404
rect 34701 24395 34759 24401
rect 34701 24392 34713 24395
rect 34480 24364 34713 24392
rect 34480 24352 34486 24364
rect 34701 24361 34713 24364
rect 34747 24361 34759 24395
rect 34701 24355 34759 24361
rect 35158 24352 35164 24404
rect 35216 24392 35222 24404
rect 35802 24392 35808 24404
rect 35216 24364 35808 24392
rect 35216 24352 35222 24364
rect 35802 24352 35808 24364
rect 35860 24352 35866 24404
rect 35345 24327 35403 24333
rect 35345 24324 35357 24327
rect 33704 24296 35357 24324
rect 33597 24287 33655 24293
rect 35345 24293 35357 24296
rect 35391 24324 35403 24327
rect 36354 24324 36360 24336
rect 35391 24296 36360 24324
rect 35391 24293 35403 24296
rect 35345 24287 35403 24293
rect 14292 24228 15332 24256
rect 15396 24228 16620 24256
rect 14292 24200 14320 24228
rect 13035 24160 13124 24188
rect 13219 24191 13277 24197
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13219 24157 13231 24191
rect 13265 24188 13277 24191
rect 13630 24188 13636 24200
rect 13265 24160 13636 24188
rect 13265 24157 13277 24160
rect 13219 24151 13277 24157
rect 12820 24120 12848 24151
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 14274 24148 14280 24200
rect 14332 24148 14338 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 14642 24148 14648 24200
rect 14700 24148 14706 24200
rect 15304 24188 15332 24228
rect 16592 24197 16620 24228
rect 18138 24216 18144 24268
rect 18196 24256 18202 24268
rect 19058 24256 19064 24268
rect 18196 24228 19064 24256
rect 18196 24216 18202 24228
rect 19058 24216 19064 24228
rect 19116 24256 19122 24268
rect 22557 24259 22615 24265
rect 22557 24256 22569 24259
rect 19116 24228 22569 24256
rect 19116 24216 19122 24228
rect 22557 24225 22569 24228
rect 22603 24225 22615 24259
rect 22557 24219 22615 24225
rect 22925 24259 22983 24265
rect 22925 24225 22937 24259
rect 22971 24256 22983 24259
rect 23290 24256 23296 24268
rect 22971 24228 23296 24256
rect 22971 24225 22983 24228
rect 22925 24219 22983 24225
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 27338 24216 27344 24268
rect 27396 24256 27402 24268
rect 32858 24256 32864 24268
rect 27396 24228 28994 24256
rect 27396 24216 27402 24228
rect 16393 24191 16451 24197
rect 16393 24188 16405 24191
rect 15304 24160 16405 24188
rect 16393 24157 16405 24160
rect 16439 24157 16451 24191
rect 16393 24151 16451 24157
rect 16577 24191 16635 24197
rect 16577 24157 16589 24191
rect 16623 24157 16635 24191
rect 16577 24151 16635 24157
rect 12636 24092 12848 24120
rect 13081 24123 13139 24129
rect 12529 24083 12587 24089
rect 13081 24089 13093 24123
rect 13127 24120 13139 24123
rect 13814 24120 13820 24132
rect 13127 24092 13820 24120
rect 13127 24089 13139 24092
rect 13081 24083 13139 24089
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 14369 24123 14427 24129
rect 14369 24089 14381 24123
rect 14415 24120 14427 24123
rect 15010 24120 15016 24132
rect 14415 24092 15016 24120
rect 14415 24089 14427 24092
rect 14369 24083 14427 24089
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 16114 24080 16120 24132
rect 16172 24080 16178 24132
rect 12032 24024 12112 24052
rect 12329 24055 12387 24061
rect 12032 24012 12038 24024
rect 12329 24021 12341 24055
rect 12375 24052 12387 24055
rect 12710 24052 12716 24064
rect 12375 24024 12716 24052
rect 12375 24021 12387 24024
rect 12329 24015 12387 24021
rect 12710 24012 12716 24024
rect 12768 24052 12774 24064
rect 12894 24052 12900 24064
rect 12768 24024 12900 24052
rect 12768 24012 12774 24024
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 13170 24012 13176 24064
rect 13228 24052 13234 24064
rect 13357 24055 13415 24061
rect 13357 24052 13369 24055
rect 13228 24024 13369 24052
rect 13228 24012 13234 24024
rect 13357 24021 13369 24024
rect 13403 24021 13415 24055
rect 13357 24015 13415 24021
rect 15933 24055 15991 24061
rect 15933 24021 15945 24055
rect 15979 24052 15991 24055
rect 16022 24052 16028 24064
rect 15979 24024 16028 24052
rect 15979 24021 15991 24024
rect 15933 24015 15991 24021
rect 16022 24012 16028 24024
rect 16080 24012 16086 24064
rect 16408 24052 16436 24151
rect 16758 24148 16764 24200
rect 16816 24148 16822 24200
rect 17218 24148 17224 24200
rect 17276 24188 17282 24200
rect 17678 24188 17684 24200
rect 17276 24160 17684 24188
rect 17276 24148 17282 24160
rect 17678 24148 17684 24160
rect 17736 24188 17742 24200
rect 19610 24188 19616 24200
rect 17736 24160 19616 24188
rect 17736 24148 17742 24160
rect 19610 24148 19616 24160
rect 19668 24148 19674 24200
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24188 20039 24191
rect 20346 24188 20352 24200
rect 20027 24160 20352 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 16485 24123 16543 24129
rect 16485 24089 16497 24123
rect 16531 24120 16543 24123
rect 17586 24120 17592 24132
rect 16531 24092 17592 24120
rect 16531 24089 16543 24092
rect 16485 24083 16543 24089
rect 17586 24080 17592 24092
rect 17644 24120 17650 24132
rect 19426 24120 19432 24132
rect 17644 24092 19432 24120
rect 17644 24080 17650 24092
rect 19426 24080 19432 24092
rect 19484 24080 19490 24132
rect 19720 24120 19748 24151
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 22738 24148 22744 24200
rect 22796 24148 22802 24200
rect 22833 24191 22891 24197
rect 22833 24157 22845 24191
rect 22879 24157 22891 24191
rect 22833 24151 22891 24157
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 19720 24092 20085 24120
rect 20073 24089 20085 24092
rect 20119 24120 20131 24123
rect 20622 24120 20628 24132
rect 20119 24092 20628 24120
rect 20119 24089 20131 24092
rect 20073 24083 20131 24089
rect 20622 24080 20628 24092
rect 20680 24080 20686 24132
rect 22848 24120 22876 24151
rect 23014 24148 23020 24200
rect 23072 24188 23078 24200
rect 24489 24191 24547 24197
rect 24489 24188 24501 24191
rect 23072 24160 24501 24188
rect 23072 24148 23078 24160
rect 24489 24157 24501 24160
rect 24535 24157 24547 24191
rect 24489 24151 24547 24157
rect 24670 24148 24676 24200
rect 24728 24148 24734 24200
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24188 24823 24191
rect 24854 24188 24860 24200
rect 24811 24160 24860 24188
rect 24811 24157 24823 24160
rect 24765 24151 24823 24157
rect 24854 24148 24860 24160
rect 24912 24148 24918 24200
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 25038 24148 25044 24200
rect 25096 24148 25102 24200
rect 25130 24148 25136 24200
rect 25188 24148 25194 24200
rect 25317 24191 25375 24197
rect 25317 24157 25329 24191
rect 25363 24188 25375 24191
rect 25774 24188 25780 24200
rect 25363 24160 25780 24188
rect 25363 24157 25375 24160
rect 25317 24151 25375 24157
rect 25774 24148 25780 24160
rect 25832 24148 25838 24200
rect 25866 24148 25872 24200
rect 25924 24148 25930 24200
rect 26326 24148 26332 24200
rect 26384 24148 26390 24200
rect 27154 24148 27160 24200
rect 27212 24188 27218 24200
rect 27249 24191 27307 24197
rect 27249 24188 27261 24191
rect 27212 24160 27261 24188
rect 27212 24148 27218 24160
rect 27249 24157 27261 24160
rect 27295 24157 27307 24191
rect 27249 24151 27307 24157
rect 28166 24148 28172 24200
rect 28224 24148 28230 24200
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24188 28595 24191
rect 28718 24188 28724 24200
rect 28583 24160 28724 24188
rect 28583 24157 28595 24160
rect 28537 24151 28595 24157
rect 28718 24148 28724 24160
rect 28776 24148 28782 24200
rect 22922 24120 22928 24132
rect 22848 24092 22928 24120
rect 22922 24080 22928 24092
rect 22980 24080 22986 24132
rect 23569 24123 23627 24129
rect 23569 24089 23581 24123
rect 23615 24120 23627 24123
rect 23750 24120 23756 24132
rect 23615 24092 23756 24120
rect 23615 24089 23627 24092
rect 23569 24083 23627 24089
rect 23750 24080 23756 24092
rect 23808 24080 23814 24132
rect 25498 24080 25504 24132
rect 25556 24080 25562 24132
rect 27617 24123 27675 24129
rect 27617 24089 27629 24123
rect 27663 24120 27675 24123
rect 27706 24120 27712 24132
rect 27663 24092 27712 24120
rect 27663 24089 27675 24092
rect 27617 24083 27675 24089
rect 27706 24080 27712 24092
rect 27764 24080 27770 24132
rect 28445 24123 28503 24129
rect 28445 24089 28457 24123
rect 28491 24089 28503 24123
rect 28445 24083 28503 24089
rect 28859 24123 28917 24129
rect 28859 24089 28871 24123
rect 28905 24120 28917 24123
rect 28966 24120 28994 24228
rect 32692 24228 32864 24256
rect 29270 24148 29276 24200
rect 29328 24188 29334 24200
rect 31021 24191 31079 24197
rect 31021 24188 31033 24191
rect 29328 24160 31033 24188
rect 29328 24148 29334 24160
rect 31021 24157 31033 24160
rect 31067 24188 31079 24191
rect 31110 24188 31116 24200
rect 31067 24160 31116 24188
rect 31067 24157 31079 24160
rect 31021 24151 31079 24157
rect 31110 24148 31116 24160
rect 31168 24148 31174 24200
rect 32490 24148 32496 24200
rect 32548 24148 32554 24200
rect 32692 24197 32720 24228
rect 32858 24216 32864 24228
rect 32916 24256 32922 24268
rect 33612 24256 33640 24287
rect 36354 24284 36360 24296
rect 36412 24284 36418 24336
rect 32916 24228 33640 24256
rect 32916 24216 32922 24228
rect 33870 24216 33876 24268
rect 33928 24216 33934 24268
rect 36170 24256 36176 24268
rect 34992 24228 36176 24256
rect 34992 24200 35020 24228
rect 36170 24216 36176 24228
rect 36228 24216 36234 24268
rect 32677 24191 32735 24197
rect 32677 24157 32689 24191
rect 32723 24157 32735 24191
rect 32677 24151 32735 24157
rect 32766 24148 32772 24200
rect 32824 24148 32830 24200
rect 33060 24197 33364 24198
rect 33045 24191 33364 24197
rect 33045 24157 33057 24191
rect 33091 24188 33364 24191
rect 33965 24191 34023 24197
rect 33091 24170 33916 24188
rect 33091 24157 33103 24170
rect 33336 24160 33916 24170
rect 33045 24151 33103 24157
rect 28905 24092 28994 24120
rect 29029 24123 29087 24129
rect 28905 24089 28917 24092
rect 28859 24083 28917 24089
rect 29029 24089 29041 24123
rect 29075 24120 29087 24123
rect 29730 24120 29736 24132
rect 29075 24092 29736 24120
rect 29075 24089 29087 24092
rect 29029 24083 29087 24089
rect 17310 24052 17316 24064
rect 16408 24024 17316 24052
rect 17310 24012 17316 24024
rect 17368 24012 17374 24064
rect 19518 24012 19524 24064
rect 19576 24052 19582 24064
rect 19794 24052 19800 24064
rect 19576 24024 19800 24052
rect 19576 24012 19582 24024
rect 19794 24012 19800 24024
rect 19852 24012 19858 24064
rect 19889 24055 19947 24061
rect 19889 24021 19901 24055
rect 19935 24052 19947 24055
rect 20162 24052 20168 24064
rect 19935 24024 20168 24052
rect 19935 24021 19947 24024
rect 19889 24015 19947 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 20257 24055 20315 24061
rect 20257 24021 20269 24055
rect 20303 24052 20315 24055
rect 21818 24052 21824 24064
rect 20303 24024 21824 24052
rect 20303 24021 20315 24024
rect 20257 24015 20315 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 22462 24012 22468 24064
rect 22520 24052 22526 24064
rect 23201 24055 23259 24061
rect 23201 24052 23213 24055
rect 22520 24024 23213 24052
rect 22520 24012 22526 24024
rect 23201 24021 23213 24024
rect 23247 24021 23259 24055
rect 23201 24015 23259 24021
rect 23369 24055 23427 24061
rect 23369 24021 23381 24055
rect 23415 24052 23427 24055
rect 23658 24052 23664 24064
rect 23415 24024 23664 24052
rect 23415 24021 23427 24024
rect 23369 24015 23427 24021
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 25516 24052 25544 24080
rect 25188 24024 25544 24052
rect 25188 24012 25194 24024
rect 25590 24012 25596 24064
rect 25648 24052 25654 24064
rect 26237 24055 26295 24061
rect 26237 24052 26249 24055
rect 25648 24024 26249 24052
rect 25648 24012 25654 24024
rect 26237 24021 26249 24024
rect 26283 24021 26295 24055
rect 26237 24015 26295 24021
rect 27801 24055 27859 24061
rect 27801 24021 27813 24055
rect 27847 24052 27859 24055
rect 28074 24052 28080 24064
rect 27847 24024 28080 24052
rect 27847 24021 27859 24024
rect 27801 24015 27859 24021
rect 28074 24012 28080 24024
rect 28132 24012 28138 24064
rect 28166 24012 28172 24064
rect 28224 24052 28230 24064
rect 28460 24052 28488 24083
rect 29730 24080 29736 24092
rect 29788 24080 29794 24132
rect 31754 24120 31760 24132
rect 31220 24092 31760 24120
rect 28224 24024 28488 24052
rect 28224 24012 28230 24024
rect 28718 24012 28724 24064
rect 28776 24052 28782 24064
rect 29914 24052 29920 24064
rect 28776 24024 29920 24052
rect 28776 24012 28782 24024
rect 29914 24012 29920 24024
rect 29972 24012 29978 24064
rect 31220 24061 31248 24092
rect 31754 24080 31760 24092
rect 31812 24080 31818 24132
rect 31938 24080 31944 24132
rect 31996 24120 32002 24132
rect 32582 24120 32588 24132
rect 31996 24092 32588 24120
rect 31996 24080 32002 24092
rect 32582 24080 32588 24092
rect 32640 24080 32646 24132
rect 32784 24120 32812 24148
rect 33888 24132 33916 24160
rect 33965 24157 33977 24191
rect 34011 24188 34023 24191
rect 34011 24160 34376 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 33410 24129 33416 24132
rect 33163 24123 33221 24129
rect 33163 24120 33175 24123
rect 32784 24092 33175 24120
rect 31205 24055 31263 24061
rect 31205 24021 31217 24055
rect 31251 24021 31263 24055
rect 31205 24015 31263 24021
rect 31662 24012 31668 24064
rect 31720 24052 31726 24064
rect 32766 24052 32772 24064
rect 31720 24024 32772 24052
rect 31720 24012 31726 24024
rect 32766 24012 32772 24024
rect 32824 24012 32830 24064
rect 32876 24061 32904 24092
rect 33163 24089 33175 24092
rect 33209 24089 33221 24123
rect 33163 24083 33221 24089
rect 33353 24123 33416 24129
rect 33353 24089 33365 24123
rect 33399 24089 33416 24123
rect 33353 24083 33416 24089
rect 33410 24080 33416 24083
rect 33468 24080 33474 24132
rect 33778 24120 33784 24132
rect 33520 24092 33784 24120
rect 33520 24061 33548 24092
rect 33778 24080 33784 24092
rect 33836 24080 33842 24132
rect 33870 24080 33876 24132
rect 33928 24080 33934 24132
rect 32861 24055 32919 24061
rect 32861 24021 32873 24055
rect 32907 24021 32919 24055
rect 32861 24015 32919 24021
rect 33505 24055 33563 24061
rect 33505 24021 33517 24055
rect 33551 24021 33563 24055
rect 33505 24015 33563 24021
rect 33594 24012 33600 24064
rect 33652 24052 33658 24064
rect 34238 24052 34244 24064
rect 33652 24024 34244 24052
rect 33652 24012 33658 24024
rect 34238 24012 34244 24024
rect 34296 24012 34302 24064
rect 34348 24052 34376 24160
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34848 24160 34897 24188
rect 34848 24148 34854 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 34974 24148 34980 24200
rect 35032 24148 35038 24200
rect 35250 24148 35256 24200
rect 35308 24148 35314 24200
rect 36078 24148 36084 24200
rect 36136 24148 36142 24200
rect 34606 24080 34612 24132
rect 34664 24120 34670 24132
rect 35069 24123 35127 24129
rect 35069 24120 35081 24123
rect 34664 24092 35081 24120
rect 34664 24080 34670 24092
rect 35069 24089 35081 24092
rect 35115 24089 35127 24123
rect 35069 24083 35127 24089
rect 35526 24080 35532 24132
rect 35584 24080 35590 24132
rect 35342 24052 35348 24064
rect 34348 24024 35348 24052
rect 35342 24012 35348 24024
rect 35400 24012 35406 24064
rect 1104 23962 36524 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 36524 23962
rect 1104 23888 36524 23910
rect 2314 23808 2320 23860
rect 2372 23808 2378 23860
rect 4062 23848 4068 23860
rect 3436 23820 4068 23848
rect 3142 23740 3148 23792
rect 3200 23780 3206 23792
rect 3436 23780 3464 23820
rect 4062 23808 4068 23820
rect 4120 23808 4126 23860
rect 4522 23808 4528 23860
rect 4580 23808 4586 23860
rect 5166 23808 5172 23860
rect 5224 23848 5230 23860
rect 5442 23848 5448 23860
rect 5224 23820 5448 23848
rect 5224 23808 5230 23820
rect 5442 23808 5448 23820
rect 5500 23808 5506 23860
rect 5994 23848 6000 23860
rect 5552 23820 6000 23848
rect 4540 23780 4568 23808
rect 5552 23789 5580 23820
rect 5994 23808 6000 23820
rect 6052 23848 6058 23860
rect 8662 23848 8668 23860
rect 6052 23820 8668 23848
rect 6052 23808 6058 23820
rect 8662 23808 8668 23820
rect 8720 23808 8726 23860
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 10045 23851 10103 23857
rect 10045 23848 10057 23851
rect 9732 23820 10057 23848
rect 9732 23808 9738 23820
rect 10045 23817 10057 23820
rect 10091 23817 10103 23851
rect 10045 23811 10103 23817
rect 10134 23808 10140 23860
rect 10192 23848 10198 23860
rect 10229 23851 10287 23857
rect 10229 23848 10241 23851
rect 10192 23820 10241 23848
rect 10192 23808 10198 23820
rect 10229 23817 10241 23820
rect 10275 23817 10287 23851
rect 10229 23811 10287 23817
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 14274 23848 14280 23860
rect 10376 23820 12388 23848
rect 10376 23808 10382 23820
rect 5537 23783 5595 23789
rect 3200 23752 3542 23780
rect 4540 23752 5304 23780
rect 3200 23740 3206 23752
rect 2682 23672 2688 23724
rect 2740 23712 2746 23724
rect 2774 23712 2780 23724
rect 2740 23684 2780 23712
rect 2740 23672 2746 23684
rect 2774 23672 2780 23684
rect 2832 23672 2838 23724
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 5276 23721 5304 23752
rect 5537 23749 5549 23783
rect 5583 23749 5595 23783
rect 6638 23780 6644 23792
rect 5537 23743 5595 23749
rect 5690 23752 6644 23780
rect 5262 23715 5320 23721
rect 5262 23681 5274 23715
rect 5308 23681 5320 23715
rect 5262 23675 5320 23681
rect 5350 23672 5356 23724
rect 5408 23712 5414 23724
rect 5690 23721 5718 23752
rect 6638 23740 6644 23752
rect 6696 23740 6702 23792
rect 7098 23740 7104 23792
rect 7156 23740 7162 23792
rect 9214 23740 9220 23792
rect 9272 23740 9278 23792
rect 12360 23789 12388 23820
rect 13740 23820 14280 23848
rect 12345 23783 12403 23789
rect 12345 23749 12357 23783
rect 12391 23749 12403 23783
rect 12345 23743 12403 23749
rect 5445 23715 5503 23721
rect 5445 23712 5457 23715
rect 5408 23684 5457 23712
rect 5408 23672 5414 23684
rect 5445 23681 5457 23684
rect 5491 23681 5503 23715
rect 5445 23675 5503 23681
rect 5675 23715 5733 23721
rect 5675 23681 5687 23715
rect 5721 23681 5733 23715
rect 5675 23675 5733 23681
rect 8941 23715 8999 23721
rect 8941 23681 8953 23715
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 2314 23604 2320 23656
rect 2372 23644 2378 23656
rect 2409 23647 2467 23653
rect 2409 23644 2421 23647
rect 2372 23616 2421 23644
rect 2372 23604 2378 23616
rect 2409 23613 2421 23616
rect 2455 23613 2467 23647
rect 2409 23607 2467 23613
rect 2590 23604 2596 23656
rect 2648 23604 2654 23656
rect 3050 23604 3056 23656
rect 3108 23604 3114 23656
rect 4706 23604 4712 23656
rect 4764 23644 4770 23656
rect 6365 23647 6423 23653
rect 6365 23644 6377 23647
rect 4764 23616 6377 23644
rect 4764 23604 4770 23616
rect 6365 23613 6377 23616
rect 6411 23613 6423 23647
rect 6365 23607 6423 23613
rect 6641 23647 6699 23653
rect 6641 23613 6653 23647
rect 6687 23644 6699 23647
rect 7006 23644 7012 23656
rect 6687 23616 7012 23644
rect 6687 23613 6699 23616
rect 6641 23607 6699 23613
rect 7006 23604 7012 23616
rect 7064 23604 7070 23656
rect 8113 23647 8171 23653
rect 8113 23613 8125 23647
rect 8159 23644 8171 23647
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 8159 23616 8769 23644
rect 8159 23613 8171 23616
rect 8113 23607 8171 23613
rect 8757 23613 8769 23616
rect 8803 23644 8815 23647
rect 8956 23644 8984 23675
rect 9122 23672 9128 23724
rect 9180 23672 9186 23724
rect 9314 23715 9372 23721
rect 9314 23681 9326 23715
rect 9360 23681 9372 23715
rect 9314 23675 9372 23681
rect 10104 23715 10162 23721
rect 10104 23681 10116 23715
rect 10150 23712 10162 23715
rect 10594 23712 10600 23724
rect 10150 23684 10600 23712
rect 10150 23681 10162 23684
rect 10104 23675 10162 23681
rect 8803 23616 8984 23644
rect 8803 23613 8815 23616
rect 8757 23607 8815 23613
rect 9214 23604 9220 23656
rect 9272 23644 9278 23656
rect 9329 23644 9357 23675
rect 10594 23672 10600 23684
rect 10652 23672 10658 23724
rect 11333 23715 11391 23721
rect 11333 23681 11345 23715
rect 11379 23712 11391 23715
rect 11422 23712 11428 23724
rect 11379 23684 11428 23712
rect 11379 23681 11391 23684
rect 11333 23675 11391 23681
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11882 23672 11888 23724
rect 11940 23672 11946 23724
rect 12434 23672 12440 23724
rect 12492 23712 12498 23724
rect 12529 23715 12587 23721
rect 12529 23712 12541 23715
rect 12492 23684 12541 23712
rect 12492 23672 12498 23684
rect 12529 23681 12541 23684
rect 12575 23681 12587 23715
rect 12529 23675 12587 23681
rect 12713 23715 12771 23721
rect 12713 23681 12725 23715
rect 12759 23712 12771 23715
rect 12894 23712 12900 23724
rect 12759 23684 12900 23712
rect 12759 23681 12771 23684
rect 12713 23675 12771 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 9272 23616 9357 23644
rect 9585 23647 9643 23653
rect 9272 23604 9278 23616
rect 9585 23613 9597 23647
rect 9631 23644 9643 23647
rect 10410 23644 10416 23656
rect 9631 23616 10416 23644
rect 9631 23613 9643 23616
rect 9585 23607 9643 23613
rect 10410 23604 10416 23616
rect 10468 23604 10474 23656
rect 11773 23647 11831 23653
rect 11773 23613 11785 23647
rect 11819 23644 11831 23647
rect 12066 23644 12072 23656
rect 11819 23616 12072 23644
rect 11819 23613 11831 23616
rect 11773 23607 11831 23613
rect 12066 23604 12072 23616
rect 12124 23604 12130 23656
rect 12158 23604 12164 23656
rect 12216 23604 12222 23656
rect 12253 23647 12311 23653
rect 12253 23613 12265 23647
rect 12299 23644 12311 23647
rect 13096 23644 13124 23675
rect 13170 23672 13176 23724
rect 13228 23672 13234 23724
rect 13354 23672 13360 23724
rect 13412 23672 13418 23724
rect 13740 23721 13768 23820
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 15933 23851 15991 23857
rect 15933 23848 15945 23851
rect 15712 23820 15945 23848
rect 15712 23808 15718 23820
rect 15933 23817 15945 23820
rect 15979 23817 15991 23851
rect 15933 23811 15991 23817
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 16448 23820 16712 23848
rect 16448 23808 16454 23820
rect 13814 23740 13820 23792
rect 13872 23740 13878 23792
rect 13909 23783 13967 23789
rect 13909 23749 13921 23783
rect 13955 23780 13967 23783
rect 14458 23780 14464 23792
rect 13955 23752 14464 23780
rect 13955 23749 13967 23752
rect 13909 23743 13967 23749
rect 14458 23740 14464 23752
rect 14516 23740 14522 23792
rect 16114 23740 16120 23792
rect 16172 23780 16178 23792
rect 16684 23789 16712 23820
rect 16942 23808 16948 23860
rect 17000 23848 17006 23860
rect 17405 23851 17463 23857
rect 17405 23848 17417 23851
rect 17000 23820 17417 23848
rect 17000 23808 17006 23820
rect 17405 23817 17417 23820
rect 17451 23817 17463 23851
rect 17405 23811 17463 23817
rect 17954 23808 17960 23860
rect 18012 23848 18018 23860
rect 18049 23851 18107 23857
rect 18049 23848 18061 23851
rect 18012 23820 18061 23848
rect 18012 23808 18018 23820
rect 18049 23817 18061 23820
rect 18095 23817 18107 23851
rect 18049 23811 18107 23817
rect 19706 23851 19764 23857
rect 19706 23817 19718 23851
rect 19752 23817 19764 23851
rect 21542 23848 21548 23860
rect 19706 23814 19764 23817
rect 19904 23820 21548 23848
rect 19904 23814 19932 23820
rect 19706 23811 19932 23814
rect 16669 23783 16727 23789
rect 16172 23752 16620 23780
rect 16172 23740 16178 23752
rect 13725 23715 13783 23721
rect 13725 23681 13737 23715
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 14090 23672 14096 23724
rect 14148 23672 14154 23724
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15381 23715 15439 23721
rect 15381 23712 15393 23715
rect 15252 23684 15393 23712
rect 15252 23672 15258 23684
rect 15381 23681 15393 23684
rect 15427 23681 15439 23715
rect 15381 23675 15439 23681
rect 15654 23672 15660 23724
rect 15712 23712 15718 23724
rect 15933 23715 15991 23721
rect 15933 23712 15945 23715
rect 15712 23684 15945 23712
rect 15712 23672 15718 23684
rect 15933 23681 15945 23684
rect 15979 23681 15991 23715
rect 15933 23675 15991 23681
rect 16298 23672 16304 23724
rect 16356 23672 16362 23724
rect 16390 23672 16396 23724
rect 16448 23712 16454 23724
rect 16485 23715 16543 23721
rect 16485 23712 16497 23715
rect 16448 23684 16497 23712
rect 16448 23672 16454 23684
rect 16485 23681 16497 23684
rect 16531 23681 16543 23715
rect 16592 23712 16620 23752
rect 16669 23749 16681 23783
rect 16715 23749 16727 23783
rect 17046 23783 17104 23789
rect 17046 23780 17058 23783
rect 16669 23743 16727 23749
rect 16960 23752 17058 23780
rect 16960 23724 16988 23752
rect 17046 23749 17058 23752
rect 17092 23749 17104 23783
rect 19150 23780 19156 23792
rect 17046 23743 17104 23749
rect 18524 23752 19156 23780
rect 16942 23712 16948 23724
rect 16592 23684 16948 23712
rect 16485 23675 16543 23681
rect 16942 23672 16948 23684
rect 17000 23672 17006 23724
rect 17310 23672 17316 23724
rect 17368 23672 17374 23724
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23712 17647 23715
rect 18046 23712 18052 23724
rect 17635 23684 18052 23712
rect 17635 23681 17647 23684
rect 17589 23675 17647 23681
rect 18046 23672 18052 23684
rect 18104 23672 18110 23724
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23712 18291 23715
rect 18322 23712 18328 23724
rect 18279 23684 18328 23712
rect 18279 23681 18291 23684
rect 18233 23675 18291 23681
rect 18322 23672 18328 23684
rect 18380 23672 18386 23724
rect 18524 23721 18552 23752
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 19720 23786 19932 23811
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 21634 23808 21640 23860
rect 21692 23848 21698 23860
rect 21821 23851 21879 23857
rect 21821 23848 21833 23851
rect 21692 23820 21833 23848
rect 21692 23808 21698 23820
rect 21821 23817 21833 23820
rect 21867 23817 21879 23851
rect 25682 23848 25688 23860
rect 21821 23811 21879 23817
rect 23032 23820 25688 23848
rect 22002 23780 22008 23792
rect 21560 23752 22008 23780
rect 21560 23724 21588 23752
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 18509 23715 18567 23721
rect 18509 23681 18521 23715
rect 18555 23681 18567 23715
rect 18509 23675 18567 23681
rect 18690 23672 18696 23724
rect 18748 23672 18754 23724
rect 18782 23672 18788 23724
rect 18840 23712 18846 23724
rect 19646 23715 19704 23721
rect 19646 23712 19658 23715
rect 18840 23684 19658 23712
rect 18840 23672 18846 23684
rect 19646 23681 19658 23684
rect 19692 23681 19704 23715
rect 19646 23675 19704 23681
rect 21542 23672 21548 23724
rect 21600 23672 21606 23724
rect 21634 23672 21640 23724
rect 21692 23712 21698 23724
rect 22097 23715 22155 23721
rect 22097 23712 22109 23715
rect 21692 23684 22109 23712
rect 21692 23672 21698 23684
rect 22097 23681 22109 23684
rect 22143 23712 22155 23715
rect 22370 23712 22376 23724
rect 22143 23684 22376 23712
rect 22143 23681 22155 23684
rect 22097 23675 22155 23681
rect 22370 23672 22376 23684
rect 22428 23672 22434 23724
rect 22554 23672 22560 23724
rect 22612 23712 22618 23724
rect 23032 23721 23060 23820
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 26510 23808 26516 23860
rect 26568 23848 26574 23860
rect 28166 23848 28172 23860
rect 26568 23820 28172 23848
rect 26568 23808 26574 23820
rect 28166 23808 28172 23820
rect 28224 23808 28230 23860
rect 28261 23851 28319 23857
rect 28261 23817 28273 23851
rect 28307 23848 28319 23851
rect 28534 23848 28540 23860
rect 28307 23820 28540 23848
rect 28307 23817 28319 23820
rect 28261 23811 28319 23817
rect 28534 23808 28540 23820
rect 28592 23808 28598 23860
rect 30190 23808 30196 23860
rect 30248 23848 30254 23860
rect 30453 23851 30511 23857
rect 30453 23848 30465 23851
rect 30248 23820 30465 23848
rect 30248 23808 30254 23820
rect 30453 23817 30465 23820
rect 30499 23848 30511 23851
rect 31037 23851 31095 23857
rect 31037 23848 31049 23851
rect 30499 23820 31049 23848
rect 30499 23817 30511 23820
rect 30453 23811 30511 23817
rect 31037 23817 31049 23820
rect 31083 23817 31095 23851
rect 33318 23848 33324 23860
rect 31037 23811 31095 23817
rect 31128 23820 33324 23848
rect 23290 23740 23296 23792
rect 23348 23780 23354 23792
rect 23750 23780 23756 23792
rect 23348 23752 23756 23780
rect 23348 23740 23354 23752
rect 23750 23740 23756 23752
rect 23808 23740 23814 23792
rect 24486 23740 24492 23792
rect 24544 23740 24550 23792
rect 25498 23780 25504 23792
rect 24872 23752 25504 23780
rect 24872 23724 24900 23752
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 22612 23684 23029 23712
rect 22612 23672 22618 23684
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 23382 23672 23388 23724
rect 23440 23672 23446 23724
rect 24670 23672 24676 23724
rect 24728 23672 24734 23724
rect 24765 23715 24823 23721
rect 24765 23681 24777 23715
rect 24811 23712 24823 23715
rect 24854 23712 24860 23724
rect 24811 23684 24860 23712
rect 24811 23681 24823 23684
rect 24765 23675 24823 23681
rect 24854 23672 24860 23684
rect 24912 23672 24918 23724
rect 24946 23672 24952 23724
rect 25004 23672 25010 23724
rect 25041 23715 25099 23721
rect 25041 23681 25053 23715
rect 25087 23712 25099 23715
rect 25222 23712 25228 23724
rect 25087 23684 25228 23712
rect 25087 23681 25099 23684
rect 25041 23675 25099 23681
rect 25222 23672 25228 23684
rect 25280 23672 25286 23724
rect 25314 23672 25320 23724
rect 25372 23672 25378 23724
rect 25424 23721 25452 23752
rect 25498 23740 25504 23752
rect 25556 23780 25562 23792
rect 25869 23783 25927 23789
rect 25869 23780 25881 23783
rect 25556 23752 25881 23780
rect 25556 23740 25562 23752
rect 25869 23749 25881 23752
rect 25915 23749 25927 23783
rect 25869 23743 25927 23749
rect 27246 23740 27252 23792
rect 27304 23780 27310 23792
rect 27304 23752 28994 23780
rect 27304 23740 27310 23752
rect 25409 23715 25467 23721
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25590 23672 25596 23724
rect 25648 23672 25654 23724
rect 25682 23672 25688 23724
rect 25740 23672 25746 23724
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23681 25835 23715
rect 25777 23675 25835 23681
rect 15286 23644 15292 23656
rect 12299 23616 12375 23644
rect 13096 23616 15292 23644
rect 12299 23613 12311 23616
rect 12253 23607 12311 23613
rect 7742 23536 7748 23588
rect 7800 23576 7806 23588
rect 8941 23579 8999 23585
rect 8941 23576 8953 23579
rect 7800 23548 8953 23576
rect 7800 23536 7806 23548
rect 8941 23545 8953 23548
rect 8987 23545 8999 23579
rect 8941 23539 8999 23545
rect 9677 23579 9735 23585
rect 9677 23545 9689 23579
rect 9723 23576 9735 23579
rect 9858 23576 9864 23588
rect 9723 23548 9864 23576
rect 9723 23545 9735 23548
rect 9677 23539 9735 23545
rect 9858 23536 9864 23548
rect 9916 23536 9922 23588
rect 10134 23536 10140 23588
rect 10192 23576 10198 23588
rect 11054 23576 11060 23588
rect 10192 23548 11060 23576
rect 10192 23536 10198 23548
rect 11054 23536 11060 23548
rect 11112 23536 11118 23588
rect 11241 23579 11299 23585
rect 11241 23545 11253 23579
rect 11287 23576 11299 23579
rect 12176 23576 12204 23604
rect 11287 23548 12204 23576
rect 11287 23545 11299 23548
rect 11241 23539 11299 23545
rect 12347 23520 12375 23616
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 15470 23604 15476 23656
rect 15528 23604 15534 23656
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 15838 23644 15844 23656
rect 15620 23616 15844 23644
rect 15620 23604 15626 23616
rect 15838 23604 15844 23616
rect 15896 23604 15902 23656
rect 17678 23604 17684 23656
rect 17736 23604 17742 23656
rect 17773 23647 17831 23653
rect 17773 23613 17785 23647
rect 17819 23613 17831 23647
rect 17773 23607 17831 23613
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 17911 23616 18644 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 13265 23579 13323 23585
rect 13265 23545 13277 23579
rect 13311 23576 13323 23579
rect 13541 23579 13599 23585
rect 13541 23576 13553 23579
rect 13311 23548 13553 23576
rect 13311 23545 13323 23548
rect 13265 23539 13323 23545
rect 13541 23545 13553 23548
rect 13587 23545 13599 23579
rect 13541 23539 13599 23545
rect 15930 23536 15936 23588
rect 15988 23576 15994 23588
rect 16298 23576 16304 23588
rect 15988 23548 16304 23576
rect 15988 23536 15994 23548
rect 16298 23536 16304 23548
rect 16356 23536 16362 23588
rect 1670 23468 1676 23520
rect 1728 23508 1734 23520
rect 1949 23511 2007 23517
rect 1949 23508 1961 23511
rect 1728 23480 1961 23508
rect 1728 23468 1734 23480
rect 1949 23477 1961 23480
rect 1995 23477 2007 23511
rect 1949 23471 2007 23477
rect 3234 23468 3240 23520
rect 3292 23508 3298 23520
rect 4982 23508 4988 23520
rect 3292 23480 4988 23508
rect 3292 23468 3298 23480
rect 4982 23468 4988 23480
rect 5040 23468 5046 23520
rect 5813 23511 5871 23517
rect 5813 23477 5825 23511
rect 5859 23508 5871 23511
rect 5994 23508 6000 23520
rect 5859 23480 6000 23508
rect 5859 23477 5871 23480
rect 5813 23471 5871 23477
rect 5994 23468 6000 23480
rect 6052 23468 6058 23520
rect 7190 23468 7196 23520
rect 7248 23508 7254 23520
rect 8018 23508 8024 23520
rect 7248 23480 8024 23508
rect 7248 23468 7254 23480
rect 8018 23468 8024 23480
rect 8076 23468 8082 23520
rect 8202 23468 8208 23520
rect 8260 23468 8266 23520
rect 8386 23468 8392 23520
rect 8444 23508 8450 23520
rect 11609 23511 11667 23517
rect 11609 23508 11621 23511
rect 8444 23480 11621 23508
rect 8444 23468 8450 23480
rect 11609 23477 11621 23480
rect 11655 23477 11667 23511
rect 11609 23471 11667 23477
rect 11790 23468 11796 23520
rect 11848 23508 11854 23520
rect 12342 23508 12348 23520
rect 11848 23480 12348 23508
rect 11848 23468 11854 23480
rect 12342 23468 12348 23480
rect 12400 23508 12406 23520
rect 12897 23511 12955 23517
rect 12897 23508 12909 23511
rect 12400 23480 12909 23508
rect 12400 23468 12406 23480
rect 12897 23477 12909 23480
rect 12943 23477 12955 23511
rect 12897 23471 12955 23477
rect 16022 23468 16028 23520
rect 16080 23508 16086 23520
rect 17037 23511 17095 23517
rect 17037 23508 17049 23511
rect 16080 23480 17049 23508
rect 16080 23468 16086 23480
rect 17037 23477 17049 23480
rect 17083 23477 17095 23511
rect 17788 23508 17816 23607
rect 18616 23588 18644 23616
rect 18966 23604 18972 23656
rect 19024 23604 19030 23656
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23644 19119 23647
rect 19242 23644 19248 23656
rect 19107 23616 19248 23644
rect 19107 23613 19119 23616
rect 19061 23607 19119 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 19429 23647 19487 23653
rect 19429 23613 19441 23647
rect 19475 23613 19487 23647
rect 19429 23607 19487 23613
rect 18598 23536 18604 23588
rect 18656 23536 18662 23588
rect 19444 23576 19472 23607
rect 19794 23604 19800 23656
rect 19852 23644 19858 23656
rect 20165 23647 20223 23653
rect 20165 23644 20177 23647
rect 19852 23616 20177 23644
rect 19852 23604 19858 23616
rect 20165 23613 20177 23616
rect 20211 23613 20223 23647
rect 20165 23607 20223 23613
rect 21818 23604 21824 23656
rect 21876 23644 21882 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 21876 23616 22017 23644
rect 21876 23604 21882 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22186 23604 22192 23656
rect 22244 23604 22250 23656
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 24688 23644 24716 23672
rect 25332 23644 25360 23672
rect 25792 23644 25820 23675
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 28074 23672 28080 23724
rect 28132 23672 28138 23724
rect 28166 23672 28172 23724
rect 28224 23712 28230 23724
rect 28534 23712 28540 23724
rect 28224 23684 28540 23712
rect 28224 23672 28230 23684
rect 28534 23672 28540 23684
rect 28592 23712 28598 23724
rect 28629 23715 28687 23721
rect 28629 23712 28641 23715
rect 28592 23684 28641 23712
rect 28592 23672 28598 23684
rect 28629 23681 28641 23684
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23681 28779 23715
rect 28966 23712 28994 23752
rect 29086 23740 29092 23792
rect 29144 23780 29150 23792
rect 30653 23783 30711 23789
rect 30653 23780 30665 23783
rect 29144 23752 30665 23780
rect 29144 23740 29150 23752
rect 30653 23749 30665 23752
rect 30699 23780 30711 23783
rect 30837 23783 30895 23789
rect 30837 23780 30849 23783
rect 30699 23752 30849 23780
rect 30699 23749 30711 23752
rect 30653 23743 30711 23749
rect 30837 23749 30849 23752
rect 30883 23780 30895 23783
rect 31128 23780 31156 23820
rect 33318 23808 33324 23820
rect 33376 23808 33382 23860
rect 33965 23851 34023 23857
rect 33965 23817 33977 23851
rect 34011 23848 34023 23851
rect 34514 23848 34520 23860
rect 34011 23820 34520 23848
rect 34011 23817 34023 23820
rect 33965 23811 34023 23817
rect 34514 23808 34520 23820
rect 34572 23848 34578 23860
rect 35250 23848 35256 23860
rect 34572 23820 35256 23848
rect 34572 23808 34578 23820
rect 35250 23808 35256 23820
rect 35308 23808 35314 23860
rect 30883 23752 31156 23780
rect 31220 23752 31524 23780
rect 30883 23749 30895 23752
rect 30837 23743 30895 23749
rect 31220 23712 31248 23752
rect 28966 23684 31248 23712
rect 28721 23675 28779 23681
rect 24688 23616 25820 23644
rect 27798 23604 27804 23656
rect 27856 23644 27862 23656
rect 27893 23647 27951 23653
rect 27893 23644 27905 23647
rect 27856 23616 27905 23644
rect 27856 23604 27862 23616
rect 27893 23613 27905 23616
rect 27939 23613 27951 23647
rect 27893 23607 27951 23613
rect 19886 23576 19892 23588
rect 19444 23548 19892 23576
rect 19886 23536 19892 23548
rect 19944 23536 19950 23588
rect 20254 23536 20260 23588
rect 20312 23576 20318 23588
rect 25133 23579 25191 23585
rect 25133 23576 25145 23579
rect 20312 23548 25145 23576
rect 20312 23536 20318 23548
rect 25133 23545 25145 23548
rect 25179 23545 25191 23579
rect 25133 23539 25191 23545
rect 26053 23579 26111 23585
rect 26053 23545 26065 23579
rect 26099 23576 26111 23579
rect 28736 23576 28764 23675
rect 31294 23672 31300 23724
rect 31352 23672 31358 23724
rect 31390 23715 31448 23721
rect 31390 23681 31402 23715
rect 31436 23681 31448 23715
rect 31496 23712 31524 23752
rect 31570 23740 31576 23792
rect 31628 23740 31634 23792
rect 31665 23715 31723 23721
rect 31665 23712 31677 23715
rect 31496 23684 31677 23712
rect 31390 23675 31448 23681
rect 31665 23681 31677 23684
rect 31711 23681 31723 23715
rect 31665 23675 31723 23681
rect 31803 23715 31861 23721
rect 31803 23681 31815 23715
rect 31849 23712 31861 23715
rect 32306 23712 32312 23724
rect 31849 23684 32312 23712
rect 31849 23681 31861 23684
rect 31803 23675 31861 23681
rect 31405 23644 31433 23675
rect 32306 23672 32312 23684
rect 32364 23672 32370 23724
rect 33045 23715 33103 23721
rect 33045 23681 33057 23715
rect 33091 23712 33103 23715
rect 33091 23684 33732 23712
rect 33091 23681 33103 23684
rect 33045 23675 33103 23681
rect 31220 23616 31433 23644
rect 26099 23548 28764 23576
rect 26099 23545 26111 23548
rect 26053 23539 26111 23545
rect 28810 23536 28816 23588
rect 28868 23576 28874 23588
rect 29730 23576 29736 23588
rect 28868 23548 29736 23576
rect 28868 23536 28874 23548
rect 29730 23536 29736 23548
rect 29788 23576 29794 23588
rect 31220 23585 31248 23616
rect 31205 23579 31263 23585
rect 29788 23548 30512 23576
rect 29788 23536 29794 23548
rect 18414 23508 18420 23520
rect 17788 23480 18420 23508
rect 17037 23471 17095 23477
rect 18414 23468 18420 23480
rect 18472 23468 18478 23520
rect 18690 23468 18696 23520
rect 18748 23508 18754 23520
rect 18785 23511 18843 23517
rect 18785 23508 18797 23511
rect 18748 23480 18797 23508
rect 18748 23468 18754 23480
rect 18785 23477 18797 23480
rect 18831 23477 18843 23511
rect 18785 23471 18843 23477
rect 19150 23468 19156 23520
rect 19208 23508 19214 23520
rect 19334 23508 19340 23520
rect 19208 23480 19340 23508
rect 19208 23468 19214 23480
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 19521 23511 19579 23517
rect 19521 23477 19533 23511
rect 19567 23508 19579 23511
rect 19610 23508 19616 23520
rect 19567 23480 19616 23508
rect 19567 23477 19579 23480
rect 19521 23471 19579 23477
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 20073 23511 20131 23517
rect 20073 23477 20085 23511
rect 20119 23508 20131 23511
rect 20346 23508 20352 23520
rect 20119 23480 20352 23508
rect 20119 23477 20131 23480
rect 20073 23471 20131 23477
rect 20346 23468 20352 23480
rect 20404 23468 20410 23520
rect 22002 23468 22008 23520
rect 22060 23508 22066 23520
rect 22278 23508 22284 23520
rect 22060 23480 22284 23508
rect 22060 23468 22066 23480
rect 22278 23468 22284 23480
rect 22336 23508 22342 23520
rect 22833 23511 22891 23517
rect 22833 23508 22845 23511
rect 22336 23480 22845 23508
rect 22336 23468 22342 23480
rect 22833 23477 22845 23480
rect 22879 23508 22891 23511
rect 27982 23508 27988 23520
rect 22879 23480 27988 23508
rect 22879 23477 22891 23480
rect 22833 23471 22891 23477
rect 27982 23468 27988 23480
rect 28040 23468 28046 23520
rect 28442 23468 28448 23520
rect 28500 23468 28506 23520
rect 28534 23468 28540 23520
rect 28592 23508 28598 23520
rect 28905 23511 28963 23517
rect 28905 23508 28917 23511
rect 28592 23480 28917 23508
rect 28592 23468 28598 23480
rect 28905 23477 28917 23480
rect 28951 23477 28963 23511
rect 28905 23471 28963 23477
rect 30282 23468 30288 23520
rect 30340 23468 30346 23520
rect 30484 23517 30512 23548
rect 31205 23545 31217 23579
rect 31251 23576 31263 23579
rect 31386 23576 31392 23588
rect 31251 23548 31392 23576
rect 31251 23545 31263 23548
rect 31205 23539 31263 23545
rect 31386 23536 31392 23548
rect 31444 23576 31450 23588
rect 31662 23576 31668 23588
rect 31444 23548 31668 23576
rect 31444 23536 31450 23548
rect 31662 23536 31668 23548
rect 31720 23536 31726 23588
rect 32324 23576 32352 23672
rect 33594 23604 33600 23656
rect 33652 23604 33658 23656
rect 33704 23644 33732 23684
rect 33778 23672 33784 23724
rect 33836 23672 33842 23724
rect 35161 23715 35219 23721
rect 35161 23681 35173 23715
rect 35207 23712 35219 23715
rect 35342 23712 35348 23724
rect 35207 23684 35348 23712
rect 35207 23681 35219 23684
rect 35161 23675 35219 23681
rect 35342 23672 35348 23684
rect 35400 23672 35406 23724
rect 36170 23672 36176 23724
rect 36228 23672 36234 23724
rect 33870 23644 33876 23656
rect 33704 23616 33876 23644
rect 33870 23604 33876 23616
rect 33928 23644 33934 23656
rect 35253 23647 35311 23653
rect 35253 23644 35265 23647
rect 33928 23616 35265 23644
rect 33928 23604 33934 23616
rect 35253 23613 35265 23616
rect 35299 23613 35311 23647
rect 35253 23607 35311 23613
rect 33226 23576 33232 23588
rect 32324 23548 33232 23576
rect 33226 23536 33232 23548
rect 33284 23536 33290 23588
rect 33410 23536 33416 23588
rect 33468 23576 33474 23588
rect 33962 23576 33968 23588
rect 33468 23548 33968 23576
rect 33468 23536 33474 23548
rect 33962 23536 33968 23548
rect 34020 23536 34026 23588
rect 35268 23576 35296 23607
rect 35989 23579 36047 23585
rect 35989 23576 36001 23579
rect 35268 23548 36001 23576
rect 35989 23545 36001 23548
rect 36035 23545 36047 23579
rect 35989 23539 36047 23545
rect 30469 23511 30527 23517
rect 30469 23477 30481 23511
rect 30515 23477 30527 23511
rect 30469 23471 30527 23477
rect 30558 23468 30564 23520
rect 30616 23508 30622 23520
rect 31021 23511 31079 23517
rect 31021 23508 31033 23511
rect 30616 23480 31033 23508
rect 30616 23468 30622 23480
rect 31021 23477 31033 23480
rect 31067 23508 31079 23511
rect 31110 23508 31116 23520
rect 31067 23480 31116 23508
rect 31067 23477 31079 23480
rect 31021 23471 31079 23477
rect 31110 23468 31116 23480
rect 31168 23468 31174 23520
rect 31941 23511 31999 23517
rect 31941 23477 31953 23511
rect 31987 23508 31999 23511
rect 32030 23508 32036 23520
rect 31987 23480 32036 23508
rect 31987 23477 31999 23480
rect 31941 23471 31999 23477
rect 32030 23468 32036 23480
rect 32088 23508 32094 23520
rect 32582 23508 32588 23520
rect 32088 23480 32588 23508
rect 32088 23468 32094 23480
rect 32582 23468 32588 23480
rect 32640 23468 32646 23520
rect 33505 23511 33563 23517
rect 33505 23477 33517 23511
rect 33551 23508 33563 23511
rect 33870 23508 33876 23520
rect 33551 23480 33876 23508
rect 33551 23477 33563 23480
rect 33505 23471 33563 23477
rect 33870 23468 33876 23480
rect 33928 23468 33934 23520
rect 35158 23468 35164 23520
rect 35216 23468 35222 23520
rect 35342 23468 35348 23520
rect 35400 23508 35406 23520
rect 35529 23511 35587 23517
rect 35529 23508 35541 23511
rect 35400 23480 35541 23508
rect 35400 23468 35406 23480
rect 35529 23477 35541 23480
rect 35575 23477 35587 23511
rect 35529 23471 35587 23477
rect 1104 23418 36524 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 36524 23418
rect 1104 23344 36524 23366
rect 3050 23264 3056 23316
rect 3108 23304 3114 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 3108 23276 3801 23304
rect 3108 23264 3114 23276
rect 3789 23273 3801 23276
rect 3835 23273 3847 23307
rect 3789 23267 3847 23273
rect 3970 23264 3976 23316
rect 4028 23304 4034 23316
rect 9125 23307 9183 23313
rect 9125 23304 9137 23307
rect 4028 23276 9137 23304
rect 4028 23264 4034 23276
rect 9125 23273 9137 23276
rect 9171 23273 9183 23307
rect 9125 23267 9183 23273
rect 9674 23264 9680 23316
rect 9732 23264 9738 23316
rect 9766 23264 9772 23316
rect 9824 23304 9830 23316
rect 12066 23304 12072 23316
rect 9824 23276 12072 23304
rect 9824 23264 9830 23276
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 13538 23304 13544 23316
rect 12176 23276 13544 23304
rect 3145 23239 3203 23245
rect 3145 23205 3157 23239
rect 3191 23236 3203 23239
rect 3418 23236 3424 23248
rect 3191 23208 3424 23236
rect 3191 23205 3203 23208
rect 3145 23199 3203 23205
rect 3418 23196 3424 23208
rect 3476 23236 3482 23248
rect 4706 23236 4712 23248
rect 3476 23208 4712 23236
rect 3476 23196 3482 23208
rect 4706 23196 4712 23208
rect 4764 23196 4770 23248
rect 4890 23196 4896 23248
rect 4948 23236 4954 23248
rect 5350 23236 5356 23248
rect 4948 23208 5356 23236
rect 4948 23196 4954 23208
rect 5350 23196 5356 23208
rect 5408 23196 5414 23248
rect 7101 23239 7159 23245
rect 7101 23205 7113 23239
rect 7147 23205 7159 23239
rect 7101 23199 7159 23205
rect 7392 23208 7788 23236
rect 1394 23128 1400 23180
rect 1452 23128 1458 23180
rect 1670 23128 1676 23180
rect 1728 23128 1734 23180
rect 4062 23128 4068 23180
rect 4120 23168 4126 23180
rect 4341 23171 4399 23177
rect 4341 23168 4353 23171
rect 4120 23140 4353 23168
rect 4120 23128 4126 23140
rect 4341 23137 4353 23140
rect 4387 23137 4399 23171
rect 6270 23168 6276 23180
rect 4341 23131 4399 23137
rect 4632 23140 6276 23168
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23100 4215 23103
rect 4522 23100 4528 23112
rect 4203 23072 4528 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 4522 23060 4528 23072
rect 4580 23060 4586 23112
rect 4632 23109 4660 23140
rect 6270 23128 6276 23140
rect 6328 23128 6334 23180
rect 7006 23128 7012 23180
rect 7064 23168 7070 23180
rect 7116 23168 7144 23199
rect 7064 23140 7144 23168
rect 7064 23128 7070 23140
rect 4617 23103 4675 23109
rect 4617 23069 4629 23103
rect 4663 23069 4675 23103
rect 4617 23063 4675 23069
rect 4706 23060 4712 23112
rect 4764 23060 4770 23112
rect 4890 23060 4896 23112
rect 4948 23060 4954 23112
rect 5121 23103 5179 23109
rect 5121 23069 5133 23103
rect 5167 23100 5179 23103
rect 5810 23100 5816 23112
rect 5167 23072 5816 23100
rect 5167 23069 5179 23072
rect 5121 23063 5179 23069
rect 5810 23060 5816 23072
rect 5868 23100 5874 23112
rect 5868 23072 6040 23100
rect 5868 23060 5874 23072
rect 3142 23032 3148 23044
rect 2898 23004 3148 23032
rect 3142 22992 3148 23004
rect 3200 22992 3206 23044
rect 3418 22992 3424 23044
rect 3476 23032 3482 23044
rect 3970 23032 3976 23044
rect 3476 23004 3976 23032
rect 3476 22992 3482 23004
rect 3970 22992 3976 23004
rect 4028 23032 4034 23044
rect 4249 23035 4307 23041
rect 4249 23032 4261 23035
rect 4028 23004 4261 23032
rect 4028 22992 4034 23004
rect 4249 23001 4261 23004
rect 4295 23001 4307 23035
rect 4249 22995 4307 23001
rect 4982 22992 4988 23044
rect 5040 22992 5046 23044
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 5261 22967 5319 22973
rect 5261 22964 5273 22967
rect 4672 22936 5273 22964
rect 4672 22924 4678 22936
rect 5261 22933 5273 22936
rect 5307 22933 5319 22967
rect 6012 22964 6040 23072
rect 6454 23060 6460 23112
rect 6512 23100 6518 23112
rect 7392 23100 7420 23208
rect 7558 23128 7564 23180
rect 7616 23168 7622 23180
rect 7653 23171 7711 23177
rect 7653 23168 7665 23171
rect 7616 23140 7665 23168
rect 7616 23128 7622 23140
rect 7653 23137 7665 23140
rect 7699 23137 7711 23171
rect 7760 23168 7788 23208
rect 8018 23196 8024 23248
rect 8076 23196 8082 23248
rect 8846 23168 8852 23180
rect 7760 23140 8852 23168
rect 7653 23131 7711 23137
rect 8846 23128 8852 23140
rect 8904 23128 8910 23180
rect 9048 23140 9536 23168
rect 6512 23072 7420 23100
rect 7469 23103 7527 23109
rect 6512 23060 6518 23072
rect 7469 23069 7481 23103
rect 7515 23100 7527 23103
rect 8202 23100 8208 23112
rect 7515 23072 8208 23100
rect 7515 23069 7527 23072
rect 7469 23063 7527 23069
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 9048 23109 9076 23140
rect 9033 23103 9091 23109
rect 9033 23069 9045 23103
rect 9079 23069 9091 23103
rect 9033 23063 9091 23069
rect 9398 23060 9404 23112
rect 9456 23060 9462 23112
rect 7561 23035 7619 23041
rect 7561 23001 7573 23035
rect 7607 23032 7619 23035
rect 8297 23035 8355 23041
rect 7607 23004 8248 23032
rect 7607 23001 7619 23004
rect 7561 22995 7619 23001
rect 8018 22964 8024 22976
rect 6012 22936 8024 22964
rect 5261 22927 5319 22933
rect 8018 22924 8024 22936
rect 8076 22924 8082 22976
rect 8220 22964 8248 23004
rect 8297 23001 8309 23035
rect 8343 23032 8355 23035
rect 9306 23032 9312 23044
rect 8343 23004 9312 23032
rect 8343 23001 8355 23004
rect 8297 22995 8355 23001
rect 9306 22992 9312 23004
rect 9364 22992 9370 23044
rect 9508 23032 9536 23140
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 9784 23100 9812 23264
rect 10134 23196 10140 23248
rect 10192 23196 10198 23248
rect 11974 23196 11980 23248
rect 12032 23236 12038 23248
rect 12176 23236 12204 23276
rect 13538 23264 13544 23276
rect 13596 23304 13602 23316
rect 13725 23307 13783 23313
rect 13725 23304 13737 23307
rect 13596 23276 13737 23304
rect 13596 23264 13602 23276
rect 13725 23273 13737 23276
rect 13771 23273 13783 23307
rect 13725 23267 13783 23273
rect 14737 23307 14795 23313
rect 14737 23273 14749 23307
rect 14783 23304 14795 23307
rect 15470 23304 15476 23316
rect 14783 23276 15476 23304
rect 14783 23273 14795 23276
rect 14737 23267 14795 23273
rect 15470 23264 15476 23276
rect 15528 23264 15534 23316
rect 15654 23264 15660 23316
rect 15712 23304 15718 23316
rect 17313 23307 17371 23313
rect 15712 23276 17172 23304
rect 15712 23264 15718 23276
rect 12526 23236 12532 23248
rect 12032 23208 12204 23236
rect 12268 23208 12532 23236
rect 12032 23196 12038 23208
rect 10042 23128 10048 23180
rect 10100 23128 10106 23180
rect 10152 23168 10180 23196
rect 10597 23176 10655 23177
rect 10520 23171 10655 23176
rect 10520 23168 10609 23171
rect 10152 23140 10364 23168
rect 9631 23072 9812 23100
rect 9861 23103 9919 23109
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 9861 23069 9873 23103
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 9876 23032 9904 23063
rect 10134 23060 10140 23112
rect 10192 23060 10198 23112
rect 10226 23060 10232 23112
rect 10284 23060 10290 23112
rect 10042 23032 10048 23044
rect 9508 23004 10048 23032
rect 10042 22992 10048 23004
rect 10100 22992 10106 23044
rect 10336 23032 10364 23140
rect 10428 23148 10609 23168
rect 10428 23140 10548 23148
rect 10428 23109 10456 23140
rect 10597 23137 10609 23148
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 11790 23168 11796 23180
rect 11664 23140 11796 23168
rect 11664 23128 11670 23140
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23069 10471 23103
rect 10413 23063 10471 23069
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23069 10563 23103
rect 10505 23063 10563 23069
rect 10689 23103 10747 23109
rect 10689 23069 10701 23103
rect 10735 23102 10747 23103
rect 10778 23102 10784 23112
rect 10735 23074 10784 23102
rect 10735 23069 10747 23074
rect 10689 23063 10747 23069
rect 10520 23032 10548 23063
rect 10778 23060 10784 23074
rect 10836 23060 10842 23112
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 11333 23103 11391 23109
rect 11333 23100 11345 23103
rect 11296 23072 11345 23100
rect 11296 23060 11302 23072
rect 11333 23069 11345 23072
rect 11379 23069 11391 23103
rect 11333 23063 11391 23069
rect 11422 23060 11428 23112
rect 11480 23100 11486 23112
rect 12268 23109 12296 23208
rect 12526 23196 12532 23208
rect 12584 23236 12590 23248
rect 12897 23239 12955 23245
rect 12897 23236 12909 23239
rect 12584 23208 12909 23236
rect 12584 23196 12590 23208
rect 12897 23205 12909 23208
rect 12943 23205 12955 23239
rect 15102 23236 15108 23248
rect 12897 23199 12955 23205
rect 14108 23208 15108 23236
rect 12802 23168 12808 23180
rect 12452 23140 12808 23168
rect 12452 23109 12480 23140
rect 12802 23128 12808 23140
rect 12860 23128 12866 23180
rect 12912 23168 12940 23199
rect 13354 23168 13360 23180
rect 12912 23140 13360 23168
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 11480 23072 11529 23100
rect 11480 23060 11486 23072
rect 11517 23069 11529 23072
rect 11563 23100 11575 23103
rect 12253 23103 12311 23109
rect 11563 23072 12112 23100
rect 11563 23069 11575 23072
rect 11517 23063 11575 23069
rect 10336 23004 10548 23032
rect 11701 23035 11759 23041
rect 11701 23001 11713 23035
rect 11747 23032 11759 23035
rect 12084 23032 12112 23072
rect 12253 23069 12265 23103
rect 12299 23069 12311 23103
rect 12253 23063 12311 23069
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 12713 23103 12771 23109
rect 12713 23069 12725 23103
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 12728 23032 12756 23063
rect 12986 23060 12992 23112
rect 13044 23060 13050 23112
rect 13188 23109 13216 23140
rect 13354 23128 13360 23140
rect 13412 23128 13418 23180
rect 13173 23103 13231 23109
rect 13173 23069 13185 23103
rect 13219 23069 13231 23103
rect 13173 23063 13231 23069
rect 13906 23060 13912 23112
rect 13964 23060 13970 23112
rect 14108 23109 14136 23208
rect 15102 23196 15108 23208
rect 15160 23236 15166 23248
rect 15930 23236 15936 23248
rect 15160 23208 15936 23236
rect 15160 23196 15166 23208
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 16390 23196 16396 23248
rect 16448 23236 16454 23248
rect 16448 23208 16804 23236
rect 16448 23196 16454 23208
rect 14645 23171 14703 23177
rect 14645 23137 14657 23171
rect 14691 23168 14703 23171
rect 15194 23168 15200 23180
rect 14691 23140 15200 23168
rect 14691 23137 14703 23140
rect 14645 23131 14703 23137
rect 15194 23128 15200 23140
rect 15252 23128 15258 23180
rect 16408 23140 16712 23168
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23100 14335 23103
rect 14366 23100 14372 23112
rect 14323 23072 14372 23100
rect 14323 23069 14335 23072
rect 14277 23063 14335 23069
rect 14366 23060 14372 23072
rect 14424 23060 14430 23112
rect 14737 23103 14795 23109
rect 14737 23069 14749 23103
rect 14783 23100 14795 23103
rect 15654 23100 15660 23112
rect 14783 23072 15660 23100
rect 14783 23069 14795 23072
rect 14737 23063 14795 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 15746 23060 15752 23112
rect 15804 23060 15810 23112
rect 16025 23103 16083 23109
rect 16025 23069 16037 23103
rect 16071 23069 16083 23103
rect 16025 23063 16083 23069
rect 11747 23004 11836 23032
rect 12084 23004 12480 23032
rect 12728 23004 14412 23032
rect 11747 23001 11759 23004
rect 11701 22995 11759 23001
rect 8386 22964 8392 22976
rect 8220 22936 8392 22964
rect 8386 22924 8392 22936
rect 8444 22964 8450 22976
rect 8662 22964 8668 22976
rect 8444 22936 8668 22964
rect 8444 22924 8450 22936
rect 8662 22924 8668 22936
rect 8720 22924 8726 22976
rect 10226 22924 10232 22976
rect 10284 22964 10290 22976
rect 11606 22964 11612 22976
rect 10284 22936 11612 22964
rect 10284 22924 10290 22936
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 11808 22964 11836 23004
rect 12452 22976 12480 23004
rect 11882 22964 11888 22976
rect 11808 22936 11888 22964
rect 11882 22924 11888 22936
rect 11940 22964 11946 22976
rect 12253 22967 12311 22973
rect 12253 22964 12265 22967
rect 11940 22936 12265 22964
rect 11940 22924 11946 22936
rect 12253 22933 12265 22936
rect 12299 22933 12311 22967
rect 12253 22927 12311 22933
rect 12434 22924 12440 22976
rect 12492 22924 12498 22976
rect 12986 22924 12992 22976
rect 13044 22924 13050 22976
rect 14185 22967 14243 22973
rect 14185 22933 14197 22967
rect 14231 22964 14243 22967
rect 14274 22964 14280 22976
rect 14231 22936 14280 22964
rect 14231 22933 14243 22936
rect 14185 22927 14243 22933
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14384 22964 14412 23004
rect 14458 22992 14464 23044
rect 14516 22992 14522 23044
rect 15105 23035 15163 23041
rect 15105 23001 15117 23035
rect 15151 23032 15163 23035
rect 15378 23032 15384 23044
rect 15151 23004 15384 23032
rect 15151 23001 15163 23004
rect 15105 22995 15163 23001
rect 15378 22992 15384 23004
rect 15436 22992 15442 23044
rect 15838 22992 15844 23044
rect 15896 23032 15902 23044
rect 16040 23032 16068 23063
rect 16114 23060 16120 23112
rect 16172 23100 16178 23112
rect 16408 23109 16436 23140
rect 16684 23109 16712 23140
rect 16776 23109 16804 23208
rect 17144 23177 17172 23276
rect 17313 23273 17325 23307
rect 17359 23304 17371 23307
rect 17862 23304 17868 23316
rect 17359 23276 17868 23304
rect 17359 23273 17371 23276
rect 17313 23267 17371 23273
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 18966 23264 18972 23316
rect 19024 23304 19030 23316
rect 19024 23276 22784 23304
rect 19024 23264 19030 23276
rect 18598 23196 18604 23248
rect 18656 23236 18662 23248
rect 18656 23208 20760 23236
rect 18656 23196 18662 23208
rect 17129 23171 17187 23177
rect 17129 23137 17141 23171
rect 17175 23137 17187 23171
rect 18138 23168 18144 23180
rect 17129 23131 17187 23137
rect 17512 23140 18144 23168
rect 16393 23103 16451 23109
rect 16393 23100 16405 23103
rect 16172 23072 16405 23100
rect 16172 23060 16178 23072
rect 16393 23069 16405 23072
rect 16439 23069 16451 23103
rect 16393 23063 16451 23069
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23069 16543 23103
rect 16485 23063 16543 23069
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 16669 23063 16727 23069
rect 16761 23103 16819 23109
rect 16761 23069 16773 23103
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 16298 23032 16304 23044
rect 15896 23004 16304 23032
rect 15896 22992 15902 23004
rect 16298 22992 16304 23004
rect 16356 22992 16362 23044
rect 14918 22964 14924 22976
rect 14384 22936 14924 22964
rect 14918 22924 14924 22936
rect 14976 22924 14982 22976
rect 15010 22924 15016 22976
rect 15068 22964 15074 22976
rect 16500 22964 16528 23063
rect 16684 23032 16712 23063
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17512 23109 17540 23140
rect 18138 23128 18144 23140
rect 18196 23128 18202 23180
rect 19242 23128 19248 23180
rect 19300 23128 19306 23180
rect 19886 23168 19892 23180
rect 19352 23140 19892 23168
rect 17497 23103 17555 23109
rect 16908 23072 16953 23100
rect 16908 23060 16914 23072
rect 17497 23069 17509 23103
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23069 17647 23103
rect 17589 23063 17647 23069
rect 17604 23032 17632 23063
rect 17678 23060 17684 23112
rect 17736 23060 17742 23112
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23100 18935 23103
rect 18966 23100 18972 23112
rect 18923 23072 18972 23100
rect 18923 23069 18935 23072
rect 18877 23063 18935 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19061 23103 19119 23109
rect 19061 23069 19073 23103
rect 19107 23100 19119 23103
rect 19352 23100 19380 23140
rect 19107 23072 19380 23100
rect 19107 23069 19119 23072
rect 19061 23063 19119 23069
rect 19426 23060 19432 23112
rect 19484 23060 19490 23112
rect 19518 23060 19524 23112
rect 19576 23060 19582 23112
rect 19628 23109 19656 23140
rect 19886 23128 19892 23140
rect 19944 23128 19950 23180
rect 20530 23128 20536 23180
rect 20588 23128 20594 23180
rect 19613 23103 19671 23109
rect 19613 23069 19625 23103
rect 19659 23069 19671 23103
rect 19613 23063 19671 23069
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23100 19855 23103
rect 20070 23100 20076 23112
rect 19843 23072 20076 23100
rect 19843 23069 19855 23072
rect 19797 23063 19855 23069
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 20346 23060 20352 23112
rect 20404 23100 20410 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20404 23072 20453 23100
rect 20404 23060 20410 23072
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 17770 23032 17776 23044
rect 16684 23004 16988 23032
rect 17604 23004 17776 23032
rect 16758 22964 16764 22976
rect 15068 22936 16764 22964
rect 15068 22924 15074 22936
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 16960 22964 16988 23004
rect 17770 22992 17776 23004
rect 17828 22992 17834 23044
rect 19150 23032 19156 23044
rect 17880 23004 19156 23032
rect 17880 22964 17908 23004
rect 19150 22992 19156 23004
rect 19208 22992 19214 23044
rect 20088 23032 20116 23060
rect 20640 23032 20668 23063
rect 20088 23004 20668 23032
rect 20732 23032 20760 23208
rect 21174 23196 21180 23248
rect 21232 23245 21238 23248
rect 21232 23239 21281 23245
rect 21232 23205 21235 23239
rect 21269 23205 21281 23239
rect 21910 23236 21916 23248
rect 21232 23199 21281 23205
rect 21376 23208 21916 23236
rect 21232 23196 21238 23199
rect 20898 23060 20904 23112
rect 20956 23060 20962 23112
rect 21085 23103 21143 23109
rect 21085 23069 21097 23103
rect 21131 23100 21143 23103
rect 21266 23100 21272 23112
rect 21131 23072 21272 23100
rect 21131 23069 21143 23072
rect 21085 23063 21143 23069
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 21376 23109 21404 23208
rect 21910 23196 21916 23208
rect 21968 23196 21974 23248
rect 22002 23196 22008 23248
rect 22060 23236 22066 23248
rect 22060 23208 22232 23236
rect 22060 23196 22066 23208
rect 21634 23128 21640 23180
rect 21692 23128 21698 23180
rect 22204 23177 22232 23208
rect 22462 23196 22468 23248
rect 22520 23236 22526 23248
rect 22756 23236 22784 23276
rect 22830 23264 22836 23316
rect 22888 23264 22894 23316
rect 23382 23264 23388 23316
rect 23440 23304 23446 23316
rect 24857 23307 24915 23313
rect 24857 23304 24869 23307
rect 23440 23276 24869 23304
rect 23440 23264 23446 23276
rect 24857 23273 24869 23276
rect 24903 23273 24915 23307
rect 24857 23267 24915 23273
rect 26142 23264 26148 23316
rect 26200 23264 26206 23316
rect 26326 23264 26332 23316
rect 26384 23304 26390 23316
rect 26605 23307 26663 23313
rect 26605 23304 26617 23307
rect 26384 23276 26617 23304
rect 26384 23264 26390 23276
rect 26605 23273 26617 23276
rect 26651 23273 26663 23307
rect 26605 23267 26663 23273
rect 27065 23307 27123 23313
rect 27065 23273 27077 23307
rect 27111 23304 27123 23307
rect 27157 23307 27215 23313
rect 27157 23304 27169 23307
rect 27111 23276 27169 23304
rect 27111 23273 27123 23276
rect 27065 23267 27123 23273
rect 27157 23273 27169 23276
rect 27203 23273 27215 23307
rect 27157 23267 27215 23273
rect 27338 23264 27344 23316
rect 27396 23264 27402 23316
rect 28169 23307 28227 23313
rect 28169 23273 28181 23307
rect 28215 23273 28227 23307
rect 28169 23267 28227 23273
rect 23109 23239 23167 23245
rect 22520 23208 22717 23236
rect 22756 23208 22876 23236
rect 22520 23196 22526 23208
rect 22189 23171 22247 23177
rect 22189 23137 22201 23171
rect 22235 23137 22247 23171
rect 22189 23131 22247 23137
rect 22370 23128 22376 23180
rect 22428 23168 22434 23180
rect 22689 23177 22717 23208
rect 22557 23171 22615 23177
rect 22557 23168 22569 23171
rect 22428 23140 22569 23168
rect 22428 23128 22434 23140
rect 22557 23137 22569 23140
rect 22603 23137 22615 23171
rect 22557 23131 22615 23137
rect 22674 23171 22732 23177
rect 22674 23137 22686 23171
rect 22720 23137 22732 23171
rect 22848 23168 22876 23208
rect 23109 23205 23121 23239
rect 23155 23236 23167 23239
rect 23474 23236 23480 23248
rect 23155 23208 23480 23236
rect 23155 23205 23167 23208
rect 23109 23199 23167 23205
rect 23474 23196 23480 23208
rect 23532 23196 23538 23248
rect 25130 23196 25136 23248
rect 25188 23236 25194 23248
rect 25590 23236 25596 23248
rect 25188 23208 25596 23236
rect 25188 23196 25194 23208
rect 25590 23196 25596 23208
rect 25648 23196 25654 23248
rect 26160 23236 26188 23264
rect 25976 23208 26188 23236
rect 25976 23177 26004 23208
rect 25961 23171 26019 23177
rect 22848 23140 25820 23168
rect 22674 23131 22732 23137
rect 21361 23103 21419 23109
rect 21361 23069 21373 23103
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23069 21787 23103
rect 21729 23063 21787 23069
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22097 23103 22155 23109
rect 22097 23069 22109 23103
rect 22143 23100 22155 23103
rect 22143 23072 22227 23100
rect 22143 23069 22155 23072
rect 22097 23063 22155 23069
rect 21744 23032 21772 23063
rect 20732 23004 21772 23032
rect 21836 23032 21864 23063
rect 22199 23032 22227 23072
rect 22278 23060 22284 23112
rect 22336 23100 22342 23112
rect 23268 23103 23326 23109
rect 23268 23100 23280 23103
rect 22336 23072 23280 23100
rect 22336 23060 22342 23072
rect 23268 23069 23280 23072
rect 23314 23069 23326 23103
rect 23268 23063 23326 23069
rect 23750 23060 23756 23112
rect 23808 23060 23814 23112
rect 25038 23060 25044 23112
rect 25096 23060 25102 23112
rect 25314 23060 25320 23112
rect 25372 23100 25378 23112
rect 25682 23100 25688 23112
rect 25372 23072 25688 23100
rect 25372 23060 25378 23072
rect 25682 23060 25688 23072
rect 25740 23060 25746 23112
rect 25792 23100 25820 23140
rect 25961 23137 25973 23171
rect 26007 23137 26019 23171
rect 28184 23168 28212 23267
rect 28534 23264 28540 23316
rect 28592 23304 28598 23316
rect 28629 23307 28687 23313
rect 28629 23304 28641 23307
rect 28592 23276 28641 23304
rect 28592 23264 28598 23276
rect 28629 23273 28641 23276
rect 28675 23304 28687 23307
rect 29086 23304 29092 23316
rect 28675 23276 29092 23304
rect 28675 23273 28687 23276
rect 28629 23267 28687 23273
rect 29086 23264 29092 23276
rect 29144 23304 29150 23316
rect 29144 23276 29684 23304
rect 29144 23264 29150 23276
rect 28350 23196 28356 23248
rect 28408 23196 28414 23248
rect 29656 23245 29684 23276
rect 30006 23264 30012 23316
rect 30064 23304 30070 23316
rect 31570 23304 31576 23316
rect 30064 23276 31576 23304
rect 30064 23264 30070 23276
rect 31570 23264 31576 23276
rect 31628 23264 31634 23316
rect 33226 23264 33232 23316
rect 33284 23304 33290 23316
rect 34790 23304 34796 23316
rect 33284 23276 34796 23304
rect 33284 23264 33290 23276
rect 34790 23264 34796 23276
rect 34848 23264 34854 23316
rect 29641 23239 29699 23245
rect 29641 23205 29653 23239
rect 29687 23205 29699 23239
rect 29641 23199 29699 23205
rect 30374 23196 30380 23248
rect 30432 23236 30438 23248
rect 31110 23236 31116 23248
rect 30432 23208 31116 23236
rect 30432 23196 30438 23208
rect 31110 23196 31116 23208
rect 31168 23196 31174 23248
rect 32030 23236 32036 23248
rect 31405 23208 32036 23236
rect 28810 23168 28816 23180
rect 28184 23140 28816 23168
rect 25961 23131 26019 23137
rect 28810 23128 28816 23140
rect 28868 23168 28874 23180
rect 28868 23140 29868 23168
rect 28868 23128 28874 23140
rect 25792 23072 26004 23100
rect 22370 23032 22376 23044
rect 21836 23004 22140 23032
rect 22199 23004 22376 23032
rect 16960 22936 17908 22964
rect 18046 22924 18052 22976
rect 18104 22964 18110 22976
rect 18877 22967 18935 22973
rect 18877 22964 18889 22967
rect 18104 22936 18889 22964
rect 18104 22924 18110 22936
rect 18877 22933 18889 22936
rect 18923 22933 18935 22967
rect 18877 22927 18935 22933
rect 19242 22924 19248 22976
rect 19300 22924 19306 22976
rect 19702 22924 19708 22976
rect 19760 22924 19766 22976
rect 19794 22924 19800 22976
rect 19852 22964 19858 22976
rect 20901 22967 20959 22973
rect 20901 22964 20913 22967
rect 19852 22936 20913 22964
rect 19852 22924 19858 22936
rect 20901 22933 20913 22936
rect 20947 22933 20959 22967
rect 20901 22927 20959 22933
rect 20990 22924 20996 22976
rect 21048 22964 21054 22976
rect 21358 22964 21364 22976
rect 21048 22936 21364 22964
rect 21048 22924 21054 22936
rect 21358 22924 21364 22936
rect 21416 22964 21422 22976
rect 22005 22967 22063 22973
rect 22005 22964 22017 22967
rect 21416 22936 22017 22964
rect 21416 22924 21422 22936
rect 22005 22933 22017 22936
rect 22051 22933 22063 22967
rect 22112 22964 22140 23004
rect 22370 22992 22376 23004
rect 22428 22992 22434 23044
rect 22465 23035 22523 23041
rect 22465 23001 22477 23035
rect 22511 23032 22523 23035
rect 22830 23032 22836 23044
rect 22511 23004 22836 23032
rect 22511 23001 22523 23004
rect 22465 22995 22523 23001
rect 22830 22992 22836 23004
rect 22888 23032 22894 23044
rect 23566 23032 23572 23044
rect 22888 23004 23572 23032
rect 22888 22992 22894 23004
rect 23566 22992 23572 23004
rect 23624 23032 23630 23044
rect 25130 23032 25136 23044
rect 23624 23004 25136 23032
rect 23624 22992 23630 23004
rect 25130 22992 25136 23004
rect 25188 22992 25194 23044
rect 25225 23035 25283 23041
rect 25225 23001 25237 23035
rect 25271 23032 25283 23035
rect 25498 23032 25504 23044
rect 25271 23004 25504 23032
rect 25271 23001 25283 23004
rect 25225 22995 25283 23001
rect 25498 22992 25504 23004
rect 25556 22992 25562 23044
rect 25976 23041 26004 23072
rect 26142 23060 26148 23112
rect 26200 23060 26206 23112
rect 26237 23103 26295 23109
rect 26237 23069 26249 23103
rect 26283 23100 26295 23103
rect 26418 23100 26424 23112
rect 26283 23072 26424 23100
rect 26283 23069 26295 23072
rect 26237 23063 26295 23069
rect 26418 23060 26424 23072
rect 26476 23100 26482 23112
rect 26694 23100 26700 23112
rect 26476 23072 26700 23100
rect 26476 23060 26482 23072
rect 26694 23060 26700 23072
rect 26752 23060 26758 23112
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 26881 23103 26939 23109
rect 26881 23069 26893 23103
rect 26927 23100 26939 23103
rect 26970 23100 26976 23112
rect 26927 23072 26976 23100
rect 26927 23069 26939 23072
rect 26881 23063 26939 23069
rect 25961 23035 26019 23041
rect 25961 23001 25973 23035
rect 26007 23001 26019 23035
rect 25961 22995 26019 23001
rect 22738 22964 22744 22976
rect 22112 22936 22744 22964
rect 22005 22927 22063 22933
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 23382 22924 23388 22976
rect 23440 22924 23446 22976
rect 23474 22924 23480 22976
rect 23532 22924 23538 22976
rect 25314 22924 25320 22976
rect 25372 22964 25378 22976
rect 26804 22964 26832 23063
rect 26970 23060 26976 23072
rect 27028 23060 27034 23112
rect 28442 23060 28448 23112
rect 28500 23060 28506 23112
rect 29840 23109 29868 23140
rect 30484 23140 30972 23168
rect 29825 23103 29883 23109
rect 29825 23069 29837 23103
rect 29871 23069 29883 23103
rect 29825 23063 29883 23069
rect 30009 23103 30067 23109
rect 30009 23069 30021 23103
rect 30055 23100 30067 23103
rect 30190 23100 30196 23112
rect 30055 23072 30196 23100
rect 30055 23069 30067 23072
rect 30009 23063 30067 23069
rect 27065 23035 27123 23041
rect 27065 23001 27077 23035
rect 27111 23001 27123 23035
rect 27065 22995 27123 23001
rect 25372 22936 26832 22964
rect 25372 22924 25378 22936
rect 26878 22924 26884 22976
rect 26936 22964 26942 22976
rect 27080 22964 27108 22995
rect 27154 22992 27160 23044
rect 27212 23032 27218 23044
rect 27522 23032 27528 23044
rect 27212 23004 27528 23032
rect 27212 22992 27218 23004
rect 27522 22992 27528 23004
rect 27580 22992 27586 23044
rect 27985 23035 28043 23041
rect 27985 23001 27997 23035
rect 28031 23032 28043 23035
rect 28534 23032 28540 23044
rect 28031 23004 28540 23032
rect 28031 23001 28043 23004
rect 27985 22995 28043 23001
rect 28534 22992 28540 23004
rect 28592 22992 28598 23044
rect 29178 22992 29184 23044
rect 29236 23032 29242 23044
rect 30024 23032 30052 23063
rect 30190 23060 30196 23072
rect 30248 23060 30254 23112
rect 30282 23060 30288 23112
rect 30340 23060 30346 23112
rect 30374 23060 30380 23112
rect 30432 23060 30438 23112
rect 30484 23032 30512 23140
rect 30558 23060 30564 23112
rect 30616 23060 30622 23112
rect 30653 23103 30711 23109
rect 30653 23069 30665 23103
rect 30699 23100 30711 23103
rect 30834 23100 30840 23112
rect 30699 23072 30840 23100
rect 30699 23069 30711 23072
rect 30653 23063 30711 23069
rect 30834 23060 30840 23072
rect 30892 23060 30898 23112
rect 30944 23100 30972 23140
rect 30944 23072 31156 23100
rect 31021 23035 31079 23041
rect 31021 23032 31033 23035
rect 29236 23004 30052 23032
rect 30116 23004 30512 23032
rect 30668 23004 31033 23032
rect 29236 22992 29242 23004
rect 26936 22936 27108 22964
rect 27325 22967 27383 22973
rect 26936 22924 26942 22936
rect 27325 22933 27337 22967
rect 27371 22964 27383 22967
rect 27890 22964 27896 22976
rect 27371 22936 27896 22964
rect 27371 22933 27383 22936
rect 27325 22927 27383 22933
rect 27890 22924 27896 22936
rect 27948 22924 27954 22976
rect 28195 22967 28253 22973
rect 28195 22933 28207 22967
rect 28241 22964 28253 22967
rect 29086 22964 29092 22976
rect 28241 22936 29092 22964
rect 28241 22933 28253 22936
rect 28195 22927 28253 22933
rect 29086 22924 29092 22936
rect 29144 22964 29150 22976
rect 29546 22964 29552 22976
rect 29144 22936 29552 22964
rect 29144 22924 29150 22936
rect 29546 22924 29552 22936
rect 29604 22924 29610 22976
rect 29822 22924 29828 22976
rect 29880 22964 29886 22976
rect 29917 22967 29975 22973
rect 29917 22964 29929 22967
rect 29880 22936 29929 22964
rect 29880 22924 29886 22936
rect 29917 22933 29929 22936
rect 29963 22933 29975 22967
rect 29917 22927 29975 22933
rect 30006 22924 30012 22976
rect 30064 22964 30070 22976
rect 30116 22964 30144 23004
rect 30668 22976 30696 23004
rect 31021 23001 31033 23004
rect 31067 23001 31079 23035
rect 31128 23032 31156 23072
rect 31202 23060 31208 23112
rect 31260 23060 31266 23112
rect 31405 23109 31433 23208
rect 32030 23196 32036 23208
rect 32088 23196 32094 23248
rect 31662 23128 31668 23180
rect 31720 23128 31726 23180
rect 31389 23103 31447 23109
rect 31389 23069 31401 23103
rect 31435 23069 31447 23103
rect 31389 23063 31447 23069
rect 31478 23060 31484 23112
rect 31536 23109 31542 23112
rect 31536 23103 31565 23109
rect 31553 23069 31565 23103
rect 31536 23063 31565 23069
rect 31536 23060 31542 23063
rect 31754 23060 31760 23112
rect 31812 23060 31818 23112
rect 32306 23060 32312 23112
rect 32364 23060 32370 23112
rect 35250 23060 35256 23112
rect 35308 23060 35314 23112
rect 31297 23035 31355 23041
rect 31297 23032 31309 23035
rect 31128 23004 31309 23032
rect 31021 22995 31079 23001
rect 31297 23001 31309 23004
rect 31343 23032 31355 23035
rect 31343 23004 32168 23032
rect 31343 23001 31355 23004
rect 31297 22995 31355 23001
rect 30064 22936 30144 22964
rect 30064 22924 30070 22936
rect 30190 22924 30196 22976
rect 30248 22924 30254 22976
rect 30650 22924 30656 22976
rect 30708 22924 30714 22976
rect 30837 22967 30895 22973
rect 30837 22933 30849 22967
rect 30883 22964 30895 22967
rect 30926 22964 30932 22976
rect 30883 22936 30932 22964
rect 30883 22933 30895 22936
rect 30837 22927 30895 22933
rect 30926 22924 30932 22936
rect 30984 22924 30990 22976
rect 31202 22924 31208 22976
rect 31260 22964 31266 22976
rect 32140 22973 32168 23004
rect 32490 22992 32496 23044
rect 32548 23032 32554 23044
rect 33042 23032 33048 23044
rect 32548 23004 33048 23032
rect 32548 22992 32554 23004
rect 33042 22992 33048 23004
rect 33100 22992 33106 23044
rect 35066 22992 35072 23044
rect 35124 22992 35130 23044
rect 31941 22967 31999 22973
rect 31941 22964 31953 22967
rect 31260 22936 31953 22964
rect 31260 22924 31266 22936
rect 31941 22933 31953 22936
rect 31987 22933 31999 22967
rect 31941 22927 31999 22933
rect 32125 22967 32183 22973
rect 32125 22933 32137 22967
rect 32171 22933 32183 22967
rect 32125 22927 32183 22933
rect 32950 22924 32956 22976
rect 33008 22964 33014 22976
rect 34422 22964 34428 22976
rect 33008 22936 34428 22964
rect 33008 22924 33014 22936
rect 34422 22924 34428 22936
rect 34480 22924 34486 22976
rect 34790 22924 34796 22976
rect 34848 22964 34854 22976
rect 35437 22967 35495 22973
rect 35437 22964 35449 22967
rect 34848 22936 35449 22964
rect 34848 22924 34854 22936
rect 35437 22933 35449 22936
rect 35483 22933 35495 22967
rect 35437 22927 35495 22933
rect 1104 22874 36524 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 36524 22874
rect 1104 22800 36524 22822
rect 2961 22763 3019 22769
rect 2961 22729 2973 22763
rect 3007 22760 3019 22763
rect 3234 22760 3240 22772
rect 3007 22732 3240 22760
rect 3007 22729 3019 22732
rect 2961 22723 3019 22729
rect 3234 22720 3240 22732
rect 3292 22760 3298 22772
rect 3602 22760 3608 22772
rect 3292 22732 3608 22760
rect 3292 22720 3298 22732
rect 3602 22720 3608 22732
rect 3660 22720 3666 22772
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 7558 22760 7564 22772
rect 7340 22732 7564 22760
rect 7340 22720 7346 22732
rect 7558 22720 7564 22732
rect 7616 22720 7622 22772
rect 8110 22760 8116 22772
rect 7668 22732 8116 22760
rect 7668 22704 7696 22732
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 8938 22760 8944 22772
rect 8352 22732 8944 22760
rect 8352 22720 8358 22732
rect 8938 22720 8944 22732
rect 8996 22720 9002 22772
rect 9398 22720 9404 22772
rect 9456 22760 9462 22772
rect 9953 22763 10011 22769
rect 9953 22760 9965 22763
rect 9456 22732 9965 22760
rect 9456 22720 9462 22732
rect 9953 22729 9965 22732
rect 9999 22729 10011 22763
rect 9953 22723 10011 22729
rect 10045 22763 10103 22769
rect 10045 22729 10057 22763
rect 10091 22760 10103 22763
rect 10594 22760 10600 22772
rect 10091 22732 10600 22760
rect 10091 22729 10103 22732
rect 10045 22723 10103 22729
rect 10594 22720 10600 22732
rect 10652 22720 10658 22772
rect 12250 22760 12256 22772
rect 10704 22732 12256 22760
rect 5534 22692 5540 22704
rect 4540 22664 4844 22692
rect 2869 22627 2927 22633
rect 2869 22593 2881 22627
rect 2915 22624 2927 22627
rect 3329 22627 3387 22633
rect 3329 22624 3341 22627
rect 2915 22596 3341 22624
rect 2915 22593 2927 22596
rect 2869 22587 2927 22593
rect 3329 22593 3341 22596
rect 3375 22593 3387 22627
rect 3329 22587 3387 22593
rect 3878 22584 3884 22636
rect 3936 22624 3942 22636
rect 4341 22627 4399 22633
rect 4341 22624 4353 22627
rect 3936 22596 4353 22624
rect 3936 22584 3942 22596
rect 4341 22593 4353 22596
rect 4387 22593 4399 22627
rect 4341 22587 4399 22593
rect 4430 22584 4436 22636
rect 4488 22584 4494 22636
rect 2590 22516 2596 22568
rect 2648 22556 2654 22568
rect 3145 22559 3203 22565
rect 3145 22556 3157 22559
rect 2648 22528 3157 22556
rect 2648 22516 2654 22528
rect 3145 22525 3157 22528
rect 3191 22525 3203 22559
rect 3145 22519 3203 22525
rect 3160 22488 3188 22519
rect 3970 22516 3976 22568
rect 4028 22516 4034 22568
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 4540 22556 4568 22664
rect 4617 22627 4675 22633
rect 4617 22593 4629 22627
rect 4663 22593 4675 22627
rect 4617 22587 4675 22593
rect 4203 22528 4568 22556
rect 4632 22556 4660 22587
rect 4706 22584 4712 22636
rect 4764 22584 4770 22636
rect 4816 22633 4844 22664
rect 5000 22664 5540 22692
rect 5000 22633 5028 22664
rect 5534 22652 5540 22664
rect 5592 22692 5598 22704
rect 6822 22692 6828 22704
rect 5592 22664 6828 22692
rect 5592 22652 5598 22664
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22593 5043 22627
rect 4985 22587 5043 22593
rect 5166 22584 5172 22636
rect 5224 22584 5230 22636
rect 5350 22584 5356 22636
rect 5408 22584 5414 22636
rect 5442 22584 5448 22636
rect 5500 22584 5506 22636
rect 5626 22584 5632 22636
rect 5684 22584 5690 22636
rect 5810 22584 5816 22636
rect 5868 22584 5874 22636
rect 6196 22633 6224 22664
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 7650 22652 7656 22704
rect 7708 22652 7714 22704
rect 7926 22652 7932 22704
rect 7984 22652 7990 22704
rect 8478 22652 8484 22704
rect 8536 22692 8542 22704
rect 10704 22692 10732 22732
rect 12250 22720 12256 22732
rect 12308 22760 12314 22772
rect 12526 22760 12532 22772
rect 12308 22732 12532 22760
rect 12308 22720 12314 22732
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 12989 22763 13047 22769
rect 12989 22760 13001 22763
rect 12768 22732 13001 22760
rect 12768 22720 12774 22732
rect 12989 22729 13001 22732
rect 13035 22729 13047 22763
rect 12989 22723 13047 22729
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 15252 22732 15301 22760
rect 15252 22720 15258 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 17678 22720 17684 22772
rect 17736 22760 17742 22772
rect 18782 22760 18788 22772
rect 17736 22732 18788 22760
rect 17736 22720 17742 22732
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 19150 22720 19156 22772
rect 19208 22760 19214 22772
rect 19429 22763 19487 22769
rect 19429 22760 19441 22763
rect 19208 22732 19441 22760
rect 19208 22720 19214 22732
rect 19429 22729 19441 22732
rect 19475 22729 19487 22763
rect 19429 22723 19487 22729
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 22189 22763 22247 22769
rect 22189 22760 22201 22763
rect 20956 22732 22201 22760
rect 20956 22720 20962 22732
rect 22189 22729 22201 22732
rect 22235 22729 22247 22763
rect 22646 22760 22652 22772
rect 22189 22723 22247 22729
rect 22480 22732 22652 22760
rect 8536 22664 10732 22692
rect 11333 22695 11391 22701
rect 8536 22652 8542 22664
rect 11333 22661 11345 22695
rect 11379 22692 11391 22695
rect 11882 22692 11888 22704
rect 11379 22664 11888 22692
rect 11379 22661 11391 22664
rect 11333 22655 11391 22661
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 13624 22695 13682 22701
rect 13624 22661 13636 22695
rect 13670 22692 13682 22695
rect 19242 22692 19248 22704
rect 13670 22664 14504 22692
rect 13670 22661 13682 22664
rect 13624 22655 13682 22661
rect 6181 22627 6239 22633
rect 6181 22593 6193 22627
rect 6227 22593 6239 22627
rect 6638 22624 6644 22636
rect 6181 22587 6239 22593
rect 6472 22596 6644 22624
rect 5184 22556 5212 22584
rect 4632 22528 5212 22556
rect 5368 22556 5396 22584
rect 5368 22528 5672 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 5644 22500 5672 22528
rect 5718 22516 5724 22568
rect 5776 22556 5782 22568
rect 6472 22556 6500 22596
rect 6638 22584 6644 22596
rect 6696 22624 6702 22636
rect 7837 22627 7895 22633
rect 7837 22624 7849 22627
rect 6696 22596 7849 22624
rect 6696 22584 6702 22596
rect 7837 22593 7849 22596
rect 7883 22593 7895 22627
rect 8018 22624 8024 22636
rect 8076 22633 8082 22636
rect 7984 22596 8024 22624
rect 7837 22587 7895 22593
rect 8018 22584 8024 22596
rect 8076 22587 8084 22633
rect 9769 22627 9827 22633
rect 9769 22624 9781 22627
rect 9416 22596 9781 22624
rect 8076 22584 8082 22587
rect 5776 22528 6500 22556
rect 5776 22516 5782 22528
rect 6730 22516 6736 22568
rect 6788 22556 6794 22568
rect 9416 22556 9444 22596
rect 9769 22593 9781 22596
rect 9815 22624 9827 22627
rect 10226 22624 10232 22636
rect 9815 22596 10232 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 10226 22584 10232 22596
rect 10284 22624 10290 22636
rect 10965 22627 11023 22633
rect 10965 22624 10977 22627
rect 10284 22596 10977 22624
rect 10284 22584 10290 22596
rect 10965 22593 10977 22596
rect 11011 22593 11023 22627
rect 10965 22587 11023 22593
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22624 12035 22627
rect 12158 22624 12164 22636
rect 12023 22596 12164 22624
rect 12023 22593 12035 22596
rect 11977 22587 12035 22593
rect 12158 22584 12164 22596
rect 12216 22584 12222 22636
rect 12434 22584 12440 22636
rect 12492 22584 12498 22636
rect 12526 22584 12532 22636
rect 12584 22584 12590 22636
rect 12618 22584 12624 22636
rect 12676 22584 12682 22636
rect 13048 22627 13106 22633
rect 13048 22593 13060 22627
rect 13094 22624 13106 22627
rect 13354 22624 13360 22636
rect 13094 22596 13360 22624
rect 13094 22593 13106 22596
rect 13048 22587 13106 22593
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 13906 22584 13912 22636
rect 13964 22624 13970 22636
rect 14001 22627 14059 22633
rect 14001 22624 14013 22627
rect 13964 22596 14013 22624
rect 13964 22584 13970 22596
rect 14001 22593 14013 22596
rect 14047 22593 14059 22627
rect 14001 22587 14059 22593
rect 14182 22584 14188 22636
rect 14240 22624 14246 22636
rect 14369 22627 14427 22633
rect 14369 22624 14381 22627
rect 14240 22596 14381 22624
rect 14240 22584 14246 22596
rect 14369 22593 14381 22596
rect 14415 22593 14427 22627
rect 14369 22587 14427 22593
rect 6788 22528 9444 22556
rect 9585 22559 9643 22565
rect 6788 22516 6794 22528
rect 9585 22525 9597 22559
rect 9631 22556 9643 22559
rect 9858 22556 9864 22568
rect 9631 22528 9864 22556
rect 9631 22525 9643 22528
rect 9585 22519 9643 22525
rect 9858 22516 9864 22528
rect 9916 22516 9922 22568
rect 10137 22559 10195 22565
rect 10137 22525 10149 22559
rect 10183 22556 10195 22559
rect 11054 22556 11060 22568
rect 10183 22528 11060 22556
rect 10183 22525 10195 22528
rect 10137 22519 10195 22525
rect 11054 22516 11060 22528
rect 11112 22516 11118 22568
rect 11149 22559 11207 22565
rect 11149 22525 11161 22559
rect 11195 22525 11207 22559
rect 11149 22519 11207 22525
rect 11885 22559 11943 22565
rect 11885 22525 11897 22559
rect 11931 22556 11943 22559
rect 12066 22556 12072 22568
rect 11931 22528 12072 22556
rect 11931 22525 11943 22528
rect 11885 22519 11943 22525
rect 4062 22488 4068 22500
rect 3160 22460 4068 22488
rect 4062 22448 4068 22460
rect 4120 22448 4126 22500
rect 4430 22448 4436 22500
rect 4488 22488 4494 22500
rect 5350 22488 5356 22500
rect 4488 22460 5356 22488
rect 4488 22448 4494 22460
rect 5350 22448 5356 22460
rect 5408 22448 5414 22500
rect 5626 22448 5632 22500
rect 5684 22448 5690 22500
rect 6089 22491 6147 22497
rect 6089 22457 6101 22491
rect 6135 22488 6147 22491
rect 7466 22488 7472 22500
rect 6135 22460 7472 22488
rect 6135 22457 6147 22460
rect 6089 22451 6147 22457
rect 7466 22448 7472 22460
rect 7524 22448 7530 22500
rect 10686 22488 10692 22500
rect 7576 22460 10692 22488
rect 1670 22380 1676 22432
rect 1728 22420 1734 22432
rect 2501 22423 2559 22429
rect 2501 22420 2513 22423
rect 1728 22392 2513 22420
rect 1728 22380 1734 22392
rect 2501 22389 2513 22392
rect 2547 22389 2559 22423
rect 2501 22383 2559 22389
rect 4893 22423 4951 22429
rect 4893 22389 4905 22423
rect 4939 22420 4951 22423
rect 7576 22420 7604 22460
rect 10686 22448 10692 22460
rect 10744 22488 10750 22500
rect 10962 22488 10968 22500
rect 10744 22460 10968 22488
rect 10744 22448 10750 22460
rect 10962 22448 10968 22460
rect 11020 22448 11026 22500
rect 11164 22488 11192 22519
rect 12066 22516 12072 22528
rect 12124 22516 12130 22568
rect 12250 22488 12256 22500
rect 11164 22460 12256 22488
rect 12250 22448 12256 22460
rect 12308 22488 12314 22500
rect 12308 22460 12434 22488
rect 12308 22448 12314 22460
rect 4939 22392 7604 22420
rect 4939 22389 4951 22392
rect 4893 22383 4951 22389
rect 7650 22380 7656 22432
rect 7708 22380 7714 22432
rect 7926 22380 7932 22432
rect 7984 22420 7990 22432
rect 10318 22420 10324 22432
rect 7984 22392 10324 22420
rect 7984 22380 7990 22392
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 11054 22420 11060 22432
rect 10836 22392 11060 22420
rect 10836 22380 10842 22392
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 11241 22423 11299 22429
rect 11241 22389 11253 22423
rect 11287 22420 11299 22423
rect 11698 22420 11704 22432
rect 11287 22392 11704 22420
rect 11287 22389 11299 22392
rect 11241 22383 11299 22389
rect 11698 22380 11704 22392
rect 11756 22380 11762 22432
rect 12406 22420 12434 22460
rect 12636 22420 12664 22584
rect 14476 22556 14504 22664
rect 14568 22664 19248 22692
rect 14568 22633 14596 22664
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 20530 22692 20536 22704
rect 20364 22664 20536 22692
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 14645 22627 14703 22633
rect 14645 22593 14657 22627
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 14660 22556 14688 22587
rect 15562 22584 15568 22636
rect 15620 22584 15626 22636
rect 15746 22584 15752 22636
rect 15804 22584 15810 22636
rect 15930 22584 15936 22636
rect 15988 22624 15994 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 15988 22596 16129 22624
rect 15988 22584 15994 22596
rect 16117 22593 16129 22596
rect 16163 22624 16175 22627
rect 16850 22624 16856 22636
rect 16163 22596 16856 22624
rect 16163 22593 16175 22596
rect 16117 22587 16175 22593
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 17218 22624 17224 22636
rect 17175 22596 17224 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17218 22584 17224 22596
rect 17276 22584 17282 22636
rect 17586 22584 17592 22636
rect 17644 22584 17650 22636
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 17681 22587 17739 22593
rect 15838 22556 15844 22568
rect 14476 22528 14596 22556
rect 14660 22528 15844 22556
rect 14568 22500 14596 22528
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 16666 22516 16672 22568
rect 16724 22556 16730 22568
rect 17313 22559 17371 22565
rect 17313 22556 17325 22559
rect 16724 22528 17325 22556
rect 16724 22516 16730 22528
rect 17313 22525 17325 22528
rect 17359 22525 17371 22559
rect 17696 22556 17724 22587
rect 17770 22584 17776 22636
rect 17828 22584 17834 22636
rect 17957 22627 18015 22633
rect 17957 22593 17969 22627
rect 18003 22624 18015 22627
rect 18322 22624 18328 22636
rect 18003 22596 18328 22624
rect 18003 22593 18015 22596
rect 17957 22587 18015 22593
rect 18322 22584 18328 22596
rect 18380 22584 18386 22636
rect 18966 22584 18972 22636
rect 19024 22624 19030 22636
rect 19153 22627 19211 22633
rect 19153 22624 19165 22627
rect 19024 22596 19165 22624
rect 19024 22584 19030 22596
rect 19153 22593 19165 22596
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22624 19395 22627
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19383 22596 19625 22624
rect 19383 22593 19395 22596
rect 19337 22587 19395 22593
rect 19613 22593 19625 22596
rect 19659 22624 19671 22627
rect 19794 22624 19800 22636
rect 19659 22596 19800 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 19886 22584 19892 22636
rect 19944 22584 19950 22636
rect 20070 22584 20076 22636
rect 20128 22584 20134 22636
rect 20162 22584 20168 22636
rect 20220 22584 20226 22636
rect 20364 22633 20392 22664
rect 20530 22652 20536 22664
rect 20588 22692 20594 22704
rect 21266 22692 21272 22704
rect 20588 22664 21272 22692
rect 20588 22652 20594 22664
rect 21266 22652 21272 22664
rect 21324 22652 21330 22704
rect 22002 22652 22008 22704
rect 22060 22652 22066 22704
rect 22480 22692 22508 22732
rect 22646 22720 22652 22732
rect 22704 22720 22710 22772
rect 23109 22763 23167 22769
rect 23109 22729 23121 22763
rect 23155 22760 23167 22763
rect 23382 22760 23388 22772
rect 23155 22732 23388 22760
rect 23155 22729 23167 22732
rect 23109 22723 23167 22729
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 25225 22763 25283 22769
rect 25225 22729 25237 22763
rect 25271 22760 25283 22763
rect 25498 22760 25504 22772
rect 25271 22732 25504 22760
rect 25271 22729 25283 22732
rect 25225 22723 25283 22729
rect 25498 22720 25504 22732
rect 25556 22720 25562 22772
rect 26142 22720 26148 22772
rect 26200 22760 26206 22772
rect 26878 22760 26884 22772
rect 26200 22732 26884 22760
rect 26200 22720 26206 22732
rect 26878 22720 26884 22732
rect 26936 22720 26942 22772
rect 26970 22720 26976 22772
rect 27028 22720 27034 22772
rect 27985 22763 28043 22769
rect 27985 22729 27997 22763
rect 28031 22760 28043 22763
rect 30558 22760 30564 22772
rect 28031 22732 30564 22760
rect 28031 22729 28043 22732
rect 27985 22723 28043 22729
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 30834 22720 30840 22772
rect 30892 22760 30898 22772
rect 30929 22763 30987 22769
rect 30929 22760 30941 22763
rect 30892 22732 30941 22760
rect 30892 22720 30898 22732
rect 30929 22729 30941 22732
rect 30975 22729 30987 22763
rect 30929 22723 30987 22729
rect 31478 22720 31484 22772
rect 31536 22760 31542 22772
rect 31536 22732 34284 22760
rect 31536 22720 31542 22732
rect 22112 22664 22508 22692
rect 22557 22695 22615 22701
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 20990 22584 20996 22636
rect 21048 22584 21054 22636
rect 21174 22584 21180 22636
rect 21232 22584 21238 22636
rect 21361 22627 21419 22633
rect 21361 22593 21373 22627
rect 21407 22624 21419 22627
rect 21450 22624 21456 22636
rect 21407 22596 21456 22624
rect 21407 22593 21419 22596
rect 21361 22587 21419 22593
rect 21450 22584 21456 22596
rect 21508 22624 21514 22636
rect 21726 22624 21732 22636
rect 21508 22596 21732 22624
rect 21508 22584 21514 22596
rect 21726 22584 21732 22596
rect 21784 22584 21790 22636
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22624 21879 22627
rect 21910 22624 21916 22636
rect 21867 22596 21916 22624
rect 21867 22593 21879 22596
rect 21821 22587 21879 22593
rect 21910 22584 21916 22596
rect 21968 22584 21974 22636
rect 22112 22633 22140 22664
rect 22557 22661 22569 22695
rect 22603 22692 22615 22695
rect 22603 22664 26556 22692
rect 22603 22661 22615 22664
rect 22557 22655 22615 22661
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22593 22155 22627
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 22097 22587 22155 22593
rect 22204 22596 22385 22624
rect 18138 22556 18144 22568
rect 17696 22528 18144 22556
rect 17313 22519 17371 22525
rect 18138 22516 18144 22528
rect 18196 22556 18202 22568
rect 18196 22528 19196 22556
rect 18196 22516 18202 22528
rect 19168 22500 19196 22528
rect 19242 22516 19248 22568
rect 19300 22516 19306 22568
rect 12802 22448 12808 22500
rect 12860 22488 12866 22500
rect 13078 22488 13084 22500
rect 12860 22460 13084 22488
rect 12860 22448 12866 22460
rect 13078 22448 13084 22460
rect 13136 22488 13142 22500
rect 13449 22491 13507 22497
rect 13449 22488 13461 22491
rect 13136 22460 13461 22488
rect 13136 22448 13142 22460
rect 13449 22457 13461 22460
rect 13495 22457 13507 22491
rect 14274 22488 14280 22500
rect 13449 22451 13507 22457
rect 13648 22460 14280 22488
rect 12406 22392 12664 22420
rect 12710 22380 12716 22432
rect 12768 22420 12774 22432
rect 13648 22429 13676 22460
rect 14274 22448 14280 22460
rect 14332 22448 14338 22500
rect 14550 22448 14556 22500
rect 14608 22448 14614 22500
rect 16298 22448 16304 22500
rect 16356 22488 16362 22500
rect 18506 22488 18512 22500
rect 16356 22460 18512 22488
rect 16356 22448 16362 22460
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 18782 22448 18788 22500
rect 18840 22488 18846 22500
rect 19058 22488 19064 22500
rect 18840 22460 19064 22488
rect 18840 22448 18846 22460
rect 19058 22448 19064 22460
rect 19116 22448 19122 22500
rect 19150 22448 19156 22500
rect 19208 22448 19214 22500
rect 21821 22491 21879 22497
rect 21821 22457 21833 22491
rect 21867 22488 21879 22491
rect 22094 22488 22100 22500
rect 21867 22460 22100 22488
rect 21867 22457 21879 22460
rect 21821 22451 21879 22457
rect 22094 22448 22100 22460
rect 22152 22448 22158 22500
rect 13173 22423 13231 22429
rect 13173 22420 13185 22423
rect 12768 22392 13185 22420
rect 12768 22380 12774 22392
rect 13173 22389 13185 22392
rect 13219 22389 13231 22423
rect 13173 22383 13231 22389
rect 13633 22423 13691 22429
rect 13633 22389 13645 22423
rect 13679 22389 13691 22423
rect 13633 22383 13691 22389
rect 14182 22380 14188 22432
rect 14240 22380 14246 22432
rect 18138 22380 18144 22432
rect 18196 22420 18202 22432
rect 19610 22420 19616 22432
rect 18196 22392 19616 22420
rect 18196 22380 18202 22392
rect 19610 22380 19616 22392
rect 19668 22380 19674 22432
rect 20254 22380 20260 22432
rect 20312 22380 20318 22432
rect 20622 22380 20628 22432
rect 20680 22420 20686 22432
rect 22204 22420 22232 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 22646 22584 22652 22636
rect 22704 22584 22710 22636
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22624 23167 22627
rect 23198 22624 23204 22636
rect 23155 22596 23204 22624
rect 23155 22593 23167 22596
rect 23109 22587 23167 22593
rect 23198 22584 23204 22596
rect 23256 22584 23262 22636
rect 24118 22584 24124 22636
rect 24176 22584 24182 22636
rect 24210 22584 24216 22636
rect 24268 22624 24274 22636
rect 24305 22627 24363 22633
rect 24305 22624 24317 22627
rect 24268 22596 24317 22624
rect 24268 22584 24274 22596
rect 24305 22593 24317 22596
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24394 22584 24400 22636
rect 24452 22584 24458 22636
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22624 24547 22627
rect 24670 22624 24676 22636
rect 24535 22596 24676 22624
rect 24535 22593 24547 22596
rect 24489 22587 24547 22593
rect 24670 22584 24676 22596
rect 24728 22624 24734 22636
rect 25317 22627 25375 22633
rect 25317 22624 25329 22627
rect 24728 22596 25329 22624
rect 24728 22584 24734 22596
rect 25317 22593 25329 22596
rect 25363 22593 25375 22627
rect 25317 22587 25375 22593
rect 22738 22516 22744 22568
rect 22796 22516 22802 22568
rect 23293 22559 23351 22565
rect 23293 22525 23305 22559
rect 23339 22556 23351 22559
rect 23339 22528 25360 22556
rect 23339 22525 23351 22528
rect 23293 22519 23351 22525
rect 22370 22448 22376 22500
rect 22428 22488 22434 22500
rect 23308 22488 23336 22519
rect 22428 22460 23336 22488
rect 22428 22448 22434 22460
rect 24118 22420 24124 22432
rect 20680 22392 24124 22420
rect 20680 22380 20686 22392
rect 24118 22380 24124 22392
rect 24176 22420 24182 22432
rect 24486 22420 24492 22432
rect 24176 22392 24492 22420
rect 24176 22380 24182 22392
rect 24486 22380 24492 22392
rect 24544 22380 24550 22432
rect 24762 22380 24768 22432
rect 24820 22380 24826 22432
rect 25332 22420 25360 22528
rect 26528 22488 26556 22664
rect 27062 22652 27068 22704
rect 27120 22692 27126 22704
rect 28261 22695 28319 22701
rect 28261 22692 28273 22695
rect 27120 22664 28273 22692
rect 27120 22652 27126 22664
rect 28261 22661 28273 22664
rect 28307 22661 28319 22695
rect 28261 22655 28319 22661
rect 28350 22652 28356 22704
rect 28408 22652 28414 22704
rect 28460 22664 29500 22692
rect 26970 22584 26976 22636
rect 27028 22624 27034 22636
rect 27249 22627 27307 22633
rect 27249 22624 27261 22627
rect 27028 22596 27261 22624
rect 27028 22584 27034 22596
rect 27249 22593 27261 22596
rect 27295 22593 27307 22627
rect 27249 22587 27307 22593
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 27433 22627 27491 22633
rect 27433 22593 27445 22627
rect 27479 22593 27491 22627
rect 27433 22587 27491 22593
rect 26602 22516 26608 22568
rect 26660 22556 26666 22568
rect 27154 22556 27160 22568
rect 26660 22528 27160 22556
rect 26660 22516 26666 22528
rect 27154 22516 27160 22528
rect 27212 22516 27218 22568
rect 27448 22488 27476 22587
rect 27522 22584 27528 22636
rect 27580 22624 27586 22636
rect 27617 22627 27675 22633
rect 27617 22624 27629 22627
rect 27580 22596 27629 22624
rect 27580 22584 27586 22596
rect 27617 22593 27629 22596
rect 27663 22593 27675 22627
rect 27617 22587 27675 22593
rect 28164 22627 28222 22633
rect 28164 22593 28176 22627
rect 28210 22593 28222 22627
rect 28164 22587 28222 22593
rect 27522 22488 27528 22500
rect 26528 22460 27528 22488
rect 27522 22448 27528 22460
rect 27580 22448 27586 22500
rect 28179 22488 28207 22587
rect 28460 22488 28488 22664
rect 28536 22627 28594 22633
rect 28536 22593 28548 22627
rect 28582 22593 28594 22627
rect 28536 22587 28594 22593
rect 28629 22627 28687 22633
rect 28629 22593 28641 22627
rect 28675 22624 28687 22627
rect 28675 22596 29224 22624
rect 28675 22593 28687 22596
rect 28629 22587 28687 22593
rect 28552 22500 28580 22587
rect 29196 22565 29224 22596
rect 29362 22584 29368 22636
rect 29420 22584 29426 22636
rect 29472 22633 29500 22664
rect 29546 22652 29552 22704
rect 29604 22692 29610 22704
rect 31110 22692 31116 22704
rect 29604 22664 30696 22692
rect 29604 22652 29610 22664
rect 29457 22627 29515 22633
rect 29457 22593 29469 22627
rect 29503 22624 29515 22627
rect 29914 22624 29920 22636
rect 29503 22596 29920 22624
rect 29503 22593 29515 22596
rect 29457 22587 29515 22593
rect 29914 22584 29920 22596
rect 29972 22584 29978 22636
rect 30006 22584 30012 22636
rect 30064 22584 30070 22636
rect 30190 22584 30196 22636
rect 30248 22584 30254 22636
rect 30282 22584 30288 22636
rect 30340 22624 30346 22636
rect 30668 22633 30696 22664
rect 31052 22664 31116 22692
rect 30377 22627 30435 22633
rect 30377 22624 30389 22627
rect 30340 22596 30389 22624
rect 30340 22584 30346 22596
rect 30377 22593 30389 22596
rect 30423 22593 30435 22627
rect 30377 22587 30435 22593
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22593 30527 22627
rect 30469 22587 30527 22593
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 30653 22587 30711 22593
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22624 30803 22627
rect 30834 22624 30840 22636
rect 30791 22596 30840 22624
rect 30791 22593 30803 22596
rect 30745 22587 30803 22593
rect 29181 22559 29239 22565
rect 29181 22525 29193 22559
rect 29227 22525 29239 22559
rect 29181 22519 29239 22525
rect 28179 22460 28488 22488
rect 28534 22448 28540 22500
rect 28592 22448 28598 22500
rect 29196 22488 29224 22519
rect 29270 22516 29276 22568
rect 29328 22516 29334 22568
rect 30101 22559 30159 22565
rect 30101 22525 30113 22559
rect 30147 22525 30159 22559
rect 30101 22519 30159 22525
rect 29733 22491 29791 22497
rect 29733 22488 29745 22491
rect 29196 22460 29745 22488
rect 29733 22457 29745 22460
rect 29779 22457 29791 22491
rect 30116 22488 30144 22519
rect 30190 22488 30196 22500
rect 30116 22460 30196 22488
rect 29733 22451 29791 22457
rect 30190 22448 30196 22460
rect 30248 22448 30254 22500
rect 26878 22420 26884 22432
rect 25332 22392 26884 22420
rect 26878 22380 26884 22392
rect 26936 22380 26942 22432
rect 28074 22380 28080 22432
rect 28132 22420 28138 22432
rect 28902 22420 28908 22432
rect 28132 22392 28908 22420
rect 28132 22380 28138 22392
rect 28902 22380 28908 22392
rect 28960 22420 28966 22432
rect 29546 22420 29552 22432
rect 28960 22392 29552 22420
rect 28960 22380 28966 22392
rect 29546 22380 29552 22392
rect 29604 22380 29610 22432
rect 29641 22423 29699 22429
rect 29641 22389 29653 22423
rect 29687 22420 29699 22423
rect 30484 22420 30512 22587
rect 30834 22584 30840 22596
rect 30892 22584 30898 22636
rect 31052 22488 31080 22664
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 31846 22652 31852 22704
rect 31904 22692 31910 22704
rect 32125 22695 32183 22701
rect 32125 22692 32137 22695
rect 31904 22664 32137 22692
rect 31904 22652 31910 22664
rect 32125 22661 32137 22664
rect 32171 22661 32183 22695
rect 32769 22695 32827 22701
rect 32125 22655 32183 22661
rect 32232 22664 32536 22692
rect 31205 22630 31263 22633
rect 31205 22627 31432 22630
rect 31205 22593 31217 22627
rect 31251 22624 31432 22627
rect 31570 22624 31576 22636
rect 31251 22602 31576 22624
rect 31251 22593 31263 22602
rect 31404 22596 31576 22602
rect 31205 22587 31263 22593
rect 31570 22584 31576 22596
rect 31628 22624 31634 22636
rect 32232 22624 32260 22664
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 31628 22596 32260 22624
rect 32324 22596 32413 22624
rect 31628 22584 31634 22596
rect 31110 22516 31116 22568
rect 31168 22516 31174 22568
rect 31297 22559 31355 22565
rect 31297 22525 31309 22559
rect 31343 22525 31355 22559
rect 31297 22519 31355 22525
rect 31312 22488 31340 22519
rect 31386 22516 31392 22568
rect 31444 22516 31450 22568
rect 32214 22516 32220 22568
rect 32272 22516 32278 22568
rect 31052 22460 31340 22488
rect 32324 22488 32352 22596
rect 32401 22593 32413 22596
rect 32447 22593 32459 22627
rect 32508 22624 32536 22664
rect 32769 22661 32781 22695
rect 32815 22692 32827 22695
rect 32950 22692 32956 22704
rect 32815 22664 32956 22692
rect 32815 22661 32827 22664
rect 32769 22655 32827 22661
rect 32950 22652 32956 22664
rect 33008 22692 33014 22704
rect 34256 22701 34284 22732
rect 34422 22720 34428 22772
rect 34480 22720 34486 22772
rect 33137 22695 33195 22701
rect 33137 22692 33149 22695
rect 33008 22664 33149 22692
rect 33008 22652 33014 22664
rect 33137 22661 33149 22664
rect 33183 22661 33195 22695
rect 33137 22655 33195 22661
rect 34241 22695 34299 22701
rect 34241 22661 34253 22695
rect 34287 22661 34299 22695
rect 34241 22655 34299 22661
rect 34330 22652 34336 22704
rect 34388 22652 34394 22704
rect 34440 22692 34468 22720
rect 34440 22664 34560 22692
rect 32508 22596 32812 22624
rect 32401 22587 32459 22593
rect 32784 22556 32812 22596
rect 32858 22584 32864 22636
rect 32916 22584 32922 22636
rect 33042 22584 33048 22636
rect 33100 22584 33106 22636
rect 33226 22584 33232 22636
rect 33284 22624 33290 22636
rect 34532 22633 34560 22664
rect 34149 22627 34207 22633
rect 34149 22624 34161 22627
rect 33284 22596 34161 22624
rect 33284 22584 33290 22596
rect 34149 22593 34161 22596
rect 34195 22593 34207 22627
rect 34149 22587 34207 22593
rect 34517 22627 34575 22633
rect 34517 22593 34529 22627
rect 34563 22593 34575 22627
rect 34517 22587 34575 22593
rect 34882 22584 34888 22636
rect 34940 22584 34946 22636
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22624 35219 22627
rect 35342 22624 35348 22636
rect 35207 22596 35348 22624
rect 35207 22593 35219 22596
rect 35161 22587 35219 22593
rect 35342 22584 35348 22596
rect 35400 22584 35406 22636
rect 35897 22559 35955 22565
rect 35897 22556 35909 22559
rect 32784 22528 35909 22556
rect 35897 22525 35909 22528
rect 35943 22525 35955 22559
rect 35897 22519 35955 22525
rect 36170 22516 36176 22568
rect 36228 22516 36234 22568
rect 33413 22491 33471 22497
rect 33413 22488 33425 22491
rect 32324 22460 33425 22488
rect 33413 22457 33425 22460
rect 33459 22488 33471 22491
rect 33459 22460 33548 22488
rect 33459 22457 33471 22460
rect 33413 22451 33471 22457
rect 33520 22432 33548 22460
rect 34606 22448 34612 22500
rect 34664 22488 34670 22500
rect 35161 22491 35219 22497
rect 35161 22488 35173 22491
rect 34664 22460 35173 22488
rect 34664 22448 34670 22460
rect 35161 22457 35173 22460
rect 35207 22457 35219 22491
rect 35161 22451 35219 22457
rect 29687 22392 30512 22420
rect 29687 22389 29699 22392
rect 29641 22383 29699 22389
rect 31570 22380 31576 22432
rect 31628 22380 31634 22432
rect 31662 22380 31668 22432
rect 31720 22420 31726 22432
rect 32125 22423 32183 22429
rect 32125 22420 32137 22423
rect 31720 22392 32137 22420
rect 31720 22380 31726 22392
rect 32125 22389 32137 22392
rect 32171 22389 32183 22423
rect 32125 22383 32183 22389
rect 32398 22380 32404 22432
rect 32456 22420 32462 22432
rect 32585 22423 32643 22429
rect 32585 22420 32597 22423
rect 32456 22392 32597 22420
rect 32456 22380 32462 22392
rect 32585 22389 32597 22392
rect 32631 22389 32643 22423
rect 32585 22383 32643 22389
rect 33502 22380 33508 22432
rect 33560 22380 33566 22432
rect 33962 22380 33968 22432
rect 34020 22380 34026 22432
rect 1104 22330 36524 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 36524 22330
rect 1104 22256 36524 22278
rect 1670 22225 1676 22228
rect 1660 22219 1676 22225
rect 1660 22185 1672 22219
rect 1660 22179 1676 22185
rect 1670 22176 1676 22179
rect 1728 22176 1734 22228
rect 3694 22176 3700 22228
rect 3752 22176 3758 22228
rect 3970 22176 3976 22228
rect 4028 22216 4034 22228
rect 4617 22219 4675 22225
rect 4028 22188 4476 22216
rect 4028 22176 4034 22188
rect 2774 22108 2780 22160
rect 2832 22148 2838 22160
rect 3712 22148 3740 22176
rect 2832 22120 4292 22148
rect 2832 22108 2838 22120
rect 1394 22040 1400 22092
rect 1452 22080 1458 22092
rect 2682 22080 2688 22092
rect 1452 22052 2688 22080
rect 1452 22040 1458 22052
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 3145 22083 3203 22089
rect 3145 22049 3157 22083
rect 3191 22080 3203 22083
rect 3970 22080 3976 22092
rect 3191 22052 3976 22080
rect 3191 22049 3203 22052
rect 3145 22043 3203 22049
rect 3970 22040 3976 22052
rect 4028 22040 4034 22092
rect 4264 22089 4292 22120
rect 4249 22083 4307 22089
rect 4249 22049 4261 22083
rect 4295 22049 4307 22083
rect 4249 22043 4307 22049
rect 4338 22040 4344 22092
rect 4396 22040 4402 22092
rect 4448 22080 4476 22188
rect 4617 22185 4629 22219
rect 4663 22216 4675 22219
rect 4706 22216 4712 22228
rect 4663 22188 4712 22216
rect 4663 22185 4675 22188
rect 4617 22179 4675 22185
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 8018 22176 8024 22228
rect 8076 22216 8082 22228
rect 8113 22219 8171 22225
rect 8113 22216 8125 22219
rect 8076 22188 8125 22216
rect 8076 22176 8082 22188
rect 8113 22185 8125 22188
rect 8159 22185 8171 22219
rect 8113 22179 8171 22185
rect 8294 22176 8300 22228
rect 8352 22216 8358 22228
rect 9582 22216 9588 22228
rect 8352 22188 9588 22216
rect 8352 22176 8358 22188
rect 9582 22176 9588 22188
rect 9640 22216 9646 22228
rect 14182 22216 14188 22228
rect 9640 22188 14188 22216
rect 9640 22176 9646 22188
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 14274 22176 14280 22228
rect 14332 22176 14338 22228
rect 15470 22176 15476 22228
rect 15528 22176 15534 22228
rect 20254 22216 20260 22228
rect 15580 22188 20260 22216
rect 5166 22108 5172 22160
rect 5224 22148 5230 22160
rect 5224 22120 6132 22148
rect 5224 22108 5230 22120
rect 5626 22080 5632 22092
rect 4448 22052 5396 22080
rect 4796 22015 4854 22021
rect 4796 21981 4808 22015
rect 4842 22012 4854 22015
rect 5074 22012 5080 22024
rect 4842 21984 5080 22012
rect 4842 21981 4854 21984
rect 4796 21975 4854 21981
rect 5074 21972 5080 21984
rect 5132 21972 5138 22024
rect 5166 21972 5172 22024
rect 5224 21972 5230 22024
rect 5258 21972 5264 22024
rect 5316 21972 5322 22024
rect 5368 22021 5396 22052
rect 5552 22052 5632 22080
rect 5552 22021 5580 22052
rect 5626 22040 5632 22052
rect 5684 22040 5690 22092
rect 6104 22024 6132 22120
rect 6638 22108 6644 22160
rect 6696 22108 6702 22160
rect 7466 22108 7472 22160
rect 7524 22148 7530 22160
rect 8478 22148 8484 22160
rect 7524 22120 8484 22148
rect 7524 22108 7530 22120
rect 8478 22108 8484 22120
rect 8536 22108 8542 22160
rect 8941 22151 8999 22157
rect 8941 22117 8953 22151
rect 8987 22148 8999 22151
rect 9306 22148 9312 22160
rect 8987 22120 9312 22148
rect 8987 22117 8999 22120
rect 8941 22111 8999 22117
rect 9306 22108 9312 22120
rect 9364 22108 9370 22160
rect 9858 22108 9864 22160
rect 9916 22148 9922 22160
rect 11701 22151 11759 22157
rect 11701 22148 11713 22151
rect 9916 22120 11713 22148
rect 9916 22108 9922 22120
rect 11701 22117 11713 22120
rect 11747 22117 11759 22151
rect 12158 22148 12164 22160
rect 11701 22111 11759 22117
rect 11808 22120 12164 22148
rect 6656 22080 6684 22108
rect 6380 22052 6684 22080
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 21981 5411 22015
rect 5353 21975 5411 21981
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 2958 21944 2964 21956
rect 2898 21916 2964 21944
rect 2958 21904 2964 21916
rect 3016 21904 3022 21956
rect 4614 21944 4620 21956
rect 3712 21916 4620 21944
rect 2406 21836 2412 21888
rect 2464 21876 2470 21888
rect 3712 21876 3740 21916
rect 4614 21904 4620 21916
rect 4672 21944 4678 21956
rect 4893 21947 4951 21953
rect 4893 21944 4905 21947
rect 4672 21916 4905 21944
rect 4672 21904 4678 21916
rect 4893 21913 4905 21916
rect 4939 21913 4951 21947
rect 4893 21907 4951 21913
rect 4985 21947 5043 21953
rect 4985 21913 4997 21947
rect 5031 21944 5043 21947
rect 5552 21944 5580 21975
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 6086 21972 6092 22024
rect 6144 21972 6150 22024
rect 6178 21972 6184 22024
rect 6236 22012 6242 22024
rect 6380 22021 6408 22052
rect 6730 22040 6736 22092
rect 6788 22040 6794 22092
rect 7650 22040 7656 22092
rect 7708 22040 7714 22092
rect 7742 22040 7748 22092
rect 7800 22040 7806 22092
rect 10888 22052 11376 22080
rect 10888 22024 10916 22052
rect 6273 22015 6331 22021
rect 6273 22012 6285 22015
rect 6236 21984 6285 22012
rect 6236 21972 6242 21984
rect 6273 21981 6285 21984
rect 6319 21981 6331 22015
rect 6273 21975 6331 21981
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 6549 22015 6607 22021
rect 6549 21981 6561 22015
rect 6595 22012 6607 22015
rect 6641 22015 6699 22021
rect 6641 22012 6653 22015
rect 6595 21984 6653 22012
rect 6595 21981 6607 21984
rect 6549 21975 6607 21981
rect 6641 21981 6653 21984
rect 6687 21981 6699 22015
rect 6641 21975 6699 21981
rect 6822 21972 6828 22024
rect 6880 21972 6886 22024
rect 7466 21972 7472 22024
rect 7524 21972 7530 22024
rect 7558 21972 7564 22024
rect 7616 21972 7622 22024
rect 8665 22015 8723 22021
rect 8665 21981 8677 22015
rect 8711 22012 8723 22015
rect 8754 22012 8760 22024
rect 8711 21984 8760 22012
rect 8711 21981 8723 21984
rect 8665 21975 8723 21981
rect 8754 21972 8760 21984
rect 8812 21972 8818 22024
rect 9309 22015 9367 22021
rect 9216 21993 9274 21999
rect 9216 21959 9228 21993
rect 9262 21959 9274 21993
rect 9309 21981 9321 22015
rect 9355 21981 9367 22015
rect 9309 21975 9367 21981
rect 9216 21956 9274 21959
rect 5031 21916 5580 21944
rect 5629 21947 5687 21953
rect 5031 21913 5043 21916
rect 4985 21907 5043 21913
rect 5629 21913 5641 21947
rect 5675 21944 5687 21947
rect 6454 21944 6460 21956
rect 5675 21916 6460 21944
rect 5675 21913 5687 21916
rect 5629 21907 5687 21913
rect 2464 21848 3740 21876
rect 2464 21836 2470 21848
rect 3786 21836 3792 21888
rect 3844 21836 3850 21888
rect 4157 21879 4215 21885
rect 4157 21845 4169 21879
rect 4203 21876 4215 21879
rect 4430 21876 4436 21888
rect 4203 21848 4436 21876
rect 4203 21845 4215 21848
rect 4157 21839 4215 21845
rect 4430 21836 4436 21848
rect 4488 21836 4494 21888
rect 4706 21836 4712 21888
rect 4764 21876 4770 21888
rect 5000 21876 5028 21907
rect 6288 21888 6316 21916
rect 6454 21904 6460 21916
rect 6512 21904 6518 21956
rect 8288 21947 8346 21953
rect 8288 21913 8300 21947
rect 8334 21944 8346 21947
rect 9214 21944 9220 21956
rect 8334 21916 9220 21944
rect 8334 21913 8346 21916
rect 8288 21907 8346 21913
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 9329 21944 9357 21975
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 9582 21972 9588 22024
rect 9640 21972 9646 22024
rect 9858 21972 9864 22024
rect 9916 21972 9922 22024
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10137 22015 10195 22021
rect 10137 22012 10149 22015
rect 10100 21984 10149 22012
rect 10100 21972 10106 21984
rect 10137 21981 10149 21984
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 11054 21972 11060 22024
rect 11112 21972 11118 22024
rect 11146 21972 11152 22024
rect 11204 21972 11210 22024
rect 11348 22021 11376 22052
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 11808 22012 11836 22120
rect 12158 22108 12164 22120
rect 12216 22108 12222 22160
rect 14366 22148 14372 22160
rect 13648 22120 14372 22148
rect 12802 22080 12808 22092
rect 11900 22052 12808 22080
rect 11900 22021 11928 22052
rect 12802 22040 12808 22052
rect 12860 22040 12866 22092
rect 13648 22080 13676 22120
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 14550 22108 14556 22160
rect 14608 22148 14614 22160
rect 15580 22148 15608 22188
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 24854 22176 24860 22228
rect 24912 22216 24918 22228
rect 27154 22216 27160 22228
rect 24912 22188 27160 22216
rect 24912 22176 24918 22188
rect 27154 22176 27160 22188
rect 27212 22176 27218 22228
rect 29362 22176 29368 22228
rect 29420 22216 29426 22228
rect 29917 22219 29975 22225
rect 29917 22216 29929 22219
rect 29420 22188 29929 22216
rect 29420 22176 29426 22188
rect 29917 22185 29929 22188
rect 29963 22185 29975 22219
rect 29917 22179 29975 22185
rect 30006 22176 30012 22228
rect 30064 22176 30070 22228
rect 30101 22219 30159 22225
rect 30101 22185 30113 22219
rect 30147 22216 30159 22219
rect 30374 22216 30380 22228
rect 30147 22188 30380 22216
rect 30147 22185 30159 22188
rect 30101 22179 30159 22185
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 30837 22219 30895 22225
rect 30837 22185 30849 22219
rect 30883 22185 30895 22219
rect 30837 22179 30895 22185
rect 31021 22219 31079 22225
rect 31021 22185 31033 22219
rect 31067 22216 31079 22219
rect 31110 22216 31116 22228
rect 31067 22188 31116 22216
rect 31067 22185 31079 22188
rect 31021 22179 31079 22185
rect 14608 22120 15608 22148
rect 14608 22108 14614 22120
rect 15746 22108 15752 22160
rect 15804 22148 15810 22160
rect 15804 22120 16620 22148
rect 15804 22108 15810 22120
rect 15856 22089 15884 22120
rect 15841 22083 15899 22089
rect 13004 22052 13676 22080
rect 14384 22052 15792 22080
rect 11379 21984 11836 22012
rect 11885 22015 11943 22021
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 11885 21981 11897 22015
rect 11931 21981 11943 22015
rect 11885 21975 11943 21981
rect 9876 21944 9904 21972
rect 9329 21916 9904 21944
rect 10594 21904 10600 21956
rect 10652 21944 10658 21956
rect 11900 21944 11928 21975
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 13004 22012 13032 22052
rect 12207 21984 13032 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 13078 21972 13084 22024
rect 13136 21972 13142 22024
rect 13265 22015 13323 22021
rect 13265 21981 13277 22015
rect 13311 22012 13323 22015
rect 13311 21984 13492 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 10652 21916 11928 21944
rect 10652 21904 10658 21916
rect 12434 21904 12440 21956
rect 12492 21944 12498 21956
rect 12897 21947 12955 21953
rect 12897 21944 12909 21947
rect 12492 21916 12909 21944
rect 12492 21904 12498 21916
rect 12897 21913 12909 21916
rect 12943 21913 12955 21947
rect 12897 21907 12955 21913
rect 4764 21848 5028 21876
rect 4764 21836 4770 21848
rect 5442 21836 5448 21888
rect 5500 21876 5506 21888
rect 5905 21879 5963 21885
rect 5905 21876 5917 21879
rect 5500 21848 5917 21876
rect 5500 21836 5506 21848
rect 5905 21845 5917 21848
rect 5951 21845 5963 21879
rect 5905 21839 5963 21845
rect 6270 21836 6276 21888
rect 6328 21836 6334 21888
rect 7926 21836 7932 21888
rect 7984 21836 7990 21888
rect 8754 21836 8760 21888
rect 8812 21876 8818 21888
rect 9398 21876 9404 21888
rect 8812 21848 9404 21876
rect 8812 21836 8818 21848
rect 9398 21836 9404 21848
rect 9456 21876 9462 21888
rect 9677 21879 9735 21885
rect 9677 21876 9689 21879
rect 9456 21848 9689 21876
rect 9456 21836 9462 21848
rect 9677 21845 9689 21848
rect 9723 21845 9735 21879
rect 9677 21839 9735 21845
rect 10045 21879 10103 21885
rect 10045 21845 10057 21879
rect 10091 21876 10103 21879
rect 10134 21876 10140 21888
rect 10091 21848 10140 21876
rect 10091 21845 10103 21848
rect 10045 21839 10103 21845
rect 10134 21836 10140 21848
rect 10192 21836 10198 21888
rect 10965 21879 11023 21885
rect 10965 21845 10977 21879
rect 11011 21876 11023 21879
rect 11054 21876 11060 21888
rect 11011 21848 11060 21876
rect 11011 21845 11023 21848
rect 10965 21839 11023 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 11241 21879 11299 21885
rect 11241 21876 11253 21879
rect 11204 21848 11253 21876
rect 11204 21836 11210 21848
rect 11241 21845 11253 21848
rect 11287 21845 11299 21879
rect 11241 21839 11299 21845
rect 11606 21836 11612 21888
rect 11664 21876 11670 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 11664 21848 13369 21876
rect 11664 21836 11670 21848
rect 13357 21845 13369 21848
rect 13403 21845 13415 21879
rect 13464 21876 13492 21984
rect 13538 21972 13544 22024
rect 13596 21972 13602 22024
rect 13817 22015 13875 22021
rect 13817 22012 13829 22015
rect 13648 21984 13829 22012
rect 13648 21876 13676 21984
rect 13817 21981 13829 21984
rect 13863 22012 13875 22015
rect 13906 22012 13912 22024
rect 13863 21984 13912 22012
rect 13863 21981 13875 21984
rect 13817 21975 13875 21981
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14384 22021 14412 22052
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 22012 14519 22015
rect 14550 22012 14556 22024
rect 14507 21984 14556 22012
rect 14507 21981 14519 21984
rect 14461 21975 14519 21981
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 15657 22015 15715 22021
rect 15657 21981 15669 22015
rect 15703 21981 15715 22015
rect 15764 22012 15792 22052
rect 15841 22049 15853 22083
rect 15887 22049 15899 22083
rect 15841 22043 15899 22049
rect 16022 22040 16028 22092
rect 16080 22040 16086 22092
rect 15930 22012 15936 22024
rect 15764 21984 15936 22012
rect 15657 21975 15715 21981
rect 13725 21947 13783 21953
rect 13725 21913 13737 21947
rect 13771 21944 13783 21947
rect 15672 21944 15700 21975
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 16040 21944 16068 22040
rect 16114 21972 16120 22024
rect 16172 21972 16178 22024
rect 16592 22012 16620 22120
rect 16758 22108 16764 22160
rect 16816 22148 16822 22160
rect 18138 22148 18144 22160
rect 16816 22120 18144 22148
rect 16816 22108 16822 22120
rect 18138 22108 18144 22120
rect 18196 22148 18202 22160
rect 18233 22151 18291 22157
rect 18233 22148 18245 22151
rect 18196 22120 18245 22148
rect 18196 22108 18202 22120
rect 18233 22117 18245 22120
rect 18279 22117 18291 22151
rect 18233 22111 18291 22117
rect 18417 22151 18475 22157
rect 18417 22117 18429 22151
rect 18463 22117 18475 22151
rect 18417 22111 18475 22117
rect 16850 22040 16856 22092
rect 16908 22080 16914 22092
rect 17402 22080 17408 22092
rect 16908 22052 17408 22080
rect 16908 22040 16914 22052
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 18432 22080 18460 22111
rect 18966 22108 18972 22160
rect 19024 22148 19030 22160
rect 19337 22151 19395 22157
rect 19337 22148 19349 22151
rect 19024 22120 19349 22148
rect 19024 22108 19030 22120
rect 19337 22117 19349 22120
rect 19383 22117 19395 22151
rect 19337 22111 19395 22117
rect 23661 22151 23719 22157
rect 23661 22117 23673 22151
rect 23707 22148 23719 22151
rect 26234 22148 26240 22160
rect 23707 22120 23741 22148
rect 24688 22120 26240 22148
rect 23707 22117 23719 22120
rect 23661 22111 23719 22117
rect 20622 22080 20628 22092
rect 17603 22052 18460 22080
rect 18708 22052 20628 22080
rect 16942 22012 16948 22024
rect 16592 21984 16948 22012
rect 16942 21972 16948 21984
rect 17000 22012 17006 22024
rect 17603 22012 17631 22052
rect 17000 21984 17631 22012
rect 17000 21972 17006 21984
rect 17954 21972 17960 22024
rect 18012 21972 18018 22024
rect 18046 21972 18052 22024
rect 18104 21972 18110 22024
rect 18138 21972 18144 22024
rect 18196 22012 18202 22024
rect 18549 22015 18607 22021
rect 18549 22012 18561 22015
rect 18196 21984 18561 22012
rect 18196 21972 18202 21984
rect 18549 21981 18561 21984
rect 18595 21981 18607 22015
rect 18549 21975 18607 21981
rect 13771 21916 15608 21944
rect 15672 21916 16068 21944
rect 13771 21913 13783 21916
rect 13725 21907 13783 21913
rect 13464 21848 13676 21876
rect 13357 21839 13415 21845
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 13872 21848 14105 21876
rect 13872 21836 13878 21848
rect 14093 21845 14105 21848
rect 14139 21845 14151 21879
rect 15580 21876 15608 21916
rect 16298 21904 16304 21956
rect 16356 21944 16362 21956
rect 18708 21953 18736 22052
rect 20622 22040 20628 22052
rect 20680 22040 20686 22092
rect 23676 22080 23704 22111
rect 23753 22083 23811 22089
rect 23753 22080 23765 22083
rect 22848 22052 23765 22080
rect 18782 21972 18788 22024
rect 18840 21972 18846 22024
rect 18969 22015 19027 22021
rect 18969 21981 18981 22015
rect 19015 21981 19027 22015
rect 18969 21975 19027 21981
rect 17497 21947 17555 21953
rect 17497 21944 17509 21947
rect 16356 21916 17509 21944
rect 16356 21904 16362 21916
rect 17497 21913 17509 21916
rect 17543 21913 17555 21947
rect 18693 21947 18751 21953
rect 18693 21944 18705 21947
rect 17497 21907 17555 21913
rect 17696 21916 18705 21944
rect 17696 21876 17724 21916
rect 18693 21913 18705 21916
rect 18739 21913 18751 21947
rect 18693 21907 18751 21913
rect 15580 21848 17724 21876
rect 14093 21839 14151 21845
rect 18598 21836 18604 21888
rect 18656 21876 18662 21888
rect 18984 21876 19012 21975
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19521 22015 19579 22021
rect 19521 22012 19533 22015
rect 19484 21984 19533 22012
rect 19484 21972 19490 21984
rect 19521 21981 19533 21984
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 22002 21904 22008 21956
rect 22060 21944 22066 21956
rect 22848 21944 22876 22052
rect 23753 22049 23765 22052
rect 23799 22049 23811 22083
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 23753 22043 23811 22049
rect 23860 22052 24409 22080
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23385 22015 23443 22021
rect 23385 22012 23397 22015
rect 22980 21984 23397 22012
rect 22980 21972 22986 21984
rect 23385 21981 23397 21984
rect 23431 21981 23443 22015
rect 23385 21975 23443 21981
rect 23661 22015 23719 22021
rect 23661 21981 23673 22015
rect 23707 22012 23719 22015
rect 23860 22012 23888 22052
rect 24397 22049 24409 22052
rect 24443 22049 24455 22083
rect 24397 22043 24455 22049
rect 24578 22040 24584 22092
rect 24636 22080 24642 22092
rect 24688 22080 24716 22120
rect 26234 22108 26240 22120
rect 26292 22108 26298 22160
rect 27338 22148 27344 22160
rect 26620 22120 27344 22148
rect 24636 22052 24716 22080
rect 24780 22052 26096 22080
rect 24636 22040 24642 22052
rect 23707 21984 23888 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 24026 21972 24032 22024
rect 24084 21972 24090 22024
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 24780 22021 24808 22052
rect 24213 22015 24271 22021
rect 24213 22012 24225 22015
rect 24176 21984 24225 22012
rect 24176 21972 24182 21984
rect 24213 21981 24225 21984
rect 24259 21981 24271 22015
rect 24213 21975 24271 21981
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 22060 21916 22876 21944
rect 22060 21904 22066 21916
rect 23842 21904 23848 21956
rect 23900 21944 23906 21956
rect 24044 21944 24072 21972
rect 23900 21916 24072 21944
rect 24688 21944 24716 21975
rect 24854 21972 24860 22024
rect 24912 21972 24918 22024
rect 25038 21972 25044 22024
rect 25096 21972 25102 22024
rect 25317 22015 25375 22021
rect 25317 21981 25329 22015
rect 25363 21981 25375 22015
rect 25317 21975 25375 21981
rect 24946 21944 24952 21956
rect 24688 21916 24952 21944
rect 23900 21904 23906 21916
rect 24946 21904 24952 21916
rect 25004 21904 25010 21956
rect 18656 21848 19012 21876
rect 18656 21836 18662 21848
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 20070 21876 20076 21888
rect 19392 21848 20076 21876
rect 19392 21836 19398 21848
rect 20070 21836 20076 21848
rect 20128 21876 20134 21888
rect 20254 21876 20260 21888
rect 20128 21848 20260 21876
rect 20128 21836 20134 21848
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 23477 21879 23535 21885
rect 23477 21845 23489 21879
rect 23523 21876 23535 21879
rect 23566 21876 23572 21888
rect 23523 21848 23572 21876
rect 23523 21845 23535 21848
rect 23477 21839 23535 21845
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 24026 21836 24032 21888
rect 24084 21836 24090 21888
rect 24121 21879 24179 21885
rect 24121 21845 24133 21879
rect 24167 21876 24179 21879
rect 24302 21876 24308 21888
rect 24167 21848 24308 21876
rect 24167 21845 24179 21848
rect 24121 21839 24179 21845
rect 24302 21836 24308 21848
rect 24360 21836 24366 21888
rect 24394 21836 24400 21888
rect 24452 21876 24458 21888
rect 25332 21876 25360 21975
rect 25682 21972 25688 22024
rect 25740 21972 25746 22024
rect 26068 22012 26096 22052
rect 26142 22040 26148 22092
rect 26200 22040 26206 22092
rect 26620 22080 26648 22120
rect 27338 22108 27344 22120
rect 27396 22148 27402 22160
rect 30024 22148 30052 22176
rect 27396 22120 30052 22148
rect 27396 22108 27402 22120
rect 30190 22108 30196 22160
rect 30248 22148 30254 22160
rect 30852 22148 30880 22179
rect 31110 22176 31116 22188
rect 31168 22176 31174 22228
rect 32214 22176 32220 22228
rect 32272 22216 32278 22228
rect 32766 22216 32772 22228
rect 32272 22188 32772 22216
rect 32272 22176 32278 22188
rect 32766 22176 32772 22188
rect 32824 22176 32830 22228
rect 33134 22176 33140 22228
rect 33192 22216 33198 22228
rect 36170 22216 36176 22228
rect 33192 22188 36176 22216
rect 33192 22176 33198 22188
rect 36170 22176 36176 22188
rect 36228 22176 36234 22228
rect 30248 22120 30880 22148
rect 30248 22108 30254 22120
rect 26344 22052 26648 22080
rect 26344 22012 26372 22052
rect 26878 22040 26884 22092
rect 26936 22040 26942 22092
rect 26988 22052 30796 22080
rect 26068 21984 26372 22012
rect 26421 22015 26479 22021
rect 26421 21981 26433 22015
rect 26467 21981 26479 22015
rect 26421 21975 26479 21981
rect 26436 21944 26464 21975
rect 26510 21972 26516 22024
rect 26568 21972 26574 22024
rect 26602 21972 26608 22024
rect 26660 21972 26666 22024
rect 26789 22015 26847 22021
rect 26789 21981 26801 22015
rect 26835 22012 26847 22015
rect 26988 22012 27016 22052
rect 26835 21984 27016 22012
rect 27065 22015 27123 22021
rect 26835 21981 26847 21984
rect 26789 21975 26847 21981
rect 27065 21981 27077 22015
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 26878 21944 26884 21956
rect 26436 21916 26884 21944
rect 26878 21904 26884 21916
rect 26936 21944 26942 21956
rect 27080 21944 27108 21975
rect 27154 21972 27160 22024
rect 27212 21972 27218 22024
rect 27525 22015 27583 22021
rect 27525 21981 27537 22015
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27540 21944 27568 21975
rect 27614 21972 27620 22024
rect 27672 22012 27678 22024
rect 28718 22012 28724 22024
rect 27672 21984 28724 22012
rect 27672 21972 27678 21984
rect 28718 21972 28724 21984
rect 28776 22012 28782 22024
rect 30190 22012 30196 22024
rect 28776 21984 30196 22012
rect 28776 21972 28782 21984
rect 30190 21972 30196 21984
rect 30248 21972 30254 22024
rect 26936 21916 27568 21944
rect 26936 21904 26942 21916
rect 29362 21904 29368 21956
rect 29420 21944 29426 21956
rect 29733 21947 29791 21953
rect 29733 21944 29745 21947
rect 29420 21916 29745 21944
rect 29420 21904 29426 21916
rect 29733 21913 29745 21916
rect 29779 21913 29791 21947
rect 29733 21907 29791 21913
rect 30558 21904 30564 21956
rect 30616 21944 30622 21956
rect 30653 21947 30711 21953
rect 30653 21944 30665 21947
rect 30616 21916 30665 21944
rect 30616 21904 30622 21916
rect 30653 21913 30665 21916
rect 30699 21913 30711 21947
rect 30768 21944 30796 22052
rect 30834 22040 30840 22092
rect 30892 22080 30898 22092
rect 34606 22080 34612 22092
rect 30892 22052 34612 22080
rect 30892 22040 30898 22052
rect 34606 22040 34612 22052
rect 34664 22040 34670 22092
rect 30926 21972 30932 22024
rect 30984 22012 30990 22024
rect 31202 22012 31208 22024
rect 30984 21984 31208 22012
rect 30984 21972 30990 21984
rect 31202 21972 31208 21984
rect 31260 21972 31266 22024
rect 32030 21972 32036 22024
rect 32088 22012 32094 22024
rect 35986 22012 35992 22024
rect 32088 21984 35992 22012
rect 32088 21972 32094 21984
rect 35986 21972 35992 21984
rect 36044 21972 36050 22024
rect 32048 21944 32076 21972
rect 30768 21916 32076 21944
rect 30653 21907 30711 21913
rect 24452 21848 25360 21876
rect 24452 21836 24458 21848
rect 26050 21836 26056 21888
rect 26108 21876 26114 21888
rect 26602 21876 26608 21888
rect 26108 21848 26608 21876
rect 26108 21836 26114 21848
rect 26602 21836 26608 21848
rect 26660 21836 26666 21888
rect 26786 21836 26792 21888
rect 26844 21876 26850 21888
rect 27341 21879 27399 21885
rect 27341 21876 27353 21879
rect 26844 21848 27353 21876
rect 26844 21836 26850 21848
rect 27341 21845 27353 21848
rect 27387 21845 27399 21879
rect 27341 21839 27399 21845
rect 28166 21836 28172 21888
rect 28224 21876 28230 21888
rect 28350 21876 28356 21888
rect 28224 21848 28356 21876
rect 28224 21836 28230 21848
rect 28350 21836 28356 21848
rect 28408 21836 28414 21888
rect 28994 21836 29000 21888
rect 29052 21876 29058 21888
rect 29914 21876 29920 21888
rect 29972 21885 29978 21888
rect 29972 21879 29991 21885
rect 29052 21848 29920 21876
rect 29052 21836 29058 21848
rect 29914 21836 29920 21848
rect 29979 21876 29991 21879
rect 30282 21876 30288 21888
rect 29979 21848 30288 21876
rect 29979 21845 29991 21848
rect 29972 21839 29991 21845
rect 29972 21836 29978 21839
rect 30282 21836 30288 21848
rect 30340 21876 30346 21888
rect 30853 21879 30911 21885
rect 30853 21876 30865 21879
rect 30340 21848 30865 21876
rect 30340 21836 30346 21848
rect 30853 21845 30865 21848
rect 30899 21876 30911 21879
rect 31110 21876 31116 21888
rect 30899 21848 31116 21876
rect 30899 21845 30911 21848
rect 30853 21839 30911 21845
rect 31110 21836 31116 21848
rect 31168 21836 31174 21888
rect 1104 21786 36524 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 36524 21786
rect 1104 21712 36524 21734
rect 3786 21672 3792 21684
rect 1780 21644 3792 21672
rect 1780 21613 1808 21644
rect 3786 21632 3792 21644
rect 3844 21632 3850 21684
rect 4430 21632 4436 21684
rect 4488 21632 4494 21684
rect 4614 21632 4620 21684
rect 4672 21672 4678 21684
rect 6362 21672 6368 21684
rect 4672 21644 6368 21672
rect 4672 21632 4678 21644
rect 6362 21632 6368 21644
rect 6420 21632 6426 21684
rect 7926 21632 7932 21684
rect 7984 21672 7990 21684
rect 9766 21672 9772 21684
rect 7984 21644 9772 21672
rect 7984 21632 7990 21644
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 10686 21632 10692 21684
rect 10744 21672 10750 21684
rect 12066 21672 12072 21684
rect 10744 21644 12072 21672
rect 10744 21632 10750 21644
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 12250 21632 12256 21684
rect 12308 21632 12314 21684
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 15565 21675 15623 21681
rect 15565 21672 15577 21675
rect 14424 21644 15577 21672
rect 14424 21632 14430 21644
rect 15565 21641 15577 21644
rect 15611 21641 15623 21675
rect 15565 21635 15623 21641
rect 15838 21632 15844 21684
rect 15896 21672 15902 21684
rect 16482 21672 16488 21684
rect 15896 21644 16488 21672
rect 15896 21632 15902 21644
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 17313 21675 17371 21681
rect 17313 21641 17325 21675
rect 17359 21672 17371 21675
rect 19426 21672 19432 21684
rect 17359 21644 19432 21672
rect 17359 21641 17371 21644
rect 17313 21635 17371 21641
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 19521 21675 19579 21681
rect 19521 21641 19533 21675
rect 19567 21672 19579 21675
rect 19610 21672 19616 21684
rect 19567 21644 19616 21672
rect 19567 21641 19579 21644
rect 19521 21635 19579 21641
rect 19610 21632 19616 21644
rect 19668 21632 19674 21684
rect 20533 21675 20591 21681
rect 20533 21641 20545 21675
rect 20579 21672 20591 21675
rect 20714 21672 20720 21684
rect 20579 21644 20720 21672
rect 20579 21641 20591 21644
rect 20533 21635 20591 21641
rect 20714 21632 20720 21644
rect 20772 21632 20778 21684
rect 21818 21632 21824 21684
rect 21876 21632 21882 21684
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 22573 21675 22631 21681
rect 22573 21672 22585 21675
rect 22336 21644 22585 21672
rect 22336 21632 22342 21644
rect 22573 21641 22585 21644
rect 22619 21641 22631 21675
rect 22573 21635 22631 21641
rect 22738 21632 22744 21684
rect 22796 21632 22802 21684
rect 24213 21675 24271 21681
rect 24213 21641 24225 21675
rect 24259 21672 24271 21675
rect 24486 21672 24492 21684
rect 24259 21644 24492 21672
rect 24259 21641 24271 21644
rect 24213 21635 24271 21641
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 25025 21675 25083 21681
rect 25025 21672 25037 21675
rect 24964 21644 25037 21672
rect 1765 21607 1823 21613
rect 1765 21573 1777 21607
rect 1811 21573 1823 21607
rect 5258 21604 5264 21616
rect 1765 21567 1823 21573
rect 3896 21576 5264 21604
rect 1394 21496 1400 21548
rect 1452 21536 1458 21548
rect 3896 21545 3924 21576
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 9122 21604 9128 21616
rect 7944 21576 9128 21604
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 1452 21508 1501 21536
rect 1452 21496 1458 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 3881 21539 3939 21545
rect 3881 21536 3893 21539
rect 2898 21508 3004 21536
rect 1489 21499 1547 21505
rect 2976 21480 3004 21508
rect 3252 21508 3893 21536
rect 2958 21428 2964 21480
rect 3016 21428 3022 21480
rect 3252 21477 3280 21508
rect 3881 21505 3893 21508
rect 3927 21505 3939 21539
rect 3881 21499 3939 21505
rect 4522 21496 4528 21548
rect 4580 21496 4586 21548
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 4893 21539 4951 21545
rect 4893 21505 4905 21539
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 5077 21539 5135 21545
rect 5077 21505 5089 21539
rect 5123 21536 5135 21539
rect 5169 21539 5227 21545
rect 5169 21536 5181 21539
rect 5123 21508 5181 21536
rect 5123 21505 5135 21508
rect 5077 21499 5135 21505
rect 5169 21505 5181 21508
rect 5215 21505 5227 21539
rect 5169 21499 5227 21505
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21536 5411 21539
rect 5534 21536 5540 21548
rect 5399 21508 5540 21536
rect 5399 21505 5411 21508
rect 5353 21499 5411 21505
rect 3237 21471 3295 21477
rect 3237 21437 3249 21471
rect 3283 21437 3295 21471
rect 3237 21431 3295 21437
rect 3326 21428 3332 21480
rect 3384 21468 3390 21480
rect 4816 21468 4844 21499
rect 3384 21440 4844 21468
rect 3384 21428 3390 21440
rect 3878 21360 3884 21412
rect 3936 21400 3942 21412
rect 4908 21400 4936 21499
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 5626 21496 5632 21548
rect 5684 21536 5690 21548
rect 7098 21536 7104 21548
rect 5684 21508 7104 21536
rect 5684 21496 5690 21508
rect 7098 21496 7104 21508
rect 7156 21536 7162 21548
rect 7944 21545 7972 21576
rect 9122 21564 9128 21576
rect 9180 21564 9186 21616
rect 9950 21604 9956 21616
rect 9784 21576 9956 21604
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7156 21508 7941 21536
rect 7156 21496 7162 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 8294 21496 8300 21548
rect 8352 21536 8358 21548
rect 8481 21539 8539 21545
rect 8481 21536 8493 21539
rect 8352 21508 8493 21536
rect 8352 21496 8358 21508
rect 8481 21505 8493 21508
rect 8527 21505 8539 21539
rect 8481 21499 8539 21505
rect 8754 21496 8760 21548
rect 8812 21496 8818 21548
rect 9214 21496 9220 21548
rect 9272 21496 9278 21548
rect 9306 21496 9312 21548
rect 9364 21536 9370 21548
rect 9539 21539 9597 21545
rect 9539 21536 9551 21539
rect 9364 21508 9551 21536
rect 9364 21496 9370 21508
rect 9539 21505 9551 21508
rect 9585 21505 9597 21539
rect 9539 21499 9597 21505
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21468 5319 21471
rect 9784 21468 9812 21576
rect 9950 21564 9956 21576
rect 10008 21564 10014 21616
rect 10870 21604 10876 21616
rect 10704 21576 10876 21604
rect 9861 21539 9919 21545
rect 9861 21505 9873 21539
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 5307 21440 9812 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 6638 21400 6644 21412
rect 3936 21372 6644 21400
rect 3936 21360 3942 21372
rect 6638 21360 6644 21372
rect 6696 21400 6702 21412
rect 9309 21403 9367 21409
rect 9309 21400 9321 21403
rect 6696 21372 9321 21400
rect 6696 21360 6702 21372
rect 9309 21369 9321 21372
rect 9355 21369 9367 21403
rect 9309 21363 9367 21369
rect 9582 21360 9588 21412
rect 9640 21400 9646 21412
rect 9876 21400 9904 21499
rect 9968 21468 9996 21564
rect 10413 21539 10471 21545
rect 10413 21505 10425 21539
rect 10459 21536 10471 21539
rect 10594 21536 10600 21548
rect 10459 21508 10600 21536
rect 10459 21505 10471 21508
rect 10413 21499 10471 21505
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 10704 21545 10732 21576
rect 10870 21564 10876 21576
rect 10928 21604 10934 21616
rect 13725 21607 13783 21613
rect 13725 21604 13737 21607
rect 10928 21576 11192 21604
rect 10928 21564 10934 21576
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 11054 21496 11060 21548
rect 11112 21496 11118 21548
rect 11164 21545 11192 21576
rect 11256 21576 13737 21604
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21505 11207 21539
rect 11149 21499 11207 21505
rect 10505 21471 10563 21477
rect 10505 21468 10517 21471
rect 9968 21440 10517 21468
rect 10505 21437 10517 21440
rect 10551 21437 10563 21471
rect 10612 21468 10640 21496
rect 11256 21468 11284 21576
rect 13725 21573 13737 21576
rect 13771 21573 13783 21607
rect 16942 21604 16948 21616
rect 13725 21567 13783 21573
rect 14384 21576 16948 21604
rect 11330 21545 11336 21546
rect 11327 21499 11336 21545
rect 11330 21494 11336 21499
rect 11388 21494 11394 21546
rect 11885 21539 11943 21545
rect 11885 21505 11897 21539
rect 11931 21536 11943 21539
rect 12158 21536 12164 21548
rect 11931 21508 12164 21536
rect 11931 21505 11943 21508
rect 11885 21499 11943 21505
rect 12158 21496 12164 21508
rect 12216 21496 12222 21548
rect 14001 21539 14059 21545
rect 14001 21505 14013 21539
rect 14047 21536 14059 21539
rect 14090 21536 14096 21548
rect 14047 21508 14096 21536
rect 14047 21505 14059 21508
rect 14001 21499 14059 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 11517 21471 11575 21477
rect 11517 21468 11529 21471
rect 10612 21440 11284 21468
rect 11440 21440 11529 21468
rect 10505 21431 10563 21437
rect 9640 21372 9904 21400
rect 9640 21360 9646 21372
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 10965 21403 11023 21409
rect 10965 21400 10977 21403
rect 10652 21372 10977 21400
rect 10652 21360 10658 21372
rect 10965 21369 10977 21372
rect 11011 21369 11023 21403
rect 10965 21363 11023 21369
rect 11333 21403 11391 21409
rect 11333 21369 11345 21403
rect 11379 21400 11391 21403
rect 11440 21400 11468 21440
rect 11517 21437 11529 21440
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 12066 21428 12072 21480
rect 12124 21428 12130 21480
rect 11379 21372 11468 21400
rect 11379 21369 11391 21372
rect 11333 21363 11391 21369
rect 11606 21360 11612 21412
rect 11664 21360 11670 21412
rect 12176 21400 12204 21496
rect 14384 21480 14412 21576
rect 16942 21564 16948 21576
rect 17000 21564 17006 21616
rect 17034 21564 17040 21616
rect 17092 21564 17098 21616
rect 17402 21564 17408 21616
rect 17460 21604 17466 21616
rect 18417 21607 18475 21613
rect 17460 21576 17632 21604
rect 17460 21564 17466 21576
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 14550 21536 14556 21548
rect 14507 21508 14556 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 14550 21496 14556 21508
rect 14608 21496 14614 21548
rect 14829 21539 14887 21545
rect 14829 21505 14841 21539
rect 14875 21536 14887 21539
rect 15102 21536 15108 21548
rect 14875 21508 15108 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15102 21496 15108 21508
rect 15160 21496 15166 21548
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21536 15623 21539
rect 16206 21536 16212 21548
rect 15611 21508 16212 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 16206 21496 16212 21508
rect 16264 21496 16270 21548
rect 16666 21496 16672 21548
rect 16724 21536 16730 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16724 21508 16865 21536
rect 16724 21496 16730 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 17218 21496 17224 21548
rect 17276 21496 17282 21548
rect 17310 21496 17316 21548
rect 17368 21536 17374 21548
rect 17604 21545 17632 21576
rect 17696 21576 18092 21604
rect 17696 21545 17724 21576
rect 18064 21548 18092 21576
rect 18417 21573 18429 21607
rect 18463 21604 18475 21607
rect 19242 21604 19248 21616
rect 18463 21576 19248 21604
rect 18463 21573 18475 21576
rect 18417 21567 18475 21573
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 19337 21607 19395 21613
rect 19337 21573 19349 21607
rect 19383 21604 19395 21607
rect 20073 21607 20131 21613
rect 19383 21576 19472 21604
rect 19383 21573 19395 21576
rect 19337 21567 19395 21573
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17368 21508 17509 21536
rect 17368 21496 17374 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 17589 21539 17647 21545
rect 17589 21505 17601 21539
rect 17635 21505 17647 21539
rect 17589 21499 17647 21505
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 17957 21539 18015 21545
rect 17957 21536 17969 21539
rect 17920 21508 17969 21536
rect 17920 21496 17926 21508
rect 17957 21505 17969 21508
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18046 21496 18052 21548
rect 18104 21496 18110 21548
rect 18230 21496 18236 21548
rect 18288 21496 18294 21548
rect 18782 21496 18788 21548
rect 18840 21536 18846 21548
rect 19061 21539 19119 21545
rect 18840 21534 19012 21536
rect 19061 21534 19073 21539
rect 18840 21508 19073 21534
rect 18840 21496 18846 21508
rect 18984 21506 19073 21508
rect 19061 21505 19073 21506
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 13078 21428 13084 21480
rect 13136 21468 13142 21480
rect 14366 21468 14372 21480
rect 13136 21440 14372 21468
rect 13136 21428 13142 21440
rect 14366 21428 14372 21440
rect 14424 21428 14430 21480
rect 15286 21428 15292 21480
rect 15344 21428 15350 21480
rect 15473 21471 15531 21477
rect 15473 21437 15485 21471
rect 15519 21468 15531 21471
rect 17773 21471 17831 21477
rect 15519 21440 17448 21468
rect 15519 21437 15531 21440
rect 15473 21431 15531 21437
rect 16298 21400 16304 21412
rect 12176 21372 16304 21400
rect 16298 21360 16304 21372
rect 16356 21360 16362 21412
rect 17034 21360 17040 21412
rect 17092 21400 17098 21412
rect 17310 21400 17316 21412
rect 17092 21372 17316 21400
rect 17092 21360 17098 21372
rect 17310 21360 17316 21372
rect 17368 21360 17374 21412
rect 17420 21400 17448 21440
rect 17773 21437 17785 21471
rect 17819 21468 17831 21471
rect 18414 21468 18420 21480
rect 17819 21440 18420 21468
rect 17819 21437 17831 21440
rect 17773 21431 17831 21437
rect 18414 21428 18420 21440
rect 18472 21428 18478 21480
rect 19245 21471 19303 21477
rect 19245 21437 19257 21471
rect 19291 21468 19303 21471
rect 19444 21468 19472 21576
rect 20073 21573 20085 21607
rect 20119 21604 20131 21607
rect 20625 21607 20683 21613
rect 20625 21604 20637 21607
rect 20119 21576 20637 21604
rect 20119 21573 20131 21576
rect 20073 21567 20131 21573
rect 20548 21548 20576 21576
rect 20625 21573 20637 21576
rect 20671 21573 20683 21607
rect 20625 21567 20683 21573
rect 21266 21564 21272 21616
rect 21324 21604 21330 21616
rect 21973 21607 22031 21613
rect 21973 21604 21985 21607
rect 21324 21576 21985 21604
rect 21324 21564 21330 21576
rect 21973 21573 21985 21576
rect 22019 21573 22031 21607
rect 21973 21567 22031 21573
rect 22186 21564 22192 21616
rect 22244 21564 22250 21616
rect 22373 21607 22431 21613
rect 22373 21573 22385 21607
rect 22419 21604 22431 21607
rect 22419 21576 22600 21604
rect 22419 21573 22431 21576
rect 22373 21567 22431 21573
rect 22572 21548 22600 21576
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 23842 21604 23848 21616
rect 23624 21576 23848 21604
rect 23624 21564 23630 21576
rect 23842 21564 23848 21576
rect 23900 21564 23906 21616
rect 24964 21604 24992 21644
rect 25025 21641 25037 21644
rect 25071 21672 25083 21675
rect 25590 21672 25596 21684
rect 25071 21644 25596 21672
rect 25071 21641 25083 21644
rect 25025 21635 25083 21641
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 28626 21672 28632 21684
rect 28552 21644 28632 21672
rect 24136 21576 24992 21604
rect 25225 21607 25283 21613
rect 20346 21496 20352 21548
rect 20404 21496 20410 21548
rect 20530 21496 20536 21548
rect 20588 21496 20594 21548
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21536 20959 21539
rect 20990 21536 20996 21548
rect 20947 21508 20996 21536
rect 20947 21505 20959 21508
rect 20901 21499 20959 21505
rect 20990 21496 20996 21508
rect 21048 21496 21054 21548
rect 22554 21496 22560 21548
rect 22612 21496 22618 21548
rect 24136 21545 24164 21576
rect 25225 21573 25237 21607
rect 25271 21604 25283 21607
rect 25271 21576 26556 21604
rect 25271 21573 25283 21576
rect 25225 21567 25283 21573
rect 24121 21539 24179 21545
rect 24121 21505 24133 21539
rect 24167 21536 24179 21539
rect 24210 21536 24216 21548
rect 24167 21508 24216 21536
rect 24167 21505 24179 21508
rect 24121 21499 24179 21505
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 24302 21496 24308 21548
rect 24360 21496 24366 21548
rect 24581 21539 24639 21545
rect 24581 21505 24593 21539
rect 24627 21536 24639 21539
rect 24670 21536 24676 21548
rect 24627 21508 24676 21536
rect 24627 21505 24639 21508
rect 24581 21499 24639 21505
rect 24670 21496 24676 21508
rect 24728 21536 24734 21548
rect 25240 21536 25268 21567
rect 24728 21508 25268 21536
rect 24728 21496 24734 21508
rect 19518 21468 19524 21480
rect 19291 21440 19524 21468
rect 19291 21437 19303 21440
rect 19245 21431 19303 21437
rect 19518 21428 19524 21440
rect 19576 21428 19582 21480
rect 20165 21471 20223 21477
rect 20165 21437 20177 21471
rect 20211 21468 20223 21471
rect 20211 21440 20245 21468
rect 20211 21437 20223 21440
rect 20165 21431 20223 21437
rect 18877 21403 18935 21409
rect 18877 21400 18889 21403
rect 17420 21372 18889 21400
rect 18877 21369 18889 21372
rect 18923 21400 18935 21403
rect 19705 21403 19763 21409
rect 18923 21372 19656 21400
rect 18923 21369 18935 21372
rect 18877 21363 18935 21369
rect 10226 21292 10232 21344
rect 10284 21332 10290 21344
rect 14918 21332 14924 21344
rect 10284 21304 14924 21332
rect 10284 21292 10290 21304
rect 14918 21292 14924 21304
rect 14976 21292 14982 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 15712 21304 16681 21332
rect 15712 21292 15718 21304
rect 16669 21301 16681 21304
rect 16715 21301 16727 21335
rect 16669 21295 16727 21301
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 18322 21332 18328 21344
rect 17000 21304 18328 21332
rect 17000 21292 17006 21304
rect 18322 21292 18328 21304
rect 18380 21292 18386 21344
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 19150 21332 19156 21344
rect 18840 21304 19156 21332
rect 18840 21292 18846 21304
rect 19150 21292 19156 21304
rect 19208 21292 19214 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19484 21304 19533 21332
rect 19484 21292 19490 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19628 21332 19656 21372
rect 19705 21369 19717 21403
rect 19751 21400 19763 21403
rect 20180 21400 20208 21431
rect 19751 21372 20208 21400
rect 20364 21400 20392 21496
rect 20438 21428 20444 21480
rect 20496 21468 20502 21480
rect 20717 21471 20775 21477
rect 20717 21468 20729 21471
rect 20496 21440 20729 21468
rect 20496 21428 20502 21440
rect 20717 21437 20729 21440
rect 20763 21437 20775 21471
rect 20717 21431 20775 21437
rect 21008 21440 23799 21468
rect 21008 21400 21036 21440
rect 20364 21372 21036 21400
rect 21085 21403 21143 21409
rect 19751 21369 19763 21372
rect 19705 21363 19763 21369
rect 20073 21335 20131 21341
rect 20073 21332 20085 21335
rect 19628 21304 20085 21332
rect 19521 21295 19579 21301
rect 20073 21301 20085 21304
rect 20119 21301 20131 21335
rect 20180 21332 20208 21372
rect 21085 21369 21097 21403
rect 21131 21400 21143 21403
rect 23106 21400 23112 21412
rect 21131 21372 23112 21400
rect 21131 21369 21143 21372
rect 21085 21363 21143 21369
rect 23106 21360 23112 21372
rect 23164 21360 23170 21412
rect 23771 21400 23799 21440
rect 23842 21428 23848 21480
rect 23900 21428 23906 21480
rect 25222 21400 25228 21412
rect 23771 21372 25228 21400
rect 20346 21332 20352 21344
rect 20180 21304 20352 21332
rect 20073 21295 20131 21301
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 20438 21292 20444 21344
rect 20496 21332 20502 21344
rect 20622 21332 20628 21344
rect 20496 21304 20628 21332
rect 20496 21292 20502 21304
rect 20622 21292 20628 21304
rect 20680 21332 20686 21344
rect 20717 21335 20775 21341
rect 20717 21332 20729 21335
rect 20680 21304 20729 21332
rect 20680 21292 20686 21304
rect 20717 21301 20729 21304
rect 20763 21301 20775 21335
rect 20717 21295 20775 21301
rect 22005 21335 22063 21341
rect 22005 21301 22017 21335
rect 22051 21332 22063 21335
rect 22557 21335 22615 21341
rect 22557 21332 22569 21335
rect 22051 21304 22569 21332
rect 22051 21301 22063 21304
rect 22005 21295 22063 21301
rect 22557 21301 22569 21304
rect 22603 21332 22615 21335
rect 24026 21332 24032 21344
rect 22603 21304 24032 21332
rect 22603 21301 22615 21304
rect 22557 21295 22615 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24486 21292 24492 21344
rect 24544 21292 24550 21344
rect 24857 21335 24915 21341
rect 24857 21301 24869 21335
rect 24903 21332 24915 21335
rect 24946 21332 24952 21344
rect 24903 21304 24952 21332
rect 24903 21301 24915 21304
rect 24857 21295 24915 21301
rect 24946 21292 24952 21304
rect 25004 21292 25010 21344
rect 25056 21341 25084 21372
rect 25222 21360 25228 21372
rect 25280 21360 25286 21412
rect 26528 21400 26556 21576
rect 27338 21564 27344 21616
rect 27396 21564 27402 21616
rect 28074 21564 28080 21616
rect 28132 21604 28138 21616
rect 28552 21613 28580 21644
rect 28626 21632 28632 21644
rect 28684 21672 28690 21684
rect 28684 21644 28994 21672
rect 28684 21632 28690 21644
rect 28307 21607 28365 21613
rect 28307 21604 28319 21607
rect 28132 21576 28319 21604
rect 28132 21564 28138 21576
rect 28307 21573 28319 21576
rect 28353 21573 28365 21607
rect 28307 21567 28365 21573
rect 28537 21607 28595 21613
rect 28537 21573 28549 21607
rect 28583 21573 28595 21607
rect 28966 21604 28994 21644
rect 30282 21632 30288 21684
rect 30340 21672 30346 21684
rect 31754 21672 31760 21684
rect 30340 21644 31760 21672
rect 30340 21632 30346 21644
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 30558 21604 30564 21616
rect 28966 21576 30564 21604
rect 28537 21567 28595 21573
rect 30558 21564 30564 21576
rect 30616 21564 30622 21616
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21536 27215 21539
rect 27356 21536 27384 21564
rect 27203 21508 27384 21536
rect 27203 21505 27215 21508
rect 27157 21499 27215 21505
rect 28166 21496 28172 21548
rect 28224 21496 28230 21548
rect 28445 21539 28503 21545
rect 28445 21505 28457 21539
rect 28491 21505 28503 21539
rect 28445 21499 28503 21505
rect 28629 21539 28687 21545
rect 28629 21505 28641 21539
rect 28675 21536 28687 21539
rect 28994 21536 29000 21548
rect 28675 21508 29000 21536
rect 28675 21505 28687 21508
rect 28629 21499 28687 21505
rect 27246 21428 27252 21480
rect 27304 21468 27310 21480
rect 27341 21471 27399 21477
rect 27341 21468 27353 21471
rect 27304 21440 27353 21468
rect 27304 21428 27310 21440
rect 27341 21437 27353 21440
rect 27387 21468 27399 21471
rect 27430 21468 27436 21480
rect 27387 21440 27436 21468
rect 27387 21437 27399 21440
rect 27341 21431 27399 21437
rect 27430 21428 27436 21440
rect 27488 21468 27494 21480
rect 28460 21468 28488 21499
rect 28994 21496 29000 21508
rect 29052 21496 29058 21548
rect 29178 21496 29184 21548
rect 29236 21536 29242 21548
rect 29914 21536 29920 21548
rect 29236 21508 29920 21536
rect 29236 21496 29242 21508
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 35526 21536 35532 21548
rect 30024 21508 35532 21536
rect 30024 21468 30052 21508
rect 35526 21496 35532 21508
rect 35584 21496 35590 21548
rect 27488 21440 28488 21468
rect 28966 21440 30052 21468
rect 27488 21428 27494 21440
rect 28966 21400 28994 21440
rect 30650 21428 30656 21480
rect 30708 21468 30714 21480
rect 31386 21468 31392 21480
rect 30708 21440 31392 21468
rect 30708 21428 30714 21440
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 26528 21372 28994 21400
rect 29546 21360 29552 21412
rect 29604 21400 29610 21412
rect 30834 21400 30840 21412
rect 29604 21372 30840 21400
rect 29604 21360 29610 21372
rect 30834 21360 30840 21372
rect 30892 21360 30898 21412
rect 31018 21360 31024 21412
rect 31076 21400 31082 21412
rect 31294 21400 31300 21412
rect 31076 21372 31300 21400
rect 31076 21360 31082 21372
rect 31294 21360 31300 21372
rect 31352 21400 31358 21412
rect 33410 21400 33416 21412
rect 31352 21372 33416 21400
rect 31352 21360 31358 21372
rect 33410 21360 33416 21372
rect 33468 21360 33474 21412
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21301 25099 21335
rect 25041 21295 25099 21301
rect 26970 21292 26976 21344
rect 27028 21292 27034 21344
rect 28813 21335 28871 21341
rect 28813 21301 28825 21335
rect 28859 21332 28871 21335
rect 31110 21332 31116 21344
rect 28859 21304 31116 21332
rect 28859 21301 28871 21304
rect 28813 21295 28871 21301
rect 31110 21292 31116 21304
rect 31168 21292 31174 21344
rect 32030 21292 32036 21344
rect 32088 21332 32094 21344
rect 32858 21332 32864 21344
rect 32088 21304 32864 21332
rect 32088 21292 32094 21304
rect 32858 21292 32864 21304
rect 32916 21292 32922 21344
rect 35342 21292 35348 21344
rect 35400 21332 35406 21344
rect 35710 21332 35716 21344
rect 35400 21304 35716 21332
rect 35400 21292 35406 21304
rect 35710 21292 35716 21304
rect 35768 21292 35774 21344
rect 1104 21242 36524 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 36524 21242
rect 1104 21168 36524 21190
rect 5718 21088 5724 21140
rect 5776 21088 5782 21140
rect 7006 21088 7012 21140
rect 7064 21128 7070 21140
rect 7466 21128 7472 21140
rect 7064 21100 7472 21128
rect 7064 21088 7070 21100
rect 7466 21088 7472 21100
rect 7524 21128 7530 21140
rect 7524 21100 7880 21128
rect 7524 21088 7530 21100
rect 4890 21060 4896 21072
rect 4816 21032 4896 21060
rect 3145 20995 3203 21001
rect 3145 20961 3157 20995
rect 3191 20992 3203 20995
rect 4062 20992 4068 21004
rect 3191 20964 4068 20992
rect 3191 20961 3203 20964
rect 3145 20955 3203 20961
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 2866 20884 2872 20936
rect 2924 20924 2930 20936
rect 2924 20896 3004 20924
rect 2924 20884 2930 20896
rect 1670 20748 1676 20800
rect 1728 20788 1734 20800
rect 2501 20791 2559 20797
rect 2501 20788 2513 20791
rect 1728 20760 2513 20788
rect 1728 20748 1734 20760
rect 2501 20757 2513 20760
rect 2547 20757 2559 20791
rect 2501 20751 2559 20757
rect 2866 20748 2872 20800
rect 2924 20748 2930 20800
rect 2976 20797 3004 20896
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 4525 20927 4583 20933
rect 4525 20893 4537 20927
rect 4571 20924 4583 20927
rect 4614 20924 4620 20936
rect 4571 20896 4620 20924
rect 4571 20893 4583 20896
rect 4525 20887 4583 20893
rect 4614 20884 4620 20896
rect 4672 20884 4678 20936
rect 4706 20884 4712 20936
rect 4764 20884 4770 20936
rect 4816 20933 4844 21032
rect 4890 21020 4896 21032
rect 4948 21060 4954 21072
rect 6546 21060 6552 21072
rect 4948 21032 6552 21060
rect 4948 21020 4954 21032
rect 6546 21020 6552 21032
rect 6604 21020 6610 21072
rect 7116 21032 7788 21060
rect 7116 21001 7144 21032
rect 7760 21004 7788 21032
rect 7101 20995 7159 21001
rect 5461 20964 5856 20992
rect 4801 20927 4859 20933
rect 4801 20893 4813 20927
rect 4847 20893 4859 20927
rect 4801 20887 4859 20893
rect 4893 20927 4951 20933
rect 4893 20893 4905 20927
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 4908 20856 4936 20887
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5461 20924 5489 20964
rect 5828 20936 5856 20964
rect 7101 20961 7113 20995
rect 7147 20961 7159 20995
rect 7101 20955 7159 20961
rect 7285 20995 7343 21001
rect 7285 20961 7297 20995
rect 7331 20992 7343 20995
rect 7374 20992 7380 21004
rect 7331 20964 7380 20992
rect 7331 20961 7343 20964
rect 7285 20955 7343 20961
rect 7374 20952 7380 20964
rect 7432 20992 7438 21004
rect 7432 20964 7604 20992
rect 7432 20952 7438 20964
rect 5534 20924 5540 20936
rect 5461 20896 5540 20924
rect 5534 20884 5540 20896
rect 5592 20884 5598 20936
rect 5626 20884 5632 20936
rect 5684 20884 5690 20936
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 7006 20884 7012 20936
rect 7064 20884 7070 20936
rect 7190 20884 7196 20936
rect 7248 20884 7254 20936
rect 7576 20933 7604 20964
rect 7742 20952 7748 21004
rect 7800 20952 7806 21004
rect 7561 20927 7619 20933
rect 7561 20893 7573 20927
rect 7607 20893 7619 20927
rect 7852 20924 7880 21100
rect 8018 21088 8024 21140
rect 8076 21128 8082 21140
rect 10502 21128 10508 21140
rect 8076 21100 10508 21128
rect 8076 21088 8082 21100
rect 10502 21088 10508 21100
rect 10560 21088 10566 21140
rect 11054 21088 11060 21140
rect 11112 21128 11118 21140
rect 11606 21128 11612 21140
rect 11112 21100 11612 21128
rect 11112 21088 11118 21100
rect 11606 21088 11612 21100
rect 11664 21088 11670 21140
rect 13173 21131 13231 21137
rect 13173 21097 13185 21131
rect 13219 21128 13231 21131
rect 13354 21128 13360 21140
rect 13219 21100 13360 21128
rect 13219 21097 13231 21100
rect 13173 21091 13231 21097
rect 13354 21088 13360 21100
rect 13412 21088 13418 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 15657 21131 15715 21137
rect 15657 21128 15669 21131
rect 15620 21100 15669 21128
rect 15620 21088 15626 21100
rect 15657 21097 15669 21100
rect 15703 21097 15715 21131
rect 17770 21128 17776 21140
rect 15657 21091 15715 21097
rect 15764 21100 17776 21128
rect 7929 21063 7987 21069
rect 7929 21029 7941 21063
rect 7975 21060 7987 21063
rect 7975 21032 11468 21060
rect 7975 21029 7987 21032
rect 7929 21023 7987 21029
rect 8294 20952 8300 21004
rect 8352 20992 8358 21004
rect 8481 20995 8539 21001
rect 8481 20992 8493 20995
rect 8352 20964 8493 20992
rect 8352 20952 8358 20964
rect 8481 20961 8493 20964
rect 8527 20961 8539 20995
rect 8481 20955 8539 20961
rect 8665 20995 8723 21001
rect 8665 20961 8677 20995
rect 8711 20992 8723 20995
rect 8754 20992 8760 21004
rect 8711 20964 8760 20992
rect 8711 20961 8723 20964
rect 8665 20955 8723 20961
rect 8754 20952 8760 20964
rect 8812 20952 8818 21004
rect 9030 20992 9036 21004
rect 8864 20964 9036 20992
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7852 20896 7941 20924
rect 7561 20887 7619 20893
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 8864 20924 8892 20964
rect 9030 20952 9036 20964
rect 9088 20952 9094 21004
rect 10226 20952 10232 21004
rect 10284 20952 10290 21004
rect 10502 20952 10508 21004
rect 10560 20992 10566 21004
rect 10597 20995 10655 21001
rect 10597 20992 10609 20995
rect 10560 20964 10609 20992
rect 10560 20952 10566 20964
rect 10597 20961 10609 20964
rect 10643 20961 10655 20995
rect 10597 20955 10655 20961
rect 11146 20952 11152 21004
rect 11204 20952 11210 21004
rect 11440 21001 11468 21032
rect 11514 21020 11520 21072
rect 11572 21060 11578 21072
rect 11885 21063 11943 21069
rect 11885 21060 11897 21063
rect 11572 21032 11897 21060
rect 11572 21020 11578 21032
rect 11885 21029 11897 21032
rect 11931 21029 11943 21063
rect 11885 21023 11943 21029
rect 12250 21020 12256 21072
rect 12308 21020 12314 21072
rect 13446 21020 13452 21072
rect 13504 21060 13510 21072
rect 15764 21060 15792 21100
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 17865 21131 17923 21137
rect 17865 21097 17877 21131
rect 17911 21128 17923 21131
rect 18138 21128 18144 21140
rect 17911 21100 18144 21128
rect 17911 21097 17923 21100
rect 17865 21091 17923 21097
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 18322 21088 18328 21140
rect 18380 21088 18386 21140
rect 18693 21131 18751 21137
rect 18693 21097 18705 21131
rect 18739 21128 18751 21131
rect 18874 21128 18880 21140
rect 18739 21100 18880 21128
rect 18739 21097 18751 21100
rect 18693 21091 18751 21097
rect 18874 21088 18880 21100
rect 18932 21088 18938 21140
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 19794 21128 19800 21140
rect 19576 21100 19800 21128
rect 19576 21088 19582 21100
rect 19794 21088 19800 21100
rect 19852 21088 19858 21140
rect 20530 21088 20536 21140
rect 20588 21088 20594 21140
rect 22646 21128 22652 21140
rect 20732 21100 22652 21128
rect 16393 21063 16451 21069
rect 16393 21060 16405 21063
rect 13504 21032 15792 21060
rect 15856 21032 16405 21060
rect 13504 21020 13510 21032
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20961 11483 20995
rect 11425 20955 11483 20961
rect 12161 20995 12219 21001
rect 12161 20961 12173 20995
rect 12207 20992 12219 20995
rect 12268 20992 12296 21020
rect 12207 20964 12296 20992
rect 13081 20995 13139 21001
rect 12207 20961 12219 20964
rect 12161 20955 12219 20961
rect 13081 20961 13093 20995
rect 13127 20992 13139 20995
rect 13998 20992 14004 21004
rect 13127 20964 14004 20992
rect 13127 20961 13139 20964
rect 13081 20955 13139 20961
rect 7929 20887 7987 20893
rect 8286 20896 8892 20924
rect 8941 20927 8999 20933
rect 5902 20856 5908 20868
rect 4908 20828 5908 20856
rect 5902 20816 5908 20828
rect 5960 20816 5966 20868
rect 7208 20856 7236 20884
rect 7653 20859 7711 20865
rect 7653 20856 7665 20859
rect 7208 20828 7665 20856
rect 7653 20825 7665 20828
rect 7699 20825 7711 20859
rect 8286 20856 8314 20896
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9214 20924 9220 20936
rect 8987 20896 9220 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 7653 20819 7711 20825
rect 7944 20828 8314 20856
rect 8389 20859 8447 20865
rect 2961 20791 3019 20797
rect 2961 20757 2973 20791
rect 3007 20788 3019 20791
rect 3510 20788 3516 20800
rect 3007 20760 3516 20788
rect 3007 20757 3019 20760
rect 2961 20751 3019 20757
rect 3510 20748 3516 20760
rect 3568 20748 3574 20800
rect 3786 20748 3792 20800
rect 3844 20748 3850 20800
rect 5077 20791 5135 20797
rect 5077 20757 5089 20791
rect 5123 20788 5135 20791
rect 5258 20788 5264 20800
rect 5123 20760 5264 20788
rect 5123 20757 5135 20760
rect 5077 20751 5135 20757
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 7374 20788 7380 20800
rect 5583 20760 7380 20788
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 7374 20748 7380 20760
rect 7432 20748 7438 20800
rect 7469 20791 7527 20797
rect 7469 20757 7481 20791
rect 7515 20788 7527 20791
rect 7944 20788 7972 20828
rect 8389 20825 8401 20859
rect 8435 20856 8447 20859
rect 8754 20856 8760 20868
rect 8435 20828 8760 20856
rect 8435 20825 8447 20828
rect 8389 20819 8447 20825
rect 8754 20816 8760 20828
rect 8812 20856 8818 20868
rect 8956 20856 8984 20887
rect 9214 20884 9220 20896
rect 9272 20884 9278 20936
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 9858 20924 9864 20936
rect 9723 20896 9864 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 10042 20884 10048 20936
rect 10100 20884 10106 20936
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20924 10839 20927
rect 10870 20924 10876 20936
rect 10827 20896 10876 20924
rect 10827 20893 10839 20896
rect 10781 20887 10839 20893
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20924 11391 20927
rect 11606 20924 11612 20936
rect 11379 20896 11612 20924
rect 11379 20893 11391 20896
rect 11333 20887 11391 20893
rect 11606 20884 11612 20896
rect 11664 20924 11670 20936
rect 12176 20924 12204 20955
rect 13998 20952 14004 20964
rect 14056 20992 14062 21004
rect 14645 20995 14703 21001
rect 14645 20992 14657 20995
rect 14056 20964 14657 20992
rect 14056 20952 14062 20964
rect 14645 20961 14657 20964
rect 14691 20961 14703 20995
rect 14645 20955 14703 20961
rect 11664 20896 12204 20924
rect 12253 20927 12311 20933
rect 11664 20884 11670 20896
rect 12253 20893 12265 20927
rect 12299 20893 12311 20927
rect 12253 20887 12311 20893
rect 12621 20927 12679 20933
rect 12621 20893 12633 20927
rect 12667 20924 12679 20927
rect 12986 20924 12992 20936
rect 12667 20896 12992 20924
rect 12667 20893 12679 20896
rect 12621 20887 12679 20893
rect 8812 20828 8984 20856
rect 8812 20816 8818 20828
rect 10410 20816 10416 20868
rect 10468 20856 10474 20868
rect 12268 20856 12296 20887
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20924 13231 20927
rect 13262 20924 13268 20936
rect 13219 20896 13268 20924
rect 13219 20893 13231 20896
rect 13173 20887 13231 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 13354 20884 13360 20936
rect 13412 20924 13418 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 13412 20896 14473 20924
rect 13412 20884 13418 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 15470 20884 15476 20936
rect 15528 20884 15534 20936
rect 15856 20933 15884 21032
rect 16393 21029 16405 21032
rect 16439 21060 16451 21063
rect 16439 21032 18184 21060
rect 16439 21029 16451 21032
rect 16393 21023 16451 21029
rect 16206 20952 16212 21004
rect 16264 20952 16270 21004
rect 18046 20992 18052 21004
rect 17420 20964 18052 20992
rect 15749 20927 15807 20933
rect 15749 20893 15761 20927
rect 15795 20893 15807 20927
rect 15749 20887 15807 20893
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 10468 20828 12296 20856
rect 12529 20859 12587 20865
rect 10468 20816 10474 20828
rect 12529 20825 12541 20859
rect 12575 20856 12587 20859
rect 13078 20856 13084 20868
rect 12575 20828 13084 20856
rect 12575 20825 12587 20828
rect 12529 20819 12587 20825
rect 13078 20816 13084 20828
rect 13136 20816 13142 20868
rect 14277 20859 14335 20865
rect 14277 20825 14289 20859
rect 14323 20856 14335 20859
rect 14918 20856 14924 20868
rect 14323 20828 14924 20856
rect 14323 20825 14335 20828
rect 14277 20819 14335 20825
rect 14918 20816 14924 20828
rect 14976 20816 14982 20868
rect 15562 20816 15568 20868
rect 15620 20816 15626 20868
rect 15764 20856 15792 20887
rect 16114 20884 16120 20936
rect 16172 20884 16178 20936
rect 16224 20856 16252 20952
rect 17420 20949 17448 20964
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20924 16359 20927
rect 17218 20924 17224 20936
rect 16347 20896 17224 20924
rect 16347 20893 16359 20896
rect 16301 20887 16359 20893
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 17329 20933 17448 20949
rect 18156 20936 18184 21032
rect 18340 20992 18368 21088
rect 18414 21020 18420 21072
rect 18472 21060 18478 21072
rect 20732 21060 20760 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 22741 21131 22799 21137
rect 22741 21097 22753 21131
rect 22787 21128 22799 21131
rect 22830 21128 22836 21140
rect 22787 21100 22836 21128
rect 22787 21097 22799 21100
rect 22741 21091 22799 21097
rect 22830 21088 22836 21100
rect 22888 21088 22894 21140
rect 23385 21131 23443 21137
rect 23385 21097 23397 21131
rect 23431 21128 23443 21131
rect 23474 21128 23480 21140
rect 23431 21100 23480 21128
rect 23431 21097 23443 21100
rect 23385 21091 23443 21097
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 24118 21088 24124 21140
rect 24176 21128 24182 21140
rect 26970 21128 26976 21140
rect 24176 21100 26976 21128
rect 24176 21088 24182 21100
rect 26970 21088 26976 21100
rect 27028 21088 27034 21140
rect 28718 21088 28724 21140
rect 28776 21128 28782 21140
rect 30193 21131 30251 21137
rect 28776 21100 29868 21128
rect 28776 21088 28782 21100
rect 18472 21032 20760 21060
rect 18472 21020 18478 21032
rect 20806 21020 20812 21072
rect 20864 21060 20870 21072
rect 20864 21032 23244 21060
rect 20864 21020 20870 21032
rect 18340 20964 18460 20992
rect 17314 20927 17448 20933
rect 17314 20893 17326 20927
rect 17360 20921 17448 20927
rect 17727 20927 17785 20933
rect 17360 20893 17372 20921
rect 17314 20887 17372 20893
rect 17727 20893 17739 20927
rect 17773 20924 17785 20927
rect 17957 20927 18015 20933
rect 17773 20896 17908 20924
rect 17773 20893 17785 20896
rect 17727 20887 17785 20893
rect 15764 20828 16252 20856
rect 17494 20816 17500 20868
rect 17552 20816 17558 20868
rect 17586 20816 17592 20868
rect 17644 20816 17650 20868
rect 17880 20800 17908 20896
rect 17957 20893 17969 20927
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 17972 20856 18000 20887
rect 18138 20884 18144 20936
rect 18196 20884 18202 20936
rect 18230 20884 18236 20936
rect 18288 20884 18294 20936
rect 18322 20884 18328 20936
rect 18380 20884 18386 20936
rect 18432 20933 18460 20964
rect 19242 20952 19248 21004
rect 19300 20952 19306 21004
rect 20622 20992 20628 21004
rect 19904 20964 20628 20992
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20924 18475 20927
rect 18966 20924 18972 20936
rect 18463 20896 18972 20924
rect 18463 20893 18475 20896
rect 18417 20887 18475 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19518 20884 19524 20936
rect 19576 20884 19582 20936
rect 19610 20884 19616 20936
rect 19668 20884 19674 20936
rect 19702 20884 19708 20936
rect 19760 20884 19766 20936
rect 19904 20933 19932 20964
rect 20622 20952 20628 20964
rect 20680 20952 20686 21004
rect 21634 20992 21640 21004
rect 20824 20964 21640 20992
rect 20070 20933 20076 20936
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 20037 20927 20076 20933
rect 20037 20893 20049 20927
rect 20037 20887 20076 20893
rect 20070 20884 20076 20887
rect 20128 20884 20134 20936
rect 20395 20927 20453 20933
rect 20395 20893 20407 20927
rect 20441 20924 20453 20927
rect 20824 20924 20852 20964
rect 21634 20952 21640 20964
rect 21692 20952 21698 21004
rect 22002 20952 22008 21004
rect 22060 20952 22066 21004
rect 20441 20896 20852 20924
rect 20441 20893 20453 20896
rect 20395 20887 20453 20893
rect 20898 20884 20904 20936
rect 20956 20924 20962 20936
rect 21545 20927 21603 20933
rect 21545 20924 21557 20927
rect 20956 20896 21557 20924
rect 20956 20884 20962 20896
rect 21545 20893 21557 20896
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 21910 20884 21916 20936
rect 21968 20924 21974 20936
rect 22097 20927 22155 20933
rect 22097 20924 22109 20927
rect 21968 20896 22109 20924
rect 21968 20884 21974 20896
rect 22097 20893 22109 20896
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 22370 20884 22376 20936
rect 22428 20924 22434 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22428 20896 22477 20924
rect 22428 20884 22434 20896
rect 22465 20893 22477 20896
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22554 20884 22560 20936
rect 22612 20933 22618 20936
rect 23216 20933 23244 21032
rect 26510 21020 26516 21072
rect 26568 21060 26574 21072
rect 29178 21060 29184 21072
rect 26568 21032 29184 21060
rect 26568 21020 26574 21032
rect 22612 20927 22640 20933
rect 22628 20924 22640 20927
rect 23201 20927 23259 20933
rect 22628 20896 23060 20924
rect 22628 20893 22640 20896
rect 22612 20887 22640 20893
rect 22612 20884 22618 20887
rect 18782 20856 18788 20868
rect 17972 20828 18788 20856
rect 18782 20816 18788 20828
rect 18840 20856 18846 20868
rect 18840 20828 19334 20856
rect 18840 20816 18846 20828
rect 7515 20760 7972 20788
rect 7515 20757 7527 20760
rect 7469 20751 7527 20757
rect 8018 20748 8024 20800
rect 8076 20748 8082 20800
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 9125 20791 9183 20797
rect 9125 20788 9137 20791
rect 8260 20760 9137 20788
rect 8260 20748 8266 20760
rect 9125 20757 9137 20760
rect 9171 20757 9183 20791
rect 9125 20751 9183 20757
rect 9306 20748 9312 20800
rect 9364 20788 9370 20800
rect 9490 20788 9496 20800
rect 9364 20760 9496 20788
rect 9364 20748 9370 20760
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 9582 20748 9588 20800
rect 9640 20788 9646 20800
rect 9861 20791 9919 20797
rect 9861 20788 9873 20791
rect 9640 20760 9873 20788
rect 9640 20748 9646 20760
rect 9861 20757 9873 20760
rect 9907 20757 9919 20791
rect 9861 20751 9919 20757
rect 11057 20791 11115 20797
rect 11057 20757 11069 20791
rect 11103 20788 11115 20791
rect 11146 20788 11152 20800
rect 11103 20760 11152 20788
rect 11103 20757 11115 20760
rect 11057 20751 11115 20757
rect 11146 20748 11152 20760
rect 11204 20748 11210 20800
rect 11425 20791 11483 20797
rect 11425 20757 11437 20791
rect 11471 20788 11483 20791
rect 11790 20788 11796 20800
rect 11471 20760 11796 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 12805 20791 12863 20797
rect 12805 20757 12817 20791
rect 12851 20788 12863 20791
rect 13630 20788 13636 20800
rect 12851 20760 13636 20788
rect 12851 20757 12863 20760
rect 12805 20751 12863 20757
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 14093 20791 14151 20797
rect 14093 20757 14105 20791
rect 14139 20788 14151 20791
rect 14182 20788 14188 20800
rect 14139 20760 14188 20788
rect 14139 20757 14151 20760
rect 14093 20751 14151 20757
rect 14182 20748 14188 20760
rect 14240 20748 14246 20800
rect 14366 20748 14372 20800
rect 14424 20788 14430 20800
rect 14826 20788 14832 20800
rect 14424 20760 14832 20788
rect 14424 20748 14430 20760
rect 14826 20748 14832 20760
rect 14884 20748 14890 20800
rect 15194 20748 15200 20800
rect 15252 20788 15258 20800
rect 15289 20791 15347 20797
rect 15289 20788 15301 20791
rect 15252 20760 15301 20788
rect 15252 20748 15258 20760
rect 15289 20757 15301 20760
rect 15335 20788 15347 20791
rect 15746 20788 15752 20800
rect 15335 20760 15752 20788
rect 15335 20757 15347 20760
rect 15289 20751 15347 20757
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 16022 20748 16028 20800
rect 16080 20748 16086 20800
rect 16390 20748 16396 20800
rect 16448 20748 16454 20800
rect 17862 20748 17868 20800
rect 17920 20748 17926 20800
rect 19306 20788 19334 20828
rect 20162 20816 20168 20868
rect 20220 20816 20226 20868
rect 20257 20859 20315 20865
rect 20257 20825 20269 20859
rect 20303 20856 20315 20859
rect 21174 20856 21180 20868
rect 20303 20828 21180 20856
rect 20303 20825 20315 20828
rect 20257 20819 20315 20825
rect 21174 20816 21180 20828
rect 21232 20816 21238 20868
rect 22833 20859 22891 20865
rect 22833 20825 22845 20859
rect 22879 20825 22891 20859
rect 22833 20819 22891 20825
rect 20346 20788 20352 20800
rect 19306 20760 20352 20788
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 21729 20791 21787 20797
rect 21729 20757 21741 20791
rect 21775 20788 21787 20791
rect 22373 20791 22431 20797
rect 22373 20788 22385 20791
rect 21775 20760 22385 20788
rect 21775 20757 21787 20760
rect 21729 20751 21787 20757
rect 22373 20757 22385 20760
rect 22419 20788 22431 20791
rect 22848 20788 22876 20819
rect 23032 20800 23060 20896
rect 23201 20893 23213 20927
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 27890 20884 27896 20936
rect 27948 20924 27954 20936
rect 28277 20933 28305 21032
rect 29178 21020 29184 21032
rect 29236 21020 29242 21072
rect 28442 20952 28448 21004
rect 28500 20992 28506 21004
rect 28629 20995 28687 21001
rect 28629 20992 28641 20995
rect 28500 20964 28641 20992
rect 28500 20952 28506 20964
rect 28629 20961 28641 20964
rect 28675 20961 28687 20995
rect 28629 20955 28687 20961
rect 28261 20927 28319 20933
rect 28169 20924 28227 20927
rect 27948 20921 28227 20924
rect 27948 20896 28181 20921
rect 27948 20884 27954 20896
rect 28169 20887 28181 20896
rect 28215 20887 28227 20921
rect 28261 20893 28273 20927
rect 28307 20893 28319 20927
rect 28261 20887 28319 20893
rect 28169 20881 28227 20887
rect 28350 20884 28356 20936
rect 28408 20884 28414 20936
rect 28718 20884 28724 20936
rect 28776 20924 28782 20936
rect 28994 20924 29000 20936
rect 28776 20896 29000 20924
rect 28776 20884 28782 20896
rect 28994 20884 29000 20896
rect 29052 20884 29058 20936
rect 29546 20884 29552 20936
rect 29604 20884 29610 20936
rect 29730 20933 29736 20936
rect 29707 20927 29736 20933
rect 29707 20893 29719 20927
rect 29707 20887 29736 20893
rect 29722 20884 29736 20887
rect 29788 20884 29794 20936
rect 29840 20924 29868 21100
rect 30193 21097 30205 21131
rect 30239 21128 30251 21131
rect 31018 21128 31024 21140
rect 30239 21100 31024 21128
rect 30239 21097 30251 21100
rect 30193 21091 30251 21097
rect 31018 21088 31024 21100
rect 31076 21088 31082 21140
rect 31386 21088 31392 21140
rect 31444 21128 31450 21140
rect 33321 21131 33379 21137
rect 33321 21128 33333 21131
rect 31444 21100 33333 21128
rect 31444 21088 31450 21100
rect 33321 21097 33333 21100
rect 33367 21097 33379 21131
rect 33321 21091 33379 21097
rect 33410 21088 33416 21140
rect 33468 21128 33474 21140
rect 34885 21131 34943 21137
rect 34885 21128 34897 21131
rect 33468 21100 34897 21128
rect 33468 21088 33474 21100
rect 34885 21097 34897 21100
rect 34931 21097 34943 21131
rect 34885 21091 34943 21097
rect 29914 21020 29920 21072
rect 29972 21060 29978 21072
rect 30929 21063 30987 21069
rect 29972 21032 30512 21060
rect 29972 21020 29978 21032
rect 30300 21001 30328 21032
rect 30285 20995 30343 21001
rect 30285 20961 30297 20995
rect 30331 20961 30343 20995
rect 30285 20955 30343 20961
rect 30374 20952 30380 21004
rect 30432 20952 30438 21004
rect 30484 20992 30512 21032
rect 30929 21029 30941 21063
rect 30975 21060 30987 21063
rect 33686 21060 33692 21072
rect 30975 21032 32536 21060
rect 30975 21029 30987 21032
rect 30929 21023 30987 21029
rect 31478 20992 31484 21004
rect 30484 20964 31484 20992
rect 31478 20952 31484 20964
rect 31536 20952 31542 21004
rect 29917 20927 29975 20933
rect 29917 20924 29929 20927
rect 29840 20896 29929 20924
rect 29917 20893 29929 20896
rect 29963 20893 29975 20927
rect 29917 20887 29975 20893
rect 30009 20927 30067 20933
rect 30009 20893 30021 20927
rect 30055 20924 30067 20927
rect 30392 20924 30420 20952
rect 30745 20927 30803 20933
rect 30745 20924 30757 20927
rect 30055 20896 30757 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 30745 20893 30757 20896
rect 30791 20893 30803 20927
rect 30745 20887 30803 20893
rect 28442 20816 28448 20868
rect 28500 20865 28506 20868
rect 28500 20859 28529 20865
rect 28517 20856 28529 20859
rect 29722 20856 29750 20884
rect 28517 20828 29750 20856
rect 29825 20859 29883 20865
rect 28517 20825 28529 20828
rect 28500 20819 28529 20825
rect 29825 20825 29837 20859
rect 29871 20825 29883 20859
rect 29825 20819 29883 20825
rect 28500 20816 28506 20819
rect 22419 20760 22876 20788
rect 22419 20757 22431 20760
rect 22373 20751 22431 20757
rect 23014 20748 23020 20800
rect 23072 20748 23078 20800
rect 23106 20748 23112 20800
rect 23164 20748 23170 20800
rect 27982 20748 27988 20800
rect 28040 20748 28046 20800
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 29840 20788 29868 20819
rect 29420 20760 29868 20788
rect 29932 20788 29960 20887
rect 31110 20884 31116 20936
rect 31168 20884 31174 20936
rect 31297 20927 31355 20933
rect 31297 20893 31309 20927
rect 31343 20924 31355 20927
rect 31570 20924 31576 20936
rect 31343 20896 31576 20924
rect 31343 20893 31355 20896
rect 31297 20887 31355 20893
rect 30190 20816 30196 20868
rect 30248 20856 30254 20868
rect 30423 20859 30481 20865
rect 30423 20856 30435 20859
rect 30248 20828 30435 20856
rect 30248 20816 30254 20828
rect 30423 20825 30435 20828
rect 30469 20825 30481 20859
rect 30423 20819 30481 20825
rect 30558 20816 30564 20868
rect 30616 20816 30622 20868
rect 30653 20859 30711 20865
rect 30653 20825 30665 20859
rect 30699 20825 30711 20859
rect 30653 20819 30711 20825
rect 30668 20788 30696 20819
rect 30834 20816 30840 20868
rect 30892 20856 30898 20868
rect 31312 20856 31340 20887
rect 31570 20884 31576 20896
rect 31628 20884 31634 20936
rect 31754 20884 31760 20936
rect 31812 20924 31818 20936
rect 31849 20927 31907 20933
rect 31849 20924 31861 20927
rect 31812 20896 31861 20924
rect 31812 20884 31818 20896
rect 31849 20893 31861 20896
rect 31895 20893 31907 20927
rect 31849 20887 31907 20893
rect 32122 20856 32128 20868
rect 30892 20828 31340 20856
rect 31404 20828 32128 20856
rect 30892 20816 30898 20828
rect 29932 20760 30696 20788
rect 29420 20748 29426 20760
rect 31018 20748 31024 20800
rect 31076 20788 31082 20800
rect 31404 20788 31432 20828
rect 32122 20816 32128 20828
rect 32180 20816 32186 20868
rect 32508 20856 32536 21032
rect 32600 21032 33692 21060
rect 32600 21001 32628 21032
rect 33686 21020 33692 21032
rect 33744 21060 33750 21072
rect 35529 21063 35587 21069
rect 35529 21060 35541 21063
rect 33744 21032 35541 21060
rect 33744 21020 33750 21032
rect 35529 21029 35541 21032
rect 35575 21029 35587 21063
rect 35529 21023 35587 21029
rect 32585 20995 32643 21001
rect 32585 20961 32597 20995
rect 32631 20961 32643 20995
rect 32585 20955 32643 20961
rect 32674 20952 32680 21004
rect 32732 20992 32738 21004
rect 32769 20995 32827 21001
rect 32769 20992 32781 20995
rect 32732 20964 32781 20992
rect 32732 20952 32738 20964
rect 32769 20961 32781 20964
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 33410 20952 33416 21004
rect 33468 20992 33474 21004
rect 33778 20992 33784 21004
rect 33468 20964 33784 20992
rect 33468 20952 33474 20964
rect 33778 20952 33784 20964
rect 33836 20952 33842 21004
rect 34238 20952 34244 21004
rect 34296 20992 34302 21004
rect 34514 20992 34520 21004
rect 34296 20964 34520 20992
rect 34296 20952 34302 20964
rect 34514 20952 34520 20964
rect 34572 20952 34578 21004
rect 34790 20952 34796 21004
rect 34848 20992 34854 21004
rect 34848 20964 34928 20992
rect 34848 20952 34854 20964
rect 33226 20884 33232 20936
rect 33284 20924 33290 20936
rect 34900 20933 34928 20964
rect 35342 20952 35348 21004
rect 35400 20992 35406 21004
rect 35400 20964 35848 20992
rect 35400 20952 35406 20964
rect 33505 20927 33563 20933
rect 33505 20924 33517 20927
rect 33284 20896 33517 20924
rect 33284 20884 33290 20896
rect 33505 20893 33517 20896
rect 33551 20893 33563 20927
rect 33505 20887 33563 20893
rect 33597 20927 33655 20933
rect 33597 20893 33609 20927
rect 33643 20924 33655 20927
rect 34885 20927 34943 20933
rect 34885 20924 34897 20927
rect 33643 20896 34897 20924
rect 33643 20893 33655 20896
rect 33597 20887 33655 20893
rect 34885 20893 34897 20896
rect 34931 20893 34943 20927
rect 34885 20887 34943 20893
rect 34974 20884 34980 20936
rect 35032 20884 35038 20936
rect 35437 20927 35495 20933
rect 35437 20924 35449 20927
rect 35084 20896 35449 20924
rect 33134 20856 33140 20868
rect 32508 20828 33140 20856
rect 33134 20816 33140 20828
rect 33192 20816 33198 20868
rect 33321 20859 33379 20865
rect 33321 20825 33333 20859
rect 33367 20825 33379 20859
rect 33321 20819 33379 20825
rect 31076 20760 31432 20788
rect 31481 20791 31539 20797
rect 31076 20748 31082 20760
rect 31481 20757 31493 20791
rect 31527 20788 31539 20791
rect 31570 20788 31576 20800
rect 31527 20760 31576 20788
rect 31527 20757 31539 20760
rect 31481 20751 31539 20757
rect 31570 20748 31576 20760
rect 31628 20748 31634 20800
rect 31662 20748 31668 20800
rect 31720 20748 31726 20800
rect 32858 20748 32864 20800
rect 32916 20748 32922 20800
rect 33229 20791 33287 20797
rect 33229 20757 33241 20791
rect 33275 20788 33287 20791
rect 33336 20788 33364 20819
rect 34514 20816 34520 20868
rect 34572 20856 34578 20868
rect 35084 20856 35112 20896
rect 35437 20893 35449 20896
rect 35483 20893 35495 20927
rect 35437 20887 35495 20893
rect 35710 20884 35716 20936
rect 35768 20884 35774 20936
rect 35820 20933 35848 20964
rect 35805 20927 35863 20933
rect 35805 20893 35817 20927
rect 35851 20893 35863 20927
rect 35805 20887 35863 20893
rect 34572 20828 35112 20856
rect 35345 20859 35403 20865
rect 34572 20816 34578 20828
rect 35345 20825 35357 20859
rect 35391 20856 35403 20859
rect 35391 20828 35480 20856
rect 35391 20825 35403 20828
rect 35345 20819 35403 20825
rect 35452 20800 35480 20828
rect 33275 20760 33364 20788
rect 33275 20757 33287 20760
rect 33229 20751 33287 20757
rect 33594 20748 33600 20800
rect 33652 20788 33658 20800
rect 33781 20791 33839 20797
rect 33781 20788 33793 20791
rect 33652 20760 33793 20788
rect 33652 20748 33658 20760
rect 33781 20757 33793 20760
rect 33827 20757 33839 20791
rect 33781 20751 33839 20757
rect 34698 20748 34704 20800
rect 34756 20748 34762 20800
rect 35434 20748 35440 20800
rect 35492 20788 35498 20800
rect 35989 20791 36047 20797
rect 35989 20788 36001 20791
rect 35492 20760 36001 20788
rect 35492 20748 35498 20760
rect 35989 20757 36001 20760
rect 36035 20757 36047 20791
rect 35989 20751 36047 20757
rect 1104 20698 36524 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 36524 20698
rect 1104 20624 36524 20646
rect 2498 20544 2504 20596
rect 2556 20584 2562 20596
rect 2556 20556 3740 20584
rect 2556 20544 2562 20556
rect 3712 20516 3740 20556
rect 3786 20544 3792 20596
rect 3844 20544 3850 20596
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 5074 20584 5080 20596
rect 4396 20556 5080 20584
rect 4396 20544 4402 20556
rect 5074 20544 5080 20556
rect 5132 20544 5138 20596
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5626 20584 5632 20596
rect 5307 20556 5632 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 5810 20544 5816 20596
rect 5868 20584 5874 20596
rect 6457 20587 6515 20593
rect 6457 20584 6469 20587
rect 5868 20556 6469 20584
rect 5868 20544 5874 20556
rect 6457 20553 6469 20556
rect 6503 20553 6515 20587
rect 6457 20547 6515 20553
rect 7558 20544 7564 20596
rect 7616 20584 7622 20596
rect 7745 20587 7803 20593
rect 7745 20584 7757 20587
rect 7616 20556 7757 20584
rect 7616 20544 7622 20556
rect 7745 20553 7757 20556
rect 7791 20553 7803 20587
rect 7745 20547 7803 20553
rect 8018 20544 8024 20596
rect 8076 20584 8082 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 8076 20556 8217 20584
rect 8076 20544 8082 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 15194 20584 15200 20596
rect 8205 20547 8263 20553
rect 14660 20556 15200 20584
rect 3712 20488 5396 20516
rect 1394 20408 1400 20460
rect 1452 20448 1458 20460
rect 1581 20451 1639 20457
rect 1581 20448 1593 20451
rect 1452 20420 1593 20448
rect 1452 20408 1458 20420
rect 1581 20417 1593 20420
rect 1627 20417 1639 20451
rect 1581 20411 1639 20417
rect 2958 20408 2964 20460
rect 3016 20408 3022 20460
rect 4525 20451 4583 20457
rect 4525 20417 4537 20451
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 1903 20352 3464 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 3436 20321 3464 20352
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 4062 20340 4068 20392
rect 4120 20340 4126 20392
rect 4540 20380 4568 20411
rect 4706 20408 4712 20460
rect 4764 20408 4770 20460
rect 4798 20408 4804 20460
rect 4856 20448 4862 20460
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 4856 20420 4905 20448
rect 4856 20408 4862 20420
rect 4893 20417 4905 20420
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 4985 20451 5043 20457
rect 4985 20417 4997 20451
rect 5031 20448 5043 20451
rect 5258 20448 5264 20460
rect 5031 20420 5264 20448
rect 5031 20417 5043 20420
rect 4985 20411 5043 20417
rect 5258 20408 5264 20420
rect 5316 20408 5322 20460
rect 5368 20457 5396 20488
rect 5718 20476 5724 20528
rect 5776 20516 5782 20528
rect 6546 20516 6552 20528
rect 5776 20488 6552 20516
rect 5776 20476 5782 20488
rect 6546 20476 6552 20488
rect 6604 20476 6610 20528
rect 6730 20476 6736 20528
rect 6788 20516 6794 20528
rect 7098 20516 7104 20528
rect 6788 20488 7104 20516
rect 6788 20476 6794 20488
rect 7098 20476 7104 20488
rect 7156 20476 7162 20528
rect 7193 20519 7251 20525
rect 7193 20485 7205 20519
rect 7239 20516 7251 20519
rect 7466 20516 7472 20528
rect 7239 20488 7472 20516
rect 7239 20485 7251 20488
rect 7193 20479 7251 20485
rect 7466 20476 7472 20488
rect 7524 20476 7530 20528
rect 8294 20476 8300 20528
rect 8352 20516 8358 20528
rect 9490 20516 9496 20528
rect 8352 20488 9496 20516
rect 8352 20476 8358 20488
rect 5902 20457 5908 20460
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 5446 20451 5504 20457
rect 5446 20417 5458 20451
rect 5492 20417 5504 20451
rect 5446 20411 5504 20417
rect 5629 20451 5687 20457
rect 5629 20417 5641 20451
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 5859 20451 5908 20457
rect 5859 20417 5871 20451
rect 5905 20417 5908 20451
rect 5859 20411 5908 20417
rect 4540 20352 4936 20380
rect 4908 20324 4936 20352
rect 5074 20340 5080 20392
rect 5132 20380 5138 20392
rect 5460 20380 5488 20411
rect 5132 20352 5488 20380
rect 5132 20340 5138 20352
rect 3421 20315 3479 20321
rect 3421 20281 3433 20315
rect 3467 20281 3479 20315
rect 3421 20275 3479 20281
rect 4890 20272 4896 20324
rect 4948 20272 4954 20324
rect 5644 20312 5672 20411
rect 5874 20408 5908 20411
rect 5960 20408 5966 20460
rect 6638 20408 6644 20460
rect 6696 20408 6702 20460
rect 6822 20408 6828 20460
rect 6880 20408 6886 20460
rect 6914 20408 6920 20460
rect 6972 20408 6978 20460
rect 7305 20451 7363 20457
rect 7305 20417 7317 20451
rect 7351 20417 7363 20451
rect 7305 20411 7363 20417
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8570 20448 8576 20460
rect 8159 20420 8576 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 5874 20380 5902 20408
rect 7320 20380 7348 20411
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 8754 20408 8760 20460
rect 8812 20408 8818 20460
rect 8956 20457 8984 20488
rect 9490 20476 9496 20488
rect 9548 20476 9554 20528
rect 13262 20476 13268 20528
rect 13320 20476 13326 20528
rect 13722 20476 13728 20528
rect 13780 20516 13786 20528
rect 14660 20516 14688 20556
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 16209 20587 16267 20593
rect 16209 20584 16221 20587
rect 15620 20556 16221 20584
rect 15620 20544 15626 20556
rect 16209 20553 16221 20556
rect 16255 20553 16267 20587
rect 16209 20547 16267 20553
rect 17034 20544 17040 20596
rect 17092 20544 17098 20596
rect 17586 20544 17592 20596
rect 17644 20584 17650 20596
rect 17644 20556 17724 20584
rect 17644 20544 17650 20556
rect 13780 20488 14766 20516
rect 13780 20476 13786 20488
rect 16298 20476 16304 20528
rect 16356 20516 16362 20528
rect 17696 20525 17724 20556
rect 17770 20544 17776 20596
rect 17828 20544 17834 20596
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 18693 20587 18751 20593
rect 18693 20584 18705 20587
rect 18288 20556 18705 20584
rect 18288 20544 18294 20556
rect 18693 20553 18705 20556
rect 18739 20553 18751 20587
rect 18693 20547 18751 20553
rect 20806 20544 20812 20596
rect 20864 20544 20870 20596
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 22186 20584 22192 20596
rect 22143 20556 22192 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 23017 20587 23075 20593
rect 23017 20584 23029 20587
rect 22296 20556 23029 20584
rect 16853 20519 16911 20525
rect 16853 20516 16865 20519
rect 16356 20488 16865 20516
rect 16356 20476 16362 20488
rect 16853 20485 16865 20488
rect 16899 20485 16911 20519
rect 16853 20479 16911 20485
rect 17681 20519 17739 20525
rect 17681 20485 17693 20519
rect 17727 20485 17739 20519
rect 17681 20479 17739 20485
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 10962 20448 10968 20460
rect 9824 20420 10968 20448
rect 9824 20408 9830 20420
rect 10962 20408 10968 20420
rect 11020 20448 11026 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11020 20420 11529 20448
rect 11020 20408 11026 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 11606 20408 11612 20460
rect 11664 20448 11670 20460
rect 11701 20451 11759 20457
rect 11701 20448 11713 20451
rect 11664 20420 11713 20448
rect 11664 20408 11670 20420
rect 11701 20417 11713 20420
rect 11747 20417 11759 20451
rect 11701 20411 11759 20417
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 13357 20451 13415 20457
rect 13357 20448 13369 20451
rect 13219 20420 13369 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 13357 20417 13369 20420
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 13630 20408 13636 20460
rect 13688 20408 13694 20460
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 16022 20448 16028 20460
rect 15620 20420 16028 20448
rect 15620 20408 15626 20420
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 16114 20408 16120 20460
rect 16172 20448 16178 20460
rect 17788 20457 17816 20544
rect 18325 20519 18383 20525
rect 18325 20485 18337 20519
rect 18371 20485 18383 20519
rect 18325 20479 18383 20485
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16172 20420 16681 20448
rect 16172 20408 16178 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20428 17647 20451
rect 17773 20451 17831 20457
rect 17635 20417 17724 20428
rect 17589 20411 17724 20417
rect 17773 20417 17785 20451
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20448 18015 20451
rect 18046 20448 18052 20460
rect 18003 20420 18052 20448
rect 18003 20417 18015 20420
rect 17957 20411 18015 20417
rect 8202 20380 8208 20392
rect 5874 20352 8208 20380
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 8389 20383 8447 20389
rect 8389 20349 8401 20383
rect 8435 20349 8447 20383
rect 8389 20343 8447 20349
rect 6730 20312 6736 20324
rect 5644 20284 6736 20312
rect 6730 20272 6736 20284
rect 6788 20272 6794 20324
rect 6917 20315 6975 20321
rect 6917 20281 6929 20315
rect 6963 20312 6975 20315
rect 7190 20312 7196 20324
rect 6963 20284 7196 20312
rect 6963 20281 6975 20284
rect 6917 20275 6975 20281
rect 7190 20272 7196 20284
rect 7248 20272 7254 20324
rect 8110 20272 8116 20324
rect 8168 20312 8174 20324
rect 8404 20312 8432 20343
rect 12526 20340 12532 20392
rect 12584 20340 12590 20392
rect 13725 20383 13783 20389
rect 13725 20349 13737 20383
rect 13771 20380 13783 20383
rect 13814 20380 13820 20392
rect 13771 20352 13820 20380
rect 13771 20349 13783 20352
rect 13725 20343 13783 20349
rect 13814 20340 13820 20352
rect 13872 20340 13878 20392
rect 13998 20340 14004 20392
rect 14056 20340 14062 20392
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 14642 20380 14648 20392
rect 14323 20352 14648 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 15746 20340 15752 20392
rect 15804 20380 15810 20392
rect 15841 20383 15899 20389
rect 15841 20380 15853 20383
rect 15804 20352 15853 20380
rect 15804 20340 15810 20352
rect 15841 20349 15853 20352
rect 15887 20380 15899 20383
rect 16132 20380 16160 20408
rect 17604 20400 17724 20411
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 18340 20448 18368 20479
rect 18506 20476 18512 20528
rect 18564 20525 18570 20528
rect 18564 20519 18583 20525
rect 18571 20485 18583 20519
rect 18564 20479 18583 20485
rect 18564 20476 18570 20479
rect 18782 20476 18788 20528
rect 18840 20476 18846 20528
rect 20162 20476 20168 20528
rect 20220 20516 20226 20528
rect 21453 20519 21511 20525
rect 21453 20516 21465 20519
rect 20220 20488 20760 20516
rect 20220 20476 20226 20488
rect 19058 20448 19064 20460
rect 18340 20420 19064 20448
rect 19058 20408 19064 20420
rect 19116 20448 19122 20460
rect 20070 20448 20076 20460
rect 19116 20420 20076 20448
rect 19116 20408 19122 20420
rect 20070 20408 20076 20420
rect 20128 20448 20134 20460
rect 20346 20448 20352 20460
rect 20128 20420 20352 20448
rect 20128 20408 20134 20420
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20622 20408 20628 20460
rect 20680 20408 20686 20460
rect 20732 20457 20760 20488
rect 20824 20488 21465 20516
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 15887 20352 16160 20380
rect 15887 20349 15899 20352
rect 15841 20343 15899 20349
rect 8573 20315 8631 20321
rect 8573 20312 8585 20315
rect 8168 20284 8585 20312
rect 8168 20272 8174 20284
rect 8573 20281 8585 20284
rect 8619 20281 8631 20315
rect 8573 20275 8631 20281
rect 17218 20272 17224 20324
rect 17276 20312 17282 20324
rect 17405 20315 17463 20321
rect 17405 20312 17417 20315
rect 17276 20284 17417 20312
rect 17276 20272 17282 20284
rect 17405 20281 17417 20284
rect 17451 20281 17463 20315
rect 17696 20312 17724 20400
rect 19702 20340 19708 20392
rect 19760 20380 19766 20392
rect 20824 20380 20852 20488
rect 21453 20485 21465 20488
rect 21499 20516 21511 20519
rect 21499 20488 22232 20516
rect 21499 20485 21511 20488
rect 21453 20479 21511 20485
rect 20898 20408 20904 20460
rect 20956 20408 20962 20460
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 19760 20352 20852 20380
rect 19760 20340 19766 20352
rect 18782 20312 18788 20324
rect 17696 20284 17748 20312
rect 17405 20275 17463 20281
rect 3329 20247 3387 20253
rect 3329 20213 3341 20247
rect 3375 20244 3387 20247
rect 4338 20244 4344 20256
rect 3375 20216 4344 20244
rect 3375 20213 3387 20216
rect 3329 20207 3387 20213
rect 4338 20204 4344 20216
rect 4396 20204 4402 20256
rect 4522 20204 4528 20256
rect 4580 20244 4586 20256
rect 4798 20244 4804 20256
rect 4580 20216 4804 20244
rect 4580 20204 4586 20216
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5994 20204 6000 20256
rect 6052 20204 6058 20256
rect 6825 20247 6883 20253
rect 6825 20213 6837 20247
rect 6871 20244 6883 20247
rect 7098 20244 7104 20256
rect 6871 20216 7104 20244
rect 6871 20213 6883 20216
rect 6825 20207 6883 20213
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 8941 20247 8999 20253
rect 8941 20213 8953 20247
rect 8987 20244 8999 20247
rect 9582 20244 9588 20256
rect 8987 20216 9588 20244
rect 8987 20213 8999 20216
rect 8941 20207 8999 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 11422 20204 11428 20256
rect 11480 20244 11486 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11480 20216 11529 20244
rect 11480 20204 11486 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 13630 20204 13636 20256
rect 13688 20244 13694 20256
rect 13909 20247 13967 20253
rect 13909 20244 13921 20247
rect 13688 20216 13921 20244
rect 13688 20204 13694 20216
rect 13909 20213 13921 20216
rect 13955 20213 13967 20247
rect 13909 20207 13967 20213
rect 15746 20204 15752 20256
rect 15804 20204 15810 20256
rect 17720 20244 17748 20284
rect 17926 20284 18788 20312
rect 17926 20244 17954 20284
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 20714 20272 20720 20324
rect 20772 20312 20778 20324
rect 21008 20312 21036 20411
rect 21100 20380 21128 20411
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21269 20451 21327 20457
rect 21269 20448 21281 20451
rect 21232 20420 21281 20448
rect 21232 20408 21238 20420
rect 21269 20417 21281 20420
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21542 20408 21548 20460
rect 21600 20448 21606 20460
rect 22002 20448 22008 20460
rect 21600 20420 22008 20448
rect 21600 20408 21606 20420
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 21634 20380 21640 20392
rect 21100 20352 21640 20380
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 22204 20380 22232 20488
rect 22296 20457 22324 20556
rect 23017 20553 23029 20556
rect 23063 20584 23075 20587
rect 23106 20584 23112 20596
rect 23063 20556 23112 20584
rect 23063 20553 23075 20556
rect 23017 20547 23075 20553
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 26329 20587 26387 20593
rect 26329 20553 26341 20587
rect 26375 20553 26387 20587
rect 26329 20547 26387 20553
rect 26497 20587 26555 20593
rect 26497 20553 26509 20587
rect 26543 20584 26555 20587
rect 26602 20584 26608 20596
rect 26543 20556 26608 20584
rect 26543 20553 26555 20556
rect 26497 20547 26555 20553
rect 22830 20516 22836 20528
rect 22388 20488 22836 20516
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22388 20380 22416 20488
rect 22830 20476 22836 20488
rect 22888 20516 22894 20528
rect 23290 20516 23296 20528
rect 22888 20488 23296 20516
rect 22888 20476 22894 20488
rect 23290 20476 23296 20488
rect 23348 20476 23354 20528
rect 23569 20519 23627 20525
rect 23569 20516 23581 20519
rect 23416 20488 23581 20516
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22704 20420 22937 20448
rect 22704 20408 22710 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23121 20451 23179 20457
rect 23121 20417 23133 20451
rect 23167 20448 23179 20451
rect 23416 20448 23444 20488
rect 23569 20485 23581 20488
rect 23615 20516 23627 20519
rect 23615 20488 25912 20516
rect 23615 20485 23627 20488
rect 23569 20479 23627 20485
rect 23167 20420 23444 20448
rect 23167 20417 23179 20420
rect 23121 20411 23179 20417
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 23532 20420 23888 20448
rect 23532 20408 23538 20420
rect 22204 20352 22416 20380
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20380 22523 20383
rect 23014 20380 23020 20392
rect 22511 20352 23020 20380
rect 22511 20349 22523 20352
rect 22465 20343 22523 20349
rect 23014 20340 23020 20352
rect 23072 20340 23078 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23860 20389 23888 20420
rect 23934 20408 23940 20460
rect 23992 20408 23998 20460
rect 24762 20408 24768 20460
rect 24820 20408 24826 20460
rect 25038 20408 25044 20460
rect 25096 20408 25102 20460
rect 25884 20457 25912 20488
rect 25869 20451 25927 20457
rect 25869 20417 25881 20451
rect 25915 20448 25927 20451
rect 26344 20448 26372 20547
rect 26602 20544 26608 20556
rect 26660 20544 26666 20596
rect 27890 20544 27896 20596
rect 27948 20584 27954 20596
rect 28718 20584 28724 20596
rect 27948 20556 28724 20584
rect 27948 20544 27954 20556
rect 28718 20544 28724 20556
rect 28776 20544 28782 20596
rect 28920 20556 33640 20584
rect 26697 20519 26755 20525
rect 26697 20485 26709 20519
rect 26743 20516 26755 20519
rect 26878 20516 26884 20528
rect 26743 20488 26884 20516
rect 26743 20485 26755 20488
rect 26697 20479 26755 20485
rect 26878 20476 26884 20488
rect 26936 20476 26942 20528
rect 28258 20516 28264 20528
rect 28000 20488 28264 20516
rect 25915 20420 26372 20448
rect 25915 20417 25927 20420
rect 25869 20411 25927 20417
rect 26602 20408 26608 20460
rect 26660 20448 26666 20460
rect 27249 20451 27307 20457
rect 27249 20448 27261 20451
rect 26660 20420 27261 20448
rect 26660 20408 26666 20420
rect 27249 20417 27261 20420
rect 27295 20417 27307 20451
rect 27249 20411 27307 20417
rect 27338 20408 27344 20460
rect 27396 20448 27402 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 27396 20420 27537 20448
rect 27396 20408 27402 20420
rect 27525 20417 27537 20420
rect 27571 20417 27583 20451
rect 27525 20411 27583 20417
rect 27709 20451 27767 20457
rect 27709 20417 27721 20451
rect 27755 20448 27767 20451
rect 27890 20448 27896 20460
rect 27755 20420 27896 20448
rect 27755 20417 27767 20420
rect 27709 20411 27767 20417
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28000 20457 28028 20488
rect 28258 20476 28264 20488
rect 28316 20476 28322 20528
rect 27985 20451 28043 20457
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28169 20451 28227 20457
rect 28169 20417 28181 20451
rect 28215 20448 28227 20451
rect 28718 20448 28724 20460
rect 28215 20420 28724 20448
rect 28215 20417 28227 20420
rect 28169 20411 28227 20417
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 23753 20383 23811 20389
rect 23753 20380 23765 20383
rect 23348 20352 23765 20380
rect 23348 20340 23354 20352
rect 23753 20349 23765 20352
rect 23799 20349 23811 20383
rect 23753 20343 23811 20349
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 24210 20380 24216 20392
rect 23891 20352 24216 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 24210 20340 24216 20352
rect 24268 20340 24274 20392
rect 24949 20383 25007 20389
rect 24949 20349 24961 20383
rect 24995 20349 25007 20383
rect 24949 20343 25007 20349
rect 21082 20312 21088 20324
rect 20772 20284 21088 20312
rect 20772 20272 20778 20284
rect 21082 20272 21088 20284
rect 21140 20272 21146 20324
rect 21266 20272 21272 20324
rect 21324 20272 21330 20324
rect 21450 20272 21456 20324
rect 21508 20312 21514 20324
rect 21508 20284 23980 20312
rect 21508 20272 21514 20284
rect 17720 20216 17954 20244
rect 18509 20247 18567 20253
rect 18509 20213 18521 20247
rect 18555 20244 18567 20247
rect 19426 20244 19432 20256
rect 18555 20216 19432 20244
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 20070 20204 20076 20256
rect 20128 20204 20134 20256
rect 23290 20204 23296 20256
rect 23348 20244 23354 20256
rect 23474 20244 23480 20256
rect 23348 20216 23480 20244
rect 23348 20204 23354 20216
rect 23474 20204 23480 20216
rect 23532 20204 23538 20256
rect 23658 20204 23664 20256
rect 23716 20244 23722 20256
rect 23753 20247 23811 20253
rect 23753 20244 23765 20247
rect 23716 20216 23765 20244
rect 23716 20204 23722 20216
rect 23753 20213 23765 20216
rect 23799 20213 23811 20247
rect 23952 20244 23980 20284
rect 24026 20272 24032 20324
rect 24084 20312 24090 20324
rect 24964 20312 24992 20343
rect 25314 20340 25320 20392
rect 25372 20380 25378 20392
rect 25593 20383 25651 20389
rect 25593 20380 25605 20383
rect 25372 20352 25605 20380
rect 25372 20340 25378 20352
rect 25593 20349 25605 20352
rect 25639 20349 25651 20383
rect 25593 20343 25651 20349
rect 27430 20340 27436 20392
rect 27488 20340 27494 20392
rect 28077 20383 28135 20389
rect 28077 20349 28089 20383
rect 28123 20380 28135 20383
rect 28626 20380 28632 20392
rect 28123 20352 28632 20380
rect 28123 20349 28135 20352
rect 28077 20343 28135 20349
rect 28626 20340 28632 20352
rect 28684 20380 28690 20392
rect 28920 20380 28948 20556
rect 29638 20476 29644 20528
rect 29696 20516 29702 20528
rect 29733 20519 29791 20525
rect 29733 20516 29745 20519
rect 29696 20488 29745 20516
rect 29696 20476 29702 20488
rect 29733 20485 29745 20488
rect 29779 20485 29791 20519
rect 30282 20516 30288 20528
rect 29733 20479 29791 20485
rect 29932 20488 30288 20516
rect 29086 20408 29092 20460
rect 29144 20448 29150 20460
rect 29549 20451 29607 20457
rect 29549 20448 29561 20451
rect 29144 20420 29561 20448
rect 29144 20408 29150 20420
rect 29549 20417 29561 20420
rect 29595 20417 29607 20451
rect 29549 20411 29607 20417
rect 28684 20352 28948 20380
rect 29564 20380 29592 20411
rect 29822 20408 29828 20460
rect 29880 20408 29886 20460
rect 29932 20457 29960 20488
rect 30282 20476 30288 20488
rect 30340 20476 30346 20528
rect 31389 20519 31447 20525
rect 31389 20485 31401 20519
rect 31435 20516 31447 20519
rect 33226 20516 33232 20528
rect 31435 20488 31708 20516
rect 31435 20485 31447 20488
rect 31389 20479 31447 20485
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20417 29975 20451
rect 29917 20411 29975 20417
rect 30190 20408 30196 20460
rect 30248 20448 30254 20460
rect 30653 20451 30711 20457
rect 30653 20448 30665 20451
rect 30248 20420 30665 20448
rect 30248 20408 30254 20420
rect 30653 20417 30665 20420
rect 30699 20417 30711 20451
rect 30653 20411 30711 20417
rect 30834 20408 30840 20460
rect 30892 20408 30898 20460
rect 31271 20451 31329 20457
rect 31271 20417 31283 20451
rect 31317 20417 31329 20451
rect 31271 20411 31329 20417
rect 31481 20451 31539 20457
rect 31481 20417 31493 20451
rect 31527 20417 31539 20451
rect 31481 20411 31539 20417
rect 31573 20451 31631 20457
rect 31573 20417 31585 20451
rect 31619 20417 31631 20451
rect 31573 20411 31631 20417
rect 30282 20380 30288 20392
rect 29564 20352 30288 20380
rect 28684 20340 28690 20352
rect 30282 20340 30288 20352
rect 30340 20340 30346 20392
rect 30742 20340 30748 20392
rect 30800 20380 30806 20392
rect 31110 20380 31116 20392
rect 30800 20352 31116 20380
rect 30800 20340 30806 20352
rect 31110 20340 31116 20352
rect 31168 20340 31174 20392
rect 31286 20380 31314 20411
rect 31386 20380 31392 20392
rect 31286 20352 31392 20380
rect 31386 20340 31392 20352
rect 31444 20340 31450 20392
rect 24084 20284 24992 20312
rect 24084 20272 24090 20284
rect 25130 20272 25136 20324
rect 25188 20272 25194 20324
rect 25774 20272 25780 20324
rect 25832 20312 25838 20324
rect 27065 20315 27123 20321
rect 27065 20312 27077 20315
rect 25832 20284 27077 20312
rect 25832 20272 25838 20284
rect 27065 20281 27077 20284
rect 27111 20312 27123 20315
rect 28810 20312 28816 20324
rect 27111 20284 28816 20312
rect 27111 20281 27123 20284
rect 27065 20275 27123 20281
rect 28810 20272 28816 20284
rect 28868 20272 28874 20324
rect 29086 20272 29092 20324
rect 29144 20312 29150 20324
rect 29822 20312 29828 20324
rect 29144 20284 29828 20312
rect 29144 20272 29150 20284
rect 29822 20272 29828 20284
rect 29880 20272 29886 20324
rect 30834 20312 30840 20324
rect 30024 20284 30840 20312
rect 24581 20247 24639 20253
rect 24581 20244 24593 20247
rect 23952 20216 24593 20244
rect 23753 20207 23811 20213
rect 24581 20213 24593 20216
rect 24627 20244 24639 20247
rect 24854 20244 24860 20256
rect 24627 20216 24860 20244
rect 24627 20213 24639 20216
rect 24581 20207 24639 20213
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 26234 20204 26240 20256
rect 26292 20244 26298 20256
rect 26513 20247 26571 20253
rect 26513 20244 26525 20247
rect 26292 20216 26525 20244
rect 26292 20204 26298 20216
rect 26513 20213 26525 20216
rect 26559 20213 26571 20247
rect 26513 20207 26571 20213
rect 27614 20204 27620 20256
rect 27672 20204 27678 20256
rect 27798 20204 27804 20256
rect 27856 20244 27862 20256
rect 28442 20244 28448 20256
rect 27856 20216 28448 20244
rect 27856 20204 27862 20216
rect 28442 20204 28448 20216
rect 28500 20204 28506 20256
rect 29178 20204 29184 20256
rect 29236 20244 29242 20256
rect 30024 20244 30052 20284
rect 30834 20272 30840 20284
rect 30892 20312 30898 20324
rect 31496 20312 31524 20411
rect 30892 20284 31524 20312
rect 30892 20272 30898 20284
rect 29236 20216 30052 20244
rect 29236 20204 29242 20216
rect 30098 20204 30104 20256
rect 30156 20204 30162 20256
rect 30650 20204 30656 20256
rect 30708 20204 30714 20256
rect 31021 20247 31079 20253
rect 31021 20213 31033 20247
rect 31067 20244 31079 20247
rect 31478 20244 31484 20256
rect 31067 20216 31484 20244
rect 31067 20213 31079 20216
rect 31021 20207 31079 20213
rect 31478 20204 31484 20216
rect 31536 20204 31542 20256
rect 31588 20244 31616 20411
rect 31680 20392 31708 20488
rect 32600 20488 33232 20516
rect 32306 20408 32312 20460
rect 32364 20448 32370 20460
rect 32600 20457 32628 20488
rect 33226 20476 33232 20488
rect 33284 20476 33290 20528
rect 32585 20451 32643 20457
rect 32585 20448 32597 20451
rect 32364 20420 32597 20448
rect 32364 20408 32370 20420
rect 32585 20417 32597 20420
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 32858 20408 32864 20460
rect 32916 20408 32922 20460
rect 33612 20457 33640 20556
rect 33505 20451 33563 20457
rect 33505 20417 33517 20451
rect 33551 20417 33563 20451
rect 33505 20411 33563 20417
rect 33597 20451 33655 20457
rect 33597 20417 33609 20451
rect 33643 20417 33655 20451
rect 33597 20411 33655 20417
rect 31662 20340 31668 20392
rect 31720 20340 31726 20392
rect 32769 20383 32827 20389
rect 32769 20349 32781 20383
rect 32815 20380 32827 20383
rect 33321 20383 33379 20389
rect 33321 20380 33333 20383
rect 32815 20352 33333 20380
rect 32815 20349 32827 20352
rect 32769 20343 32827 20349
rect 33321 20349 33333 20352
rect 33367 20349 33379 20383
rect 33520 20380 33548 20411
rect 33686 20408 33692 20460
rect 33744 20448 33750 20460
rect 33781 20451 33839 20457
rect 33781 20448 33793 20451
rect 33744 20420 33793 20448
rect 33744 20408 33750 20420
rect 33781 20417 33793 20420
rect 33827 20417 33839 20451
rect 33781 20411 33839 20417
rect 33870 20408 33876 20460
rect 33928 20408 33934 20460
rect 34422 20408 34428 20460
rect 34480 20448 34486 20460
rect 34609 20451 34667 20457
rect 34609 20448 34621 20451
rect 34480 20420 34621 20448
rect 34480 20408 34486 20420
rect 34609 20417 34621 20420
rect 34655 20417 34667 20451
rect 34609 20411 34667 20417
rect 34790 20408 34796 20460
rect 34848 20408 34854 20460
rect 35250 20380 35256 20392
rect 33520 20352 35256 20380
rect 33321 20343 33379 20349
rect 35250 20340 35256 20352
rect 35308 20380 35314 20392
rect 35526 20380 35532 20392
rect 35308 20352 35532 20380
rect 35308 20340 35314 20352
rect 35526 20340 35532 20352
rect 35584 20340 35590 20392
rect 33134 20272 33140 20324
rect 33192 20312 33198 20324
rect 33686 20312 33692 20324
rect 33192 20284 33692 20312
rect 33192 20272 33198 20284
rect 33686 20272 33692 20284
rect 33744 20272 33750 20324
rect 31662 20244 31668 20256
rect 31588 20216 31668 20244
rect 31662 20204 31668 20216
rect 31720 20204 31726 20256
rect 31757 20247 31815 20253
rect 31757 20213 31769 20247
rect 31803 20244 31815 20247
rect 31846 20244 31852 20256
rect 31803 20216 31852 20244
rect 31803 20213 31815 20216
rect 31757 20207 31815 20213
rect 31846 20204 31852 20216
rect 31904 20204 31910 20256
rect 32398 20204 32404 20256
rect 32456 20204 32462 20256
rect 32582 20204 32588 20256
rect 32640 20204 32646 20256
rect 34698 20204 34704 20256
rect 34756 20244 34762 20256
rect 35342 20244 35348 20256
rect 34756 20216 35348 20244
rect 34756 20204 34762 20216
rect 35342 20204 35348 20216
rect 35400 20204 35406 20256
rect 1104 20154 36524 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 36524 20154
rect 1104 20080 36524 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 2924 20012 3801 20040
rect 2924 20000 2930 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 4614 20040 4620 20052
rect 3789 20003 3847 20009
rect 4448 20012 4620 20040
rect 3145 19975 3203 19981
rect 3145 19941 3157 19975
rect 3191 19972 3203 19975
rect 4448 19972 4476 20012
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 5077 20043 5135 20049
rect 5077 20009 5089 20043
rect 5123 20040 5135 20043
rect 5350 20040 5356 20052
rect 5123 20012 5356 20040
rect 5123 20009 5135 20012
rect 5077 20003 5135 20009
rect 5350 20000 5356 20012
rect 5408 20000 5414 20052
rect 5537 20043 5595 20049
rect 5537 20009 5549 20043
rect 5583 20040 5595 20043
rect 5902 20040 5908 20052
rect 5583 20012 5908 20040
rect 5583 20009 5595 20012
rect 5537 20003 5595 20009
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 7101 20043 7159 20049
rect 7101 20040 7113 20043
rect 7064 20012 7113 20040
rect 7064 20000 7070 20012
rect 7101 20009 7113 20012
rect 7147 20009 7159 20043
rect 7101 20003 7159 20009
rect 7469 20043 7527 20049
rect 7469 20009 7481 20043
rect 7515 20040 7527 20043
rect 7742 20040 7748 20052
rect 7515 20012 7748 20040
rect 7515 20009 7527 20012
rect 7469 20003 7527 20009
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 12161 20043 12219 20049
rect 12161 20009 12173 20043
rect 12207 20040 12219 20043
rect 12526 20040 12532 20052
rect 12207 20012 12532 20040
rect 12207 20009 12219 20012
rect 12161 20003 12219 20009
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 13262 20000 13268 20052
rect 13320 20040 13326 20052
rect 13320 20012 14412 20040
rect 13320 20000 13326 20012
rect 4798 19972 4804 19984
rect 3191 19944 4476 19972
rect 3191 19941 3203 19944
rect 3145 19935 3203 19941
rect 1394 19864 1400 19916
rect 1452 19864 1458 19916
rect 1670 19864 1676 19916
rect 1728 19864 1734 19916
rect 4448 19913 4476 19944
rect 4632 19944 4804 19972
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 4522 19796 4528 19848
rect 4580 19796 4586 19848
rect 4632 19845 4660 19944
rect 4798 19932 4804 19944
rect 4856 19972 4862 19984
rect 6086 19972 6092 19984
rect 4856 19944 6092 19972
rect 4856 19932 4862 19944
rect 6086 19932 6092 19944
rect 6144 19972 6150 19984
rect 6181 19975 6239 19981
rect 6181 19972 6193 19975
rect 6144 19944 6193 19972
rect 6144 19932 6150 19944
rect 6181 19941 6193 19944
rect 6227 19941 6239 19975
rect 6181 19935 6239 19941
rect 6270 19932 6276 19984
rect 6328 19972 6334 19984
rect 9674 19972 9680 19984
rect 6328 19944 9680 19972
rect 6328 19932 6334 19944
rect 9674 19932 9680 19944
rect 9732 19932 9738 19984
rect 14384 19972 14412 20012
rect 14642 20000 14648 20052
rect 14700 20000 14706 20052
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 15344 20012 15485 20040
rect 15344 20000 15350 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 17126 20000 17132 20052
rect 17184 20040 17190 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 17184 20012 17233 20040
rect 17184 20000 17190 20012
rect 17221 20009 17233 20012
rect 17267 20009 17279 20043
rect 17221 20003 17279 20009
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18506 20040 18512 20052
rect 18104 20012 18512 20040
rect 18104 20000 18110 20012
rect 18506 20000 18512 20012
rect 18564 20000 18570 20052
rect 19610 20000 19616 20052
rect 19668 20000 19674 20052
rect 20162 20000 20168 20052
rect 20220 20040 20226 20052
rect 20441 20043 20499 20049
rect 20441 20040 20453 20043
rect 20220 20012 20453 20040
rect 20220 20000 20226 20012
rect 20441 20009 20453 20012
rect 20487 20009 20499 20043
rect 20441 20003 20499 20009
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24213 20043 24271 20049
rect 24213 20040 24225 20043
rect 23992 20012 24225 20040
rect 23992 20000 23998 20012
rect 24213 20009 24225 20012
rect 24259 20040 24271 20043
rect 24854 20040 24860 20052
rect 24259 20012 24860 20040
rect 24259 20009 24271 20012
rect 24213 20003 24271 20009
rect 24854 20000 24860 20012
rect 24912 20000 24918 20052
rect 29822 20040 29828 20052
rect 27908 20012 29828 20040
rect 14829 19975 14887 19981
rect 14829 19972 14841 19975
rect 14384 19944 14841 19972
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4724 19876 5181 19904
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 2958 19768 2964 19780
rect 2898 19740 2964 19768
rect 2958 19728 2964 19740
rect 3016 19728 3022 19780
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 4724 19768 4752 19876
rect 5169 19873 5181 19876
rect 5215 19873 5227 19907
rect 7098 19904 7104 19916
rect 5169 19867 5227 19873
rect 6288 19876 7104 19904
rect 4798 19796 4804 19848
rect 4856 19796 4862 19848
rect 4890 19796 4896 19848
rect 4948 19796 4954 19848
rect 6288 19845 6316 19876
rect 7098 19864 7104 19876
rect 7156 19904 7162 19916
rect 7193 19907 7251 19913
rect 7193 19904 7205 19907
rect 7156 19876 7205 19904
rect 7156 19864 7162 19876
rect 7193 19873 7205 19876
rect 7239 19904 7251 19907
rect 7929 19907 7987 19913
rect 7929 19904 7941 19907
rect 7239 19876 7941 19904
rect 7239 19873 7251 19876
rect 7193 19867 7251 19873
rect 7929 19873 7941 19876
rect 7975 19904 7987 19907
rect 8018 19904 8024 19916
rect 7975 19876 8024 19904
rect 7975 19873 7987 19876
rect 7929 19867 7987 19873
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 8110 19864 8116 19916
rect 8168 19864 8174 19916
rect 11238 19864 11244 19916
rect 11296 19864 11302 19916
rect 13630 19864 13636 19916
rect 13688 19864 13694 19916
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19805 6331 19839
rect 6273 19799 6331 19805
rect 6457 19839 6515 19845
rect 6457 19805 6469 19839
rect 6503 19805 6515 19839
rect 6457 19799 6515 19805
rect 4304 19740 4752 19768
rect 4908 19768 4936 19796
rect 5368 19768 5396 19799
rect 6472 19768 6500 19799
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 7285 19839 7343 19845
rect 7285 19836 7297 19839
rect 6880 19808 7297 19836
rect 6880 19796 6886 19808
rect 7285 19805 7297 19808
rect 7331 19836 7343 19839
rect 10410 19836 10416 19848
rect 7331 19808 10416 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19836 11575 19839
rect 12342 19836 12348 19848
rect 11563 19808 12348 19836
rect 11563 19805 11575 19808
rect 11517 19799 11575 19805
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 13998 19836 14004 19848
rect 13955 19808 14004 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 13998 19796 14004 19808
rect 14056 19796 14062 19848
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 6638 19768 6644 19780
rect 4908 19740 6644 19768
rect 4304 19728 4310 19740
rect 6638 19728 6644 19740
rect 6696 19768 6702 19780
rect 7009 19771 7067 19777
rect 7009 19768 7021 19771
rect 6696 19740 7021 19768
rect 6696 19728 6702 19740
rect 7009 19737 7021 19740
rect 7055 19737 7067 19771
rect 7009 19731 7067 19737
rect 7837 19771 7895 19777
rect 7837 19737 7849 19771
rect 7883 19768 7895 19771
rect 8294 19768 8300 19780
rect 7883 19740 8300 19768
rect 7883 19737 7895 19740
rect 7837 19731 7895 19737
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 9030 19728 9036 19780
rect 9088 19768 9094 19780
rect 9769 19771 9827 19777
rect 9769 19768 9781 19771
rect 9088 19740 9781 19768
rect 9088 19728 9094 19740
rect 9769 19737 9781 19740
rect 9815 19737 9827 19771
rect 13722 19768 13728 19780
rect 13202 19740 13728 19768
rect 9769 19731 9827 19737
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 14108 19768 14136 19799
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14240 19808 14289 19836
rect 14240 19796 14246 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14384 19836 14412 19944
rect 14829 19941 14841 19944
rect 14875 19941 14887 19975
rect 14829 19935 14887 19941
rect 14918 19932 14924 19984
rect 14976 19972 14982 19984
rect 16666 19972 16672 19984
rect 14976 19944 16672 19972
rect 14976 19932 14982 19944
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 17954 19932 17960 19984
rect 18012 19972 18018 19984
rect 18138 19972 18144 19984
rect 18012 19944 18144 19972
rect 18012 19932 18018 19944
rect 18138 19932 18144 19944
rect 18196 19972 18202 19984
rect 19429 19975 19487 19981
rect 19429 19972 19441 19975
rect 18196 19944 19441 19972
rect 18196 19932 18202 19944
rect 19429 19941 19441 19944
rect 19475 19972 19487 19975
rect 20530 19972 20536 19984
rect 19475 19944 20536 19972
rect 19475 19941 19487 19944
rect 19429 19935 19487 19941
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 20622 19932 20628 19984
rect 20680 19972 20686 19984
rect 21174 19972 21180 19984
rect 20680 19944 21180 19972
rect 20680 19932 20686 19944
rect 21174 19932 21180 19944
rect 21232 19932 21238 19984
rect 23658 19932 23664 19984
rect 23716 19972 23722 19984
rect 25866 19972 25872 19984
rect 23716 19944 25872 19972
rect 23716 19932 23722 19944
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 14384 19808 14473 19836
rect 14277 19799 14335 19805
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 14737 19839 14795 19845
rect 14737 19836 14749 19839
rect 14700 19808 14749 19836
rect 14700 19796 14706 19808
rect 14737 19805 14749 19808
rect 14783 19836 14795 19839
rect 14826 19836 14832 19848
rect 14783 19808 14832 19836
rect 14783 19805 14795 19808
rect 14737 19799 14795 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 14936 19845 14964 19932
rect 16393 19907 16451 19913
rect 15212 19876 15700 19904
rect 15212 19848 15240 19876
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 15562 19836 15568 19848
rect 15335 19808 15568 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15672 19836 15700 19876
rect 16393 19873 16405 19907
rect 16439 19904 16451 19907
rect 16439 19876 23796 19904
rect 16439 19873 16451 19876
rect 16393 19867 16451 19873
rect 16298 19845 16304 19848
rect 16289 19839 16304 19845
rect 16289 19836 16301 19839
rect 15672 19808 16301 19836
rect 16289 19805 16301 19808
rect 16289 19799 16304 19805
rect 16298 19796 16304 19799
rect 16356 19796 16362 19848
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19805 16543 19839
rect 16485 19799 16543 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 14369 19771 14427 19777
rect 14108 19740 14228 19768
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 6270 19700 6276 19712
rect 3936 19672 6276 19700
rect 3936 19660 3942 19672
rect 6270 19660 6276 19672
rect 6328 19660 6334 19712
rect 7098 19660 7104 19712
rect 7156 19700 7162 19712
rect 10042 19700 10048 19712
rect 7156 19672 10048 19700
rect 7156 19660 7162 19672
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 11241 19703 11299 19709
rect 11241 19669 11253 19703
rect 11287 19700 11299 19703
rect 11974 19700 11980 19712
rect 11287 19672 11980 19700
rect 11287 19669 11299 19672
rect 11241 19663 11299 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14200 19700 14228 19740
rect 14369 19737 14381 19771
rect 14415 19768 14427 19771
rect 15746 19768 15752 19780
rect 14415 19740 15752 19768
rect 14415 19737 14427 19740
rect 14369 19731 14427 19737
rect 15746 19728 15752 19740
rect 15804 19768 15810 19780
rect 16500 19768 16528 19799
rect 15804 19740 16528 19768
rect 17052 19768 17080 19799
rect 17218 19796 17224 19848
rect 17276 19796 17282 19848
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 17862 19836 17868 19848
rect 17552 19808 17868 19836
rect 17552 19796 17558 19808
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 23658 19836 23664 19848
rect 18564 19808 23664 19836
rect 18564 19796 18570 19808
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 23768 19845 23796 19876
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19836 23903 19839
rect 23952 19836 23980 19944
rect 25866 19932 25872 19944
rect 25924 19932 25930 19984
rect 27908 19981 27936 20012
rect 29822 20000 29828 20012
rect 29880 20000 29886 20052
rect 29914 20000 29920 20052
rect 29972 20040 29978 20052
rect 31481 20043 31539 20049
rect 31481 20040 31493 20043
rect 29972 20012 31493 20040
rect 29972 20000 29978 20012
rect 31481 20009 31493 20012
rect 31527 20040 31539 20043
rect 31662 20040 31668 20052
rect 31527 20012 31668 20040
rect 31527 20009 31539 20012
rect 31481 20003 31539 20009
rect 31662 20000 31668 20012
rect 31720 20000 31726 20052
rect 35342 20000 35348 20052
rect 35400 20040 35406 20052
rect 35526 20040 35532 20052
rect 35400 20012 35532 20040
rect 35400 20000 35406 20012
rect 35526 20000 35532 20012
rect 35584 20000 35590 20052
rect 27893 19975 27951 19981
rect 27893 19941 27905 19975
rect 27939 19941 27951 19975
rect 28258 19972 28264 19984
rect 27893 19935 27951 19941
rect 28092 19944 28264 19972
rect 25406 19864 25412 19916
rect 25464 19864 25470 19916
rect 27706 19864 27712 19916
rect 27764 19904 27770 19916
rect 28092 19913 28120 19944
rect 28258 19932 28264 19944
rect 28316 19932 28322 19984
rect 27985 19907 28043 19913
rect 27985 19904 27997 19907
rect 27764 19876 27997 19904
rect 27764 19864 27770 19876
rect 27985 19873 27997 19876
rect 28031 19873 28043 19907
rect 27985 19867 28043 19873
rect 28077 19907 28135 19913
rect 28077 19873 28089 19907
rect 28123 19873 28135 19907
rect 28077 19867 28135 19873
rect 28276 19876 31754 19904
rect 23891 19808 23980 19836
rect 24029 19839 24087 19845
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 24029 19805 24041 19839
rect 24075 19836 24087 19839
rect 24210 19836 24216 19848
rect 24075 19808 24216 19836
rect 24075 19805 24087 19808
rect 24029 19799 24087 19805
rect 18046 19768 18052 19780
rect 17052 19740 18052 19768
rect 15804 19728 15810 19740
rect 18046 19728 18052 19740
rect 18104 19728 18110 19780
rect 19794 19728 19800 19780
rect 19852 19728 19858 19780
rect 20073 19771 20131 19777
rect 20073 19737 20085 19771
rect 20119 19737 20131 19771
rect 20073 19731 20131 19737
rect 20257 19771 20315 19777
rect 20257 19737 20269 19771
rect 20303 19768 20315 19771
rect 20806 19768 20812 19780
rect 20303 19740 20812 19768
rect 20303 19737 20315 19740
rect 20257 19731 20315 19737
rect 14826 19700 14832 19712
rect 13872 19672 14832 19700
rect 13872 19660 13878 19672
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 19597 19703 19655 19709
rect 19597 19669 19609 19703
rect 19643 19700 19655 19703
rect 19702 19700 19708 19712
rect 19643 19672 19708 19700
rect 19643 19669 19655 19672
rect 19597 19663 19655 19669
rect 19702 19660 19708 19672
rect 19760 19660 19766 19712
rect 20088 19700 20116 19731
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 21174 19728 21180 19780
rect 21232 19768 21238 19780
rect 21634 19768 21640 19780
rect 21232 19740 21640 19768
rect 21232 19728 21238 19740
rect 21634 19728 21640 19740
rect 21692 19768 21698 19780
rect 23771 19768 23799 19799
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 24394 19796 24400 19848
rect 24452 19796 24458 19848
rect 24578 19796 24584 19848
rect 24636 19796 24642 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19836 24915 19839
rect 24946 19836 24952 19848
rect 24903 19808 24952 19836
rect 24903 19805 24915 19808
rect 24857 19799 24915 19805
rect 24946 19796 24952 19808
rect 25004 19796 25010 19848
rect 26234 19796 26240 19848
rect 26292 19836 26298 19848
rect 26697 19839 26755 19845
rect 26697 19836 26709 19839
rect 26292 19808 26709 19836
rect 26292 19796 26298 19808
rect 26697 19805 26709 19808
rect 26743 19805 26755 19839
rect 26697 19799 26755 19805
rect 26878 19796 26884 19848
rect 26936 19796 26942 19848
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 28276 19845 28304 19876
rect 27801 19839 27859 19845
rect 27801 19836 27813 19839
rect 27580 19808 27813 19836
rect 27580 19796 27586 19808
rect 27801 19805 27813 19808
rect 27847 19805 27859 19839
rect 27801 19799 27859 19805
rect 28261 19839 28319 19845
rect 28261 19805 28273 19839
rect 28307 19805 28319 19839
rect 28261 19799 28319 19805
rect 29730 19796 29736 19848
rect 29788 19836 29794 19848
rect 30466 19836 30472 19848
rect 29788 19808 30472 19836
rect 29788 19796 29794 19808
rect 30466 19796 30472 19808
rect 30524 19796 30530 19848
rect 31294 19796 31300 19848
rect 31352 19796 31358 19848
rect 31726 19836 31754 19876
rect 34698 19836 34704 19848
rect 31726 19808 34704 19836
rect 34698 19796 34704 19808
rect 34756 19796 34762 19848
rect 25222 19768 25228 19780
rect 21692 19740 21956 19768
rect 23771 19740 25228 19768
rect 21692 19728 21698 19740
rect 21082 19700 21088 19712
rect 20088 19672 21088 19700
rect 21082 19660 21088 19672
rect 21140 19660 21146 19712
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21818 19700 21824 19712
rect 21324 19672 21824 19700
rect 21324 19660 21330 19672
rect 21818 19660 21824 19672
rect 21876 19660 21882 19712
rect 21928 19700 21956 19740
rect 25222 19728 25228 19740
rect 25280 19728 25286 19780
rect 32674 19768 32680 19780
rect 27632 19740 32680 19768
rect 25774 19700 25780 19712
rect 21928 19672 25780 19700
rect 25774 19660 25780 19672
rect 25832 19660 25838 19712
rect 26510 19660 26516 19712
rect 26568 19660 26574 19712
rect 27632 19709 27660 19740
rect 32674 19728 32680 19740
rect 32732 19728 32738 19780
rect 27617 19703 27675 19709
rect 27617 19669 27629 19703
rect 27663 19669 27675 19703
rect 27617 19663 27675 19669
rect 28718 19660 28724 19712
rect 28776 19700 28782 19712
rect 31294 19700 31300 19712
rect 28776 19672 31300 19700
rect 28776 19660 28782 19672
rect 31294 19660 31300 19672
rect 31352 19700 31358 19712
rect 34422 19700 34428 19712
rect 31352 19672 34428 19700
rect 31352 19660 31358 19672
rect 34422 19660 34428 19672
rect 34480 19660 34486 19712
rect 1104 19610 36524 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 36524 19610
rect 1104 19536 36524 19558
rect 2682 19456 2688 19508
rect 2740 19496 2746 19508
rect 8478 19496 8484 19508
rect 2740 19468 8484 19496
rect 2740 19456 2746 19468
rect 8478 19456 8484 19468
rect 8536 19456 8542 19508
rect 9398 19456 9404 19508
rect 9456 19496 9462 19508
rect 10321 19499 10379 19505
rect 10321 19496 10333 19499
rect 9456 19468 10333 19496
rect 9456 19456 9462 19468
rect 10321 19465 10333 19468
rect 10367 19465 10379 19499
rect 10321 19459 10379 19465
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 13725 19499 13783 19505
rect 13725 19496 13737 19499
rect 10468 19468 13737 19496
rect 10468 19456 10474 19468
rect 13725 19465 13737 19468
rect 13771 19465 13783 19499
rect 13725 19459 13783 19465
rect 17218 19456 17224 19508
rect 17276 19496 17282 19508
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 17276 19468 17325 19496
rect 17276 19456 17282 19468
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 18322 19496 18328 19508
rect 17313 19459 17371 19465
rect 17788 19468 18328 19496
rect 3234 19388 3240 19440
rect 3292 19388 3298 19440
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 5166 19428 5172 19440
rect 3476 19400 5172 19428
rect 3476 19388 3482 19400
rect 5166 19388 5172 19400
rect 5224 19388 5230 19440
rect 10042 19428 10048 19440
rect 9982 19400 10048 19428
rect 10042 19388 10048 19400
rect 10100 19388 10106 19440
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 11480 19400 12173 19428
rect 11480 19388 11486 19400
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 12342 19388 12348 19440
rect 12400 19388 12406 19440
rect 13538 19388 13544 19440
rect 13596 19428 13602 19440
rect 16574 19428 16580 19440
rect 13596 19400 16580 19428
rect 13596 19388 13602 19400
rect 16574 19388 16580 19400
rect 16632 19388 16638 19440
rect 17586 19428 17592 19440
rect 17052 19400 17592 19428
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19360 3203 19363
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 3191 19332 3617 19360
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 3605 19329 3617 19332
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 4246 19320 4252 19372
rect 4304 19320 4310 19372
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5258 19360 5264 19372
rect 4764 19332 5264 19360
rect 4764 19320 4770 19332
rect 5258 19320 5264 19332
rect 5316 19360 5322 19372
rect 5353 19363 5411 19369
rect 5353 19360 5365 19363
rect 5316 19332 5365 19360
rect 5316 19320 5322 19332
rect 5353 19329 5365 19332
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 8481 19363 8539 19369
rect 8481 19360 8493 19363
rect 7064 19332 8493 19360
rect 7064 19320 7070 19332
rect 8481 19329 8493 19332
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 10744 19332 11560 19360
rect 10744 19320 10750 19332
rect 2958 19252 2964 19304
rect 3016 19292 3022 19304
rect 3329 19295 3387 19301
rect 3329 19292 3341 19295
rect 3016 19264 3341 19292
rect 3016 19252 3022 19264
rect 3329 19261 3341 19264
rect 3375 19261 3387 19295
rect 3329 19255 3387 19261
rect 8754 19252 8760 19304
rect 8812 19252 8818 19304
rect 10229 19295 10287 19301
rect 10229 19261 10241 19295
rect 10275 19292 10287 19295
rect 10318 19292 10324 19304
rect 10275 19264 10324 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 10318 19252 10324 19264
rect 10376 19292 10382 19304
rect 10873 19295 10931 19301
rect 10873 19292 10885 19295
rect 10376 19264 10885 19292
rect 10376 19252 10382 19264
rect 10873 19261 10885 19264
rect 10919 19261 10931 19295
rect 10873 19255 10931 19261
rect 3694 19184 3700 19236
rect 3752 19224 3758 19236
rect 8386 19224 8392 19236
rect 3752 19196 8392 19224
rect 3752 19184 3758 19196
rect 8386 19184 8392 19196
rect 8444 19184 8450 19236
rect 11532 19233 11560 19332
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19329 11851 19363
rect 11793 19323 11851 19329
rect 11808 19292 11836 19323
rect 11882 19320 11888 19372
rect 11940 19320 11946 19372
rect 12066 19320 12072 19372
rect 12124 19320 12130 19372
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 16482 19360 16488 19372
rect 13955 19332 16488 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 17052 19369 17080 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17037 19363 17095 19369
rect 17037 19329 17049 19363
rect 17083 19329 17095 19363
rect 17788 19360 17816 19468
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 18785 19499 18843 19505
rect 18785 19465 18797 19499
rect 18831 19496 18843 19499
rect 19426 19496 19432 19508
rect 18831 19468 19432 19496
rect 18831 19465 18843 19468
rect 18785 19459 18843 19465
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21542 19496 21548 19508
rect 20864 19468 21548 19496
rect 20864 19456 20870 19468
rect 21542 19456 21548 19468
rect 21600 19456 21606 19508
rect 23750 19456 23756 19508
rect 23808 19456 23814 19508
rect 24394 19456 24400 19508
rect 24452 19496 24458 19508
rect 24489 19499 24547 19505
rect 24489 19496 24501 19499
rect 24452 19468 24501 19496
rect 24452 19456 24458 19468
rect 24489 19465 24501 19468
rect 24535 19465 24547 19499
rect 24489 19459 24547 19465
rect 24762 19456 24768 19508
rect 24820 19496 24826 19508
rect 25041 19499 25099 19505
rect 25041 19496 25053 19499
rect 24820 19468 25053 19496
rect 24820 19456 24826 19468
rect 25041 19465 25053 19468
rect 25087 19465 25099 19499
rect 25041 19459 25099 19465
rect 27430 19456 27436 19508
rect 27488 19496 27494 19508
rect 27706 19496 27712 19508
rect 27488 19468 27712 19496
rect 27488 19456 27494 19468
rect 27706 19456 27712 19468
rect 27764 19456 27770 19508
rect 28905 19499 28963 19505
rect 28905 19465 28917 19499
rect 28951 19496 28963 19499
rect 30101 19499 30159 19505
rect 28951 19468 29868 19496
rect 28951 19465 28963 19468
rect 28905 19459 28963 19465
rect 18156 19400 19196 19428
rect 18156 19372 18184 19400
rect 17037 19323 17095 19329
rect 17604 19332 17816 19360
rect 12618 19292 12624 19304
rect 11808 19264 12624 19292
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 14093 19295 14151 19301
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14642 19292 14648 19304
rect 14139 19264 14648 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 16868 19292 16896 19323
rect 17402 19292 17408 19304
rect 16868 19264 17408 19292
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 11517 19227 11575 19233
rect 11517 19193 11529 19227
rect 11563 19193 11575 19227
rect 11517 19187 11575 19193
rect 2774 19116 2780 19168
rect 2832 19116 2838 19168
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 4672 19128 4813 19156
rect 4672 19116 4678 19128
rect 4801 19125 4813 19128
rect 4847 19125 4859 19159
rect 4801 19119 4859 19125
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 12529 19159 12587 19165
rect 12529 19156 12541 19159
rect 12216 19128 12541 19156
rect 12216 19116 12222 19128
rect 12529 19125 12541 19128
rect 12575 19125 12587 19159
rect 12529 19119 12587 19125
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17604 19165 17632 19332
rect 17862 19320 17868 19372
rect 17920 19320 17926 19372
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 18027 19332 18061 19360
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 17773 19295 17831 19301
rect 17773 19261 17785 19295
rect 17819 19292 17831 19295
rect 17954 19292 17960 19304
rect 17819 19264 17960 19292
rect 17819 19261 17831 19264
rect 17773 19255 17831 19261
rect 17954 19252 17960 19264
rect 18012 19252 18018 19304
rect 18064 19224 18092 19323
rect 18138 19320 18144 19372
rect 18196 19320 18202 19372
rect 18322 19369 18328 19372
rect 18289 19363 18328 19369
rect 18289 19329 18301 19363
rect 18289 19323 18328 19329
rect 18322 19320 18328 19323
rect 18380 19320 18386 19372
rect 18417 19363 18475 19369
rect 18417 19329 18429 19363
rect 18463 19329 18475 19363
rect 18417 19323 18475 19329
rect 18138 19224 18144 19236
rect 18064 19196 18144 19224
rect 18138 19184 18144 19196
rect 18196 19184 18202 19236
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 18432 19224 18460 19323
rect 18506 19320 18512 19372
rect 18564 19320 18570 19372
rect 18647 19363 18705 19369
rect 18647 19329 18659 19363
rect 18693 19360 18705 19363
rect 18782 19360 18788 19372
rect 18693 19332 18788 19360
rect 18693 19329 18705 19332
rect 18647 19323 18705 19329
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 18874 19320 18880 19372
rect 18932 19320 18938 19372
rect 19058 19320 19064 19372
rect 19116 19320 19122 19372
rect 19168 19369 19196 19400
rect 19242 19388 19248 19440
rect 19300 19428 19306 19440
rect 20824 19428 20852 19456
rect 19300 19400 20852 19428
rect 19300 19388 19306 19400
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19260 19304 19288 19388
rect 19518 19360 19524 19372
rect 19352 19332 19524 19360
rect 19242 19252 19248 19304
rect 19300 19252 19306 19304
rect 19352 19233 19380 19332
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 20530 19320 20536 19372
rect 20588 19320 20594 19372
rect 20824 19369 20852 19400
rect 20898 19388 20904 19440
rect 20956 19428 20962 19440
rect 21726 19428 21732 19440
rect 20956 19400 21732 19428
rect 20956 19388 20962 19400
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19329 20867 19363
rect 20809 19323 20867 19329
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19329 21051 19363
rect 21192 19360 21220 19400
rect 21726 19388 21732 19400
rect 21784 19388 21790 19440
rect 22830 19388 22836 19440
rect 22888 19428 22894 19440
rect 25314 19428 25320 19440
rect 22888 19400 25320 19428
rect 22888 19388 22894 19400
rect 24249 19372 24277 19400
rect 21252 19363 21310 19369
rect 21252 19360 21264 19363
rect 21192 19332 21264 19360
rect 20993 19323 21051 19329
rect 21252 19329 21264 19332
rect 21298 19329 21310 19363
rect 21252 19323 21310 19329
rect 21361 19363 21419 19369
rect 21361 19329 21373 19363
rect 21407 19360 21419 19363
rect 21450 19360 21456 19372
rect 21407 19332 21456 19360
rect 21407 19329 21419 19332
rect 21361 19323 21419 19329
rect 20257 19295 20315 19301
rect 20257 19261 20269 19295
rect 20303 19292 20315 19295
rect 20622 19292 20628 19304
rect 20303 19264 20628 19292
rect 20303 19261 20315 19264
rect 20257 19255 20315 19261
rect 20622 19252 20628 19264
rect 20680 19252 20686 19304
rect 18288 19196 18460 19224
rect 19337 19227 19395 19233
rect 18288 19184 18294 19196
rect 19337 19193 19349 19227
rect 19383 19193 19395 19227
rect 21008 19224 21036 19323
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 21637 19363 21695 19369
rect 21637 19329 21649 19363
rect 21683 19360 21695 19363
rect 21818 19360 21824 19372
rect 21683 19332 21824 19360
rect 21683 19329 21695 19332
rect 21637 19323 21695 19329
rect 21818 19320 21824 19332
rect 21876 19320 21882 19372
rect 23934 19320 23940 19372
rect 23992 19360 23998 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23992 19332 24041 19360
rect 23992 19320 23998 19332
rect 24029 19329 24041 19332
rect 24075 19329 24087 19363
rect 24029 19323 24087 19329
rect 24134 19363 24192 19369
rect 24134 19329 24146 19363
rect 24180 19329 24192 19363
rect 24134 19323 24192 19329
rect 24234 19366 24292 19372
rect 24234 19332 24246 19366
rect 24280 19332 24292 19366
rect 24234 19326 24292 19332
rect 24136 19292 24164 19323
rect 24394 19320 24400 19372
rect 24452 19320 24458 19372
rect 24486 19320 24492 19372
rect 24544 19320 24550 19372
rect 24688 19369 24716 19400
rect 25314 19388 25320 19400
rect 25372 19388 25378 19440
rect 25590 19388 25596 19440
rect 25648 19428 25654 19440
rect 27617 19431 27675 19437
rect 27617 19428 27629 19431
rect 25648 19400 27629 19428
rect 25648 19388 25654 19400
rect 27617 19397 27629 19400
rect 27663 19397 27675 19431
rect 27617 19391 27675 19397
rect 28276 19400 29500 19428
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19329 24731 19363
rect 24673 19323 24731 19329
rect 24854 19320 24860 19372
rect 24912 19320 24918 19372
rect 24949 19363 25007 19369
rect 24949 19329 24961 19363
rect 24995 19360 25007 19363
rect 25038 19360 25044 19372
rect 24995 19332 25044 19360
rect 24995 19329 25007 19332
rect 24949 19323 25007 19329
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 25222 19320 25228 19372
rect 25280 19320 25286 19372
rect 25406 19320 25412 19372
rect 25464 19320 25470 19372
rect 25498 19320 25504 19372
rect 25556 19320 25562 19372
rect 25774 19320 25780 19372
rect 25832 19360 25838 19372
rect 26053 19363 26111 19369
rect 26053 19360 26065 19363
rect 25832 19332 26065 19360
rect 25832 19320 25838 19332
rect 26053 19329 26065 19332
rect 26099 19329 26111 19363
rect 26053 19323 26111 19329
rect 26878 19320 26884 19372
rect 26936 19360 26942 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26936 19332 27169 19360
rect 26936 19320 26942 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 27982 19320 27988 19372
rect 28040 19360 28046 19372
rect 28276 19369 28304 19400
rect 28261 19363 28319 19369
rect 28261 19360 28273 19363
rect 28040 19332 28273 19360
rect 28040 19320 28046 19332
rect 28261 19329 28273 19332
rect 28307 19329 28319 19363
rect 28261 19323 28319 19329
rect 28350 19320 28356 19372
rect 28408 19360 28414 19372
rect 28537 19363 28595 19369
rect 28537 19360 28549 19363
rect 28408 19332 28453 19360
rect 28515 19332 28549 19360
rect 28408 19320 28414 19332
rect 28537 19329 28549 19332
rect 28583 19329 28595 19363
rect 28537 19323 28595 19329
rect 28629 19363 28687 19369
rect 28629 19329 28641 19363
rect 28675 19329 28687 19363
rect 28629 19323 28687 19329
rect 24504 19292 24532 19320
rect 24136 19264 24532 19292
rect 25130 19252 25136 19304
rect 25188 19292 25194 19304
rect 26145 19295 26203 19301
rect 26145 19292 26157 19295
rect 25188 19264 26157 19292
rect 25188 19252 25194 19264
rect 26145 19261 26157 19264
rect 26191 19261 26203 19295
rect 26145 19255 26203 19261
rect 27246 19252 27252 19304
rect 27304 19252 27310 19304
rect 27890 19252 27896 19304
rect 27948 19292 27954 19304
rect 28166 19292 28172 19304
rect 27948 19264 28172 19292
rect 27948 19252 27954 19264
rect 28166 19252 28172 19264
rect 28224 19292 28230 19304
rect 28552 19292 28580 19323
rect 28224 19264 28580 19292
rect 28224 19252 28230 19264
rect 21450 19224 21456 19236
rect 21008 19196 21456 19224
rect 19337 19187 19395 19193
rect 21450 19184 21456 19196
rect 21508 19184 21514 19236
rect 23474 19184 23480 19236
rect 23532 19224 23538 19236
rect 26234 19224 26240 19236
rect 23532 19196 26240 19224
rect 23532 19184 23538 19196
rect 26234 19184 26240 19196
rect 26292 19184 26298 19236
rect 26326 19184 26332 19236
rect 26384 19224 26390 19236
rect 26973 19227 27031 19233
rect 26973 19224 26985 19227
rect 26384 19196 26985 19224
rect 26384 19184 26390 19196
rect 26973 19193 26985 19196
rect 27019 19193 27031 19227
rect 26973 19187 27031 19193
rect 28534 19184 28540 19236
rect 28592 19224 28598 19236
rect 28644 19224 28672 19323
rect 28718 19320 28724 19372
rect 28776 19369 28782 19372
rect 29472 19369 29500 19400
rect 29730 19388 29736 19440
rect 29788 19388 29794 19440
rect 29840 19428 29868 19468
rect 30101 19465 30113 19499
rect 30147 19496 30159 19499
rect 30742 19496 30748 19508
rect 30147 19468 30748 19496
rect 30147 19465 30159 19468
rect 30101 19459 30159 19465
rect 30742 19456 30748 19468
rect 30800 19456 30806 19508
rect 30837 19499 30895 19505
rect 30837 19465 30849 19499
rect 30883 19496 30895 19499
rect 32122 19496 32128 19508
rect 30883 19468 32128 19496
rect 30883 19465 30895 19468
rect 30837 19459 30895 19465
rect 32122 19456 32128 19468
rect 32180 19456 32186 19508
rect 29840 19400 30236 19428
rect 30208 19372 30236 19400
rect 30466 19388 30472 19440
rect 30524 19388 30530 19440
rect 31294 19388 31300 19440
rect 31352 19388 31358 19440
rect 28776 19360 28784 19369
rect 29457 19363 29515 19369
rect 28776 19332 28821 19360
rect 28776 19323 28784 19332
rect 29457 19329 29469 19363
rect 29503 19329 29515 19363
rect 29457 19323 29515 19329
rect 28776 19320 28782 19323
rect 29546 19320 29552 19372
rect 29604 19360 29610 19372
rect 29825 19363 29883 19369
rect 29825 19360 29837 19363
rect 29604 19332 29649 19360
rect 29722 19332 29837 19360
rect 29604 19320 29610 19332
rect 29178 19252 29184 19304
rect 29236 19292 29242 19304
rect 29722 19292 29750 19332
rect 29825 19329 29837 19332
rect 29871 19329 29883 19363
rect 29825 19323 29883 19329
rect 29914 19320 29920 19372
rect 29972 19369 29978 19372
rect 29972 19360 29980 19369
rect 29972 19332 30017 19360
rect 29972 19323 29980 19332
rect 29972 19320 29978 19323
rect 30190 19320 30196 19372
rect 30248 19320 30254 19372
rect 30282 19320 30288 19372
rect 30340 19360 30346 19372
rect 30561 19363 30619 19369
rect 30340 19332 30385 19360
rect 30340 19320 30346 19332
rect 30561 19329 30573 19363
rect 30607 19329 30619 19363
rect 30561 19323 30619 19329
rect 30699 19363 30757 19369
rect 30699 19329 30711 19363
rect 30745 19360 30757 19363
rect 31312 19360 31340 19388
rect 30745 19332 31340 19360
rect 30745 19329 30757 19332
rect 30699 19323 30757 19329
rect 30576 19292 30604 19323
rect 29236 19264 30604 19292
rect 29236 19252 29242 19264
rect 28592 19196 28672 19224
rect 28592 19184 28598 19196
rect 32490 19184 32496 19236
rect 32548 19224 32554 19236
rect 33042 19224 33048 19236
rect 32548 19196 33048 19224
rect 32548 19184 32554 19196
rect 33042 19184 33048 19196
rect 33100 19184 33106 19236
rect 17589 19159 17647 19165
rect 17589 19156 17601 19159
rect 17000 19128 17601 19156
rect 17000 19116 17006 19128
rect 17589 19125 17601 19128
rect 17635 19125 17647 19159
rect 17589 19119 17647 19125
rect 17681 19159 17739 19165
rect 17681 19125 17693 19159
rect 17727 19156 17739 19159
rect 18322 19156 18328 19168
rect 17727 19128 18328 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 18322 19116 18328 19128
rect 18380 19156 18386 19168
rect 18877 19159 18935 19165
rect 18877 19156 18889 19159
rect 18380 19128 18889 19156
rect 18380 19116 18386 19128
rect 18877 19125 18889 19128
rect 18923 19125 18935 19159
rect 18877 19119 18935 19125
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20625 19159 20683 19165
rect 20625 19156 20637 19159
rect 20128 19128 20637 19156
rect 20128 19116 20134 19128
rect 20625 19125 20637 19128
rect 20671 19125 20683 19159
rect 20625 19119 20683 19125
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 21085 19159 21143 19165
rect 21085 19156 21097 19159
rect 20763 19128 21097 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 21085 19125 21097 19128
rect 21131 19125 21143 19159
rect 21085 19119 21143 19125
rect 21545 19159 21603 19165
rect 21545 19125 21557 19159
rect 21591 19156 21603 19159
rect 22094 19156 22100 19168
rect 21591 19128 22100 19156
rect 21591 19125 21603 19128
rect 21545 19119 21603 19125
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 24394 19116 24400 19168
rect 24452 19156 24458 19168
rect 26050 19156 26056 19168
rect 24452 19128 26056 19156
rect 24452 19116 24458 19128
rect 26050 19116 26056 19128
rect 26108 19116 26114 19168
rect 26142 19116 26148 19168
rect 26200 19116 26206 19168
rect 26418 19116 26424 19168
rect 26476 19116 26482 19168
rect 27154 19116 27160 19168
rect 27212 19156 27218 19168
rect 27522 19156 27528 19168
rect 27212 19128 27528 19156
rect 27212 19116 27218 19128
rect 27522 19116 27528 19128
rect 27580 19116 27586 19168
rect 27614 19116 27620 19168
rect 27672 19156 27678 19168
rect 34514 19156 34520 19168
rect 27672 19128 34520 19156
rect 27672 19116 27678 19128
rect 34514 19116 34520 19128
rect 34572 19116 34578 19168
rect 1104 19066 36524 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 36524 19066
rect 1104 18992 36524 19014
rect 3605 18955 3663 18961
rect 3605 18921 3617 18955
rect 3651 18952 3663 18955
rect 4062 18952 4068 18964
rect 3651 18924 4068 18952
rect 3651 18921 3663 18924
rect 3605 18915 3663 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 5534 18952 5540 18964
rect 5224 18924 5540 18952
rect 5224 18912 5230 18924
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 6549 18955 6607 18961
rect 6549 18921 6561 18955
rect 6595 18952 6607 18955
rect 6914 18952 6920 18964
rect 6595 18924 6920 18952
rect 6595 18921 6607 18924
rect 6549 18915 6607 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 7834 18912 7840 18964
rect 7892 18952 7898 18964
rect 7892 18924 8156 18952
rect 7892 18912 7898 18924
rect 6641 18887 6699 18893
rect 6641 18853 6653 18887
rect 6687 18853 6699 18887
rect 6932 18884 6960 18912
rect 8128 18884 8156 18924
rect 8294 18912 8300 18964
rect 8352 18912 8358 18964
rect 8570 18912 8576 18964
rect 8628 18912 8634 18964
rect 8754 18912 8760 18964
rect 8812 18952 8818 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8812 18924 8953 18952
rect 8812 18912 8818 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 9953 18955 10011 18961
rect 9953 18921 9965 18955
rect 9999 18952 10011 18955
rect 12066 18952 12072 18964
rect 9999 18924 12072 18952
rect 9999 18921 10011 18924
rect 9953 18915 10011 18921
rect 12066 18912 12072 18924
rect 12124 18912 12130 18964
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 17129 18955 17187 18961
rect 17129 18952 17141 18955
rect 16540 18924 17141 18952
rect 16540 18912 16546 18924
rect 17129 18921 17141 18924
rect 17175 18921 17187 18955
rect 17129 18915 17187 18921
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 18380 18924 19380 18952
rect 18380 18912 18386 18924
rect 10410 18884 10416 18896
rect 6932 18856 8064 18884
rect 8128 18856 10416 18884
rect 6641 18847 6699 18853
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 1857 18819 1915 18825
rect 1857 18816 1869 18819
rect 1452 18788 1869 18816
rect 1452 18776 1458 18788
rect 1857 18785 1869 18788
rect 1903 18816 1915 18819
rect 2682 18816 2688 18828
rect 1903 18788 2688 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 2682 18776 2688 18788
rect 2740 18816 2746 18828
rect 2740 18788 4384 18816
rect 2740 18776 2746 18788
rect 4356 18748 4384 18788
rect 4430 18776 4436 18828
rect 4488 18816 4494 18828
rect 4525 18819 4583 18825
rect 4525 18816 4537 18819
rect 4488 18788 4537 18816
rect 4488 18776 4494 18788
rect 4525 18785 4537 18788
rect 4571 18785 4583 18819
rect 4525 18779 4583 18785
rect 5077 18819 5135 18825
rect 5077 18785 5089 18819
rect 5123 18816 5135 18819
rect 6656 18816 6684 18847
rect 5123 18788 6684 18816
rect 5123 18785 5135 18788
rect 5077 18779 5135 18785
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7558 18816 7564 18828
rect 7340 18788 7564 18816
rect 7340 18776 7346 18788
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 8036 18825 8064 18856
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 16850 18844 16856 18896
rect 16908 18884 16914 18896
rect 17218 18884 17224 18896
rect 16908 18856 17224 18884
rect 16908 18844 16914 18856
rect 17218 18844 17224 18856
rect 17276 18844 17282 18896
rect 17310 18844 17316 18896
rect 17368 18884 17374 18896
rect 19245 18887 19303 18893
rect 17368 18856 18644 18884
rect 17368 18844 17374 18856
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 8444 18788 9352 18816
rect 8444 18776 8450 18788
rect 4706 18748 4712 18760
rect 4356 18720 4712 18748
rect 4706 18708 4712 18720
rect 4764 18748 4770 18760
rect 4801 18751 4859 18757
rect 4801 18748 4813 18751
rect 4764 18720 4813 18748
rect 4764 18708 4770 18720
rect 4801 18717 4813 18720
rect 4847 18717 4859 18751
rect 7098 18748 7104 18760
rect 6210 18734 7104 18748
rect 4801 18711 4859 18717
rect 6196 18720 7104 18734
rect 2133 18683 2191 18689
rect 2133 18649 2145 18683
rect 2179 18649 2191 18683
rect 3418 18680 3424 18692
rect 3358 18652 3424 18680
rect 2133 18643 2191 18649
rect 2148 18612 2176 18643
rect 3418 18640 3424 18652
rect 3476 18640 3482 18692
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 4341 18683 4399 18689
rect 3568 18652 4292 18680
rect 3568 18640 3574 18652
rect 2774 18612 2780 18624
rect 2148 18584 2780 18612
rect 2774 18572 2780 18584
rect 2832 18572 2838 18624
rect 3694 18572 3700 18624
rect 3752 18612 3758 18624
rect 3973 18615 4031 18621
rect 3973 18612 3985 18615
rect 3752 18584 3985 18612
rect 3752 18572 3758 18584
rect 3973 18581 3985 18584
rect 4019 18581 4031 18615
rect 4264 18612 4292 18652
rect 4341 18649 4353 18683
rect 4387 18680 4399 18683
rect 4614 18680 4620 18692
rect 4387 18652 4620 18680
rect 4387 18649 4399 18652
rect 4341 18643 4399 18649
rect 4614 18640 4620 18652
rect 4672 18640 4678 18692
rect 4433 18615 4491 18621
rect 4433 18612 4445 18615
rect 4264 18584 4445 18612
rect 3973 18575 4031 18581
rect 4433 18581 4445 18584
rect 4479 18612 4491 18615
rect 4522 18612 4528 18624
rect 4479 18584 4528 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 6196 18612 6224 18720
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8205 18751 8263 18757
rect 8205 18748 8217 18751
rect 8168 18720 8217 18748
rect 8168 18708 8174 18720
rect 8205 18717 8217 18720
rect 8251 18717 8263 18751
rect 8205 18711 8263 18717
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18748 8723 18751
rect 8754 18748 8760 18760
rect 8711 18720 8760 18748
rect 8711 18717 8723 18720
rect 8665 18711 8723 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 9324 18748 9352 18788
rect 9398 18776 9404 18828
rect 9456 18776 9462 18828
rect 9493 18819 9551 18825
rect 9493 18785 9505 18819
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 10965 18819 11023 18825
rect 10965 18785 10977 18819
rect 11011 18816 11023 18819
rect 11054 18816 11060 18828
rect 11011 18788 11060 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 9508 18748 9536 18779
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 11572 18788 11713 18816
rect 11572 18776 11578 18788
rect 11701 18785 11713 18788
rect 11747 18785 11759 18819
rect 11701 18779 11759 18785
rect 12250 18776 12256 18828
rect 12308 18816 12314 18828
rect 12437 18819 12495 18825
rect 12437 18816 12449 18819
rect 12308 18788 12449 18816
rect 12308 18776 12314 18788
rect 12437 18785 12449 18788
rect 12483 18785 12495 18819
rect 12437 18779 12495 18785
rect 12618 18776 12624 18828
rect 12676 18776 12682 18828
rect 17126 18776 17132 18828
rect 17184 18816 17190 18828
rect 18616 18825 18644 18856
rect 19245 18853 19257 18887
rect 19291 18853 19303 18887
rect 19245 18847 19303 18853
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 17184 18788 18061 18816
rect 17184 18776 17190 18788
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 18049 18779 18107 18785
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18966 18816 18972 18828
rect 18647 18788 18972 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18816 19119 18819
rect 19260 18816 19288 18847
rect 19107 18788 19288 18816
rect 19352 18816 19380 18924
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 19610 18912 19616 18964
rect 19668 18952 19674 18964
rect 19981 18955 20039 18961
rect 19981 18952 19993 18955
rect 19668 18924 19993 18952
rect 19668 18912 19674 18924
rect 19981 18921 19993 18924
rect 20027 18952 20039 18955
rect 22097 18955 22155 18961
rect 20027 18924 21588 18952
rect 20027 18921 20039 18924
rect 19981 18915 20039 18921
rect 20806 18844 20812 18896
rect 20864 18884 20870 18896
rect 21358 18884 21364 18896
rect 20864 18856 21364 18884
rect 20864 18844 20870 18856
rect 21358 18844 21364 18856
rect 21416 18844 21422 18896
rect 19352 18788 19656 18816
rect 19107 18785 19119 18788
rect 19061 18779 19119 18785
rect 10042 18748 10048 18760
rect 9324 18720 10048 18748
rect 10042 18708 10048 18720
rect 10100 18708 10106 18760
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18748 10287 18751
rect 10410 18748 10416 18760
rect 10275 18720 10416 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18748 10839 18751
rect 11238 18748 11244 18760
rect 10827 18720 11244 18748
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 11238 18708 11244 18720
rect 11296 18748 11302 18760
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 11296 18720 11621 18748
rect 11296 18708 11302 18720
rect 11609 18717 11621 18720
rect 11655 18748 11667 18751
rect 12066 18748 12072 18760
rect 11655 18720 12072 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 14090 18708 14096 18760
rect 14148 18708 14154 18760
rect 16574 18708 16580 18760
rect 16632 18708 16638 18760
rect 16850 18708 16856 18760
rect 16908 18708 16914 18760
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18726 17095 18751
rect 17083 18717 17172 18726
rect 17037 18711 17172 18717
rect 7009 18683 7067 18689
rect 7009 18649 7021 18683
rect 7055 18680 7067 18683
rect 7469 18683 7527 18689
rect 7469 18680 7481 18683
rect 7055 18652 7481 18680
rect 7055 18649 7067 18652
rect 7009 18643 7067 18649
rect 7469 18649 7481 18652
rect 7515 18649 7527 18683
rect 9766 18680 9772 18692
rect 7469 18643 7527 18649
rect 8312 18652 9772 18680
rect 5408 18584 6224 18612
rect 5408 18572 5414 18584
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 8312 18612 8340 18652
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 9950 18640 9956 18692
rect 10008 18640 10014 18692
rect 10689 18683 10747 18689
rect 10689 18649 10701 18683
rect 10735 18680 10747 18683
rect 11517 18683 11575 18689
rect 11517 18680 11529 18683
rect 10735 18652 11529 18680
rect 10735 18649 10747 18652
rect 10689 18643 10747 18649
rect 11517 18649 11529 18652
rect 11563 18680 11575 18683
rect 11698 18680 11704 18692
rect 11563 18652 11704 18680
rect 11563 18649 11575 18652
rect 11517 18643 11575 18649
rect 11698 18640 11704 18652
rect 11756 18640 11762 18692
rect 14366 18640 14372 18692
rect 14424 18640 14430 18692
rect 15378 18640 15384 18692
rect 15436 18640 15442 18692
rect 16592 18680 16620 18708
rect 17061 18698 17172 18711
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 17276 18720 17325 18748
rect 17276 18708 17282 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 17770 18748 17776 18760
rect 17460 18720 17776 18748
rect 17460 18708 17466 18720
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18748 18935 18751
rect 19242 18748 19248 18760
rect 18923 18720 19248 18748
rect 18923 18717 18935 18720
rect 18877 18711 18935 18717
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 15856 18652 16620 18680
rect 7156 18584 8340 18612
rect 7156 18572 7162 18584
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 8720 18584 9321 18612
rect 8720 18572 8726 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9309 18575 9367 18581
rect 10137 18615 10195 18621
rect 10137 18581 10149 18615
rect 10183 18612 10195 18615
rect 10226 18612 10232 18624
rect 10183 18584 10232 18612
rect 10183 18581 10195 18584
rect 10137 18575 10195 18581
rect 10226 18572 10232 18584
rect 10284 18572 10290 18624
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 11149 18615 11207 18621
rect 11149 18612 11161 18615
rect 10928 18584 11161 18612
rect 10928 18572 10934 18584
rect 11149 18581 11161 18584
rect 11195 18581 11207 18615
rect 11149 18575 11207 18581
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 11977 18615 12035 18621
rect 11977 18612 11989 18615
rect 11848 18584 11989 18612
rect 11848 18572 11854 18584
rect 11977 18581 11989 18584
rect 12023 18581 12035 18615
rect 11977 18575 12035 18581
rect 12342 18572 12348 18624
rect 12400 18572 12406 18624
rect 14090 18572 14096 18624
rect 14148 18612 14154 18624
rect 15010 18612 15016 18624
rect 14148 18584 15016 18612
rect 14148 18572 14154 18584
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15856 18621 15884 18652
rect 15841 18615 15899 18621
rect 15841 18581 15853 18615
rect 15887 18581 15899 18615
rect 15841 18575 15899 18581
rect 15930 18572 15936 18624
rect 15988 18572 15994 18624
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16669 18615 16727 18621
rect 16669 18612 16681 18615
rect 16080 18584 16681 18612
rect 16080 18572 16086 18584
rect 16669 18581 16681 18584
rect 16715 18581 16727 18615
rect 17144 18612 17172 18698
rect 18966 18640 18972 18692
rect 19024 18680 19030 18692
rect 19444 18680 19472 18711
rect 19518 18708 19524 18760
rect 19576 18708 19582 18760
rect 19024 18652 19472 18680
rect 19628 18680 19656 18788
rect 19702 18776 19708 18828
rect 19760 18776 19766 18828
rect 20346 18776 20352 18828
rect 20404 18816 20410 18828
rect 20622 18816 20628 18828
rect 20404 18788 20628 18816
rect 20404 18776 20410 18788
rect 20622 18776 20628 18788
rect 20680 18816 20686 18828
rect 21560 18816 21588 18924
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22186 18952 22192 18964
rect 22143 18924 22192 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 22281 18955 22339 18961
rect 22281 18921 22293 18955
rect 22327 18952 22339 18955
rect 22649 18955 22707 18961
rect 22649 18952 22661 18955
rect 22327 18924 22661 18952
rect 22327 18921 22339 18924
rect 22281 18915 22339 18921
rect 22649 18921 22661 18924
rect 22695 18921 22707 18955
rect 22649 18915 22707 18921
rect 25038 18912 25044 18964
rect 25096 18912 25102 18964
rect 25225 18955 25283 18961
rect 25225 18921 25237 18955
rect 25271 18952 25283 18955
rect 25406 18952 25412 18964
rect 25271 18924 25412 18952
rect 25271 18921 25283 18924
rect 25225 18915 25283 18921
rect 21726 18844 21732 18896
rect 21784 18884 21790 18896
rect 22741 18887 22799 18893
rect 22741 18884 22753 18887
rect 21784 18856 22753 18884
rect 21784 18844 21790 18856
rect 22741 18853 22753 18856
rect 22787 18853 22799 18887
rect 22741 18847 22799 18853
rect 20680 18788 21036 18816
rect 21560 18788 22140 18816
rect 20680 18776 20686 18788
rect 19720 18748 19748 18776
rect 19720 18723 19948 18748
rect 19720 18720 19993 18723
rect 19920 18717 19993 18720
rect 19702 18680 19708 18692
rect 19628 18652 19708 18680
rect 19024 18640 19030 18652
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 19920 18686 19947 18717
rect 19935 18683 19947 18686
rect 19981 18683 19993 18717
rect 20806 18708 20812 18760
rect 20864 18708 20870 18760
rect 21008 18757 21036 18788
rect 22112 18760 22140 18788
rect 22186 18776 22192 18828
rect 22244 18816 22250 18828
rect 22557 18819 22615 18825
rect 22557 18816 22569 18819
rect 22244 18788 22569 18816
rect 22244 18776 22250 18788
rect 22557 18785 22569 18788
rect 22603 18785 22615 18819
rect 22557 18779 22615 18785
rect 24946 18776 24952 18828
rect 25004 18816 25010 18828
rect 25240 18816 25268 18915
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 26513 18955 26571 18961
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 27614 18952 27620 18964
rect 26559 18924 27620 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 27614 18912 27620 18924
rect 27672 18912 27678 18964
rect 31202 18912 31208 18964
rect 31260 18952 31266 18964
rect 31941 18955 31999 18961
rect 31941 18952 31953 18955
rect 31260 18924 31953 18952
rect 31260 18912 31266 18924
rect 31941 18921 31953 18924
rect 31987 18921 31999 18955
rect 31941 18915 31999 18921
rect 32401 18955 32459 18961
rect 32401 18921 32413 18955
rect 32447 18952 32459 18955
rect 32493 18955 32551 18961
rect 32493 18952 32505 18955
rect 32447 18924 32505 18952
rect 32447 18921 32459 18924
rect 32401 18915 32459 18921
rect 32493 18921 32505 18924
rect 32539 18921 32551 18955
rect 32493 18915 32551 18921
rect 32858 18912 32864 18964
rect 32916 18912 32922 18964
rect 32950 18912 32956 18964
rect 33008 18952 33014 18964
rect 33321 18955 33379 18961
rect 33321 18952 33333 18955
rect 33008 18924 33333 18952
rect 33008 18912 33014 18924
rect 33321 18921 33333 18924
rect 33367 18921 33379 18955
rect 33321 18915 33379 18921
rect 34698 18912 34704 18964
rect 34756 18952 34762 18964
rect 35897 18955 35955 18961
rect 35897 18952 35909 18955
rect 34756 18924 35909 18952
rect 34756 18912 34762 18924
rect 35897 18921 35909 18924
rect 35943 18921 35955 18955
rect 35897 18915 35955 18921
rect 26881 18887 26939 18893
rect 26881 18853 26893 18887
rect 26927 18884 26939 18887
rect 28718 18884 28724 18896
rect 26927 18856 28724 18884
rect 26927 18853 26939 18856
rect 26881 18847 26939 18853
rect 28718 18844 28724 18856
rect 28776 18884 28782 18896
rect 29362 18884 29368 18896
rect 28776 18856 29368 18884
rect 28776 18844 28782 18856
rect 29362 18844 29368 18856
rect 29420 18844 29426 18896
rect 31570 18844 31576 18896
rect 31628 18884 31634 18896
rect 31628 18856 35756 18884
rect 31628 18844 31634 18856
rect 25004 18788 25268 18816
rect 25004 18776 25010 18788
rect 25866 18776 25872 18828
rect 25924 18816 25930 18828
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 25924 18788 26709 18816
rect 25924 18776 25930 18788
rect 26697 18785 26709 18788
rect 26743 18785 26755 18819
rect 26697 18779 26755 18785
rect 32125 18819 32183 18825
rect 32125 18785 32137 18819
rect 32171 18816 32183 18819
rect 32398 18816 32404 18828
rect 32171 18788 32404 18816
rect 32171 18785 32183 18788
rect 32125 18779 32183 18785
rect 32398 18776 32404 18788
rect 32456 18776 32462 18828
rect 32600 18825 32628 18856
rect 32585 18819 32643 18825
rect 32585 18785 32597 18819
rect 32631 18785 32643 18819
rect 32585 18779 32643 18785
rect 33502 18776 33508 18828
rect 33560 18776 33566 18828
rect 34146 18776 34152 18828
rect 34204 18816 34210 18828
rect 34422 18816 34428 18828
rect 34204 18788 34428 18816
rect 34204 18776 34210 18788
rect 34422 18776 34428 18788
rect 34480 18816 34486 18828
rect 34480 18788 35112 18816
rect 34480 18776 34486 18788
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18717 21051 18751
rect 20993 18711 21051 18717
rect 21082 18708 21088 18760
rect 21140 18708 21146 18760
rect 21177 18751 21235 18757
rect 21177 18717 21189 18751
rect 21223 18717 21235 18751
rect 21177 18711 21235 18717
rect 19935 18677 19993 18683
rect 20165 18683 20223 18689
rect 20165 18649 20177 18683
rect 20211 18680 20223 18683
rect 20714 18680 20720 18692
rect 20211 18652 20720 18680
rect 20211 18649 20223 18652
rect 20165 18643 20223 18649
rect 20714 18640 20720 18652
rect 20772 18640 20778 18692
rect 19426 18612 19432 18624
rect 17144 18584 19432 18612
rect 16669 18575 16727 18581
rect 19426 18572 19432 18584
rect 19484 18572 19490 18624
rect 19518 18572 19524 18624
rect 19576 18612 19582 18624
rect 19797 18615 19855 18621
rect 19797 18612 19809 18615
rect 19576 18584 19809 18612
rect 19576 18572 19582 18584
rect 19797 18581 19809 18584
rect 19843 18581 19855 18615
rect 19797 18575 19855 18581
rect 20438 18572 20444 18624
rect 20496 18612 20502 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 20496 18584 20637 18612
rect 20496 18572 20502 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 20898 18572 20904 18624
rect 20956 18612 20962 18624
rect 21192 18612 21220 18711
rect 21266 18708 21272 18760
rect 21324 18708 21330 18760
rect 21450 18708 21456 18760
rect 21508 18708 21514 18760
rect 21637 18751 21695 18757
rect 21637 18717 21649 18751
rect 21683 18748 21695 18751
rect 21726 18748 21732 18760
rect 21683 18720 21732 18748
rect 21683 18717 21695 18720
rect 21637 18711 21695 18717
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 22833 18751 22891 18757
rect 22833 18717 22845 18751
rect 22879 18748 22891 18751
rect 24394 18748 24400 18760
rect 22879 18720 24400 18748
rect 22879 18717 22891 18720
rect 22833 18711 22891 18717
rect 24394 18708 24400 18720
rect 24452 18708 24458 18760
rect 24670 18708 24676 18760
rect 24728 18748 24734 18760
rect 26145 18751 26203 18757
rect 24728 18720 25452 18748
rect 24728 18708 24734 18720
rect 21542 18640 21548 18692
rect 21600 18640 21606 18692
rect 22249 18683 22307 18689
rect 22249 18680 22261 18683
rect 21744 18652 22261 18680
rect 20956 18584 21220 18612
rect 21361 18615 21419 18621
rect 20956 18572 20962 18584
rect 21361 18581 21373 18615
rect 21407 18612 21419 18615
rect 21744 18612 21772 18652
rect 22249 18649 22261 18652
rect 22295 18649 22307 18683
rect 22249 18643 22307 18649
rect 22462 18640 22468 18692
rect 22520 18640 22526 18692
rect 22646 18640 22652 18692
rect 22704 18680 22710 18692
rect 22922 18680 22928 18692
rect 22704 18652 22928 18680
rect 22704 18640 22710 18652
rect 22922 18640 22928 18652
rect 22980 18640 22986 18692
rect 25222 18689 25228 18692
rect 25209 18683 25228 18689
rect 25209 18649 25221 18683
rect 25209 18643 25228 18649
rect 25222 18640 25228 18643
rect 25280 18640 25286 18692
rect 25424 18689 25452 18720
rect 26145 18717 26157 18751
rect 26191 18748 26203 18751
rect 26234 18748 26240 18760
rect 26191 18720 26240 18748
rect 26191 18717 26203 18720
rect 26145 18711 26203 18717
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26326 18708 26332 18760
rect 26384 18708 26390 18760
rect 26605 18751 26663 18757
rect 26605 18717 26617 18751
rect 26651 18717 26663 18751
rect 26605 18711 26663 18717
rect 25409 18683 25467 18689
rect 25409 18649 25421 18683
rect 25455 18680 25467 18683
rect 25682 18680 25688 18692
rect 25455 18652 25688 18680
rect 25455 18649 25467 18652
rect 25409 18643 25467 18649
rect 25682 18640 25688 18652
rect 25740 18640 25746 18692
rect 26418 18680 26424 18692
rect 26252 18652 26424 18680
rect 21407 18584 21772 18612
rect 21407 18581 21419 18584
rect 21361 18575 21419 18581
rect 23750 18572 23756 18624
rect 23808 18612 23814 18624
rect 24486 18612 24492 18624
rect 23808 18584 24492 18612
rect 23808 18572 23814 18584
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 25240 18612 25268 18640
rect 25498 18612 25504 18624
rect 25240 18584 25504 18612
rect 25498 18572 25504 18584
rect 25556 18612 25562 18624
rect 26252 18621 26280 18652
rect 26418 18640 26424 18652
rect 26476 18640 26482 18692
rect 25869 18615 25927 18621
rect 25869 18612 25881 18615
rect 25556 18584 25881 18612
rect 25556 18572 25562 18584
rect 25869 18581 25881 18584
rect 25915 18581 25927 18615
rect 25869 18575 25927 18581
rect 26237 18615 26295 18621
rect 26237 18581 26249 18615
rect 26283 18581 26295 18615
rect 26237 18575 26295 18581
rect 26326 18572 26332 18624
rect 26384 18612 26390 18624
rect 26620 18612 26648 18711
rect 26970 18708 26976 18760
rect 27028 18748 27034 18760
rect 29178 18748 29184 18760
rect 27028 18720 29184 18748
rect 27028 18708 27034 18720
rect 29178 18708 29184 18720
rect 29236 18708 29242 18760
rect 32214 18708 32220 18760
rect 32272 18708 32278 18760
rect 32490 18708 32496 18760
rect 32548 18708 32554 18760
rect 32674 18708 32680 18760
rect 32732 18748 32738 18760
rect 33229 18751 33287 18757
rect 33229 18748 33241 18751
rect 32732 18720 33241 18748
rect 32732 18708 32738 18720
rect 33229 18717 33241 18720
rect 33275 18717 33287 18751
rect 33229 18711 33287 18717
rect 33689 18751 33747 18757
rect 33689 18717 33701 18751
rect 33735 18748 33747 18751
rect 34698 18748 34704 18760
rect 33735 18720 34704 18748
rect 33735 18717 33747 18720
rect 33689 18711 33747 18717
rect 34698 18708 34704 18720
rect 34756 18708 34762 18760
rect 34793 18751 34851 18757
rect 34793 18717 34805 18751
rect 34839 18717 34851 18751
rect 34793 18711 34851 18717
rect 27157 18683 27215 18689
rect 27157 18649 27169 18683
rect 27203 18680 27215 18683
rect 27246 18680 27252 18692
rect 27203 18652 27252 18680
rect 27203 18649 27215 18652
rect 27157 18643 27215 18649
rect 27246 18640 27252 18652
rect 27304 18640 27310 18692
rect 29546 18640 29552 18692
rect 29604 18680 29610 18692
rect 31018 18680 31024 18692
rect 29604 18652 31024 18680
rect 29604 18640 29610 18652
rect 31018 18640 31024 18652
rect 31076 18640 31082 18692
rect 31202 18640 31208 18692
rect 31260 18680 31266 18692
rect 31941 18683 31999 18689
rect 31941 18680 31953 18683
rect 31260 18652 31953 18680
rect 31260 18640 31266 18652
rect 31941 18649 31953 18652
rect 31987 18649 31999 18683
rect 34808 18680 34836 18711
rect 34882 18708 34888 18760
rect 34940 18748 34946 18760
rect 35084 18748 35112 18788
rect 35728 18757 35756 18856
rect 35258 18751 35316 18757
rect 35258 18748 35270 18751
rect 34940 18720 34985 18748
rect 35084 18720 35270 18748
rect 34940 18708 34946 18720
rect 35258 18717 35270 18720
rect 35304 18717 35316 18751
rect 35258 18711 35316 18717
rect 35713 18751 35771 18757
rect 35713 18717 35725 18751
rect 35759 18717 35771 18751
rect 35713 18711 35771 18717
rect 31941 18643 31999 18649
rect 33336 18652 34836 18680
rect 26384 18584 26648 18612
rect 26384 18572 26390 18584
rect 30098 18572 30104 18624
rect 30156 18612 30162 18624
rect 33336 18612 33364 18652
rect 35066 18640 35072 18692
rect 35124 18640 35130 18692
rect 35161 18683 35219 18689
rect 35161 18649 35173 18683
rect 35207 18649 35219 18683
rect 35161 18643 35219 18649
rect 35529 18683 35587 18689
rect 35529 18649 35541 18683
rect 35575 18649 35587 18683
rect 35529 18643 35587 18649
rect 30156 18584 33364 18612
rect 33873 18615 33931 18621
rect 30156 18572 30162 18584
rect 33873 18581 33885 18615
rect 33919 18612 33931 18615
rect 33962 18612 33968 18624
rect 33919 18584 33968 18612
rect 33919 18581 33931 18584
rect 33873 18575 33931 18581
rect 33962 18572 33968 18584
rect 34020 18572 34026 18624
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 35176 18612 35204 18643
rect 34572 18584 35204 18612
rect 35437 18615 35495 18621
rect 34572 18572 34578 18584
rect 35437 18581 35449 18615
rect 35483 18612 35495 18615
rect 35544 18612 35572 18643
rect 35483 18584 35572 18612
rect 35483 18581 35495 18584
rect 35437 18575 35495 18581
rect 1104 18522 36524 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 36524 18522
rect 1104 18448 36524 18470
rect 3145 18411 3203 18417
rect 3145 18377 3157 18411
rect 3191 18408 3203 18411
rect 3326 18408 3332 18420
rect 3191 18380 3332 18408
rect 3191 18377 3203 18380
rect 3145 18371 3203 18377
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 5169 18411 5227 18417
rect 3476 18380 5028 18408
rect 3476 18368 3482 18380
rect 3436 18340 3464 18368
rect 2898 18312 3464 18340
rect 3694 18300 3700 18352
rect 3752 18300 3758 18352
rect 5000 18340 5028 18380
rect 5169 18377 5181 18411
rect 5215 18408 5227 18411
rect 5258 18408 5264 18420
rect 5215 18380 5264 18408
rect 5215 18377 5227 18380
rect 5169 18371 5227 18377
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 5905 18411 5963 18417
rect 5905 18377 5917 18411
rect 5951 18408 5963 18411
rect 7098 18408 7104 18420
rect 5951 18380 7104 18408
rect 5951 18377 5963 18380
rect 5905 18371 5963 18377
rect 7098 18368 7104 18380
rect 7156 18368 7162 18420
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 9309 18411 9367 18417
rect 9309 18408 9321 18411
rect 8260 18380 9321 18408
rect 8260 18368 8266 18380
rect 9309 18377 9321 18380
rect 9355 18377 9367 18411
rect 9309 18371 9367 18377
rect 9677 18411 9735 18417
rect 9677 18377 9689 18411
rect 9723 18408 9735 18411
rect 10318 18408 10324 18420
rect 9723 18380 10324 18408
rect 9723 18377 9735 18380
rect 9677 18371 9735 18377
rect 10318 18368 10324 18380
rect 10376 18368 10382 18420
rect 10870 18368 10876 18420
rect 10928 18368 10934 18420
rect 10962 18368 10968 18420
rect 11020 18368 11026 18420
rect 11882 18368 11888 18420
rect 11940 18368 11946 18420
rect 12066 18368 12072 18420
rect 12124 18368 12130 18420
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 12529 18411 12587 18417
rect 12529 18408 12541 18411
rect 12400 18380 12541 18408
rect 12400 18368 12406 18380
rect 12529 18377 12541 18380
rect 12575 18377 12587 18411
rect 12529 18371 12587 18377
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 14737 18411 14795 18417
rect 14737 18408 14749 18411
rect 14424 18380 14749 18408
rect 14424 18368 14430 18380
rect 14737 18377 14749 18380
rect 14783 18377 14795 18411
rect 14737 18371 14795 18377
rect 15105 18411 15163 18417
rect 15105 18377 15117 18411
rect 15151 18408 15163 18411
rect 15930 18408 15936 18420
rect 15151 18380 15936 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16574 18368 16580 18420
rect 16632 18408 16638 18420
rect 17494 18408 17500 18420
rect 16632 18380 17500 18408
rect 16632 18368 16638 18380
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 18874 18368 18880 18420
rect 18932 18368 18938 18420
rect 19705 18411 19763 18417
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 19978 18408 19984 18420
rect 19751 18380 19984 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 19978 18368 19984 18380
rect 20036 18368 20042 18420
rect 21085 18411 21143 18417
rect 21085 18377 21097 18411
rect 21131 18408 21143 18411
rect 21450 18408 21456 18420
rect 21131 18380 21456 18408
rect 21131 18377 21143 18380
rect 21085 18371 21143 18377
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 21726 18368 21732 18420
rect 21784 18408 21790 18420
rect 22002 18408 22008 18420
rect 21784 18380 22008 18408
rect 21784 18368 21790 18380
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 22830 18408 22836 18420
rect 22112 18380 22836 18408
rect 5350 18340 5356 18352
rect 4922 18312 5356 18340
rect 5350 18300 5356 18312
rect 5408 18300 5414 18352
rect 9030 18340 9036 18352
rect 8510 18326 9036 18340
rect 8496 18312 9036 18326
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18272 5871 18275
rect 6638 18272 6644 18284
rect 5859 18244 6644 18272
rect 5859 18241 5871 18244
rect 5813 18235 5871 18241
rect 6638 18232 6644 18244
rect 6696 18232 6702 18284
rect 7006 18232 7012 18284
rect 7064 18232 7070 18284
rect 1670 18164 1676 18216
rect 1728 18164 1734 18216
rect 2682 18164 2688 18216
rect 2740 18204 2746 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 2740 18176 3433 18204
rect 2740 18164 2746 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 4430 18204 4436 18216
rect 4120 18176 4436 18204
rect 4120 18164 4126 18176
rect 4430 18164 4436 18176
rect 4488 18204 4494 18216
rect 6089 18207 6147 18213
rect 6089 18204 6101 18207
rect 4488 18176 6101 18204
rect 4488 18164 4494 18176
rect 6089 18173 6101 18176
rect 6135 18204 6147 18207
rect 6822 18204 6828 18216
rect 6135 18176 6828 18204
rect 6135 18173 6147 18176
rect 6089 18167 6147 18173
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 7282 18164 7288 18216
rect 7340 18164 7346 18216
rect 7374 18164 7380 18216
rect 7432 18204 7438 18216
rect 8496 18204 8524 18312
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 9490 18300 9496 18352
rect 9548 18340 9554 18352
rect 9769 18343 9827 18349
rect 9769 18340 9781 18343
rect 9548 18312 9781 18340
rect 9548 18300 9554 18312
rect 9769 18309 9781 18312
rect 9815 18309 9827 18343
rect 9769 18303 9827 18309
rect 10226 18300 10232 18352
rect 10284 18340 10290 18352
rect 10284 18312 11652 18340
rect 10284 18300 10290 18312
rect 10410 18232 10416 18284
rect 10468 18272 10474 18284
rect 11422 18272 11428 18284
rect 10468 18244 11428 18272
rect 10468 18232 10474 18244
rect 11422 18232 11428 18244
rect 11480 18272 11486 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11480 18244 11529 18272
rect 11480 18232 11486 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11624 18272 11652 18312
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 13357 18343 13415 18349
rect 13357 18340 13369 18343
rect 11756 18312 13369 18340
rect 11756 18300 11762 18312
rect 13357 18309 13369 18312
rect 13403 18309 13415 18343
rect 13357 18303 13415 18309
rect 13541 18343 13599 18349
rect 13541 18309 13553 18343
rect 13587 18340 13599 18343
rect 13814 18340 13820 18352
rect 13587 18312 13820 18340
rect 13587 18309 13599 18312
rect 13541 18303 13599 18309
rect 13814 18300 13820 18312
rect 13872 18340 13878 18352
rect 15010 18340 15016 18352
rect 13872 18312 15016 18340
rect 13872 18300 13878 18312
rect 15010 18300 15016 18312
rect 15068 18300 15074 18352
rect 18138 18300 18144 18352
rect 18196 18340 18202 18352
rect 18509 18343 18567 18349
rect 18509 18340 18521 18343
rect 18196 18312 18521 18340
rect 18196 18300 18202 18312
rect 18509 18309 18521 18312
rect 18555 18340 18567 18343
rect 18555 18312 18904 18340
rect 18555 18309 18567 18312
rect 18509 18303 18567 18309
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 11624 18244 12173 18272
rect 11517 18235 11575 18241
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 7432 18176 8524 18204
rect 7432 18164 7438 18176
rect 9950 18164 9956 18216
rect 10008 18204 10014 18216
rect 11149 18207 11207 18213
rect 11149 18204 11161 18207
rect 10008 18176 11161 18204
rect 10008 18164 10014 18176
rect 11149 18173 11161 18176
rect 11195 18204 11207 18207
rect 12176 18204 12204 18235
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 13725 18275 13783 18281
rect 13725 18241 13737 18275
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 12986 18204 12992 18216
rect 11195 18176 12020 18204
rect 12176 18176 12992 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 11606 18136 11612 18148
rect 10100 18108 11612 18136
rect 10100 18096 10106 18108
rect 11606 18096 11612 18108
rect 11664 18096 11670 18148
rect 11992 18136 12020 18176
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 13078 18164 13084 18216
rect 13136 18164 13142 18216
rect 13170 18164 13176 18216
rect 13228 18204 13234 18216
rect 13740 18204 13768 18235
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18414 18281 18420 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18012 18244 18245 18272
rect 18012 18232 18018 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18381 18275 18420 18281
rect 18381 18241 18393 18275
rect 18381 18235 18420 18241
rect 18414 18232 18420 18235
rect 18472 18232 18478 18284
rect 18782 18281 18788 18284
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18739 18275 18788 18281
rect 18739 18241 18751 18275
rect 18785 18241 18788 18275
rect 18739 18235 18788 18241
rect 13228 18176 13768 18204
rect 13228 18164 13234 18176
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 14884 18176 15209 18204
rect 14884 18164 14890 18176
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18204 15439 18207
rect 15654 18204 15660 18216
rect 15427 18176 15660 18204
rect 15427 18173 15439 18176
rect 15381 18167 15439 18173
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 12618 18136 12624 18148
rect 11992 18108 12624 18136
rect 12618 18096 12624 18108
rect 12676 18096 12682 18148
rect 13096 18136 13124 18164
rect 14274 18136 14280 18148
rect 13096 18108 14280 18136
rect 14274 18096 14280 18108
rect 14332 18096 14338 18148
rect 18230 18096 18236 18148
rect 18288 18136 18294 18148
rect 18506 18136 18512 18148
rect 18288 18108 18512 18136
rect 18288 18096 18294 18108
rect 18506 18096 18512 18108
rect 18564 18136 18570 18148
rect 18616 18136 18644 18235
rect 18782 18232 18788 18235
rect 18840 18232 18846 18284
rect 18876 18272 18904 18312
rect 19150 18300 19156 18352
rect 19208 18340 19214 18352
rect 19518 18340 19524 18352
rect 19208 18312 19524 18340
rect 19208 18300 19214 18312
rect 19518 18300 19524 18312
rect 19576 18300 19582 18352
rect 20162 18340 20168 18352
rect 19628 18312 20168 18340
rect 19628 18272 19656 18312
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 22112 18340 22140 18380
rect 22830 18368 22836 18380
rect 22888 18368 22894 18420
rect 22922 18368 22928 18420
rect 22980 18408 22986 18420
rect 23201 18411 23259 18417
rect 23201 18408 23213 18411
rect 22980 18380 23213 18408
rect 22980 18368 22986 18380
rect 23201 18377 23213 18380
rect 23247 18377 23259 18411
rect 23201 18371 23259 18377
rect 23369 18411 23427 18417
rect 23369 18377 23381 18411
rect 23415 18408 23427 18411
rect 23750 18408 23756 18420
rect 23415 18380 23756 18408
rect 23415 18377 23427 18380
rect 23369 18371 23427 18377
rect 23750 18368 23756 18380
rect 23808 18368 23814 18420
rect 24486 18368 24492 18420
rect 24544 18408 24550 18420
rect 24544 18380 26188 18408
rect 24544 18368 24550 18380
rect 20732 18312 22140 18340
rect 18876 18244 19656 18272
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 20073 18275 20131 18281
rect 20073 18272 20085 18275
rect 19760 18244 20085 18272
rect 19760 18232 19766 18244
rect 20073 18241 20085 18244
rect 20119 18241 20131 18275
rect 20073 18235 20131 18241
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20272 18204 20300 18235
rect 20438 18232 20444 18284
rect 20496 18232 20502 18284
rect 20732 18281 20760 18312
rect 22462 18300 22468 18352
rect 22520 18340 22526 18352
rect 22649 18343 22707 18349
rect 22649 18340 22661 18343
rect 22520 18312 22661 18340
rect 22520 18300 22526 18312
rect 22649 18309 22661 18312
rect 22695 18309 22707 18343
rect 22649 18303 22707 18309
rect 22738 18300 22744 18352
rect 22796 18340 22802 18352
rect 23569 18343 23627 18349
rect 22796 18312 23244 18340
rect 22796 18300 22802 18312
rect 20717 18275 20775 18281
rect 20717 18241 20729 18275
rect 20763 18241 20775 18275
rect 20717 18235 20775 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 21358 18272 21364 18284
rect 21315 18244 21364 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 21450 18232 21456 18284
rect 21508 18232 21514 18284
rect 22278 18272 22284 18284
rect 21560 18244 22284 18272
rect 19352 18176 20300 18204
rect 20993 18207 21051 18213
rect 18564 18108 18644 18136
rect 18564 18096 18570 18108
rect 18782 18096 18788 18148
rect 18840 18136 18846 18148
rect 19150 18136 19156 18148
rect 18840 18108 19156 18136
rect 18840 18096 18846 18108
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 5445 18071 5503 18077
rect 5445 18037 5457 18071
rect 5491 18068 5503 18071
rect 5810 18068 5816 18080
rect 5491 18040 5816 18068
rect 5491 18037 5503 18040
rect 5445 18031 5503 18037
rect 5810 18028 5816 18040
rect 5868 18028 5874 18080
rect 8754 18028 8760 18080
rect 8812 18028 8818 18080
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10505 18071 10563 18077
rect 10505 18068 10517 18071
rect 10192 18040 10517 18068
rect 10192 18028 10198 18040
rect 10505 18037 10517 18040
rect 10551 18037 10563 18071
rect 10505 18031 10563 18037
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 19352 18068 19380 18176
rect 20993 18173 21005 18207
rect 21039 18204 21051 18207
rect 21174 18204 21180 18216
rect 21039 18176 21180 18204
rect 21039 18173 21051 18176
rect 20993 18167 21051 18173
rect 21174 18164 21180 18176
rect 21232 18164 21238 18216
rect 19426 18096 19432 18148
rect 19484 18136 19490 18148
rect 21560 18136 21588 18244
rect 22278 18232 22284 18244
rect 22336 18232 22342 18284
rect 22554 18232 22560 18284
rect 22612 18272 22618 18284
rect 23017 18275 23075 18281
rect 23017 18272 23029 18275
rect 22612 18244 23029 18272
rect 22612 18232 22618 18244
rect 23017 18241 23029 18244
rect 23063 18241 23075 18275
rect 23017 18235 23075 18241
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18241 23167 18275
rect 23216 18272 23244 18312
rect 23569 18309 23581 18343
rect 23615 18340 23627 18343
rect 23615 18312 25284 18340
rect 23615 18309 23627 18312
rect 23569 18303 23627 18309
rect 23750 18272 23756 18284
rect 23216 18244 23756 18272
rect 23109 18235 23167 18241
rect 22738 18164 22744 18216
rect 22796 18164 22802 18216
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23124 18204 23152 18235
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 23934 18232 23940 18284
rect 23992 18232 23998 18284
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 23290 18204 23296 18216
rect 22980 18176 23296 18204
rect 22980 18164 22986 18176
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 23842 18164 23848 18216
rect 23900 18204 23906 18216
rect 24136 18204 24164 18235
rect 24946 18232 24952 18284
rect 25004 18232 25010 18284
rect 25130 18232 25136 18284
rect 25188 18232 25194 18284
rect 23900 18176 24164 18204
rect 24581 18207 24639 18213
rect 23900 18164 23906 18176
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 24762 18204 24768 18216
rect 24627 18176 24768 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 19484 18108 21588 18136
rect 19484 18096 19490 18108
rect 21818 18096 21824 18148
rect 21876 18136 21882 18148
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 21876 18108 24685 18136
rect 21876 18096 21882 18108
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 25256 18136 25284 18312
rect 25314 18300 25320 18352
rect 25372 18300 25378 18352
rect 25533 18343 25591 18349
rect 25533 18309 25545 18343
rect 25579 18340 25591 18343
rect 25682 18340 25688 18352
rect 25579 18312 25688 18340
rect 25579 18309 25591 18312
rect 25533 18303 25591 18309
rect 25682 18300 25688 18312
rect 25740 18300 25746 18352
rect 26160 18340 26188 18380
rect 26234 18368 26240 18420
rect 26292 18368 26298 18420
rect 26418 18368 26424 18420
rect 26476 18408 26482 18420
rect 29362 18408 29368 18420
rect 26476 18380 28304 18408
rect 26476 18368 26482 18380
rect 28276 18352 28304 18380
rect 28368 18380 29368 18408
rect 28169 18343 28227 18349
rect 28169 18340 28181 18343
rect 26160 18312 28181 18340
rect 28169 18309 28181 18312
rect 28215 18309 28227 18343
rect 28169 18303 28227 18309
rect 25332 18204 25360 18300
rect 25869 18275 25927 18281
rect 25869 18241 25881 18275
rect 25915 18272 25927 18275
rect 26050 18272 26056 18284
rect 25915 18244 26056 18272
rect 25915 18241 25927 18244
rect 25869 18235 25927 18241
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 27798 18232 27804 18284
rect 27856 18272 27862 18284
rect 27982 18272 27988 18284
rect 27856 18244 27988 18272
rect 27856 18232 27862 18244
rect 27982 18232 27988 18244
rect 28040 18281 28046 18284
rect 28040 18275 28089 18281
rect 28040 18241 28043 18275
rect 28077 18241 28089 18275
rect 28040 18235 28089 18241
rect 28040 18232 28046 18235
rect 25961 18207 26019 18213
rect 25961 18204 25973 18207
rect 25332 18176 25973 18204
rect 25961 18173 25973 18176
rect 26007 18173 26019 18207
rect 25961 18167 26019 18173
rect 27893 18207 27951 18213
rect 27893 18173 27905 18207
rect 27939 18173 27951 18207
rect 28184 18204 28212 18303
rect 28258 18300 28264 18352
rect 28316 18300 28322 18352
rect 28368 18281 28396 18380
rect 29362 18368 29368 18380
rect 29420 18408 29426 18420
rect 29914 18408 29920 18420
rect 29420 18380 29920 18408
rect 29420 18368 29426 18380
rect 29914 18368 29920 18380
rect 29972 18368 29978 18420
rect 31202 18368 31208 18420
rect 31260 18368 31266 18420
rect 28537 18343 28595 18349
rect 28537 18309 28549 18343
rect 28583 18340 28595 18343
rect 28583 18312 30328 18340
rect 28583 18309 28595 18312
rect 28537 18303 28595 18309
rect 30300 18284 30328 18312
rect 30742 18300 30748 18352
rect 30800 18300 30806 18352
rect 28353 18275 28411 18281
rect 28353 18241 28365 18275
rect 28399 18241 28411 18275
rect 28353 18235 28411 18241
rect 28905 18275 28963 18281
rect 28905 18241 28917 18275
rect 28951 18272 28963 18275
rect 30006 18272 30012 18284
rect 28951 18244 30012 18272
rect 28951 18241 28963 18244
rect 28905 18235 28963 18241
rect 30006 18232 30012 18244
rect 30064 18232 30070 18284
rect 30282 18232 30288 18284
rect 30340 18272 30346 18284
rect 31021 18275 31079 18281
rect 31021 18272 31033 18275
rect 30340 18244 31033 18272
rect 30340 18232 30346 18244
rect 31021 18241 31033 18244
rect 31067 18241 31079 18275
rect 31021 18235 31079 18241
rect 29178 18204 29184 18216
rect 28184 18176 29184 18204
rect 27893 18167 27951 18173
rect 25314 18136 25320 18148
rect 25256 18108 25320 18136
rect 24673 18099 24731 18105
rect 25314 18096 25320 18108
rect 25372 18096 25378 18148
rect 27798 18096 27804 18148
rect 27856 18136 27862 18148
rect 27908 18136 27936 18167
rect 29178 18164 29184 18176
rect 29236 18164 29242 18216
rect 30834 18164 30840 18216
rect 30892 18164 30898 18216
rect 29454 18136 29460 18148
rect 27856 18108 29460 18136
rect 27856 18096 27862 18108
rect 29454 18096 29460 18108
rect 29512 18096 29518 18148
rect 17644 18040 19380 18068
rect 17644 18028 17650 18040
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19576 18040 19993 18068
rect 19576 18028 19582 18040
rect 19981 18037 19993 18040
rect 20027 18068 20039 18071
rect 20070 18068 20076 18080
rect 20027 18040 20076 18068
rect 20027 18037 20039 18040
rect 19981 18031 20039 18037
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 20165 18071 20223 18077
rect 20165 18037 20177 18071
rect 20211 18068 20223 18071
rect 20533 18071 20591 18077
rect 20533 18068 20545 18071
rect 20211 18040 20545 18068
rect 20211 18037 20223 18040
rect 20165 18031 20223 18037
rect 20533 18037 20545 18040
rect 20579 18037 20591 18071
rect 20533 18031 20591 18037
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 21634 18068 21640 18080
rect 20947 18040 21640 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 22646 18028 22652 18080
rect 22704 18068 22710 18080
rect 22833 18071 22891 18077
rect 22833 18068 22845 18071
rect 22704 18040 22845 18068
rect 22704 18028 22710 18040
rect 22833 18037 22845 18040
rect 22879 18037 22891 18071
rect 22833 18031 22891 18037
rect 23198 18028 23204 18080
rect 23256 18068 23262 18080
rect 23385 18071 23443 18077
rect 23385 18068 23397 18071
rect 23256 18040 23397 18068
rect 23256 18028 23262 18040
rect 23385 18037 23397 18040
rect 23431 18037 23443 18071
rect 23385 18031 23443 18037
rect 23750 18028 23756 18080
rect 23808 18028 23814 18080
rect 24210 18028 24216 18080
rect 24268 18068 24274 18080
rect 24305 18071 24363 18077
rect 24305 18068 24317 18071
rect 24268 18040 24317 18068
rect 24268 18028 24274 18040
rect 24305 18037 24317 18040
rect 24351 18037 24363 18071
rect 24305 18031 24363 18037
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 25501 18071 25559 18077
rect 25501 18068 25513 18071
rect 25280 18040 25513 18068
rect 25280 18028 25286 18040
rect 25501 18037 25513 18040
rect 25547 18037 25559 18071
rect 25501 18031 25559 18037
rect 25682 18028 25688 18080
rect 25740 18028 25746 18080
rect 26053 18071 26111 18077
rect 26053 18037 26065 18071
rect 26099 18068 26111 18071
rect 26142 18068 26148 18080
rect 26099 18040 26148 18068
rect 26099 18037 26111 18040
rect 26053 18031 26111 18037
rect 26142 18028 26148 18040
rect 26200 18028 26206 18080
rect 28258 18028 28264 18080
rect 28316 18068 28322 18080
rect 28721 18071 28779 18077
rect 28721 18068 28733 18071
rect 28316 18040 28733 18068
rect 28316 18028 28322 18040
rect 28721 18037 28733 18040
rect 28767 18037 28779 18071
rect 28721 18031 28779 18037
rect 30466 18028 30472 18080
rect 30524 18068 30530 18080
rect 30745 18071 30803 18077
rect 30745 18068 30757 18071
rect 30524 18040 30757 18068
rect 30524 18028 30530 18040
rect 30745 18037 30757 18040
rect 30791 18068 30803 18071
rect 30926 18068 30932 18080
rect 30791 18040 30932 18068
rect 30791 18037 30803 18040
rect 30745 18031 30803 18037
rect 30926 18028 30932 18040
rect 30984 18028 30990 18080
rect 34238 18028 34244 18080
rect 34296 18068 34302 18080
rect 35066 18068 35072 18080
rect 34296 18040 35072 18068
rect 34296 18028 34302 18040
rect 35066 18028 35072 18040
rect 35124 18028 35130 18080
rect 1104 17978 36524 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 36524 17978
rect 1104 17904 36524 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 1728 17836 2145 17864
rect 1728 17824 1734 17836
rect 2133 17833 2145 17836
rect 2179 17833 2191 17867
rect 2133 17827 2191 17833
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 7098 17864 7104 17876
rect 4672 17836 7104 17864
rect 4672 17824 4678 17836
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 7282 17824 7288 17876
rect 7340 17864 7346 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7340 17836 7665 17864
rect 7340 17824 7346 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 8220 17836 12848 17864
rect 2958 17796 2964 17808
rect 2700 17768 2964 17796
rect 2314 17688 2320 17740
rect 2372 17728 2378 17740
rect 2498 17728 2504 17740
rect 2372 17700 2504 17728
rect 2372 17688 2378 17700
rect 2498 17688 2504 17700
rect 2556 17728 2562 17740
rect 2700 17737 2728 17768
rect 2958 17756 2964 17768
rect 3016 17756 3022 17808
rect 6822 17756 6828 17808
rect 6880 17796 6886 17808
rect 8220 17796 8248 17836
rect 6880 17768 8248 17796
rect 12820 17796 12848 17836
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 12952 17836 13093 17864
rect 12952 17824 12958 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 15286 17824 15292 17876
rect 15344 17824 15350 17876
rect 15930 17824 15936 17876
rect 15988 17824 15994 17876
rect 21082 17864 21088 17876
rect 17236 17836 21088 17864
rect 13722 17796 13728 17808
rect 12820 17768 13728 17796
rect 6880 17756 6886 17768
rect 2593 17731 2651 17737
rect 2593 17728 2605 17731
rect 2556 17700 2605 17728
rect 2556 17688 2562 17700
rect 2593 17697 2605 17700
rect 2639 17697 2651 17731
rect 2593 17691 2651 17697
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17697 2743 17731
rect 2685 17691 2743 17697
rect 3326 17688 3332 17740
rect 3384 17728 3390 17740
rect 3513 17731 3571 17737
rect 3513 17728 3525 17731
rect 3384 17700 3525 17728
rect 3384 17688 3390 17700
rect 3513 17697 3525 17700
rect 3559 17697 3571 17731
rect 3513 17691 3571 17697
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 5537 17731 5595 17737
rect 5537 17728 5549 17731
rect 4764 17700 5549 17728
rect 4764 17688 4770 17700
rect 5537 17697 5549 17700
rect 5583 17697 5595 17731
rect 5537 17691 5595 17697
rect 5810 17688 5816 17740
rect 5868 17688 5874 17740
rect 7282 17688 7288 17740
rect 7340 17728 7346 17740
rect 8110 17728 8116 17740
rect 7340 17700 8116 17728
rect 7340 17688 7346 17700
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 8220 17737 8248 17768
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 14918 17756 14924 17808
rect 14976 17796 14982 17808
rect 16666 17796 16672 17808
rect 14976 17768 16672 17796
rect 14976 17756 14982 17768
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 8205 17731 8263 17737
rect 8205 17697 8217 17731
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 8754 17688 8760 17740
rect 8812 17728 8818 17740
rect 9493 17731 9551 17737
rect 9493 17728 9505 17731
rect 8812 17700 9505 17728
rect 8812 17688 8818 17700
rect 9493 17697 9505 17700
rect 9539 17697 9551 17731
rect 12342 17728 12348 17740
rect 9493 17691 9551 17697
rect 9600 17700 12348 17728
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2746 17632 2973 17660
rect 2501 17595 2559 17601
rect 2501 17561 2513 17595
rect 2547 17592 2559 17595
rect 2746 17592 2774 17632
rect 2961 17629 2973 17632
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 5442 17660 5448 17672
rect 4479 17632 5448 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4724 17604 4752 17632
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 9600 17660 9628 17700
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 13538 17728 13544 17740
rect 12452 17700 13544 17728
rect 7484 17632 9628 17660
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 2547 17564 2774 17592
rect 2884 17564 3801 17592
rect 2547 17561 2559 17564
rect 2501 17555 2559 17561
rect 2682 17484 2688 17536
rect 2740 17524 2746 17536
rect 2884 17524 2912 17564
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 3789 17555 3847 17561
rect 4706 17552 4712 17604
rect 4764 17552 4770 17604
rect 7190 17592 7196 17604
rect 7038 17564 7196 17592
rect 7190 17552 7196 17564
rect 7248 17592 7254 17604
rect 7374 17592 7380 17604
rect 7248 17564 7380 17592
rect 7248 17552 7254 17564
rect 7374 17552 7380 17564
rect 7432 17552 7438 17604
rect 2740 17496 2912 17524
rect 2740 17484 2746 17496
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 7484 17524 7512 17632
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11020 17632 11100 17660
rect 11020 17620 11026 17632
rect 8021 17595 8079 17601
rect 8021 17561 8033 17595
rect 8067 17592 8079 17595
rect 8941 17595 8999 17601
rect 8941 17592 8953 17595
rect 8067 17564 8953 17592
rect 8067 17561 8079 17564
rect 8021 17555 8079 17561
rect 8941 17561 8953 17564
rect 8987 17561 8999 17595
rect 11072 17592 11100 17632
rect 11146 17620 11152 17672
rect 11204 17620 11210 17672
rect 12158 17620 12164 17672
rect 12216 17660 12222 17672
rect 12452 17669 12480 17700
rect 12253 17663 12311 17669
rect 12253 17660 12265 17663
rect 12216 17632 12265 17660
rect 12216 17620 12222 17632
rect 12253 17629 12265 17632
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 13004 17669 13032 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13814 17728 13820 17740
rect 13648 17700 13820 17728
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12676 17632 12817 17660
rect 12676 17620 12682 17632
rect 12805 17629 12817 17632
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17629 13047 17663
rect 12989 17623 13047 17629
rect 12176 17592 12204 17620
rect 11072 17564 12204 17592
rect 12820 17592 12848 17623
rect 13078 17620 13084 17672
rect 13136 17620 13142 17672
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17660 13323 17663
rect 13648 17660 13676 17700
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 16390 17728 16396 17740
rect 14016 17700 16396 17728
rect 13311 17632 13676 17660
rect 13725 17663 13783 17669
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 13725 17629 13737 17663
rect 13771 17660 13783 17663
rect 13906 17660 13912 17672
rect 13771 17632 13912 17660
rect 13771 17629 13783 17632
rect 13725 17623 13783 17629
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 14016 17592 14044 17700
rect 16390 17688 16396 17700
rect 16448 17688 16454 17740
rect 16482 17688 16488 17740
rect 16540 17688 16546 17740
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14918 17660 14924 17672
rect 14507 17632 14924 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 15102 17620 15108 17672
rect 15160 17620 15166 17672
rect 15194 17620 15200 17672
rect 15252 17620 15258 17672
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17660 16083 17663
rect 16206 17660 16212 17672
rect 16071 17632 16212 17660
rect 16071 17629 16083 17632
rect 16025 17623 16083 17629
rect 12820 17564 14044 17592
rect 8941 17555 8999 17561
rect 13280 17536 13308 17564
rect 14642 17552 14648 17604
rect 14700 17552 14706 17604
rect 14829 17595 14887 17601
rect 14829 17561 14841 17595
rect 14875 17592 14887 17595
rect 15212 17592 15240 17620
rect 14875 17564 15240 17592
rect 15381 17595 15439 17601
rect 14875 17561 14887 17564
rect 14829 17555 14887 17561
rect 15381 17561 15393 17595
rect 15427 17561 15439 17595
rect 15948 17592 15976 17623
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17660 16359 17663
rect 16500 17660 16528 17688
rect 17236 17669 17264 17836
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 22370 17824 22376 17876
rect 22428 17824 22434 17876
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 22520 17836 22569 17864
rect 22520 17824 22526 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 22664 17836 23796 17864
rect 18230 17796 18236 17808
rect 17328 17768 18236 17796
rect 17328 17669 17356 17768
rect 18230 17756 18236 17768
rect 18288 17756 18294 17808
rect 18417 17799 18475 17805
rect 18417 17765 18429 17799
rect 18463 17765 18475 17799
rect 18417 17759 18475 17765
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 18138 17728 18144 17740
rect 17819 17700 18144 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 18432 17728 18460 17759
rect 18506 17756 18512 17808
rect 18564 17796 18570 17808
rect 20714 17796 20720 17808
rect 18564 17768 20720 17796
rect 18564 17756 18570 17768
rect 20714 17756 20720 17768
rect 20772 17756 20778 17808
rect 20901 17799 20959 17805
rect 20901 17765 20913 17799
rect 20947 17796 20959 17799
rect 21450 17796 21456 17808
rect 20947 17768 21456 17796
rect 20947 17765 20959 17768
rect 20901 17759 20959 17765
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 22278 17756 22284 17808
rect 22336 17796 22342 17808
rect 22664 17796 22692 17836
rect 22336 17768 22692 17796
rect 22336 17756 22342 17768
rect 23658 17756 23664 17808
rect 23716 17756 23722 17808
rect 23768 17796 23796 17836
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24213 17867 24271 17873
rect 24213 17864 24225 17867
rect 24084 17836 24225 17864
rect 24084 17824 24090 17836
rect 24213 17833 24225 17836
rect 24259 17833 24271 17867
rect 24213 17827 24271 17833
rect 25222 17824 25228 17876
rect 25280 17824 25286 17876
rect 25409 17799 25467 17805
rect 23768 17768 24072 17796
rect 18432 17700 19104 17728
rect 16347 17632 16528 17660
rect 17221 17663 17279 17669
rect 16347 17629 16359 17632
rect 16301 17623 16359 17629
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17589 17663 17647 17669
rect 17589 17629 17601 17663
rect 17635 17660 17647 17663
rect 17862 17660 17868 17672
rect 17635 17632 17868 17660
rect 17635 17629 17647 17632
rect 17589 17623 17647 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 18012 17632 18705 17660
rect 18012 17620 18018 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 18693 17623 18751 17629
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 18874 17620 18880 17672
rect 18932 17620 18938 17672
rect 19076 17669 19104 17700
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 20312 17700 23980 17728
rect 20312 17688 20318 17700
rect 19061 17663 19119 17669
rect 19061 17629 19073 17663
rect 19107 17629 19119 17663
rect 19061 17623 19119 17629
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17660 20039 17663
rect 20622 17660 20628 17672
rect 20027 17632 20628 17660
rect 20027 17629 20039 17632
rect 19981 17623 20039 17629
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 21358 17620 21364 17672
rect 21416 17620 21422 17672
rect 22646 17660 22652 17672
rect 21468 17632 22652 17660
rect 16114 17592 16120 17604
rect 15948 17564 16120 17592
rect 15381 17555 15439 17561
rect 3292 17496 7512 17524
rect 8113 17527 8171 17533
rect 3292 17484 3298 17496
rect 8113 17493 8125 17527
rect 8159 17524 8171 17527
rect 8662 17524 8668 17536
rect 8159 17496 8668 17524
rect 8159 17493 8171 17496
rect 8113 17487 8171 17493
rect 8662 17484 8668 17496
rect 8720 17524 8726 17536
rect 9582 17524 9588 17536
rect 8720 17496 9588 17524
rect 8720 17484 8726 17496
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 11054 17484 11060 17536
rect 11112 17484 11118 17536
rect 12345 17527 12403 17533
rect 12345 17493 12357 17527
rect 12391 17524 12403 17527
rect 12526 17524 12532 17536
rect 12391 17496 12532 17524
rect 12391 17493 12403 17496
rect 12345 17487 12403 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 12802 17484 12808 17536
rect 12860 17484 12866 17536
rect 13262 17484 13268 17536
rect 13320 17484 13326 17536
rect 13538 17484 13544 17536
rect 13596 17484 13602 17536
rect 14918 17484 14924 17536
rect 14976 17484 14982 17536
rect 15010 17484 15016 17536
rect 15068 17524 15074 17536
rect 15396 17524 15424 17555
rect 16114 17552 16120 17564
rect 16172 17552 16178 17604
rect 16485 17595 16543 17601
rect 16485 17561 16497 17595
rect 16531 17592 16543 17595
rect 17126 17592 17132 17604
rect 16531 17564 17132 17592
rect 16531 17561 16543 17564
rect 16485 17555 16543 17561
rect 17126 17552 17132 17564
rect 17184 17552 17190 17604
rect 17405 17595 17463 17601
rect 17405 17561 17417 17595
rect 17451 17561 17463 17595
rect 17405 17555 17463 17561
rect 15068 17496 15424 17524
rect 15068 17484 15074 17496
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15620 17496 15669 17524
rect 15620 17484 15626 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 17034 17484 17040 17536
rect 17092 17484 17098 17536
rect 17420 17524 17448 17555
rect 17494 17552 17500 17604
rect 17552 17592 17558 17604
rect 18049 17595 18107 17601
rect 18049 17592 18061 17595
rect 17552 17564 18061 17592
rect 17552 17552 17558 17564
rect 18049 17561 18061 17564
rect 18095 17561 18107 17595
rect 18049 17555 18107 17561
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 19334 17592 19340 17604
rect 18196 17564 19340 17592
rect 18196 17552 18202 17564
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 20530 17552 20536 17604
rect 20588 17592 20594 17604
rect 21085 17595 21143 17601
rect 21085 17592 21097 17595
rect 20588 17564 21097 17592
rect 20588 17552 20594 17564
rect 21085 17561 21097 17564
rect 21131 17561 21143 17595
rect 21085 17555 21143 17561
rect 21174 17552 21180 17604
rect 21232 17592 21238 17604
rect 21269 17595 21327 17601
rect 21269 17592 21281 17595
rect 21232 17564 21281 17592
rect 21232 17552 21238 17564
rect 21269 17561 21281 17564
rect 21315 17592 21327 17595
rect 21468 17592 21496 17632
rect 22646 17620 22652 17632
rect 22704 17620 22710 17672
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17660 23535 17663
rect 23566 17660 23572 17672
rect 23523 17632 23572 17660
rect 23523 17629 23535 17632
rect 23477 17623 23535 17629
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 21315 17564 21496 17592
rect 21545 17595 21603 17601
rect 21315 17561 21327 17564
rect 21269 17555 21327 17561
rect 21545 17561 21557 17595
rect 21591 17592 21603 17595
rect 21634 17592 21640 17604
rect 21591 17564 21640 17592
rect 21591 17561 21603 17564
rect 21545 17555 21603 17561
rect 21634 17552 21640 17564
rect 21692 17552 21698 17604
rect 21726 17552 21732 17604
rect 21784 17552 21790 17604
rect 22738 17552 22744 17604
rect 22796 17552 22802 17604
rect 23290 17552 23296 17604
rect 23348 17592 23354 17604
rect 23845 17595 23903 17601
rect 23845 17592 23857 17595
rect 23348 17564 23857 17592
rect 23348 17552 23354 17564
rect 23845 17561 23857 17564
rect 23891 17561 23903 17595
rect 23845 17555 23903 17561
rect 17586 17524 17592 17536
rect 17420 17496 17592 17524
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 17957 17527 18015 17533
rect 17957 17493 17969 17527
rect 18003 17524 18015 17527
rect 18414 17524 18420 17536
rect 18003 17496 18420 17524
rect 18003 17493 18015 17496
rect 17957 17487 18015 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18506 17484 18512 17536
rect 18564 17484 18570 17536
rect 19794 17484 19800 17536
rect 19852 17484 19858 17536
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 22278 17524 22284 17536
rect 20772 17496 22284 17524
rect 20772 17484 20778 17496
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 22554 17533 22560 17536
rect 22541 17527 22560 17533
rect 22541 17493 22553 17527
rect 22541 17487 22560 17493
rect 22554 17484 22560 17487
rect 22612 17484 22618 17536
rect 23952 17524 23980 17700
rect 24044 17669 24072 17768
rect 25409 17765 25421 17799
rect 25455 17765 25467 17799
rect 25409 17759 25467 17765
rect 25424 17728 25452 17759
rect 25501 17731 25559 17737
rect 25501 17728 25513 17731
rect 25424 17700 25513 17728
rect 25501 17697 25513 17700
rect 25547 17697 25559 17731
rect 25501 17691 25559 17697
rect 26234 17688 26240 17740
rect 26292 17688 26298 17740
rect 27062 17728 27068 17740
rect 26344 17700 27068 17728
rect 24029 17663 24087 17669
rect 24029 17629 24041 17663
rect 24075 17660 24087 17663
rect 24210 17660 24216 17672
rect 24075 17632 24216 17660
rect 24075 17629 24087 17632
rect 24029 17623 24087 17629
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 24946 17620 24952 17672
rect 25004 17660 25010 17672
rect 25004 17632 25544 17660
rect 25004 17620 25010 17632
rect 25038 17552 25044 17604
rect 25096 17552 25102 17604
rect 25516 17533 25544 17632
rect 25682 17620 25688 17672
rect 25740 17620 25746 17672
rect 25866 17620 25872 17672
rect 25924 17660 25930 17672
rect 26344 17669 26372 17700
rect 27062 17688 27068 17700
rect 27120 17688 27126 17740
rect 25961 17663 26019 17669
rect 25961 17660 25973 17663
rect 25924 17632 25973 17660
rect 25924 17620 25930 17632
rect 25961 17629 25973 17632
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 26329 17663 26387 17669
rect 26329 17629 26341 17663
rect 26375 17629 26387 17663
rect 26329 17623 26387 17629
rect 29638 17552 29644 17604
rect 29696 17592 29702 17604
rect 31018 17592 31024 17604
rect 29696 17564 31024 17592
rect 29696 17552 29702 17564
rect 31018 17552 31024 17564
rect 31076 17552 31082 17604
rect 32306 17552 32312 17604
rect 32364 17592 32370 17604
rect 33410 17592 33416 17604
rect 32364 17564 33416 17592
rect 32364 17552 32370 17564
rect 33410 17552 33416 17564
rect 33468 17552 33474 17604
rect 25241 17527 25299 17533
rect 25241 17524 25253 17527
rect 23952 17496 25253 17524
rect 25241 17493 25253 17496
rect 25287 17493 25299 17527
rect 25241 17487 25299 17493
rect 25501 17527 25559 17533
rect 25501 17493 25513 17527
rect 25547 17493 25559 17527
rect 25501 17487 25559 17493
rect 29178 17484 29184 17536
rect 29236 17524 29242 17536
rect 34054 17524 34060 17536
rect 29236 17496 34060 17524
rect 29236 17484 29242 17496
rect 34054 17484 34060 17496
rect 34112 17484 34118 17536
rect 36446 17484 36452 17536
rect 36504 17524 36510 17536
rect 36504 17496 36584 17524
rect 36504 17484 36510 17496
rect 1104 17434 36524 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 36524 17434
rect 1104 17360 36524 17382
rect 2682 17280 2688 17332
rect 2740 17280 2746 17332
rect 6638 17280 6644 17332
rect 6696 17280 6702 17332
rect 8757 17323 8815 17329
rect 8757 17289 8769 17323
rect 8803 17320 8815 17323
rect 8846 17320 8852 17332
rect 8803 17292 8852 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 8938 17280 8944 17332
rect 8996 17320 9002 17332
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 8996 17292 9597 17320
rect 8996 17280 9002 17292
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 9585 17283 9643 17289
rect 10137 17323 10195 17329
rect 10137 17289 10149 17323
rect 10183 17320 10195 17323
rect 10962 17320 10968 17332
rect 10183 17292 10968 17320
rect 10183 17289 10195 17292
rect 10137 17283 10195 17289
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 2777 17255 2835 17261
rect 2777 17252 2789 17255
rect 2648 17224 2789 17252
rect 2648 17212 2654 17224
rect 2777 17221 2789 17224
rect 2823 17221 2835 17255
rect 2777 17215 2835 17221
rect 2958 17212 2964 17264
rect 3016 17252 3022 17264
rect 3970 17252 3976 17264
rect 3016 17224 3976 17252
rect 3016 17212 3022 17224
rect 3970 17212 3976 17224
rect 4028 17212 4034 17264
rect 5350 17252 5356 17264
rect 5106 17224 5356 17252
rect 5350 17212 5356 17224
rect 5408 17212 5414 17264
rect 2976 17125 3004 17212
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5368 17156 6101 17184
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17085 3019 17119
rect 2961 17079 3019 17085
rect 3602 17076 3608 17128
rect 3660 17076 3666 17128
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17116 3939 17119
rect 4614 17116 4620 17128
rect 3927 17088 4620 17116
rect 3927 17085 3939 17088
rect 3881 17079 3939 17085
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 5368 17125 5396 17156
rect 6089 17153 6101 17156
rect 6135 17184 6147 17187
rect 6178 17184 6184 17196
rect 6135 17156 6184 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 7282 17144 7288 17196
rect 7340 17144 7346 17196
rect 8018 17144 8024 17196
rect 8076 17144 8082 17196
rect 8113 17187 8171 17193
rect 8113 17153 8125 17187
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 9048 17156 9904 17184
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 8128 17048 8156 17147
rect 9048 17125 9076 17156
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 5276 17020 8156 17048
rect 8297 17051 8355 17057
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 2317 16983 2375 16989
rect 2317 16980 2329 16983
rect 1728 16952 2329 16980
rect 1728 16940 1734 16952
rect 2317 16949 2329 16952
rect 2363 16949 2375 16983
rect 2317 16943 2375 16949
rect 2498 16940 2504 16992
rect 2556 16980 2562 16992
rect 5276 16980 5304 17020
rect 8297 17017 8309 17051
rect 8343 17048 8355 17051
rect 8662 17048 8668 17060
rect 8343 17020 8668 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 8864 17048 8892 17079
rect 9674 17076 9680 17128
rect 9732 17076 9738 17128
rect 9876 17125 9904 17156
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 10008 17156 10057 17184
rect 10008 17144 10014 17156
rect 10045 17153 10057 17156
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 10152 17116 10180 17283
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 12713 17323 12771 17329
rect 12713 17320 12725 17323
rect 11808 17292 12725 17320
rect 10226 17212 10232 17264
rect 10284 17252 10290 17264
rect 10870 17252 10876 17264
rect 10284 17224 10876 17252
rect 10284 17212 10290 17224
rect 10870 17212 10876 17224
rect 10928 17212 10934 17264
rect 10778 17144 10784 17196
rect 10836 17184 10842 17196
rect 11808 17193 11836 17292
rect 12713 17289 12725 17292
rect 12759 17320 12771 17323
rect 12894 17320 12900 17332
rect 12759 17292 12900 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 13630 17280 13636 17332
rect 13688 17320 13694 17332
rect 14077 17323 14135 17329
rect 13688 17292 14044 17320
rect 13688 17280 13694 17292
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 12618 17252 12624 17264
rect 12400 17224 12624 17252
rect 12400 17212 12406 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 13648 17252 13676 17280
rect 13556 17224 13676 17252
rect 14016 17252 14044 17292
rect 14077 17289 14089 17323
rect 14123 17320 14135 17323
rect 14182 17320 14188 17332
rect 14123 17292 14188 17320
rect 14123 17289 14135 17292
rect 14077 17283 14135 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14369 17323 14427 17329
rect 14369 17289 14381 17323
rect 14415 17320 14427 17323
rect 14458 17320 14464 17332
rect 14415 17292 14464 17320
rect 14415 17289 14427 17292
rect 14369 17283 14427 17289
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 15988 17292 19809 17320
rect 15988 17280 15994 17292
rect 16040 17261 16068 17292
rect 19797 17289 19809 17292
rect 19843 17289 19855 17323
rect 19797 17283 19855 17289
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17320 20867 17323
rect 21174 17320 21180 17332
rect 20855 17292 21180 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 21174 17280 21180 17292
rect 21232 17320 21238 17332
rect 21358 17320 21364 17332
rect 21232 17292 21364 17320
rect 21232 17280 21238 17292
rect 21358 17280 21364 17292
rect 21416 17280 21422 17332
rect 22554 17280 22560 17332
rect 22612 17280 22618 17332
rect 22738 17280 22744 17332
rect 22796 17280 22802 17332
rect 23290 17280 23296 17332
rect 23348 17280 23354 17332
rect 23566 17280 23572 17332
rect 23624 17320 23630 17332
rect 24762 17320 24768 17332
rect 23624 17292 24768 17320
rect 23624 17280 23630 17292
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 25222 17280 25228 17332
rect 25280 17320 25286 17332
rect 25685 17323 25743 17329
rect 25685 17320 25697 17323
rect 25280 17292 25697 17320
rect 25280 17280 25286 17292
rect 25685 17289 25697 17292
rect 25731 17289 25743 17323
rect 25685 17283 25743 17289
rect 25866 17280 25872 17332
rect 25924 17280 25930 17332
rect 27062 17280 27068 17332
rect 27120 17280 27126 17332
rect 29362 17280 29368 17332
rect 29420 17320 29426 17332
rect 29473 17323 29531 17329
rect 29473 17320 29485 17323
rect 29420 17292 29485 17320
rect 29420 17280 29426 17292
rect 29473 17289 29485 17292
rect 29519 17289 29531 17323
rect 29473 17283 29531 17289
rect 29641 17323 29699 17329
rect 29641 17289 29653 17323
rect 29687 17289 29699 17323
rect 29641 17283 29699 17289
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 14016 17224 14289 17252
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 10836 17156 11805 17184
rect 10836 17144 10842 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 11974 17144 11980 17196
rect 12032 17144 12038 17196
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17153 12863 17187
rect 12805 17147 12863 17153
rect 9907 17088 10180 17116
rect 11057 17119 11115 17125
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 11057 17085 11069 17119
rect 11103 17116 11115 17119
rect 11146 17116 11152 17128
rect 11103 17088 11152 17116
rect 11103 17085 11115 17088
rect 11057 17079 11115 17085
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 12710 17116 12716 17128
rect 12667 17088 12716 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 10413 17051 10471 17057
rect 10413 17048 10425 17051
rect 8864 17020 10425 17048
rect 10413 17017 10425 17020
rect 10459 17017 10471 17051
rect 10413 17011 10471 17017
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 12636 17048 12664 17079
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 12492 17020 12664 17048
rect 12820 17048 12848 17147
rect 13556 17116 13584 17224
rect 14277 17221 14289 17224
rect 14323 17221 14335 17255
rect 14277 17215 14335 17221
rect 16025 17255 16083 17261
rect 16025 17221 16037 17255
rect 16071 17221 16083 17255
rect 16025 17215 16083 17221
rect 16114 17212 16120 17264
rect 16172 17252 16178 17264
rect 20441 17255 20499 17261
rect 16172 17224 18368 17252
rect 16172 17212 16178 17224
rect 13630 17144 13636 17196
rect 13688 17144 13694 17196
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17184 14611 17187
rect 14734 17184 14740 17196
rect 14599 17156 14740 17184
rect 14599 17153 14611 17156
rect 14553 17147 14611 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17184 14887 17187
rect 15102 17184 15108 17196
rect 14875 17156 15108 17184
rect 14875 17153 14887 17156
rect 14829 17147 14887 17153
rect 15102 17144 15108 17156
rect 15160 17184 15166 17196
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 15160 17156 15209 17184
rect 15160 17144 15166 17156
rect 15197 17153 15209 17156
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 15378 17184 15384 17196
rect 15335 17156 15384 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15473 17187 15531 17193
rect 15473 17153 15485 17187
rect 15519 17153 15531 17187
rect 15473 17147 15531 17153
rect 13817 17119 13875 17125
rect 13817 17116 13829 17119
rect 13556 17088 13829 17116
rect 13817 17085 13829 17088
rect 13863 17085 13875 17119
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 13817 17079 13875 17085
rect 13924 17088 15025 17116
rect 12986 17048 12992 17060
rect 12820 17020 12992 17048
rect 12492 17008 12498 17020
rect 12986 17008 12992 17020
rect 13044 17048 13050 17060
rect 13924 17048 13952 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15488 17116 15516 17147
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16301 17187 16359 17193
rect 16301 17184 16313 17187
rect 15712 17156 16313 17184
rect 15712 17144 15718 17156
rect 16301 17153 16313 17156
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 16945 17187 17003 17193
rect 16945 17184 16957 17187
rect 16724 17156 16957 17184
rect 16724 17144 16730 17156
rect 16945 17153 16957 17156
rect 16991 17153 17003 17187
rect 16945 17147 17003 17153
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17184 17279 17187
rect 17310 17184 17316 17196
rect 17267 17156 17316 17184
rect 17267 17153 17279 17156
rect 17221 17147 17279 17153
rect 17310 17144 17316 17156
rect 17368 17144 17374 17196
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17184 17647 17187
rect 18230 17184 18236 17196
rect 17635 17156 18236 17184
rect 17635 17153 17647 17156
rect 17589 17147 17647 17153
rect 18230 17144 18236 17156
rect 18288 17144 18294 17196
rect 15838 17116 15844 17128
rect 15013 17079 15071 17085
rect 15120 17088 15844 17116
rect 15120 17060 15148 17088
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 16114 17076 16120 17128
rect 16172 17076 16178 17128
rect 16390 17076 16396 17128
rect 16448 17116 16454 17128
rect 16761 17119 16819 17125
rect 16761 17116 16773 17119
rect 16448 17088 16773 17116
rect 16448 17076 16454 17088
rect 16761 17085 16773 17088
rect 16807 17085 16819 17119
rect 17681 17119 17739 17125
rect 17681 17116 17693 17119
rect 16761 17079 16819 17085
rect 16868 17088 17693 17116
rect 14918 17048 14924 17060
rect 13044 17020 13952 17048
rect 14108 17020 14924 17048
rect 13044 17008 13050 17020
rect 2556 16952 5304 16980
rect 2556 16940 2562 16952
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 8389 16983 8447 16989
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 8570 16980 8576 16992
rect 8435 16952 8576 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9217 16983 9275 16989
rect 9217 16980 9229 16983
rect 9088 16952 9229 16980
rect 9088 16940 9094 16952
rect 9217 16949 9229 16952
rect 9263 16949 9275 16983
rect 9217 16943 9275 16949
rect 11514 16940 11520 16992
rect 11572 16940 11578 16992
rect 13170 16940 13176 16992
rect 13228 16940 13234 16992
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 13906 16940 13912 16992
rect 13964 16940 13970 16992
rect 14108 16989 14136 17020
rect 14918 17008 14924 17020
rect 14976 17008 14982 17060
rect 15102 17008 15108 17060
rect 15160 17008 15166 17060
rect 15378 17008 15384 17060
rect 15436 17008 15442 17060
rect 15470 17008 15476 17060
rect 15528 17048 15534 17060
rect 16868 17048 16896 17088
rect 17681 17085 17693 17088
rect 17727 17116 17739 17119
rect 17862 17116 17868 17128
rect 17727 17088 17868 17116
rect 17727 17085 17739 17088
rect 17681 17079 17739 17085
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 15528 17020 16896 17048
rect 15528 17008 15534 17020
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 17092 17020 17632 17048
rect 17092 17008 17098 17020
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16949 14151 16983
rect 14093 16943 14151 16949
rect 14734 16940 14740 16992
rect 14792 16940 14798 16992
rect 16022 16940 16028 16992
rect 16080 16940 16086 16992
rect 16485 16983 16543 16989
rect 16485 16949 16497 16983
rect 16531 16980 16543 16983
rect 17310 16980 17316 16992
rect 16531 16952 17316 16980
rect 16531 16949 16543 16952
rect 16485 16943 16543 16949
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17604 16989 17632 17020
rect 17954 17008 17960 17060
rect 18012 17008 18018 17060
rect 18340 17048 18368 17224
rect 20441 17221 20453 17255
rect 20487 17252 20499 17255
rect 20714 17252 20720 17264
rect 20487 17224 20720 17252
rect 20487 17221 20499 17224
rect 20441 17215 20499 17221
rect 20714 17212 20720 17224
rect 20772 17212 20778 17264
rect 23477 17255 23535 17261
rect 23477 17252 23489 17255
rect 22756 17224 23489 17252
rect 22756 17196 22784 17224
rect 23477 17221 23489 17224
rect 23523 17252 23535 17255
rect 23523 17224 24532 17252
rect 23523 17221 23535 17224
rect 23477 17215 23535 17221
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17184 19303 17187
rect 19334 17184 19340 17196
rect 19291 17156 19340 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 19334 17144 19340 17156
rect 19392 17144 19398 17196
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 19610 17184 19616 17196
rect 19475 17156 19616 17184
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 19610 17144 19616 17156
rect 19668 17184 19674 17196
rect 19794 17184 19800 17196
rect 19668 17156 19800 17184
rect 19668 17144 19674 17156
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20027 17156 20392 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 20070 17116 20076 17128
rect 19208 17088 20076 17116
rect 19208 17076 19214 17088
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20162 17076 20168 17128
rect 20220 17076 20226 17128
rect 20364 17116 20392 17156
rect 20622 17144 20628 17196
rect 20680 17144 20686 17196
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 21082 17193 21088 17196
rect 21049 17187 21088 17193
rect 21049 17153 21061 17187
rect 21049 17147 21088 17153
rect 21082 17144 21088 17147
rect 21140 17144 21146 17196
rect 21174 17144 21180 17196
rect 21232 17144 21238 17196
rect 21266 17144 21272 17196
rect 21324 17144 21330 17196
rect 21407 17187 21465 17193
rect 21407 17153 21419 17187
rect 21453 17184 21465 17187
rect 21542 17184 21548 17196
rect 21453 17156 21548 17184
rect 21453 17153 21465 17156
rect 21407 17147 21465 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 22278 17144 22284 17196
rect 22336 17144 22342 17196
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 22388 17156 22661 17184
rect 21726 17116 21732 17128
rect 20364 17088 21732 17116
rect 21726 17076 21732 17088
rect 21784 17076 21790 17128
rect 19702 17048 19708 17060
rect 18340 17020 19708 17048
rect 19702 17008 19708 17020
rect 19760 17008 19766 17060
rect 20180 17048 20208 17076
rect 20438 17048 20444 17060
rect 20180 17020 20444 17048
rect 20438 17008 20444 17020
rect 20496 17048 20502 17060
rect 21082 17048 21088 17060
rect 20496 17020 21088 17048
rect 20496 17008 20502 17020
rect 21082 17008 21088 17020
rect 21140 17048 21146 17060
rect 22186 17048 22192 17060
rect 21140 17020 22192 17048
rect 21140 17008 21146 17020
rect 22186 17008 22192 17020
rect 22244 17048 22250 17060
rect 22388 17048 22416 17156
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 22738 17144 22744 17196
rect 22796 17144 22802 17196
rect 22833 17187 22891 17193
rect 22833 17153 22845 17187
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 22554 17076 22560 17128
rect 22612 17076 22618 17128
rect 22848 17116 22876 17147
rect 23658 17144 23664 17196
rect 23716 17144 23722 17196
rect 24228 17193 24256 17224
rect 23937 17187 23995 17193
rect 23937 17153 23949 17187
rect 23983 17153 23995 17187
rect 23937 17147 23995 17153
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 22664 17088 22876 17116
rect 23952 17116 23980 17147
rect 24394 17144 24400 17196
rect 24452 17144 24458 17196
rect 24504 17184 24532 17224
rect 25314 17212 25320 17264
rect 25372 17252 25378 17264
rect 27706 17252 27712 17264
rect 25372 17224 27712 17252
rect 25372 17212 25378 17224
rect 27706 17212 27712 17224
rect 27764 17252 27770 17264
rect 29273 17255 29331 17261
rect 29273 17252 29285 17255
rect 27764 17224 29285 17252
rect 27764 17212 27770 17224
rect 29273 17221 29285 17224
rect 29319 17221 29331 17255
rect 29273 17215 29331 17221
rect 25682 17184 25688 17196
rect 24504 17156 25688 17184
rect 25682 17144 25688 17156
rect 25740 17144 25746 17196
rect 26142 17144 26148 17196
rect 26200 17184 26206 17196
rect 26970 17184 26976 17196
rect 26200 17156 26976 17184
rect 26200 17144 26206 17156
rect 26970 17144 26976 17156
rect 27028 17144 27034 17196
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 27522 17184 27528 17196
rect 27203 17156 27528 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 29288 17128 29316 17215
rect 29380 17128 29408 17280
rect 29656 17252 29684 17283
rect 30282 17280 30288 17332
rect 30340 17320 30346 17332
rect 30340 17292 32996 17320
rect 30340 17280 30346 17292
rect 29656 17224 32444 17252
rect 31202 17144 31208 17196
rect 31260 17184 31266 17196
rect 32030 17184 32036 17196
rect 31260 17156 32036 17184
rect 31260 17144 31266 17156
rect 32030 17144 32036 17156
rect 32088 17184 32094 17196
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 32088 17156 32137 17184
rect 32088 17144 32094 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32217 17187 32275 17193
rect 32217 17153 32229 17187
rect 32263 17184 32275 17187
rect 32306 17184 32312 17196
rect 32263 17156 32312 17184
rect 32263 17153 32275 17156
rect 32217 17147 32275 17153
rect 32306 17144 32312 17156
rect 32364 17144 32370 17196
rect 32416 17193 32444 17224
rect 32968 17193 32996 17292
rect 33226 17280 33232 17332
rect 33284 17320 33290 17332
rect 33502 17320 33508 17332
rect 33284 17292 33508 17320
rect 33284 17280 33290 17292
rect 33502 17280 33508 17292
rect 33560 17320 33566 17332
rect 33560 17292 34376 17320
rect 33560 17280 33566 17292
rect 34054 17212 34060 17264
rect 34112 17252 34118 17264
rect 34348 17261 34376 17292
rect 34241 17255 34299 17261
rect 34241 17252 34253 17255
rect 34112 17224 34253 17252
rect 34112 17212 34118 17224
rect 34241 17221 34253 17224
rect 34287 17221 34299 17255
rect 34241 17215 34299 17221
rect 34333 17255 34391 17261
rect 34333 17221 34345 17255
rect 34379 17221 34391 17255
rect 34333 17215 34391 17221
rect 34471 17255 34529 17261
rect 34471 17221 34483 17255
rect 34517 17252 34529 17255
rect 34790 17252 34796 17264
rect 34517 17224 34796 17252
rect 34517 17221 34529 17224
rect 34471 17215 34529 17221
rect 34790 17212 34796 17224
rect 34848 17212 34854 17264
rect 32401 17187 32459 17193
rect 32401 17153 32413 17187
rect 32447 17153 32459 17187
rect 32861 17187 32919 17193
rect 32861 17184 32873 17187
rect 32401 17147 32459 17153
rect 32600 17156 32873 17184
rect 26786 17116 26792 17128
rect 23952 17088 26792 17116
rect 22244 17020 22416 17048
rect 22244 17008 22250 17020
rect 22664 16992 22692 17088
rect 26786 17076 26792 17088
rect 26844 17076 26850 17128
rect 29270 17076 29276 17128
rect 29328 17076 29334 17128
rect 29362 17076 29368 17128
rect 29420 17076 29426 17128
rect 23290 17008 23296 17060
rect 23348 17048 23354 17060
rect 23348 17020 23888 17048
rect 23348 17008 23354 17020
rect 17589 16983 17647 16989
rect 17589 16949 17601 16983
rect 17635 16949 17647 16983
rect 17589 16943 17647 16949
rect 19150 16940 19156 16992
rect 19208 16940 19214 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19392 16952 19625 16980
rect 19392 16940 19398 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 20404 16952 21557 16980
rect 20404 16940 20410 16952
rect 21545 16949 21557 16952
rect 21591 16949 21603 16983
rect 21545 16943 21603 16949
rect 22373 16983 22431 16989
rect 22373 16949 22385 16983
rect 22419 16980 22431 16983
rect 22646 16980 22652 16992
rect 22419 16952 22652 16980
rect 22419 16949 22431 16952
rect 22373 16943 22431 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 23474 16940 23480 16992
rect 23532 16980 23538 16992
rect 23753 16983 23811 16989
rect 23753 16980 23765 16983
rect 23532 16952 23765 16980
rect 23532 16940 23538 16952
rect 23753 16949 23765 16952
rect 23799 16949 23811 16983
rect 23860 16980 23888 17020
rect 24026 17008 24032 17060
rect 24084 17008 24090 17060
rect 24118 17008 24124 17060
rect 24176 17008 24182 17060
rect 24581 17051 24639 17057
rect 24581 17017 24593 17051
rect 24627 17048 24639 17051
rect 24670 17048 24676 17060
rect 24627 17020 24676 17048
rect 24627 17017 24639 17020
rect 24581 17011 24639 17017
rect 24596 16980 24624 17011
rect 24670 17008 24676 17020
rect 24728 17008 24734 17060
rect 25317 17051 25375 17057
rect 25317 17017 25329 17051
rect 25363 17048 25375 17051
rect 25590 17048 25596 17060
rect 25363 17020 25596 17048
rect 25363 17017 25375 17020
rect 25317 17011 25375 17017
rect 25590 17008 25596 17020
rect 25648 17008 25654 17060
rect 32030 17008 32036 17060
rect 32088 17048 32094 17060
rect 32324 17048 32352 17144
rect 32088 17020 32352 17048
rect 32088 17008 32094 17020
rect 32600 16992 32628 17156
rect 32861 17153 32873 17156
rect 32907 17153 32919 17187
rect 32861 17147 32919 17153
rect 32953 17187 33011 17193
rect 32953 17153 32965 17187
rect 32999 17153 33011 17187
rect 32953 17147 33011 17153
rect 33137 17187 33195 17193
rect 33137 17153 33149 17187
rect 33183 17184 33195 17187
rect 33965 17187 34023 17193
rect 33965 17184 33977 17187
rect 33183 17156 33977 17184
rect 33183 17153 33195 17156
rect 33137 17147 33195 17153
rect 33965 17153 33977 17156
rect 34011 17153 34023 17187
rect 33965 17147 34023 17153
rect 34146 17144 34152 17196
rect 34204 17144 34210 17196
rect 36446 17144 36452 17196
rect 36504 17184 36510 17196
rect 36556 17184 36584 17496
rect 36504 17156 36584 17184
rect 36504 17144 36510 17156
rect 33410 17076 33416 17128
rect 33468 17116 33474 17128
rect 34609 17119 34667 17125
rect 34609 17116 34621 17119
rect 33468 17088 34621 17116
rect 33468 17076 33474 17088
rect 34609 17085 34621 17088
rect 34655 17085 34667 17119
rect 34609 17079 34667 17085
rect 23860 16952 24624 16980
rect 23753 16943 23811 16949
rect 25038 16940 25044 16992
rect 25096 16980 25102 16992
rect 25685 16983 25743 16989
rect 25685 16980 25697 16983
rect 25096 16952 25697 16980
rect 25096 16940 25102 16952
rect 25685 16949 25697 16952
rect 25731 16949 25743 16983
rect 25685 16943 25743 16949
rect 27706 16940 27712 16992
rect 27764 16980 27770 16992
rect 28994 16980 29000 16992
rect 27764 16952 29000 16980
rect 27764 16940 27770 16952
rect 28994 16940 29000 16952
rect 29052 16940 29058 16992
rect 29178 16940 29184 16992
rect 29236 16980 29242 16992
rect 29457 16983 29515 16989
rect 29457 16980 29469 16983
rect 29236 16952 29469 16980
rect 29236 16940 29242 16952
rect 29457 16949 29469 16952
rect 29503 16949 29515 16983
rect 29457 16943 29515 16949
rect 32582 16940 32588 16992
rect 32640 16940 32646 16992
rect 32674 16940 32680 16992
rect 32732 16940 32738 16992
rect 32766 16940 32772 16992
rect 32824 16980 32830 16992
rect 32861 16983 32919 16989
rect 32861 16980 32873 16983
rect 32824 16952 32873 16980
rect 32824 16940 32830 16952
rect 32861 16949 32873 16952
rect 32907 16949 32919 16983
rect 32861 16943 32919 16949
rect 1104 16890 36524 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 36524 16890
rect 1104 16816 36524 16838
rect 2120 16779 2178 16785
rect 2120 16745 2132 16779
rect 2166 16776 2178 16779
rect 2682 16776 2688 16788
rect 2166 16748 2688 16776
rect 2166 16745 2178 16748
rect 2120 16739 2178 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4614 16776 4620 16788
rect 4387 16748 4620 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 7098 16736 7104 16788
rect 7156 16776 7162 16788
rect 7929 16779 7987 16785
rect 7929 16776 7941 16779
rect 7156 16748 7941 16776
rect 7156 16736 7162 16748
rect 7929 16745 7941 16748
rect 7975 16776 7987 16779
rect 9398 16776 9404 16788
rect 7975 16748 9404 16776
rect 7975 16745 7987 16748
rect 7929 16739 7987 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 10413 16779 10471 16785
rect 10413 16776 10425 16779
rect 9732 16748 10425 16776
rect 9732 16736 9738 16748
rect 10413 16745 10425 16748
rect 10459 16745 10471 16779
rect 10413 16739 10471 16745
rect 10502 16736 10508 16788
rect 10560 16776 10566 16788
rect 10560 16748 12434 16776
rect 10560 16736 10566 16748
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 4120 16680 4936 16708
rect 4120 16668 4126 16680
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 2590 16640 2596 16652
rect 1903 16612 2596 16640
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 2682 16600 2688 16652
rect 2740 16640 2746 16652
rect 3418 16640 3424 16652
rect 2740 16612 3424 16640
rect 2740 16600 2746 16612
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 4908 16649 4936 16680
rect 8018 16668 8024 16720
rect 8076 16708 8082 16720
rect 8076 16680 9674 16708
rect 8076 16668 8082 16680
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16609 4951 16643
rect 4893 16603 4951 16609
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 6270 16640 6276 16652
rect 5951 16612 6276 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 8496 16612 9076 16640
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5442 16572 5448 16584
rect 4755 16544 5448 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 8496 16581 8524 16612
rect 8480 16575 8538 16581
rect 8036 16544 8432 16572
rect 5350 16504 5356 16516
rect 3358 16476 5356 16504
rect 3050 16396 3056 16448
rect 3108 16436 3114 16448
rect 3436 16436 3464 16476
rect 5350 16464 5356 16476
rect 5408 16504 5414 16516
rect 7913 16507 7971 16513
rect 5408 16476 6394 16504
rect 5408 16464 5414 16476
rect 7913 16473 7925 16507
rect 7959 16504 7971 16507
rect 8036 16504 8064 16544
rect 7959 16476 8064 16504
rect 8113 16507 8171 16513
rect 7959 16473 7971 16476
rect 7913 16467 7971 16473
rect 8113 16473 8125 16507
rect 8159 16473 8171 16507
rect 8404 16504 8432 16544
rect 8480 16541 8492 16575
rect 8526 16541 8538 16575
rect 8480 16535 8538 16541
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 8938 16532 8944 16584
rect 8996 16532 9002 16584
rect 8588 16504 8616 16532
rect 8404 16476 8616 16504
rect 9048 16504 9076 16612
rect 9140 16581 9168 16680
rect 9646 16584 9674 16680
rect 10042 16668 10048 16720
rect 10100 16708 10106 16720
rect 10594 16708 10600 16720
rect 10100 16680 10600 16708
rect 10100 16668 10106 16680
rect 10594 16668 10600 16680
rect 10652 16708 10658 16720
rect 12406 16708 12434 16748
rect 13998 16736 14004 16788
rect 14056 16776 14062 16788
rect 14182 16776 14188 16788
rect 14056 16748 14188 16776
rect 14056 16736 14062 16748
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 15194 16736 15200 16788
rect 15252 16776 15258 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 15252 16748 15393 16776
rect 15252 16736 15258 16748
rect 15381 16745 15393 16748
rect 15427 16745 15439 16779
rect 15381 16739 15439 16745
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 15528 16748 15669 16776
rect 15528 16736 15534 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 15657 16739 15715 16745
rect 16117 16779 16175 16785
rect 16117 16745 16129 16779
rect 16163 16776 16175 16779
rect 16206 16776 16212 16788
rect 16163 16748 16212 16776
rect 16163 16745 16175 16748
rect 16117 16739 16175 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 17126 16736 17132 16788
rect 17184 16736 17190 16788
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 17368 16748 17417 16776
rect 17368 16736 17374 16748
rect 17405 16745 17417 16748
rect 17451 16745 17463 16779
rect 17405 16739 17463 16745
rect 19242 16736 19248 16788
rect 19300 16736 19306 16788
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 21085 16779 21143 16785
rect 21085 16776 21097 16779
rect 20036 16748 21097 16776
rect 20036 16736 20042 16748
rect 21085 16745 21097 16748
rect 21131 16745 21143 16779
rect 21085 16739 21143 16745
rect 13906 16708 13912 16720
rect 10652 16680 11008 16708
rect 12406 16680 13912 16708
rect 10652 16668 10658 16680
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10502 16640 10508 16652
rect 10008 16612 10508 16640
rect 10008 16600 10014 16612
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16572 9183 16575
rect 9217 16575 9275 16581
rect 9217 16572 9229 16575
rect 9171 16544 9229 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9217 16541 9229 16544
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 9398 16532 9404 16584
rect 9456 16532 9462 16584
rect 9646 16544 9680 16584
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 10336 16581 10364 16612
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 10870 16600 10876 16652
rect 10928 16600 10934 16652
rect 10980 16649 11008 16680
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 14642 16668 14648 16720
rect 14700 16668 14706 16720
rect 15746 16708 15752 16720
rect 15488 16680 15752 16708
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 12158 16600 12164 16652
rect 12216 16640 12222 16652
rect 12805 16643 12863 16649
rect 12805 16640 12817 16643
rect 12216 16612 12817 16640
rect 12216 16600 12222 16612
rect 12805 16609 12817 16612
rect 12851 16609 12863 16643
rect 14660 16640 14688 16668
rect 14660 16612 15424 16640
rect 12805 16603 12863 16609
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9824 16544 9873 16572
rect 9824 16532 9830 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 9048 16476 9260 16504
rect 8113 16467 8171 16473
rect 3108 16408 3464 16436
rect 3605 16439 3663 16445
rect 3108 16396 3114 16408
rect 3605 16405 3617 16439
rect 3651 16436 3663 16439
rect 4706 16436 4712 16448
rect 3651 16408 4712 16436
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 4706 16396 4712 16408
rect 4764 16396 4770 16448
rect 4801 16439 4859 16445
rect 4801 16405 4813 16439
rect 4847 16436 4859 16439
rect 4890 16436 4896 16448
rect 4847 16408 4896 16436
rect 4847 16405 4859 16408
rect 4801 16399 4859 16405
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 7377 16439 7435 16445
rect 7377 16405 7389 16439
rect 7423 16436 7435 16439
rect 7466 16436 7472 16448
rect 7423 16408 7472 16436
rect 7423 16405 7435 16408
rect 7377 16399 7435 16405
rect 7466 16396 7472 16408
rect 7524 16396 7530 16448
rect 7742 16396 7748 16448
rect 7800 16396 7806 16448
rect 8018 16396 8024 16448
rect 8076 16436 8082 16448
rect 8128 16436 8156 16467
rect 9232 16448 9260 16476
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10152 16504 10180 16535
rect 10778 16532 10784 16584
rect 10836 16532 10842 16584
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11241 16575 11299 16581
rect 11241 16572 11253 16575
rect 11112 16544 11253 16572
rect 11112 16532 11118 16544
rect 11241 16541 11253 16544
rect 11287 16541 11299 16575
rect 11241 16535 11299 16541
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16572 11483 16575
rect 11514 16572 11520 16584
rect 11471 16544 11520 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 11698 16572 11704 16584
rect 11624 16544 11704 16572
rect 9640 16476 10180 16504
rect 10229 16507 10287 16513
rect 9640 16464 9646 16476
rect 10229 16473 10241 16507
rect 10275 16504 10287 16507
rect 11624 16504 11652 16544
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16572 12311 16575
rect 12526 16572 12532 16584
rect 12299 16544 12532 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 12894 16572 12900 16584
rect 12667 16544 12900 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 12894 16532 12900 16544
rect 12952 16532 12958 16584
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16572 13047 16575
rect 13170 16572 13176 16584
rect 13035 16544 13176 16572
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16541 13323 16575
rect 13265 16535 13323 16541
rect 10275 16476 11652 16504
rect 10275 16473 10287 16476
rect 10229 16467 10287 16473
rect 12710 16464 12716 16516
rect 12768 16504 12774 16516
rect 13280 16504 13308 16535
rect 13538 16532 13544 16584
rect 13596 16532 13602 16584
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13872 16544 14105 16572
rect 13872 16532 13878 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14642 16532 14648 16584
rect 14700 16532 14706 16584
rect 12768 16476 13308 16504
rect 12768 16464 12774 16476
rect 8076 16408 8156 16436
rect 8076 16396 8082 16408
rect 8202 16396 8208 16448
rect 8260 16396 8266 16448
rect 9122 16396 9128 16448
rect 9180 16396 9186 16448
rect 9214 16396 9220 16448
rect 9272 16396 9278 16448
rect 9769 16439 9827 16445
rect 9769 16405 9781 16439
rect 9815 16436 9827 16439
rect 9950 16436 9956 16448
rect 9815 16408 9956 16436
rect 9815 16405 9827 16408
rect 9769 16399 9827 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11020 16408 11897 16436
rect 11020 16396 11026 16408
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 11885 16399 11943 16405
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 14185 16439 14243 16445
rect 14185 16436 14197 16439
rect 12032 16408 14197 16436
rect 12032 16396 12038 16408
rect 14185 16405 14197 16408
rect 14231 16405 14243 16439
rect 14185 16399 14243 16405
rect 15194 16396 15200 16448
rect 15252 16396 15258 16448
rect 15396 16436 15424 16612
rect 15488 16581 15516 16680
rect 15746 16668 15752 16680
rect 15804 16668 15810 16720
rect 20346 16708 20352 16720
rect 16040 16680 20352 16708
rect 16040 16649 16068 16680
rect 20346 16668 20352 16680
rect 20404 16668 20410 16720
rect 21100 16708 21128 16739
rect 21174 16736 21180 16788
rect 21232 16776 21238 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 21232 16748 21281 16776
rect 21232 16736 21238 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 29733 16779 29791 16785
rect 29733 16776 29745 16779
rect 24084 16748 25452 16776
rect 24084 16736 24090 16748
rect 21726 16708 21732 16720
rect 21100 16680 21732 16708
rect 21726 16668 21732 16680
rect 21784 16668 21790 16720
rect 25424 16708 25452 16748
rect 27632 16748 29745 16776
rect 25869 16711 25927 16717
rect 25869 16708 25881 16711
rect 25424 16680 25881 16708
rect 25869 16677 25881 16680
rect 25915 16677 25927 16711
rect 25869 16671 25927 16677
rect 25958 16668 25964 16720
rect 26016 16708 26022 16720
rect 26053 16711 26111 16717
rect 26053 16708 26065 16711
rect 26016 16680 26065 16708
rect 26016 16668 26022 16680
rect 26053 16677 26065 16680
rect 26099 16677 26111 16711
rect 26053 16671 26111 16677
rect 16025 16643 16083 16649
rect 16025 16609 16037 16643
rect 16071 16609 16083 16643
rect 20254 16640 20260 16652
rect 16025 16603 16083 16609
rect 17604 16612 18000 16640
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16541 15531 16575
rect 15473 16535 15531 16541
rect 15562 16532 15568 16584
rect 15620 16532 15626 16584
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 15930 16572 15936 16584
rect 15887 16544 15936 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 17034 16532 17040 16584
rect 17092 16532 17098 16584
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 16114 16464 16120 16516
rect 16172 16464 16178 16516
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17144 16504 17172 16535
rect 17310 16532 17316 16584
rect 17368 16532 17374 16584
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 17604 16581 17632 16612
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 17552 16544 17601 16572
rect 17552 16532 17558 16544
rect 17589 16541 17601 16544
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 17862 16572 17868 16584
rect 17727 16544 17868 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 17972 16572 18000 16612
rect 19725 16612 20260 16640
rect 18141 16575 18199 16581
rect 18141 16572 18153 16575
rect 17972 16544 18153 16572
rect 18141 16541 18153 16544
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 18690 16532 18696 16584
rect 18748 16572 18754 16584
rect 18966 16572 18972 16584
rect 18748 16544 18972 16572
rect 18748 16532 18754 16544
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 19426 16532 19432 16584
rect 19484 16532 19490 16584
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16572 19579 16575
rect 19725 16572 19753 16612
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 25501 16643 25559 16649
rect 25501 16640 25513 16643
rect 22848 16612 25513 16640
rect 19567 16544 19753 16572
rect 19567 16541 19579 16544
rect 19521 16535 19579 16541
rect 19794 16532 19800 16584
rect 19852 16532 19858 16584
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 17000 16476 17172 16504
rect 17000 16464 17006 16476
rect 16206 16436 16212 16448
rect 15396 16408 16212 16436
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 16850 16396 16856 16448
rect 16908 16396 16914 16448
rect 17144 16436 17172 16476
rect 17405 16507 17463 16513
rect 17405 16473 17417 16507
rect 17451 16504 17463 16507
rect 17770 16504 17776 16516
rect 17451 16476 17776 16504
rect 17451 16473 17463 16476
rect 17405 16467 17463 16473
rect 17770 16464 17776 16476
rect 17828 16464 17834 16516
rect 17954 16464 17960 16516
rect 18012 16464 18018 16516
rect 18325 16507 18383 16513
rect 18325 16473 18337 16507
rect 18371 16473 18383 16507
rect 18325 16467 18383 16473
rect 17218 16436 17224 16448
rect 17144 16408 17224 16436
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 17865 16439 17923 16445
rect 17865 16436 17877 16439
rect 17736 16408 17877 16436
rect 17736 16396 17742 16408
rect 17865 16405 17877 16408
rect 17911 16405 17923 16439
rect 18340 16436 18368 16467
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 19150 16504 19156 16516
rect 18564 16476 19156 16504
rect 18564 16464 18570 16476
rect 19150 16464 19156 16476
rect 19208 16504 19214 16516
rect 19613 16507 19671 16513
rect 19613 16504 19625 16507
rect 19208 16476 19625 16504
rect 19208 16464 19214 16476
rect 19613 16473 19625 16476
rect 19659 16473 19671 16507
rect 19613 16467 19671 16473
rect 19702 16464 19708 16516
rect 19760 16504 19766 16516
rect 19904 16504 19932 16535
rect 20070 16532 20076 16584
rect 20128 16532 20134 16584
rect 20162 16532 20168 16584
rect 20220 16532 20226 16584
rect 20349 16575 20407 16581
rect 20349 16541 20361 16575
rect 20395 16572 20407 16575
rect 20622 16572 20628 16584
rect 20395 16544 20628 16572
rect 20395 16541 20407 16544
rect 20349 16535 20407 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 22848 16572 22876 16612
rect 25501 16609 25513 16612
rect 25547 16609 25559 16643
rect 26068 16640 26096 16671
rect 26068 16612 26280 16640
rect 25501 16603 25559 16609
rect 20732 16544 22876 16572
rect 20732 16504 20760 16544
rect 23290 16532 23296 16584
rect 23348 16532 23354 16584
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 19760 16476 19932 16504
rect 20456 16476 20760 16504
rect 20901 16507 20959 16513
rect 19760 16464 19766 16476
rect 20456 16436 20484 16476
rect 20901 16473 20913 16507
rect 20947 16504 20959 16507
rect 22738 16504 22744 16516
rect 20947 16476 22744 16504
rect 20947 16473 20959 16476
rect 20901 16467 20959 16473
rect 18340 16408 20484 16436
rect 17865 16399 17923 16405
rect 20530 16396 20536 16448
rect 20588 16396 20594 16448
rect 20622 16396 20628 16448
rect 20680 16436 20686 16448
rect 20916 16436 20944 16467
rect 22738 16464 22744 16476
rect 22796 16464 22802 16516
rect 23492 16504 23520 16535
rect 23566 16532 23572 16584
rect 23624 16532 23630 16584
rect 23658 16532 23664 16584
rect 23716 16532 23722 16584
rect 24854 16532 24860 16584
rect 24912 16572 24918 16584
rect 24949 16575 25007 16581
rect 24949 16572 24961 16575
rect 24912 16544 24961 16572
rect 24912 16532 24918 16544
rect 24949 16541 24961 16544
rect 24995 16541 25007 16575
rect 24949 16535 25007 16541
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 24026 16504 24032 16516
rect 23492 16476 24032 16504
rect 20680 16408 20944 16436
rect 21111 16439 21169 16445
rect 20680 16396 20686 16408
rect 21111 16405 21123 16439
rect 21157 16436 21169 16439
rect 21266 16436 21272 16448
rect 21157 16408 21272 16436
rect 21157 16405 21169 16408
rect 21111 16399 21169 16405
rect 21266 16396 21272 16408
rect 21324 16436 21330 16448
rect 21450 16436 21456 16448
rect 21324 16408 21456 16436
rect 21324 16396 21330 16408
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 21726 16396 21732 16448
rect 21784 16436 21790 16448
rect 23492 16436 23520 16476
rect 24026 16464 24032 16476
rect 24084 16464 24090 16516
rect 24394 16464 24400 16516
rect 24452 16464 24458 16516
rect 21784 16408 23520 16436
rect 23937 16439 23995 16445
rect 21784 16396 21790 16408
rect 23937 16405 23949 16439
rect 23983 16436 23995 16439
rect 25240 16436 25268 16535
rect 25406 16532 25412 16584
rect 25464 16532 25470 16584
rect 25682 16532 25688 16584
rect 25740 16532 25746 16584
rect 25958 16532 25964 16584
rect 26016 16532 26022 16584
rect 26252 16572 26280 16612
rect 27632 16584 27660 16748
rect 29733 16745 29745 16748
rect 29779 16745 29791 16779
rect 29733 16739 29791 16745
rect 32493 16779 32551 16785
rect 32493 16745 32505 16779
rect 32539 16776 32551 16779
rect 32582 16776 32588 16788
rect 32539 16748 32588 16776
rect 32539 16745 32551 16748
rect 32493 16739 32551 16745
rect 32582 16736 32588 16748
rect 32640 16736 32646 16788
rect 33410 16736 33416 16788
rect 33468 16736 33474 16788
rect 28261 16711 28319 16717
rect 28261 16677 28273 16711
rect 28307 16708 28319 16711
rect 34330 16708 34336 16720
rect 28307 16680 32536 16708
rect 28307 16677 28319 16680
rect 28261 16671 28319 16677
rect 28350 16600 28356 16652
rect 28408 16640 28414 16652
rect 28902 16640 28908 16652
rect 28408 16612 28908 16640
rect 28408 16600 28414 16612
rect 28902 16600 28908 16612
rect 28960 16640 28966 16652
rect 28960 16612 29776 16640
rect 28960 16600 28966 16612
rect 26513 16575 26571 16581
rect 26513 16572 26525 16575
rect 26252 16544 26525 16572
rect 26513 16541 26525 16544
rect 26559 16541 26571 16575
rect 26513 16535 26571 16541
rect 27614 16532 27620 16584
rect 27672 16532 27678 16584
rect 27798 16581 27804 16584
rect 27765 16575 27804 16581
rect 27765 16541 27777 16575
rect 27765 16535 27804 16541
rect 27798 16532 27804 16535
rect 27856 16532 27862 16584
rect 27890 16532 27896 16584
rect 27948 16532 27954 16584
rect 28074 16532 28080 16584
rect 28132 16581 28138 16584
rect 28132 16575 28181 16581
rect 28132 16541 28135 16575
rect 28169 16572 28181 16575
rect 29362 16572 29368 16584
rect 28169 16544 29368 16572
rect 28169 16541 28181 16544
rect 28132 16535 28181 16541
rect 28132 16532 28138 16535
rect 29362 16532 29368 16544
rect 29420 16532 29426 16584
rect 29748 16572 29776 16612
rect 29822 16600 29828 16652
rect 29880 16600 29886 16652
rect 29932 16612 32352 16640
rect 29932 16572 29960 16612
rect 29748 16544 29960 16572
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16572 30067 16575
rect 30098 16572 30104 16584
rect 30055 16544 30104 16572
rect 30055 16541 30067 16544
rect 30009 16535 30067 16541
rect 30098 16532 30104 16544
rect 30156 16532 30162 16584
rect 27430 16464 27436 16516
rect 27488 16504 27494 16516
rect 27985 16507 28043 16513
rect 27985 16504 27997 16507
rect 27488 16476 27997 16504
rect 27488 16464 27494 16476
rect 27985 16473 27997 16476
rect 28031 16473 28043 16507
rect 27985 16467 28043 16473
rect 29733 16507 29791 16513
rect 29733 16473 29745 16507
rect 29779 16504 29791 16507
rect 30282 16504 30288 16516
rect 29779 16476 30288 16504
rect 29779 16473 29791 16476
rect 29733 16467 29791 16473
rect 30282 16464 30288 16476
rect 30340 16464 30346 16516
rect 31846 16464 31852 16516
rect 31904 16504 31910 16516
rect 32217 16507 32275 16513
rect 32217 16504 32229 16507
rect 31904 16476 32229 16504
rect 31904 16464 31910 16476
rect 32217 16473 32229 16476
rect 32263 16473 32275 16507
rect 32324 16504 32352 16612
rect 32398 16600 32404 16652
rect 32456 16600 32462 16652
rect 32508 16581 32536 16680
rect 33336 16680 34336 16708
rect 33336 16640 33364 16680
rect 33060 16612 33364 16640
rect 32493 16575 32551 16581
rect 32493 16541 32505 16575
rect 32539 16572 32551 16575
rect 32950 16572 32956 16584
rect 32539 16544 32956 16572
rect 32539 16541 32551 16544
rect 32493 16535 32551 16541
rect 32950 16532 32956 16544
rect 33008 16532 33014 16584
rect 33060 16504 33088 16612
rect 33796 16581 33824 16680
rect 34330 16668 34336 16680
rect 34388 16668 34394 16720
rect 33597 16575 33655 16581
rect 33597 16572 33609 16575
rect 32324 16476 33088 16504
rect 33152 16544 33609 16572
rect 32217 16467 32275 16473
rect 23983 16408 25268 16436
rect 23983 16405 23995 16408
rect 23937 16399 23995 16405
rect 25682 16396 25688 16448
rect 25740 16436 25746 16448
rect 26329 16439 26387 16445
rect 26329 16436 26341 16439
rect 25740 16408 26341 16436
rect 25740 16396 25746 16408
rect 26329 16405 26341 16408
rect 26375 16405 26387 16439
rect 26329 16399 26387 16405
rect 30193 16439 30251 16445
rect 30193 16405 30205 16439
rect 30239 16436 30251 16439
rect 30650 16436 30656 16448
rect 30239 16408 30656 16436
rect 30239 16405 30251 16408
rect 30193 16399 30251 16405
rect 30650 16396 30656 16408
rect 30708 16396 30714 16448
rect 32490 16396 32496 16448
rect 32548 16436 32554 16448
rect 32677 16439 32735 16445
rect 32677 16436 32689 16439
rect 32548 16408 32689 16436
rect 32548 16396 32554 16408
rect 32677 16405 32689 16408
rect 32723 16405 32735 16439
rect 32677 16399 32735 16405
rect 32950 16396 32956 16448
rect 33008 16436 33014 16448
rect 33152 16436 33180 16544
rect 33597 16541 33609 16544
rect 33643 16541 33655 16575
rect 33597 16535 33655 16541
rect 33781 16575 33839 16581
rect 33781 16541 33793 16575
rect 33827 16541 33839 16575
rect 33781 16535 33839 16541
rect 34606 16532 34612 16584
rect 34664 16572 34670 16584
rect 34977 16575 35035 16581
rect 34977 16572 34989 16575
rect 34664 16544 34989 16572
rect 34664 16532 34670 16544
rect 34977 16541 34989 16544
rect 35023 16541 35035 16575
rect 35345 16575 35403 16581
rect 35345 16572 35357 16575
rect 34977 16535 35035 16541
rect 35084 16544 35357 16572
rect 33226 16464 33232 16516
rect 33284 16504 33290 16516
rect 34146 16504 34152 16516
rect 33284 16476 34152 16504
rect 33284 16464 33290 16476
rect 34146 16464 34152 16476
rect 34204 16504 34210 16516
rect 35084 16504 35112 16544
rect 35345 16541 35357 16544
rect 35391 16541 35403 16575
rect 35345 16535 35403 16541
rect 34204 16476 35112 16504
rect 34204 16464 34210 16476
rect 35158 16464 35164 16516
rect 35216 16464 35222 16516
rect 35250 16464 35256 16516
rect 35308 16464 35314 16516
rect 33008 16408 33180 16436
rect 33008 16396 33014 16408
rect 35342 16396 35348 16448
rect 35400 16436 35406 16448
rect 35529 16439 35587 16445
rect 35529 16436 35541 16439
rect 35400 16408 35541 16436
rect 35400 16396 35406 16408
rect 35529 16405 35541 16408
rect 35575 16405 35587 16439
rect 35529 16399 35587 16405
rect 1104 16346 36524 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 36524 16346
rect 1104 16272 36524 16294
rect 2590 16232 2596 16244
rect 1412 16204 2596 16232
rect 1412 16105 1440 16204
rect 2590 16192 2596 16204
rect 2648 16232 2654 16244
rect 3602 16232 3608 16244
rect 2648 16204 3608 16232
rect 2648 16192 2654 16204
rect 3602 16192 3608 16204
rect 3660 16232 3666 16244
rect 3660 16204 6224 16232
rect 3660 16192 3666 16204
rect 1670 16124 1676 16176
rect 1728 16124 1734 16176
rect 3050 16164 3056 16176
rect 2898 16136 3056 16164
rect 3050 16124 3056 16136
rect 3108 16124 3114 16176
rect 4614 16164 4620 16176
rect 3160 16136 4620 16164
rect 1397 16099 1455 16105
rect 1397 16065 1409 16099
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 3160 16037 3188 16136
rect 4614 16124 4620 16136
rect 4672 16124 4678 16176
rect 5350 16124 5356 16176
rect 5408 16124 5414 16176
rect 6196 16164 6224 16204
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 6328 16204 6377 16232
rect 6328 16192 6334 16204
rect 6365 16201 6377 16204
rect 6411 16201 6423 16235
rect 6365 16195 6423 16201
rect 6733 16235 6791 16241
rect 6733 16201 6745 16235
rect 6779 16232 6791 16235
rect 7466 16232 7472 16244
rect 6779 16204 7472 16232
rect 6779 16201 6791 16204
rect 6733 16195 6791 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 11974 16232 11980 16244
rect 7616 16204 11980 16232
rect 7616 16192 7622 16204
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 12802 16232 12808 16244
rect 12759 16204 12808 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 13814 16192 13820 16244
rect 13872 16192 13878 16244
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14366 16232 14372 16244
rect 14323 16204 14372 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 15565 16235 15623 16241
rect 15565 16201 15577 16235
rect 15611 16232 15623 16235
rect 16114 16232 16120 16244
rect 15611 16204 16120 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 17221 16235 17279 16241
rect 17221 16201 17233 16235
rect 17267 16232 17279 16235
rect 17494 16232 17500 16244
rect 17267 16204 17500 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 17678 16192 17684 16244
rect 17736 16232 17742 16244
rect 17736 16204 18828 16232
rect 17736 16192 17742 16204
rect 7006 16164 7012 16176
rect 6196 16136 7012 16164
rect 3786 16056 3792 16108
rect 3844 16056 3850 16108
rect 3878 16056 3884 16108
rect 3936 16056 3942 16108
rect 6196 16105 6224 16136
rect 7006 16124 7012 16136
rect 7064 16124 7070 16176
rect 13538 16164 13544 16176
rect 12544 16136 13544 16164
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16065 6239 16099
rect 6181 16059 6239 16065
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 7098 16096 7104 16108
rect 6871 16068 7104 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 8018 16056 8024 16108
rect 8076 16096 8082 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 8076 16068 8217 16096
rect 8076 16056 8082 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 8205 16059 8263 16065
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 8478 16096 8484 16108
rect 8435 16068 8484 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 9640 16068 10793 16096
rect 9640 16056 9646 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 3145 16031 3203 16037
rect 3145 15997 3157 16031
rect 3191 15997 3203 16031
rect 3145 15991 3203 15997
rect 4062 15988 4068 16040
rect 4120 15988 4126 16040
rect 5902 15988 5908 16040
rect 5960 15988 5966 16040
rect 6454 15988 6460 16040
rect 6512 15988 6518 16040
rect 6914 15988 6920 16040
rect 6972 15988 6978 16040
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 3418 15920 3424 15972
rect 3476 15920 3482 15972
rect 6472 15960 6500 15988
rect 7760 15960 7788 15991
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10594 16028 10600 16040
rect 9732 16000 10600 16028
rect 9732 15988 9738 16000
rect 10594 15988 10600 16000
rect 10652 16028 10658 16040
rect 10888 16028 10916 16059
rect 11054 16056 11060 16108
rect 11112 16056 11118 16108
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11514 16096 11520 16108
rect 11195 16068 11520 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 12161 16099 12219 16105
rect 12161 16065 12173 16099
rect 12207 16096 12219 16099
rect 12434 16096 12440 16108
rect 12207 16068 12440 16096
rect 12207 16065 12219 16068
rect 12161 16059 12219 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12544 16105 12572 16136
rect 13538 16124 13544 16136
rect 13596 16124 13602 16176
rect 13832 16164 13860 16192
rect 13998 16164 14004 16176
rect 13832 16136 14004 16164
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12710 16096 12716 16108
rect 12667 16068 12716 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12544 16028 12572 16059
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 13170 16096 13176 16108
rect 12943 16068 13176 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 13446 16056 13452 16108
rect 13504 16056 13510 16108
rect 13832 16105 13860 16136
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 16942 16164 16948 16176
rect 16816 16136 16948 16164
rect 16816 16124 16822 16136
rect 16942 16124 16948 16136
rect 17000 16164 17006 16176
rect 17589 16167 17647 16173
rect 17000 16136 17540 16164
rect 17000 16124 17006 16136
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 13906 16056 13912 16108
rect 13964 16096 13970 16108
rect 14093 16099 14151 16105
rect 14093 16096 14105 16099
rect 13964 16068 14105 16096
rect 13964 16056 13970 16068
rect 14093 16065 14105 16068
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 15105 16099 15163 16105
rect 15105 16065 15117 16099
rect 15151 16065 15163 16099
rect 15105 16059 15163 16065
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15562 16096 15568 16108
rect 15427 16068 15568 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 10652 16000 12572 16028
rect 12989 16031 13047 16037
rect 10652 15988 10658 16000
rect 12989 15997 13001 16031
rect 13035 16028 13047 16031
rect 13262 16028 13268 16040
rect 13035 16000 13268 16028
rect 13035 15997 13047 16000
rect 12989 15991 13047 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 6104 15932 7788 15960
rect 12069 15963 12127 15969
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 6104 15892 6132 15932
rect 12069 15929 12081 15963
rect 12115 15960 12127 15963
rect 12342 15960 12348 15972
rect 12115 15932 12348 15960
rect 12115 15929 12127 15932
rect 12069 15923 12127 15929
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 12802 15920 12808 15972
rect 12860 15960 12866 15972
rect 13357 15963 13415 15969
rect 13357 15960 13369 15963
rect 12860 15932 13369 15960
rect 12860 15920 12866 15932
rect 13357 15929 13369 15932
rect 13403 15929 13415 15963
rect 13357 15923 13415 15929
rect 14826 15920 14832 15972
rect 14884 15960 14890 15972
rect 15120 15960 15148 16059
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 16206 16056 16212 16108
rect 16264 16096 16270 16108
rect 16264 16068 17356 16096
rect 16264 16056 16270 16068
rect 15289 16031 15347 16037
rect 15289 15997 15301 16031
rect 15335 16028 15347 16031
rect 16666 16028 16672 16040
rect 15335 16000 16672 16028
rect 15335 15997 15347 16000
rect 15289 15991 15347 15997
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 17328 16028 17356 16068
rect 17402 16056 17408 16108
rect 17460 16056 17466 16108
rect 17512 16105 17540 16136
rect 17589 16133 17601 16167
rect 17635 16164 17647 16167
rect 17862 16164 17868 16176
rect 17635 16136 17868 16164
rect 17635 16133 17647 16136
rect 17589 16127 17647 16133
rect 17862 16124 17868 16136
rect 17920 16124 17926 16176
rect 18690 16124 18696 16176
rect 18748 16124 18754 16176
rect 18800 16164 18828 16204
rect 19150 16192 19156 16244
rect 19208 16192 19214 16244
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 20530 16232 20536 16244
rect 19300 16204 20536 16232
rect 19300 16192 19306 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 23382 16192 23388 16244
rect 23440 16232 23446 16244
rect 24121 16235 24179 16241
rect 24121 16232 24133 16235
rect 23440 16204 24133 16232
rect 23440 16192 23446 16204
rect 24121 16201 24133 16204
rect 24167 16201 24179 16235
rect 24121 16195 24179 16201
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 25130 16232 25136 16244
rect 24820 16204 25136 16232
rect 24820 16192 24826 16204
rect 25130 16192 25136 16204
rect 25188 16232 25194 16244
rect 25188 16204 25268 16232
rect 25188 16192 25194 16204
rect 19613 16167 19671 16173
rect 18800 16136 19564 16164
rect 17497 16099 17555 16105
rect 17497 16065 17509 16099
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16096 17831 16099
rect 17954 16096 17960 16108
rect 17819 16068 17960 16096
rect 17819 16065 17831 16068
rect 17773 16059 17831 16065
rect 17954 16056 17960 16068
rect 18012 16096 18018 16108
rect 18506 16096 18512 16108
rect 18012 16068 18512 16096
rect 18012 16056 18018 16068
rect 18506 16056 18512 16068
rect 18564 16056 18570 16108
rect 18966 16056 18972 16108
rect 19024 16056 19030 16108
rect 19426 16105 19432 16108
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19393 16099 19432 16105
rect 19393 16065 19405 16099
rect 19393 16059 19432 16065
rect 18782 16028 18788 16040
rect 17328 16000 18788 16028
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 19150 16028 19156 16040
rect 18892 16000 19156 16028
rect 18892 15960 18920 16000
rect 19150 15988 19156 16000
rect 19208 16028 19214 16040
rect 19260 16028 19288 16059
rect 19426 16056 19432 16059
rect 19484 16056 19490 16108
rect 19536 16105 19564 16136
rect 19613 16133 19625 16167
rect 19659 16164 19671 16167
rect 20070 16164 20076 16176
rect 19659 16136 20076 16164
rect 19659 16133 19671 16136
rect 19613 16127 19671 16133
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 22830 16164 22836 16176
rect 20916 16136 22836 16164
rect 19521 16099 19579 16105
rect 19521 16065 19533 16099
rect 19567 16065 19579 16099
rect 19521 16059 19579 16065
rect 19208 16000 19288 16028
rect 19536 16028 19564 16059
rect 19702 16056 19708 16108
rect 19760 16105 19766 16108
rect 19760 16096 19768 16105
rect 20916 16096 20944 16136
rect 22830 16124 22836 16136
rect 22888 16124 22894 16176
rect 25038 16173 25044 16176
rect 25025 16167 25044 16173
rect 25025 16133 25037 16167
rect 25025 16127 25044 16133
rect 23477 16121 23535 16127
rect 25038 16124 25044 16127
rect 25096 16124 25102 16176
rect 25240 16173 25268 16204
rect 25774 16192 25780 16244
rect 25832 16192 25838 16244
rect 27614 16192 27620 16244
rect 27672 16192 27678 16244
rect 27890 16232 27896 16244
rect 27724 16204 27896 16232
rect 25225 16167 25283 16173
rect 25225 16133 25237 16167
rect 25271 16133 25283 16167
rect 26237 16167 26295 16173
rect 26237 16164 26249 16167
rect 25225 16127 25283 16133
rect 25608 16136 26249 16164
rect 19760 16068 19805 16096
rect 19895 16068 20944 16096
rect 19760 16059 19768 16068
rect 19760 16056 19766 16059
rect 19895 16028 19923 16068
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21048 16068 22017 16096
rect 21048 16056 21054 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19536 16000 19923 16028
rect 19208 15988 19214 16000
rect 19980 15997 19993 16028
rect 20027 15997 20039 16031
rect 19980 15991 20039 15997
rect 19794 15960 19800 15972
rect 14884 15932 18920 15960
rect 18984 15932 19800 15960
rect 14884 15920 14890 15932
rect 4479 15864 6132 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 6454 15852 6460 15904
rect 6512 15892 6518 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 6512 15864 7205 15892
rect 6512 15852 6518 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7193 15855 7251 15861
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 10597 15895 10655 15901
rect 10597 15861 10609 15895
rect 10643 15892 10655 15895
rect 10686 15892 10692 15904
rect 10643 15864 10692 15892
rect 10643 15861 10655 15864
rect 10597 15855 10655 15861
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12986 15892 12992 15904
rect 12299 15864 12992 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 12986 15852 12992 15864
rect 13044 15852 13050 15904
rect 15378 15852 15384 15904
rect 15436 15852 15442 15904
rect 18984 15901 19012 15932
rect 19794 15920 19800 15932
rect 19852 15920 19858 15972
rect 19886 15920 19892 15972
rect 19944 15920 19950 15972
rect 18969 15895 19027 15901
rect 18969 15861 18981 15895
rect 19015 15861 19027 15895
rect 18969 15855 19027 15861
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19702 15892 19708 15904
rect 19392 15864 19708 15892
rect 19392 15852 19398 15864
rect 19702 15852 19708 15864
rect 19760 15892 19766 15904
rect 19980 15892 20008 15991
rect 20162 15988 20168 16040
rect 20220 16028 20226 16040
rect 20257 16031 20315 16037
rect 20257 16028 20269 16031
rect 20220 16000 20269 16028
rect 20220 15988 20226 16000
rect 20257 15997 20269 16000
rect 20303 15997 20315 16031
rect 20257 15991 20315 15997
rect 21818 15988 21824 16040
rect 21876 15988 21882 16040
rect 22204 16028 22232 16059
rect 22278 16056 22284 16108
rect 22336 16056 22342 16108
rect 23477 16087 23489 16121
rect 23523 16087 23535 16121
rect 23477 16081 23535 16087
rect 23492 16040 23520 16081
rect 23658 16056 23664 16108
rect 23716 16056 23722 16108
rect 24118 16056 24124 16108
rect 24176 16096 24182 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 24176 16068 24317 16096
rect 24176 16056 24182 16068
rect 24305 16065 24317 16068
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 24397 16099 24455 16105
rect 24397 16065 24409 16099
rect 24443 16065 24455 16099
rect 24397 16059 24455 16065
rect 23290 16028 23296 16040
rect 22204 16000 23296 16028
rect 23290 15988 23296 16000
rect 23348 15988 23354 16040
rect 23474 15988 23480 16040
rect 23532 15988 23538 16040
rect 22278 15920 22284 15972
rect 22336 15960 22342 15972
rect 23845 15963 23903 15969
rect 22336 15932 23612 15960
rect 22336 15920 22342 15932
rect 19760 15864 20008 15892
rect 19760 15852 19766 15864
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 23477 15895 23535 15901
rect 23477 15892 23489 15895
rect 20128 15864 23489 15892
rect 20128 15852 20134 15864
rect 23477 15861 23489 15864
rect 23523 15861 23535 15895
rect 23584 15892 23612 15932
rect 23845 15929 23857 15963
rect 23891 15960 23903 15963
rect 24302 15960 24308 15972
rect 23891 15932 24308 15960
rect 23891 15929 23903 15932
rect 23845 15923 23903 15929
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 24412 15960 24440 16059
rect 24486 16056 24492 16108
rect 24544 16056 24550 16108
rect 24578 16056 24584 16108
rect 24636 16105 24642 16108
rect 25608 16105 25636 16136
rect 26237 16133 26249 16136
rect 26283 16133 26295 16167
rect 26237 16127 26295 16133
rect 26326 16124 26332 16176
rect 26384 16164 26390 16176
rect 26384 16136 26556 16164
rect 26384 16124 26390 16136
rect 24636 16099 24665 16105
rect 24653 16065 24665 16099
rect 24636 16059 24665 16065
rect 25593 16099 25651 16105
rect 25593 16065 25605 16099
rect 25639 16065 25651 16099
rect 25593 16059 25651 16065
rect 24636 16056 24642 16059
rect 25682 16056 25688 16108
rect 25740 16096 25746 16108
rect 26528 16105 26556 16136
rect 25777 16099 25835 16105
rect 25777 16096 25789 16099
rect 25740 16068 25789 16096
rect 25740 16056 25746 16068
rect 25777 16065 25789 16068
rect 25823 16065 25835 16099
rect 25777 16059 25835 16065
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 26513 16099 26571 16105
rect 26513 16065 26525 16099
rect 26559 16096 26571 16099
rect 26602 16096 26608 16108
rect 26559 16068 26608 16096
rect 26559 16065 26571 16068
rect 26513 16059 26571 16065
rect 24765 16031 24823 16037
rect 24765 15997 24777 16031
rect 24811 16028 24823 16031
rect 24811 16000 25452 16028
rect 24811 15997 24823 16000
rect 24765 15991 24823 15997
rect 24412 15932 25084 15960
rect 25056 15901 25084 15932
rect 24857 15895 24915 15901
rect 24857 15892 24869 15895
rect 23584 15864 24869 15892
rect 23477 15855 23535 15861
rect 24857 15861 24869 15864
rect 24903 15861 24915 15895
rect 24857 15855 24915 15861
rect 25041 15895 25099 15901
rect 25041 15861 25053 15895
rect 25087 15892 25099 15895
rect 25314 15892 25320 15904
rect 25087 15864 25320 15892
rect 25087 15861 25099 15864
rect 25041 15855 25099 15861
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 25424 15892 25452 16000
rect 26142 15988 26148 16040
rect 26200 15988 26206 16040
rect 26436 16028 26464 16059
rect 26602 16056 26608 16068
rect 26660 16056 26666 16108
rect 26694 16056 26700 16108
rect 26752 16056 26758 16108
rect 26786 16056 26792 16108
rect 26844 16056 26850 16108
rect 27614 16028 27620 16040
rect 26436 16000 27620 16028
rect 27614 15988 27620 16000
rect 27672 15988 27678 16040
rect 27724 16028 27752 16204
rect 27890 16192 27896 16204
rect 27948 16232 27954 16244
rect 29457 16235 29515 16241
rect 27948 16204 29132 16232
rect 27948 16192 27954 16204
rect 28074 16164 28080 16176
rect 27816 16136 28080 16164
rect 27816 16105 27844 16136
rect 28074 16124 28080 16136
rect 28132 16124 28138 16176
rect 29104 16173 29132 16204
rect 29457 16201 29469 16235
rect 29503 16232 29515 16235
rect 29822 16232 29828 16244
rect 29503 16204 29828 16232
rect 29503 16201 29515 16204
rect 29457 16195 29515 16201
rect 29822 16192 29828 16204
rect 29880 16192 29886 16244
rect 30208 16204 31754 16232
rect 29089 16167 29147 16173
rect 29089 16133 29101 16167
rect 29135 16164 29147 16167
rect 30208 16164 30236 16204
rect 29135 16136 30236 16164
rect 29135 16133 29147 16136
rect 29089 16127 29147 16133
rect 30558 16124 30564 16176
rect 30616 16164 30622 16176
rect 30742 16164 30748 16176
rect 30616 16136 30748 16164
rect 30616 16124 30622 16136
rect 30742 16124 30748 16136
rect 30800 16164 30806 16176
rect 31297 16167 31355 16173
rect 31297 16164 31309 16167
rect 30800 16136 31309 16164
rect 30800 16124 30806 16136
rect 31297 16133 31309 16136
rect 31343 16133 31355 16167
rect 31297 16127 31355 16133
rect 27801 16099 27859 16105
rect 27801 16065 27813 16099
rect 27847 16065 27859 16099
rect 27801 16059 27859 16065
rect 27890 16056 27896 16108
rect 27948 16056 27954 16108
rect 27985 16099 28043 16105
rect 27985 16065 27997 16099
rect 28031 16065 28043 16099
rect 27985 16059 28043 16065
rect 28169 16099 28227 16105
rect 28169 16065 28181 16099
rect 28215 16096 28227 16099
rect 28442 16096 28448 16108
rect 28215 16068 28448 16096
rect 28215 16065 28227 16068
rect 28169 16059 28227 16065
rect 28000 16028 28028 16059
rect 28442 16056 28448 16068
rect 28500 16096 28506 16108
rect 28626 16096 28632 16108
rect 28500 16068 28632 16096
rect 28500 16056 28506 16068
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 28905 16099 28963 16105
rect 28905 16065 28917 16099
rect 28951 16065 28963 16099
rect 28905 16059 28963 16065
rect 27724 16000 28028 16028
rect 28920 16028 28948 16059
rect 29178 16056 29184 16108
rect 29236 16056 29242 16108
rect 29273 16099 29331 16105
rect 29273 16065 29285 16099
rect 29319 16096 29331 16099
rect 29362 16096 29368 16108
rect 29319 16068 29368 16096
rect 29319 16065 29331 16068
rect 29273 16059 29331 16065
rect 29362 16056 29368 16068
rect 29420 16056 29426 16108
rect 30374 16056 30380 16108
rect 30432 16096 30438 16108
rect 30653 16099 30711 16105
rect 30653 16096 30665 16099
rect 30432 16068 30665 16096
rect 30432 16056 30438 16068
rect 30653 16065 30665 16068
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30837 16099 30895 16105
rect 30837 16065 30849 16099
rect 30883 16096 30895 16099
rect 30926 16096 30932 16108
rect 30883 16068 30932 16096
rect 30883 16065 30895 16068
rect 30837 16059 30895 16065
rect 30926 16056 30932 16068
rect 30984 16056 30990 16108
rect 31113 16102 31171 16105
rect 31202 16102 31208 16108
rect 31113 16099 31208 16102
rect 31113 16096 31125 16099
rect 31036 16068 31125 16096
rect 29914 16028 29920 16040
rect 28920 16000 29920 16028
rect 29914 15988 29920 16000
rect 29972 16028 29978 16040
rect 30190 16028 30196 16040
rect 29972 16000 30196 16028
rect 29972 15988 29978 16000
rect 30190 15988 30196 16000
rect 30248 15988 30254 16040
rect 30558 15988 30564 16040
rect 30616 16028 30622 16040
rect 31036 16028 31064 16068
rect 31113 16065 31125 16068
rect 31159 16074 31208 16099
rect 31159 16065 31171 16074
rect 31113 16059 31171 16065
rect 31202 16056 31208 16074
rect 31260 16056 31266 16108
rect 31386 16056 31392 16108
rect 31444 16056 31450 16108
rect 31481 16099 31539 16105
rect 31481 16065 31493 16099
rect 31527 16086 31539 16099
rect 31570 16086 31576 16108
rect 31527 16065 31576 16086
rect 31481 16059 31576 16065
rect 31501 16058 31576 16059
rect 31570 16056 31576 16058
rect 31628 16056 31634 16108
rect 30616 16000 31064 16028
rect 30616 15988 30622 16000
rect 25958 15920 25964 15972
rect 26016 15960 26022 15972
rect 30098 15960 30104 15972
rect 26016 15932 30104 15960
rect 26016 15920 26022 15932
rect 30098 15920 30104 15932
rect 30156 15920 30162 15972
rect 31726 15960 31754 16204
rect 31938 16192 31944 16244
rect 31996 16232 32002 16244
rect 32766 16232 32772 16244
rect 31996 16204 32772 16232
rect 31996 16192 32002 16204
rect 32766 16192 32772 16204
rect 32824 16192 32830 16244
rect 34514 16192 34520 16244
rect 34572 16232 34578 16244
rect 34698 16232 34704 16244
rect 34572 16204 34704 16232
rect 34572 16192 34578 16204
rect 34698 16192 34704 16204
rect 34756 16192 34762 16244
rect 33318 15988 33324 16040
rect 33376 16028 33382 16040
rect 34422 16028 34428 16040
rect 33376 16000 34428 16028
rect 33376 15988 33382 16000
rect 34422 15988 34428 16000
rect 34480 15988 34486 16040
rect 35158 15960 35164 15972
rect 31726 15932 35164 15960
rect 35158 15920 35164 15932
rect 35216 15920 35222 15972
rect 28350 15892 28356 15904
rect 25424 15864 28356 15892
rect 28350 15852 28356 15864
rect 28408 15852 28414 15904
rect 30650 15852 30656 15904
rect 30708 15852 30714 15904
rect 31021 15895 31079 15901
rect 31021 15861 31033 15895
rect 31067 15892 31079 15895
rect 31570 15892 31576 15904
rect 31067 15864 31576 15892
rect 31067 15861 31079 15864
rect 31021 15855 31079 15861
rect 31570 15852 31576 15864
rect 31628 15852 31634 15904
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15892 31723 15895
rect 31846 15892 31852 15904
rect 31711 15864 31852 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 31846 15852 31852 15864
rect 31904 15852 31910 15904
rect 1104 15802 36524 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 36524 15802
rect 1104 15728 36524 15750
rect 3786 15648 3792 15700
rect 3844 15648 3850 15700
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 6089 15691 6147 15697
rect 6089 15688 6101 15691
rect 5960 15660 6101 15688
rect 5960 15648 5966 15660
rect 6089 15657 6101 15660
rect 6135 15657 6147 15691
rect 8570 15688 8576 15700
rect 6089 15651 6147 15657
rect 7668 15660 8576 15688
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4706 15552 4712 15564
rect 4479 15524 4712 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15552 6791 15555
rect 6914 15552 6920 15564
rect 6779 15524 6920 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 6914 15512 6920 15524
rect 6972 15552 6978 15564
rect 7668 15552 7696 15660
rect 8570 15648 8576 15660
rect 8628 15688 8634 15700
rect 8628 15660 12434 15688
rect 8628 15648 8634 15660
rect 8113 15623 8171 15629
rect 8113 15589 8125 15623
rect 8159 15620 8171 15623
rect 8202 15620 8208 15632
rect 8159 15592 8208 15620
rect 8159 15589 8171 15592
rect 8113 15583 8171 15589
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 10134 15620 10140 15632
rect 8444 15592 9260 15620
rect 8444 15580 8450 15592
rect 6972 15524 7696 15552
rect 6972 15512 6978 15524
rect 7742 15512 7748 15564
rect 7800 15512 7806 15564
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 8754 15552 8760 15564
rect 8619 15524 8760 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 6454 15444 6460 15496
rect 6512 15444 6518 15496
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15484 6607 15487
rect 6595 15456 8245 15484
rect 6595 15453 6607 15456
rect 6549 15447 6607 15453
rect 8217 15416 8245 15456
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 8352 15456 8493 15484
rect 8352 15444 8358 15456
rect 8481 15453 8493 15456
rect 8527 15453 8539 15487
rect 8481 15447 8539 15453
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 8846 15484 8852 15496
rect 8711 15456 8852 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 9232 15493 9260 15592
rect 9876 15592 10140 15620
rect 9398 15512 9404 15564
rect 9456 15512 9462 15564
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8996 15456 9137 15484
rect 8996 15444 9002 15456
rect 9125 15453 9137 15456
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 9674 15444 9680 15496
rect 9732 15444 9738 15496
rect 9876 15493 9904 15592
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 12406 15620 12434 15660
rect 12710 15648 12716 15700
rect 12768 15648 12774 15700
rect 12894 15648 12900 15700
rect 12952 15648 12958 15700
rect 14642 15648 14648 15700
rect 14700 15688 14706 15700
rect 15010 15688 15016 15700
rect 14700 15660 15016 15688
rect 14700 15648 14706 15660
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 15470 15648 15476 15700
rect 15528 15688 15534 15700
rect 16301 15691 16359 15697
rect 15528 15660 15976 15688
rect 15528 15648 15534 15660
rect 12618 15620 12624 15632
rect 12406 15592 12624 15620
rect 12618 15580 12624 15592
rect 12676 15580 12682 15632
rect 12728 15620 12756 15648
rect 13078 15620 13084 15632
rect 12728 15592 13084 15620
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 14734 15580 14740 15632
rect 14792 15620 14798 15632
rect 15841 15623 15899 15629
rect 15841 15620 15853 15623
rect 14792 15592 15853 15620
rect 14792 15580 14798 15592
rect 15841 15589 15853 15592
rect 15887 15589 15899 15623
rect 15948 15620 15976 15660
rect 16301 15657 16313 15691
rect 16347 15688 16359 15691
rect 16390 15688 16396 15700
rect 16347 15660 16396 15688
rect 16347 15657 16359 15660
rect 16301 15651 16359 15657
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 17126 15648 17132 15700
rect 17184 15688 17190 15700
rect 17497 15691 17555 15697
rect 17497 15688 17509 15691
rect 17184 15660 17509 15688
rect 17184 15648 17190 15660
rect 17497 15657 17509 15660
rect 17543 15657 17555 15691
rect 17497 15651 17555 15657
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 20441 15691 20499 15697
rect 20441 15688 20453 15691
rect 18840 15660 20453 15688
rect 18840 15648 18846 15660
rect 20441 15657 20453 15660
rect 20487 15688 20499 15691
rect 20898 15688 20904 15700
rect 20487 15660 20904 15688
rect 20487 15657 20499 15660
rect 20441 15651 20499 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 21729 15691 21787 15697
rect 21729 15657 21741 15691
rect 21775 15688 21787 15691
rect 21910 15688 21916 15700
rect 21775 15660 21916 15688
rect 21775 15657 21787 15660
rect 21729 15651 21787 15657
rect 21910 15648 21916 15660
rect 21968 15648 21974 15700
rect 22370 15648 22376 15700
rect 22428 15688 22434 15700
rect 22649 15691 22707 15697
rect 22649 15688 22661 15691
rect 22428 15660 22661 15688
rect 22428 15648 22434 15660
rect 22649 15657 22661 15660
rect 22695 15688 22707 15691
rect 23106 15688 23112 15700
rect 22695 15660 23112 15688
rect 22695 15657 22707 15660
rect 22649 15651 22707 15657
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 25406 15648 25412 15700
rect 25464 15688 25470 15700
rect 25961 15691 26019 15697
rect 25961 15688 25973 15691
rect 25464 15660 25973 15688
rect 25464 15648 25470 15660
rect 25961 15657 25973 15660
rect 26007 15657 26019 15691
rect 25961 15651 26019 15657
rect 26142 15648 26148 15700
rect 26200 15688 26206 15700
rect 26513 15691 26571 15697
rect 26513 15688 26525 15691
rect 26200 15660 26525 15688
rect 26200 15648 26206 15660
rect 26513 15657 26525 15660
rect 26559 15657 26571 15691
rect 26513 15651 26571 15657
rect 27249 15691 27307 15697
rect 27249 15657 27261 15691
rect 27295 15688 27307 15691
rect 27890 15688 27896 15700
rect 27295 15660 27896 15688
rect 27295 15657 27307 15660
rect 27249 15651 27307 15657
rect 16482 15620 16488 15632
rect 15948 15592 16488 15620
rect 15841 15583 15899 15589
rect 16482 15580 16488 15592
rect 16540 15580 16546 15632
rect 17034 15580 17040 15632
rect 17092 15620 17098 15632
rect 19518 15620 19524 15632
rect 17092 15592 19524 15620
rect 17092 15580 17098 15592
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 19794 15580 19800 15632
rect 19852 15620 19858 15632
rect 22278 15620 22284 15632
rect 19852 15592 22284 15620
rect 19852 15580 19858 15592
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 26329 15623 26387 15629
rect 26329 15589 26341 15623
rect 26375 15620 26387 15623
rect 27264 15620 27292 15651
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 30098 15648 30104 15700
rect 30156 15688 30162 15700
rect 31386 15688 31392 15700
rect 30156 15660 31392 15688
rect 30156 15648 30162 15660
rect 31386 15648 31392 15660
rect 31444 15648 31450 15700
rect 31478 15648 31484 15700
rect 31536 15648 31542 15700
rect 33318 15688 33324 15700
rect 31588 15660 33324 15688
rect 31588 15620 31616 15660
rect 33318 15648 33324 15660
rect 33376 15648 33382 15700
rect 26375 15592 27292 15620
rect 27356 15592 31616 15620
rect 26375 15589 26387 15592
rect 26329 15583 26387 15589
rect 10962 15552 10968 15564
rect 9968 15524 10364 15552
rect 9968 15496 9996 15524
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 9950 15444 9956 15496
rect 10008 15444 10014 15496
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10336 15493 10364 15524
rect 10520 15524 10968 15552
rect 10520 15496 10548 15524
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15552 12403 15555
rect 12713 15555 12771 15561
rect 12391 15524 12664 15552
rect 12391 15521 12403 15524
rect 12345 15515 12403 15521
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10410 15484 10416 15496
rect 10367 15456 10416 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 10502 15444 10508 15496
rect 10560 15444 10566 15496
rect 10686 15493 10692 15496
rect 10659 15487 10692 15493
rect 10659 15453 10671 15487
rect 10659 15447 10692 15453
rect 10686 15444 10692 15447
rect 10744 15444 10750 15496
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12268 15416 12296 15447
rect 12434 15444 12440 15496
rect 12492 15444 12498 15496
rect 12526 15444 12532 15496
rect 12584 15444 12590 15496
rect 12636 15484 12664 15524
rect 12713 15521 12725 15555
rect 12759 15552 12771 15555
rect 12802 15552 12808 15564
rect 12759 15524 12808 15552
rect 12759 15521 12771 15524
rect 12713 15515 12771 15521
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 16666 15552 16672 15564
rect 15335 15524 16672 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 17865 15555 17923 15561
rect 17865 15552 17877 15555
rect 17420 15524 17877 15552
rect 17420 15496 17448 15524
rect 17865 15521 17877 15524
rect 17911 15521 17923 15555
rect 17865 15515 17923 15521
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15552 18015 15555
rect 18138 15552 18144 15564
rect 18003 15524 18144 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 18138 15512 18144 15524
rect 18196 15512 18202 15564
rect 18506 15512 18512 15564
rect 18564 15552 18570 15564
rect 19426 15552 19432 15564
rect 18564 15524 19432 15552
rect 18564 15512 18570 15524
rect 19426 15512 19432 15524
rect 19484 15552 19490 15564
rect 23842 15552 23848 15564
rect 19484 15524 20208 15552
rect 19484 15512 19490 15524
rect 12636 15456 12940 15484
rect 12713 15419 12771 15425
rect 12713 15416 12725 15419
rect 8217 15388 12112 15416
rect 12268 15388 12725 15416
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 7708 15320 8217 15348
rect 7708 15308 7714 15320
rect 8205 15317 8217 15320
rect 8251 15348 8263 15351
rect 8386 15348 8392 15360
rect 8251 15320 8392 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8536 15320 8953 15348
rect 8536 15308 8542 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 9398 15308 9404 15360
rect 9456 15348 9462 15360
rect 10229 15351 10287 15357
rect 10229 15348 10241 15351
rect 9456 15320 10241 15348
rect 9456 15308 9462 15320
rect 10229 15317 10241 15320
rect 10275 15317 10287 15351
rect 10229 15311 10287 15317
rect 10870 15308 10876 15360
rect 10928 15308 10934 15360
rect 12084 15357 12112 15388
rect 12713 15385 12725 15388
rect 12759 15385 12771 15419
rect 12912 15416 12940 15456
rect 12986 15444 12992 15496
rect 13044 15444 13050 15496
rect 15378 15444 15384 15496
rect 15436 15444 15442 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 15838 15444 15844 15496
rect 15896 15484 15902 15496
rect 16025 15487 16083 15493
rect 16025 15484 16037 15487
rect 15896 15456 16037 15484
rect 15896 15444 15902 15456
rect 16025 15453 16037 15456
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 16117 15487 16175 15493
rect 16117 15453 16129 15487
rect 16163 15484 16175 15487
rect 16206 15484 16212 15496
rect 16163 15456 16212 15484
rect 16163 15453 16175 15456
rect 16117 15447 16175 15453
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 17402 15444 17408 15496
rect 17460 15444 17466 15496
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15484 17739 15487
rect 18524 15484 18552 15512
rect 17727 15456 18552 15484
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 19794 15444 19800 15496
rect 19852 15444 19858 15496
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 20180 15493 20208 15524
rect 20364 15524 23848 15552
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15484 20223 15487
rect 20254 15484 20260 15496
rect 20211 15456 20260 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 13354 15416 13360 15428
rect 12912 15388 13360 15416
rect 12713 15379 12771 15385
rect 13354 15376 13360 15388
rect 13412 15376 13418 15428
rect 15396 15416 15424 15444
rect 16298 15416 16304 15428
rect 15396 15388 16304 15416
rect 16298 15376 16304 15388
rect 16356 15376 16362 15428
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 19426 15416 19432 15428
rect 18012 15388 19432 15416
rect 18012 15376 18018 15388
rect 19426 15376 19432 15388
rect 19484 15376 19490 15428
rect 20088 15416 20116 15447
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20364 15416 20392 15524
rect 20824 15496 20852 15524
rect 23842 15512 23848 15524
rect 23900 15512 23906 15564
rect 25038 15512 25044 15564
rect 25096 15552 25102 15564
rect 27356 15552 27384 15592
rect 31662 15580 31668 15632
rect 31720 15620 31726 15632
rect 36170 15620 36176 15632
rect 31720 15592 36176 15620
rect 31720 15580 31726 15592
rect 36170 15580 36176 15592
rect 36228 15580 36234 15632
rect 28994 15552 29000 15564
rect 25096 15524 27384 15552
rect 28552 15524 29000 15552
rect 25096 15512 25102 15524
rect 20806 15444 20812 15496
rect 20864 15444 20870 15496
rect 21358 15444 21364 15496
rect 21416 15484 21422 15496
rect 21818 15484 21824 15496
rect 21416 15456 21824 15484
rect 21416 15444 21422 15456
rect 21818 15444 21824 15456
rect 21876 15484 21882 15496
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21876 15456 22017 15484
rect 21876 15444 21882 15456
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 22005 15447 22063 15453
rect 22094 15444 22100 15496
rect 22152 15444 22158 15496
rect 22186 15444 22192 15496
rect 22244 15444 22250 15496
rect 22465 15487 22523 15493
rect 22465 15453 22477 15487
rect 22511 15484 22523 15487
rect 22646 15484 22652 15496
rect 22511 15456 22652 15484
rect 22511 15453 22523 15456
rect 22465 15447 22523 15453
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 22830 15444 22836 15496
rect 22888 15484 22894 15496
rect 24762 15484 24768 15496
rect 22888 15456 24768 15484
rect 22888 15444 22894 15456
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 25682 15444 25688 15496
rect 25740 15484 25746 15496
rect 26145 15487 26203 15493
rect 26145 15484 26157 15487
rect 25740 15456 26157 15484
rect 25740 15444 25746 15456
rect 26145 15453 26157 15456
rect 26191 15453 26203 15487
rect 26145 15447 26203 15453
rect 26418 15444 26424 15496
rect 26476 15444 26482 15496
rect 26697 15487 26755 15493
rect 26697 15453 26709 15487
rect 26743 15453 26755 15487
rect 26697 15447 26755 15453
rect 20088 15388 20392 15416
rect 22738 15376 22744 15428
rect 22796 15376 22802 15428
rect 24486 15376 24492 15428
rect 24544 15416 24550 15428
rect 26712 15416 26740 15447
rect 26786 15444 26792 15496
rect 26844 15484 26850 15496
rect 26881 15487 26939 15493
rect 26881 15484 26893 15487
rect 26844 15456 26893 15484
rect 26844 15444 26850 15456
rect 26881 15453 26893 15456
rect 26927 15453 26939 15487
rect 26881 15447 26939 15453
rect 26973 15487 27031 15493
rect 26973 15453 26985 15487
rect 27019 15453 27031 15487
rect 26973 15447 27031 15453
rect 27065 15487 27123 15493
rect 27065 15453 27077 15487
rect 27111 15484 27123 15487
rect 27154 15484 27160 15496
rect 27111 15456 27160 15484
rect 27111 15453 27123 15456
rect 27065 15447 27123 15453
rect 24544 15388 26740 15416
rect 24544 15376 24550 15388
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 14366 15308 14372 15360
rect 14424 15348 14430 15360
rect 15470 15348 15476 15360
rect 14424 15320 15476 15348
rect 14424 15308 14430 15320
rect 15470 15308 15476 15320
rect 15528 15308 15534 15360
rect 15654 15308 15660 15360
rect 15712 15308 15718 15360
rect 15746 15308 15752 15360
rect 15804 15348 15810 15360
rect 16114 15348 16120 15360
rect 15804 15320 16120 15348
rect 15804 15308 15810 15320
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16206 15308 16212 15360
rect 16264 15348 16270 15360
rect 19702 15348 19708 15360
rect 16264 15320 19708 15348
rect 16264 15308 16270 15320
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 22373 15351 22431 15357
rect 22373 15348 22385 15351
rect 19852 15320 22385 15348
rect 19852 15308 19858 15320
rect 22373 15317 22385 15320
rect 22419 15348 22431 15351
rect 22922 15348 22928 15360
rect 22419 15320 22928 15348
rect 22419 15317 22431 15320
rect 22373 15311 22431 15317
rect 22922 15308 22928 15320
rect 22980 15348 22986 15360
rect 23290 15348 23296 15360
rect 22980 15320 23296 15348
rect 22980 15308 22986 15320
rect 23290 15308 23296 15320
rect 23348 15308 23354 15360
rect 25958 15308 25964 15360
rect 26016 15348 26022 15360
rect 26142 15348 26148 15360
rect 26016 15320 26148 15348
rect 26016 15308 26022 15320
rect 26142 15308 26148 15320
rect 26200 15308 26206 15360
rect 26602 15308 26608 15360
rect 26660 15348 26666 15360
rect 26988 15348 27016 15447
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27249 15487 27307 15493
rect 27249 15453 27261 15487
rect 27295 15484 27307 15487
rect 27430 15484 27436 15496
rect 27295 15456 27436 15484
rect 27295 15453 27307 15456
rect 27249 15447 27307 15453
rect 27430 15444 27436 15456
rect 27488 15444 27494 15496
rect 28552 15493 28580 15524
rect 28994 15512 29000 15524
rect 29052 15552 29058 15564
rect 29362 15552 29368 15564
rect 29052 15524 29368 15552
rect 29052 15512 29058 15524
rect 29362 15512 29368 15524
rect 29420 15512 29426 15564
rect 31018 15512 31024 15564
rect 31076 15552 31082 15564
rect 33778 15552 33784 15564
rect 31076 15524 33456 15552
rect 31076 15512 31082 15524
rect 28537 15487 28595 15493
rect 28537 15453 28549 15487
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 28626 15444 28632 15496
rect 28684 15444 28690 15496
rect 28810 15444 28816 15496
rect 28868 15484 28874 15496
rect 28905 15487 28963 15493
rect 28905 15484 28917 15487
rect 28868 15456 28917 15484
rect 28868 15444 28874 15456
rect 28905 15453 28917 15456
rect 28951 15484 28963 15487
rect 29730 15484 29736 15496
rect 28951 15456 29736 15484
rect 28951 15453 28963 15456
rect 28905 15447 28963 15453
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 30742 15444 30748 15496
rect 30800 15484 30806 15496
rect 31386 15484 31392 15496
rect 30800 15456 31392 15484
rect 30800 15444 30806 15456
rect 31386 15444 31392 15456
rect 31444 15444 31450 15496
rect 31478 15444 31484 15496
rect 31536 15444 31542 15496
rect 31570 15444 31576 15496
rect 31628 15444 31634 15496
rect 33042 15484 33048 15496
rect 32416 15456 33048 15484
rect 28718 15376 28724 15428
rect 28776 15376 28782 15428
rect 31757 15419 31815 15425
rect 31757 15385 31769 15419
rect 31803 15416 31815 15419
rect 32416 15416 32444 15456
rect 33042 15444 33048 15456
rect 33100 15444 33106 15496
rect 33226 15493 33232 15496
rect 33224 15484 33232 15493
rect 33187 15456 33232 15484
rect 33224 15447 33232 15456
rect 33226 15444 33232 15447
rect 33284 15444 33290 15496
rect 33428 15493 33456 15524
rect 33612 15524 33784 15552
rect 33612 15493 33640 15524
rect 33778 15512 33784 15524
rect 33836 15512 33842 15564
rect 33413 15487 33471 15493
rect 33413 15453 33425 15487
rect 33459 15453 33471 15487
rect 33413 15447 33471 15453
rect 33596 15487 33654 15493
rect 33596 15453 33608 15487
rect 33642 15453 33654 15487
rect 33596 15447 33654 15453
rect 33686 15444 33692 15496
rect 33744 15444 33750 15496
rect 31803 15388 32444 15416
rect 31803 15385 31815 15388
rect 31757 15379 31815 15385
rect 32858 15376 32864 15428
rect 32916 15416 32922 15428
rect 33321 15419 33379 15425
rect 33321 15416 33333 15419
rect 32916 15388 33333 15416
rect 32916 15376 32922 15388
rect 33321 15385 33333 15388
rect 33367 15385 33379 15419
rect 33321 15379 33379 15385
rect 27154 15348 27160 15360
rect 26660 15320 27160 15348
rect 26660 15308 26666 15320
rect 27154 15308 27160 15320
rect 27212 15308 27218 15360
rect 27706 15308 27712 15360
rect 27764 15348 27770 15360
rect 28258 15348 28264 15360
rect 27764 15320 28264 15348
rect 27764 15308 27770 15320
rect 28258 15308 28264 15320
rect 28316 15308 28322 15360
rect 28350 15308 28356 15360
rect 28408 15308 28414 15360
rect 31294 15308 31300 15360
rect 31352 15308 31358 15360
rect 33042 15308 33048 15360
rect 33100 15308 33106 15360
rect 1104 15258 36524 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 36524 15258
rect 1104 15184 36524 15206
rect 4614 15104 4620 15156
rect 4672 15144 4678 15156
rect 4709 15147 4767 15153
rect 4709 15144 4721 15147
rect 4672 15116 4721 15144
rect 4672 15104 4678 15116
rect 4709 15113 4721 15116
rect 4755 15144 4767 15147
rect 5258 15144 5264 15156
rect 4755 15116 5264 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 7190 15144 7196 15156
rect 6104 15116 7196 15144
rect 6104 15076 6132 15116
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 7377 15147 7435 15153
rect 7377 15113 7389 15147
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 7392 15076 7420 15107
rect 7466 15104 7472 15156
rect 7524 15144 7530 15156
rect 7742 15144 7748 15156
rect 7524 15116 7748 15144
rect 7524 15104 7530 15116
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 8754 15144 8760 15156
rect 8444 15116 8760 15144
rect 8444 15104 8450 15116
rect 8754 15104 8760 15116
rect 8812 15144 8818 15156
rect 10781 15147 10839 15153
rect 10781 15144 10793 15147
rect 8812 15116 10793 15144
rect 8812 15104 8818 15116
rect 10781 15113 10793 15116
rect 10827 15113 10839 15147
rect 10781 15107 10839 15113
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 12621 15147 12679 15153
rect 12621 15144 12633 15147
rect 12584 15116 12633 15144
rect 12584 15104 12590 15116
rect 12621 15113 12633 15116
rect 12667 15113 12679 15147
rect 12621 15107 12679 15113
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12768 15116 12817 15144
rect 12768 15104 12774 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 13541 15147 13599 15153
rect 13541 15113 13553 15147
rect 13587 15144 13599 15147
rect 13906 15144 13912 15156
rect 13587 15116 13912 15144
rect 13587 15113 13599 15116
rect 13541 15107 13599 15113
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 15654 15104 15660 15156
rect 15712 15144 15718 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15712 15116 15945 15144
rect 15712 15104 15718 15116
rect 15933 15113 15945 15116
rect 15979 15144 15991 15147
rect 16206 15144 16212 15156
rect 15979 15116 16212 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 16298 15104 16304 15156
rect 16356 15144 16362 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 16356 15116 17325 15144
rect 16356 15104 16362 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 18230 15144 18236 15156
rect 17911 15116 18236 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 19058 15153 19064 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18380 15116 18797 15144
rect 18380 15104 18386 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 18877 15147 18935 15153
rect 18877 15113 18889 15147
rect 18923 15113 18935 15147
rect 18877 15107 18935 15113
rect 19045 15147 19064 15153
rect 19045 15113 19057 15147
rect 19045 15107 19064 15113
rect 9674 15076 9680 15088
rect 4462 15062 6132 15076
rect 4448 15048 6132 15062
rect 6840 15048 7420 15076
rect 8956 15048 9680 15076
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 2961 15011 3019 15017
rect 2961 15008 2973 15011
rect 2648 14980 2973 15008
rect 2648 14968 2654 14980
rect 2961 14977 2973 14980
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 3234 14900 3240 14952
rect 3292 14900 3298 14952
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 4448 14940 4476 15048
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 5261 15011 5319 15017
rect 5261 14977 5273 15011
rect 5307 15008 5319 15011
rect 6730 15008 6736 15020
rect 5307 14980 6736 15008
rect 5307 14977 5319 14980
rect 5261 14971 5319 14977
rect 4028 14912 4476 14940
rect 5092 14940 5120 14971
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 6840 15017 6868 15048
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 7101 15011 7159 15017
rect 7101 14977 7113 15011
rect 7147 15008 7159 15011
rect 7190 15008 7196 15020
rect 7147 14980 7196 15008
rect 7147 14977 7159 14980
rect 7101 14971 7159 14977
rect 5534 14940 5540 14952
rect 5092 14912 5540 14940
rect 4028 14900 4034 14912
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 7024 14940 7052 14971
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 8956 15017 8984 15048
rect 9674 15036 9680 15048
rect 9732 15036 9738 15088
rect 10318 15036 10324 15088
rect 10376 15076 10382 15088
rect 10376 15048 11652 15076
rect 10376 15036 10382 15048
rect 8849 15011 8907 15017
rect 8849 15008 8861 15011
rect 8772 14980 8861 15008
rect 7024 14912 7144 14940
rect 7116 14872 7144 14912
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 8018 14900 8024 14952
rect 8076 14900 8082 14952
rect 7926 14872 7932 14884
rect 7116 14844 7932 14872
rect 7926 14832 7932 14844
rect 7984 14832 7990 14884
rect 8772 14872 8800 14980
rect 8849 14977 8861 14980
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 9490 14968 9496 15020
rect 9548 15008 9554 15020
rect 10339 15008 10367 15036
rect 11624 15020 11652 15048
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 14553 15079 14611 15085
rect 11756 15048 12388 15076
rect 11756 15036 11762 15048
rect 9548 14980 10367 15008
rect 9548 14968 9554 14980
rect 10410 14968 10416 15020
rect 10468 14968 10474 15020
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 10784 15011 10842 15017
rect 10784 15008 10796 15011
rect 10744 14980 10796 15008
rect 10744 14968 10750 14980
rect 10784 14977 10796 14980
rect 10830 14977 10842 15011
rect 10784 14971 10842 14977
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11664 14980 11805 15008
rect 11664 14968 11670 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 11974 14968 11980 15020
rect 12032 14968 12038 15020
rect 12360 15017 12388 15048
rect 14553 15045 14565 15079
rect 14599 15076 14611 15079
rect 14826 15076 14832 15088
rect 14599 15048 14832 15076
rect 14599 15045 14611 15048
rect 14553 15039 14611 15045
rect 14826 15036 14832 15048
rect 14884 15036 14890 15088
rect 15194 15036 15200 15088
rect 15252 15036 15258 15088
rect 16316 15076 16344 15104
rect 15764 15048 16344 15076
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 15008 12127 15011
rect 12345 15011 12403 15017
rect 12115 14980 12296 15008
rect 12115 14977 12127 14980
rect 12069 14971 12127 14977
rect 9582 14900 9588 14952
rect 9640 14940 9646 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 9640 14912 10333 14940
rect 9640 14900 9646 14912
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 11992 14940 12020 14968
rect 10321 14903 10379 14909
rect 10428 14912 12020 14940
rect 12161 14943 12219 14949
rect 10428 14872 10456 14912
rect 12161 14909 12173 14943
rect 12207 14909 12219 14943
rect 12268 14940 12296 14980
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 12746 15011 12804 15017
rect 12746 15008 12758 15011
rect 12575 14980 12758 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 12746 14977 12758 14980
rect 12792 14977 12804 15011
rect 12746 14971 12804 14977
rect 12986 14968 12992 15020
rect 13044 15008 13050 15020
rect 13265 15011 13323 15017
rect 13265 15008 13277 15011
rect 13044 14980 13277 15008
rect 13044 14968 13050 14980
rect 13265 14977 13277 14980
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14323 14980 14504 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 12894 14940 12900 14952
rect 12268 14912 12900 14940
rect 12161 14903 12219 14909
rect 8772 14844 10456 14872
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 5169 14807 5227 14813
rect 5169 14804 5181 14807
rect 4856 14776 5181 14804
rect 4856 14764 4862 14776
rect 5169 14773 5181 14776
rect 5215 14773 5227 14807
rect 5169 14767 5227 14773
rect 5258 14764 5264 14816
rect 5316 14804 5322 14816
rect 6641 14807 6699 14813
rect 6641 14804 6653 14807
rect 5316 14776 6653 14804
rect 5316 14764 5322 14776
rect 6641 14773 6653 14776
rect 6687 14773 6699 14807
rect 6641 14767 6699 14773
rect 8018 14764 8024 14816
rect 8076 14804 8082 14816
rect 8665 14807 8723 14813
rect 8665 14804 8677 14807
rect 8076 14776 8677 14804
rect 8076 14764 8082 14776
rect 8665 14773 8677 14776
rect 8711 14773 8723 14807
rect 8665 14767 8723 14773
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 8904 14776 9137 14804
rect 8904 14764 8910 14776
rect 9125 14773 9137 14776
rect 9171 14804 9183 14807
rect 9582 14804 9588 14816
rect 9171 14776 9588 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9582 14764 9588 14776
rect 9640 14804 9646 14816
rect 10226 14804 10232 14816
rect 9640 14776 10232 14804
rect 9640 14764 9646 14776
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 10836 14776 10977 14804
rect 10836 14764 10842 14776
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 10965 14767 11023 14773
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 12176 14804 12204 14903
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13357 14943 13415 14949
rect 13357 14909 13369 14943
rect 13403 14940 13415 14943
rect 13446 14940 13452 14952
rect 13403 14912 13452 14940
rect 13403 14909 13415 14912
rect 13357 14903 13415 14909
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14940 13783 14943
rect 13814 14940 13820 14952
rect 13771 14912 13820 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 14366 14900 14372 14952
rect 14424 14900 14430 14952
rect 14476 14940 14504 14980
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 14700 14980 14933 15008
rect 14700 14968 14706 14980
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15654 15008 15660 15020
rect 15059 14980 15660 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 15764 15017 15792 15048
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 18892 15076 18920 15107
rect 19058 15104 19064 15107
rect 19116 15104 19122 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 19337 15147 19395 15153
rect 19337 15144 19349 15147
rect 19208 15116 19349 15144
rect 19208 15104 19214 15116
rect 19337 15113 19349 15116
rect 19383 15113 19395 15147
rect 19337 15107 19395 15113
rect 20241 15147 20299 15153
rect 20241 15113 20253 15147
rect 20287 15144 20299 15147
rect 20898 15144 20904 15156
rect 20287 15116 20904 15144
rect 20287 15113 20299 15116
rect 20241 15107 20299 15113
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 21450 15104 21456 15156
rect 21508 15144 21514 15156
rect 22465 15147 22523 15153
rect 22465 15144 22477 15147
rect 21508 15116 22477 15144
rect 21508 15104 21514 15116
rect 22465 15113 22477 15116
rect 22511 15144 22523 15147
rect 22554 15144 22560 15156
rect 22511 15116 22560 15144
rect 22511 15113 22523 15116
rect 22465 15107 22523 15113
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 23014 15104 23020 15156
rect 23072 15144 23078 15156
rect 23566 15144 23572 15156
rect 23072 15116 23572 15144
rect 23072 15104 23078 15116
rect 23566 15104 23572 15116
rect 23624 15104 23630 15156
rect 24026 15144 24032 15156
rect 23860 15116 24032 15144
rect 19245 15079 19303 15085
rect 19245 15076 19257 15079
rect 16448 15048 19088 15076
rect 16448 15036 16454 15048
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 14977 15807 15011
rect 15749 14971 15807 14977
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16114 15008 16120 15020
rect 16071 14980 16120 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16114 14968 16120 14980
rect 16172 15008 16178 15020
rect 16758 15008 16764 15020
rect 16172 14980 16764 15008
rect 16172 14968 16178 14980
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 17497 15011 17555 15017
rect 17954 15011 17960 15020
rect 17497 14977 17509 15011
rect 17543 15008 17555 15011
rect 17788 15008 17960 15011
rect 17543 14983 17960 15008
rect 17543 14980 17816 14983
rect 17926 14980 17960 14983
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 15008 18199 15011
rect 18230 15008 18236 15020
rect 18187 14980 18236 15008
rect 18187 14977 18199 14980
rect 18141 14971 18199 14977
rect 15102 14940 15108 14952
rect 14476 14912 15108 14940
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 15289 14943 15347 14949
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 15562 14940 15568 14952
rect 15335 14912 15568 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 17773 14943 17831 14949
rect 17773 14940 17785 14943
rect 17644 14912 17785 14940
rect 17644 14900 17650 14912
rect 17773 14909 17785 14912
rect 17819 14909 17831 14943
rect 18064 14940 18092 14971
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 18325 15011 18383 15017
rect 18325 14977 18337 15011
rect 18371 14977 18383 15011
rect 18325 14971 18383 14977
rect 18340 14940 18368 14971
rect 18506 14968 18512 15020
rect 18564 14968 18570 15020
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 15008 18659 15011
rect 18782 15008 18788 15020
rect 18647 14980 18788 15008
rect 18647 14977 18659 14980
rect 18601 14971 18659 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19060 14940 19088 15048
rect 19168 15048 19257 15076
rect 19168 15020 19196 15048
rect 19245 15045 19257 15048
rect 19291 15076 19303 15079
rect 20441 15079 20499 15085
rect 19291 15048 20024 15076
rect 19291 15045 19303 15048
rect 19245 15039 19303 15045
rect 19150 14968 19156 15020
rect 19208 14968 19214 15020
rect 19518 14968 19524 15020
rect 19576 15009 19582 15020
rect 19613 15011 19671 15017
rect 19613 15009 19625 15011
rect 19576 14981 19625 15009
rect 19576 14968 19582 14981
rect 19613 14977 19625 14981
rect 19659 14977 19671 15011
rect 19613 14971 19671 14977
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 15008 19855 15011
rect 19886 15008 19892 15020
rect 19843 14980 19892 15008
rect 19843 14977 19855 14980
rect 19797 14971 19855 14977
rect 19334 14940 19340 14952
rect 18064 14912 18276 14940
rect 18340 14912 19012 14940
rect 19060 14912 19340 14940
rect 17773 14903 17831 14909
rect 12250 14832 12256 14884
rect 12308 14872 12314 14884
rect 13173 14875 13231 14881
rect 13173 14872 13185 14875
rect 12308 14844 13185 14872
rect 12308 14832 12314 14844
rect 13173 14841 13185 14844
rect 13219 14872 13231 14875
rect 13262 14872 13268 14884
rect 13219 14844 13268 14872
rect 13219 14841 13231 14844
rect 13173 14835 13231 14841
rect 13262 14832 13268 14844
rect 13320 14832 13326 14884
rect 14093 14875 14151 14881
rect 14093 14841 14105 14875
rect 14139 14872 14151 14875
rect 15378 14872 15384 14884
rect 14139 14844 15384 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 15838 14872 15844 14884
rect 15580 14844 15844 14872
rect 12124 14776 12204 14804
rect 13909 14807 13967 14813
rect 12124 14764 12130 14776
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 13998 14804 14004 14816
rect 13955 14776 14004 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14553 14807 14611 14813
rect 14553 14773 14565 14807
rect 14599 14804 14611 14807
rect 14642 14804 14648 14816
rect 14599 14776 14648 14804
rect 14599 14773 14611 14776
rect 14553 14767 14611 14773
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 14734 14764 14740 14816
rect 14792 14764 14798 14816
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 15580 14813 15608 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 17681 14875 17739 14881
rect 17681 14872 17693 14875
rect 17552 14844 17693 14872
rect 17552 14832 17558 14844
rect 17681 14841 17693 14844
rect 17727 14872 17739 14875
rect 18138 14872 18144 14884
rect 17727 14844 18144 14872
rect 17727 14841 17739 14844
rect 17681 14835 17739 14841
rect 18138 14832 18144 14844
rect 18196 14832 18202 14884
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 14884 14776 14933 14804
rect 14884 14764 14890 14776
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 14921 14767 14979 14773
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14773 15623 14807
rect 15565 14767 15623 14773
rect 15657 14807 15715 14813
rect 15657 14773 15669 14807
rect 15703 14804 15715 14807
rect 16574 14804 16580 14816
rect 15703 14776 16580 14804
rect 15703 14773 15715 14776
rect 15657 14767 15715 14773
rect 16574 14764 16580 14776
rect 16632 14764 16638 14816
rect 17770 14764 17776 14816
rect 17828 14804 17834 14816
rect 18049 14807 18107 14813
rect 18049 14804 18061 14807
rect 17828 14776 18061 14804
rect 17828 14764 17834 14776
rect 18049 14773 18061 14776
rect 18095 14773 18107 14807
rect 18248 14804 18276 14912
rect 18984 14872 19012 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19720 14940 19748 14971
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 19996 15017 20024 15048
rect 20441 15045 20453 15079
rect 20487 15076 20499 15079
rect 20714 15076 20720 15088
rect 20487 15048 20720 15076
rect 20487 15045 20499 15048
rect 20441 15039 20499 15045
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 22649 15079 22707 15085
rect 22649 15076 22661 15079
rect 22112 15048 22661 15076
rect 22112 15020 22140 15048
rect 22649 15045 22661 15048
rect 22695 15045 22707 15079
rect 22649 15039 22707 15045
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 15008 20039 15011
rect 20162 15008 20168 15020
rect 20027 14980 20168 15008
rect 20027 14977 20039 14980
rect 19981 14971 20039 14977
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 21450 15008 21456 15020
rect 21048 14980 21456 15008
rect 21048 14968 21054 14980
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 22094 14968 22100 15020
rect 22152 14968 22158 15020
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22278 15008 22284 15020
rect 22235 14980 22284 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22554 14968 22560 15020
rect 22612 14968 22618 15020
rect 22833 15011 22891 15017
rect 22833 14977 22845 15011
rect 22879 15008 22891 15011
rect 22922 15008 22928 15020
rect 22879 14980 22928 15008
rect 22879 14977 22891 14980
rect 22833 14971 22891 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 23032 15017 23060 15104
rect 23198 15036 23204 15088
rect 23256 15076 23262 15088
rect 23860 15085 23888 15116
rect 24026 15104 24032 15116
rect 24084 15104 24090 15156
rect 26326 15104 26332 15156
rect 26384 15104 26390 15156
rect 26970 15144 26976 15156
rect 26528 15116 26976 15144
rect 23753 15079 23811 15085
rect 23753 15076 23765 15079
rect 23256 15048 23765 15076
rect 23256 15036 23262 15048
rect 23753 15045 23765 15048
rect 23799 15045 23811 15079
rect 23753 15039 23811 15045
rect 23845 15079 23903 15085
rect 23845 15045 23857 15079
rect 23891 15045 23903 15079
rect 24210 15076 24216 15088
rect 23845 15039 23903 15045
rect 23952 15048 24216 15076
rect 23017 15011 23075 15017
rect 23017 14977 23029 15011
rect 23063 14977 23075 15011
rect 23017 14971 23075 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23293 15011 23351 15017
rect 23293 14977 23305 15011
rect 23339 15008 23351 15011
rect 23382 15008 23388 15020
rect 23339 14980 23388 15008
rect 23339 14977 23351 14980
rect 23293 14971 23351 14977
rect 20254 14940 20260 14952
rect 19720 14912 20260 14940
rect 20254 14900 20260 14912
rect 20312 14940 20318 14952
rect 21177 14943 21235 14949
rect 20312 14912 21128 14940
rect 20312 14900 20318 14912
rect 19242 14872 19248 14884
rect 18984 14844 19248 14872
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 20070 14832 20076 14884
rect 20128 14832 20134 14884
rect 21100 14872 21128 14912
rect 21177 14909 21189 14943
rect 21223 14940 21235 14943
rect 21634 14940 21640 14952
rect 21223 14912 21640 14940
rect 21223 14909 21235 14912
rect 21177 14903 21235 14909
rect 21634 14900 21640 14912
rect 21692 14900 21698 14952
rect 21928 14912 22968 14940
rect 21928 14872 21956 14912
rect 21100 14844 21956 14872
rect 22002 14832 22008 14884
rect 22060 14872 22066 14884
rect 22940 14881 22968 14912
rect 22925 14875 22983 14881
rect 22060 14844 22501 14872
rect 22060 14832 22066 14844
rect 18966 14804 18972 14816
rect 18248 14776 18972 14804
rect 18049 14767 18107 14773
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19061 14807 19119 14813
rect 19061 14773 19073 14807
rect 19107 14804 19119 14807
rect 19978 14804 19984 14816
rect 19107 14776 19984 14804
rect 19107 14773 19119 14776
rect 19061 14767 19119 14773
rect 19978 14764 19984 14776
rect 20036 14764 20042 14816
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 20257 14807 20315 14813
rect 20257 14804 20269 14807
rect 20220 14776 20269 14804
rect 20220 14764 20226 14776
rect 20257 14773 20269 14776
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 21174 14764 21180 14816
rect 21232 14804 21238 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 21232 14776 21281 14804
rect 21232 14764 21238 14776
rect 21269 14773 21281 14776
rect 21315 14773 21327 14807
rect 21269 14767 21327 14773
rect 21450 14764 21456 14816
rect 21508 14804 21514 14816
rect 21637 14807 21695 14813
rect 21637 14804 21649 14807
rect 21508 14776 21649 14804
rect 21508 14764 21514 14776
rect 21637 14773 21649 14776
rect 21683 14773 21695 14807
rect 21637 14767 21695 14773
rect 21818 14764 21824 14816
rect 21876 14764 21882 14816
rect 22281 14807 22339 14813
rect 22281 14773 22293 14807
rect 22327 14804 22339 14807
rect 22370 14804 22376 14816
rect 22327 14776 22376 14804
rect 22327 14773 22339 14776
rect 22281 14767 22339 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 22473 14804 22501 14844
rect 22925 14841 22937 14875
rect 22971 14841 22983 14875
rect 23124 14872 23152 14971
rect 23382 14968 23388 14980
rect 23440 14968 23446 15020
rect 23952 15017 23980 15048
rect 24210 15036 24216 15048
rect 24268 15036 24274 15088
rect 23635 15011 23693 15017
rect 23635 14977 23647 15011
rect 23681 14977 23693 15011
rect 23635 14971 23693 14977
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 24121 15011 24179 15017
rect 24121 14977 24133 15011
rect 24167 15008 24179 15011
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24167 14980 24501 15008
rect 24167 14977 24179 14980
rect 24121 14971 24179 14977
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 23474 14900 23480 14952
rect 23532 14900 23538 14952
rect 23650 14940 23678 14971
rect 24762 14968 24768 15020
rect 24820 15008 24826 15020
rect 25314 15008 25320 15020
rect 24820 14980 25320 15008
rect 24820 14968 24826 14980
rect 25314 14968 25320 14980
rect 25372 14968 25378 15020
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 26528 15008 26556 15116
rect 26970 15104 26976 15116
rect 27028 15144 27034 15156
rect 27430 15144 27436 15156
rect 27028 15116 27436 15144
rect 27028 15104 27034 15116
rect 27430 15104 27436 15116
rect 27488 15104 27494 15156
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 27709 15147 27767 15153
rect 27709 15144 27721 15147
rect 27672 15116 27721 15144
rect 27672 15104 27678 15116
rect 27709 15113 27721 15116
rect 27755 15144 27767 15147
rect 28902 15144 28908 15156
rect 27755 15116 28908 15144
rect 27755 15113 27767 15116
rect 27709 15107 27767 15113
rect 28902 15104 28908 15116
rect 28960 15104 28966 15156
rect 29181 15147 29239 15153
rect 29181 15113 29193 15147
rect 29227 15144 29239 15147
rect 29227 15116 30052 15144
rect 29227 15113 29239 15116
rect 29181 15107 29239 15113
rect 27356 15048 27752 15076
rect 27356 15020 27384 15048
rect 26467 14980 26556 15008
rect 26605 15011 26663 15017
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 26605 14977 26617 15011
rect 26651 14977 26663 15011
rect 27065 15011 27123 15017
rect 27065 15008 27077 15011
rect 26605 14971 26663 14977
rect 26712 14980 27077 15008
rect 23650 14912 23980 14940
rect 23952 14872 23980 14912
rect 24394 14900 24400 14952
rect 24452 14900 24458 14952
rect 24857 14943 24915 14949
rect 24857 14909 24869 14943
rect 24903 14940 24915 14943
rect 25038 14940 25044 14952
rect 24903 14912 25044 14940
rect 24903 14909 24915 14912
rect 24857 14903 24915 14909
rect 25038 14900 25044 14912
rect 25096 14900 25102 14952
rect 25682 14900 25688 14952
rect 25740 14940 25746 14952
rect 26620 14940 26648 14971
rect 25740 14912 26648 14940
rect 25740 14900 25746 14912
rect 25222 14872 25228 14884
rect 23124 14844 23612 14872
rect 23952 14844 25228 14872
rect 22925 14835 22983 14841
rect 23014 14804 23020 14816
rect 22473 14776 23020 14804
rect 23014 14764 23020 14776
rect 23072 14804 23078 14816
rect 23474 14804 23480 14816
rect 23072 14776 23480 14804
rect 23072 14764 23078 14776
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 23584 14804 23612 14844
rect 25222 14832 25228 14844
rect 25280 14832 25286 14884
rect 25866 14832 25872 14884
rect 25924 14872 25930 14884
rect 26712 14872 26740 14980
rect 27065 14977 27077 14980
rect 27111 14977 27123 15011
rect 27065 14971 27123 14977
rect 27338 14968 27344 15020
rect 27396 14968 27402 15020
rect 27522 14968 27528 15020
rect 27580 15008 27586 15020
rect 27724 15017 27752 15048
rect 27798 15036 27804 15088
rect 27856 15076 27862 15088
rect 27856 15048 28672 15076
rect 27856 15036 27862 15048
rect 27617 15011 27675 15017
rect 27617 15008 27629 15011
rect 27580 14980 27629 15008
rect 27580 14968 27586 14980
rect 27617 14977 27629 14980
rect 27663 14977 27675 15011
rect 27617 14971 27675 14977
rect 27709 15011 27767 15017
rect 27709 14977 27721 15011
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 28350 14968 28356 15020
rect 28408 15008 28414 15020
rect 28644 15017 28672 15048
rect 28810 15036 28816 15088
rect 28868 15036 28874 15088
rect 29270 15036 29276 15088
rect 29328 15036 29334 15088
rect 29638 15076 29644 15088
rect 29380 15048 29644 15076
rect 28537 15011 28595 15017
rect 28537 15008 28549 15011
rect 28408 14980 28549 15008
rect 28408 14968 28414 14980
rect 28537 14977 28549 14980
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 28630 15011 28688 15017
rect 28630 14977 28642 15011
rect 28676 14977 28688 15011
rect 28630 14971 28688 14977
rect 28552 14940 28580 14971
rect 28902 14968 28908 15020
rect 28960 14968 28966 15020
rect 28994 14968 29000 15020
rect 29052 15017 29058 15020
rect 29052 15008 29060 15017
rect 29052 14980 29097 15008
rect 29052 14971 29060 14980
rect 29052 14968 29058 14971
rect 28810 14940 28816 14952
rect 28552 14912 28816 14940
rect 28810 14900 28816 14912
rect 28868 14900 28874 14952
rect 29270 14900 29276 14952
rect 29328 14940 29334 14952
rect 29380 14940 29408 15048
rect 29638 15036 29644 15048
rect 29696 15036 29702 15088
rect 29549 15011 29607 15017
rect 29549 14977 29561 15011
rect 29595 15008 29607 15011
rect 29595 14980 29684 15008
rect 29595 14977 29607 14980
rect 29549 14971 29607 14977
rect 29656 14952 29684 14980
rect 29822 14968 29828 15020
rect 29880 14968 29886 15020
rect 30024 15017 30052 15116
rect 30742 15104 30748 15156
rect 30800 15144 30806 15156
rect 32950 15144 32956 15156
rect 30800 15116 32956 15144
rect 30800 15104 30806 15116
rect 32950 15104 32956 15116
rect 33008 15104 33014 15156
rect 33410 15104 33416 15156
rect 33468 15144 33474 15156
rect 33468 15116 35204 15144
rect 33468 15104 33474 15116
rect 31205 15079 31263 15085
rect 31205 15045 31217 15079
rect 31251 15076 31263 15079
rect 31754 15076 31760 15088
rect 31251 15048 31760 15076
rect 31251 15045 31263 15048
rect 31205 15039 31263 15045
rect 31754 15036 31760 15048
rect 31812 15036 31818 15088
rect 33226 15076 33232 15088
rect 32416 15048 33232 15076
rect 32416 15017 32444 15048
rect 33226 15036 33232 15048
rect 33284 15036 33290 15088
rect 35176 15085 35204 15116
rect 35161 15079 35219 15085
rect 35161 15045 35173 15079
rect 35207 15045 35219 15079
rect 35161 15039 35219 15045
rect 30009 15011 30067 15017
rect 30009 14977 30021 15011
rect 30055 14977 30067 15011
rect 31665 15011 31723 15017
rect 31665 15008 31677 15011
rect 30009 14971 30067 14977
rect 31036 14980 31677 15008
rect 29328 14912 29408 14940
rect 29328 14900 29334 14912
rect 29454 14900 29460 14952
rect 29512 14900 29518 14952
rect 29638 14900 29644 14952
rect 29696 14900 29702 14952
rect 30282 14900 30288 14952
rect 30340 14940 30346 14952
rect 31036 14949 31064 14980
rect 31665 14977 31677 14980
rect 31711 15008 31723 15011
rect 32401 15011 32459 15017
rect 31711 14980 32352 15008
rect 31711 14977 31723 14980
rect 31665 14971 31723 14977
rect 31021 14943 31079 14949
rect 31021 14940 31033 14943
rect 30340 14912 31033 14940
rect 30340 14900 30346 14912
rect 31021 14909 31033 14912
rect 31067 14909 31079 14943
rect 32214 14940 32220 14952
rect 31021 14903 31079 14909
rect 31726 14912 32220 14940
rect 25924 14844 26740 14872
rect 27065 14875 27123 14881
rect 25924 14832 25930 14844
rect 27065 14841 27077 14875
rect 27111 14841 27123 14875
rect 27065 14835 27123 14841
rect 29733 14875 29791 14881
rect 29733 14841 29745 14875
rect 29779 14872 29791 14875
rect 31726 14872 31754 14912
rect 32214 14900 32220 14912
rect 32272 14900 32278 14952
rect 32324 14940 32352 14980
rect 32401 14977 32413 15011
rect 32447 14977 32459 15011
rect 32401 14971 32459 14977
rect 32490 14968 32496 15020
rect 32548 14968 32554 15020
rect 32582 14968 32588 15020
rect 32640 14968 32646 15020
rect 32769 15011 32827 15017
rect 32769 14977 32781 15011
rect 32815 15008 32827 15011
rect 33778 15008 33784 15020
rect 32815 14980 33784 15008
rect 32815 14977 32827 14980
rect 32769 14971 32827 14977
rect 33778 14968 33784 14980
rect 33836 14968 33842 15020
rect 34931 15011 34989 15017
rect 34931 15008 34943 15011
rect 33888 14980 34943 15008
rect 32324 14912 32536 14940
rect 29779 14844 31754 14872
rect 29779 14841 29791 14844
rect 29733 14835 29791 14841
rect 24026 14804 24032 14816
rect 23584 14776 24032 14804
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 24210 14764 24216 14816
rect 24268 14764 24274 14816
rect 24762 14764 24768 14816
rect 24820 14804 24826 14816
rect 26786 14804 26792 14816
rect 24820 14776 26792 14804
rect 24820 14764 24826 14776
rect 26786 14764 26792 14776
rect 26844 14804 26850 14816
rect 27080 14804 27108 14835
rect 28534 14804 28540 14816
rect 26844 14776 28540 14804
rect 26844 14764 26850 14776
rect 28534 14764 28540 14776
rect 28592 14764 28598 14816
rect 28810 14764 28816 14816
rect 28868 14804 28874 14816
rect 29273 14807 29331 14813
rect 29273 14804 29285 14807
rect 28868 14776 29285 14804
rect 28868 14764 28874 14776
rect 29273 14773 29285 14776
rect 29319 14773 29331 14807
rect 29273 14767 29331 14773
rect 30009 14807 30067 14813
rect 30009 14773 30021 14807
rect 30055 14804 30067 14807
rect 30650 14804 30656 14816
rect 30055 14776 30656 14804
rect 30055 14773 30067 14776
rect 30009 14767 30067 14773
rect 30650 14764 30656 14776
rect 30708 14764 30714 14816
rect 31478 14764 31484 14816
rect 31536 14764 31542 14816
rect 31570 14764 31576 14816
rect 31628 14804 31634 14816
rect 31938 14804 31944 14816
rect 31628 14776 31944 14804
rect 31628 14764 31634 14776
rect 31938 14764 31944 14776
rect 31996 14764 32002 14816
rect 32217 14807 32275 14813
rect 32217 14773 32229 14807
rect 32263 14804 32275 14807
rect 32398 14804 32404 14816
rect 32263 14776 32404 14804
rect 32263 14773 32275 14776
rect 32217 14767 32275 14773
rect 32398 14764 32404 14776
rect 32456 14764 32462 14816
rect 32508 14804 32536 14912
rect 33502 14804 33508 14816
rect 32508 14776 33508 14804
rect 33502 14764 33508 14776
rect 33560 14804 33566 14816
rect 33888 14804 33916 14980
rect 34931 14977 34943 14980
rect 34977 14977 34989 15011
rect 34931 14971 34989 14977
rect 35066 14968 35072 15020
rect 35124 14968 35130 15020
rect 35289 15011 35347 15017
rect 35289 15008 35301 15011
rect 35176 14980 35301 15008
rect 34790 14900 34796 14952
rect 34848 14940 34854 14952
rect 35176 14940 35204 14980
rect 35289 14977 35301 14980
rect 35335 14977 35347 15011
rect 35289 14971 35347 14977
rect 35437 15011 35495 15017
rect 35437 14977 35449 15011
rect 35483 15008 35495 15011
rect 36170 15008 36176 15020
rect 35483 14980 36176 15008
rect 35483 14977 35495 14980
rect 35437 14971 35495 14977
rect 36170 14968 36176 14980
rect 36228 14968 36234 15020
rect 34848 14912 35204 14940
rect 34848 14900 34854 14912
rect 33560 14776 33916 14804
rect 33560 14764 33566 14776
rect 34790 14764 34796 14816
rect 34848 14764 34854 14816
rect 1104 14714 36524 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 36524 14714
rect 1104 14640 36524 14662
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3292 14572 4169 14600
rect 3292 14560 3298 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 4157 14563 4215 14569
rect 7098 14560 7104 14612
rect 7156 14560 7162 14612
rect 7834 14560 7840 14612
rect 7892 14560 7898 14612
rect 10321 14603 10379 14609
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 11054 14600 11060 14612
rect 10367 14572 11060 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12492 14572 12725 14600
rect 12492 14560 12498 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 12894 14560 12900 14612
rect 12952 14560 12958 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 14826 14600 14832 14612
rect 13504 14572 14832 14600
rect 13504 14560 13510 14572
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 16206 14600 16212 14612
rect 15528 14572 16212 14600
rect 15528 14560 15534 14572
rect 16206 14560 16212 14572
rect 16264 14600 16270 14612
rect 16301 14603 16359 14609
rect 16301 14600 16313 14603
rect 16264 14572 16313 14600
rect 16264 14560 16270 14572
rect 16301 14569 16313 14572
rect 16347 14569 16359 14603
rect 18322 14600 18328 14612
rect 16301 14563 16359 14569
rect 17696 14572 17954 14600
rect 5534 14532 5540 14544
rect 5000 14504 5540 14532
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4614 14396 4620 14408
rect 4387 14368 4620 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4709 14399 4767 14405
rect 4709 14365 4721 14399
rect 4755 14396 4767 14399
rect 4798 14396 4804 14408
rect 4755 14368 4804 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 5000 14405 5028 14504
rect 5534 14492 5540 14504
rect 5592 14532 5598 14544
rect 5592 14504 6592 14532
rect 5592 14492 5598 14504
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14464 5135 14467
rect 5350 14464 5356 14476
rect 5123 14436 5356 14464
rect 5123 14433 5135 14436
rect 5077 14427 5135 14433
rect 5350 14424 5356 14436
rect 5408 14424 5414 14476
rect 5718 14424 5724 14476
rect 5776 14424 5782 14476
rect 6564 14473 6592 14504
rect 9306 14492 9312 14544
rect 9364 14532 9370 14544
rect 9364 14504 12434 14532
rect 9364 14492 9370 14504
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 6822 14464 6828 14476
rect 6595 14436 6828 14464
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 7650 14424 7656 14476
rect 7708 14424 7714 14476
rect 8478 14464 8484 14476
rect 8036 14436 8484 14464
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 4430 14288 4436 14340
rect 4488 14288 4494 14340
rect 4522 14288 4528 14340
rect 4580 14288 4586 14340
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 4801 14263 4859 14269
rect 4801 14260 4813 14263
rect 4672 14232 4813 14260
rect 4672 14220 4678 14232
rect 4801 14229 4813 14232
rect 4847 14229 4859 14263
rect 5184 14260 5212 14359
rect 5258 14356 5264 14408
rect 5316 14356 5322 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5592 14368 5641 14396
rect 5592 14356 5598 14368
rect 5629 14365 5641 14368
rect 5675 14396 5687 14399
rect 6362 14396 6368 14408
rect 5675 14368 6368 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 8036 14405 8064 14436
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 8846 14464 8852 14476
rect 8711 14436 8852 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 8846 14424 8852 14436
rect 8904 14464 8910 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 8904 14436 9505 14464
rect 8904 14424 8910 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 10502 14464 10508 14476
rect 9493 14427 9551 14433
rect 10244 14436 10508 14464
rect 7561 14399 7619 14405
rect 7561 14365 7573 14399
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8021 14399 8079 14405
rect 8021 14365 8033 14399
rect 8067 14365 8079 14399
rect 8021 14359 8079 14365
rect 6733 14331 6791 14337
rect 6733 14328 6745 14331
rect 6012 14300 6745 14328
rect 5258 14260 5264 14272
rect 5184 14232 5264 14260
rect 4801 14223 4859 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 6012 14269 6040 14300
rect 6733 14297 6745 14300
rect 6779 14297 6791 14331
rect 6733 14291 6791 14297
rect 7466 14288 7472 14340
rect 7524 14328 7530 14340
rect 7576 14328 7604 14359
rect 8202 14356 8208 14408
rect 8260 14356 8266 14408
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8386 14396 8392 14408
rect 8343 14368 8392 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 9674 14396 9680 14408
rect 8803 14368 9680 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 7524 14300 7604 14328
rect 7524 14288 7530 14300
rect 8478 14288 8484 14340
rect 8536 14328 8542 14340
rect 8588 14328 8616 14359
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 9766 14356 9772 14408
rect 9824 14356 9830 14408
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10244 14405 10272 14436
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11388 14436 12081 14464
rect 11388 14424 11394 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12406 14464 12434 14504
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 13357 14535 13415 14541
rect 13357 14532 13369 14535
rect 12676 14504 13369 14532
rect 12676 14492 12682 14504
rect 13357 14501 13369 14504
rect 13403 14501 13415 14535
rect 13357 14495 13415 14501
rect 13464 14464 13492 14560
rect 17696 14544 17724 14572
rect 13725 14535 13783 14541
rect 13725 14501 13737 14535
rect 13771 14532 13783 14535
rect 14090 14532 14096 14544
rect 13771 14504 14096 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 14090 14492 14096 14504
rect 14148 14532 14154 14544
rect 14734 14532 14740 14544
rect 14148 14504 14740 14532
rect 14148 14492 14154 14504
rect 14734 14492 14740 14504
rect 14792 14492 14798 14544
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 16117 14535 16175 14541
rect 16117 14532 16129 14535
rect 15988 14504 16129 14532
rect 15988 14492 15994 14504
rect 16117 14501 16129 14504
rect 16163 14501 16175 14535
rect 16117 14495 16175 14501
rect 17129 14535 17187 14541
rect 17129 14501 17141 14535
rect 17175 14532 17187 14535
rect 17586 14532 17592 14544
rect 17175 14504 17592 14532
rect 17175 14501 17187 14504
rect 17129 14495 17187 14501
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 17678 14492 17684 14544
rect 17736 14492 17742 14544
rect 17926 14532 17954 14572
rect 18064 14572 18328 14600
rect 18064 14532 18092 14572
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 19058 14560 19064 14612
rect 19116 14600 19122 14612
rect 19521 14603 19579 14609
rect 19521 14600 19533 14603
rect 19116 14572 19533 14600
rect 19116 14560 19122 14572
rect 19521 14569 19533 14572
rect 19567 14569 19579 14603
rect 19521 14563 19579 14569
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 21358 14560 21364 14612
rect 21416 14560 21422 14612
rect 21450 14560 21456 14612
rect 21508 14560 21514 14612
rect 21545 14603 21603 14609
rect 21545 14569 21557 14603
rect 21591 14600 21603 14603
rect 21818 14600 21824 14612
rect 21591 14572 21824 14600
rect 21591 14569 21603 14572
rect 21545 14563 21603 14569
rect 21818 14560 21824 14572
rect 21876 14560 21882 14612
rect 22186 14560 22192 14612
rect 22244 14600 22250 14612
rect 22465 14603 22523 14609
rect 22465 14600 22477 14603
rect 22244 14572 22477 14600
rect 22244 14560 22250 14572
rect 22465 14569 22477 14572
rect 22511 14569 22523 14603
rect 22465 14563 22523 14569
rect 23658 14560 23664 14612
rect 23716 14600 23722 14612
rect 23842 14600 23848 14612
rect 23716 14572 23848 14600
rect 23716 14560 23722 14572
rect 23842 14560 23848 14572
rect 23900 14600 23906 14612
rect 24394 14600 24400 14612
rect 23900 14572 24400 14600
rect 23900 14560 23906 14572
rect 24394 14560 24400 14572
rect 24452 14560 24458 14612
rect 27614 14600 27620 14612
rect 27264 14572 27620 14600
rect 17926 14504 18092 14532
rect 18414 14492 18420 14544
rect 18472 14532 18478 14544
rect 18509 14535 18567 14541
rect 18509 14532 18521 14535
rect 18472 14504 18521 14532
rect 18472 14492 18478 14504
rect 18509 14501 18521 14504
rect 18555 14501 18567 14535
rect 19242 14532 19248 14544
rect 18509 14495 18567 14501
rect 19060 14504 19248 14532
rect 14458 14464 14464 14476
rect 12406 14436 13492 14464
rect 13556 14436 14464 14464
rect 12069 14427 12127 14433
rect 10876 14408 10928 14414
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 10008 14368 10241 14396
rect 10008 14356 10014 14368
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14396 11943 14399
rect 11931 14368 12296 14396
rect 11931 14365 11943 14368
rect 11885 14359 11943 14365
rect 10876 14350 10928 14356
rect 9398 14328 9404 14340
rect 8536 14300 9404 14328
rect 8536 14288 8542 14300
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 10781 14331 10839 14337
rect 10781 14297 10793 14331
rect 10827 14297 10839 14331
rect 12268 14328 12296 14368
rect 12434 14356 12440 14408
rect 12492 14356 12498 14408
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 12894 14396 12900 14408
rect 12584 14368 12900 14396
rect 12584 14356 12590 14368
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 13556 14405 13584 14436
rect 14458 14424 14464 14436
rect 14516 14464 14522 14476
rect 15948 14464 15976 14492
rect 14516 14436 15976 14464
rect 14516 14424 14522 14436
rect 17034 14424 17040 14476
rect 17092 14464 17098 14476
rect 17221 14467 17279 14473
rect 17221 14464 17233 14467
rect 17092 14436 17233 14464
rect 17092 14424 17098 14436
rect 17221 14433 17233 14436
rect 17267 14433 17279 14467
rect 19060 14464 19088 14504
rect 19242 14492 19248 14504
rect 19300 14532 19306 14544
rect 19889 14535 19947 14541
rect 19889 14532 19901 14535
rect 19300 14504 19901 14532
rect 19300 14492 19306 14504
rect 19889 14501 19901 14504
rect 19935 14501 19947 14535
rect 19889 14495 19947 14501
rect 20180 14504 20448 14532
rect 17221 14427 17279 14433
rect 17420 14436 18092 14464
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14365 13599 14399
rect 13541 14359 13599 14365
rect 12618 14328 12624 14340
rect 12268 14300 12624 14328
rect 10781 14291 10839 14297
rect 5997 14263 6055 14269
rect 5997 14229 6009 14263
rect 6043 14229 6055 14263
rect 5997 14223 6055 14229
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 8202 14260 8208 14272
rect 6687 14232 8208 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8386 14220 8392 14272
rect 8444 14260 8450 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8444 14232 8953 14260
rect 8444 14220 8450 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 10796 14260 10824 14291
rect 12618 14288 12624 14300
rect 12676 14328 12682 14340
rect 13004 14328 13032 14356
rect 12676 14300 13032 14328
rect 12676 14288 12682 14300
rect 11238 14260 11244 14272
rect 10796 14232 11244 14260
rect 8941 14223 8999 14229
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 11882 14260 11888 14272
rect 11664 14232 11888 14260
rect 11664 14220 11670 14232
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 12434 14220 12440 14272
rect 12492 14260 12498 14272
rect 12802 14260 12808 14272
rect 12492 14232 12808 14260
rect 12492 14220 12498 14232
rect 12802 14220 12808 14232
rect 12860 14260 12866 14272
rect 13096 14260 13124 14359
rect 13630 14356 13636 14408
rect 13688 14356 13694 14408
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 13872 14368 14657 14396
rect 13872 14356 13878 14368
rect 14645 14365 14657 14368
rect 14691 14396 14703 14399
rect 15010 14396 15016 14408
rect 14691 14368 15016 14396
rect 14691 14365 14703 14368
rect 14645 14359 14703 14365
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15194 14356 15200 14408
rect 15252 14356 15258 14408
rect 15565 14399 15623 14405
rect 15565 14365 15577 14399
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 14734 14288 14740 14340
rect 14792 14288 14798 14340
rect 15580 14328 15608 14359
rect 15654 14356 15660 14408
rect 15712 14356 15718 14408
rect 16298 14356 16304 14408
rect 16356 14356 16362 14408
rect 16390 14356 16396 14408
rect 16448 14396 16454 14408
rect 16761 14399 16819 14405
rect 16761 14396 16773 14399
rect 16448 14368 16773 14396
rect 16448 14356 16454 14368
rect 16761 14365 16773 14368
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14396 17003 14399
rect 17420 14396 17448 14436
rect 16991 14368 17448 14396
rect 17497 14399 17555 14405
rect 16991 14365 17003 14368
rect 16945 14359 17003 14365
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 15930 14328 15936 14340
rect 15580 14300 15936 14328
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 16574 14288 16580 14340
rect 16632 14288 16638 14340
rect 17512 14328 17540 14359
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18064 14405 18092 14436
rect 18616 14436 19088 14464
rect 19797 14467 19855 14473
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17644 14368 17785 14396
rect 17644 14356 17650 14368
rect 17773 14365 17785 14368
rect 17819 14365 17831 14399
rect 18049 14399 18107 14405
rect 17773 14359 17831 14365
rect 17960 14377 18018 14383
rect 17960 14343 17972 14377
rect 18006 14343 18018 14377
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 17960 14340 18018 14343
rect 17862 14328 17868 14340
rect 17512 14300 17868 14328
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 17954 14288 17960 14340
rect 18012 14288 18018 14340
rect 12860 14232 13124 14260
rect 12860 14220 12866 14232
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 15010 14260 15016 14272
rect 13504 14232 15016 14260
rect 13504 14220 13510 14232
rect 15010 14220 15016 14232
rect 15068 14260 15074 14272
rect 16114 14260 16120 14272
rect 15068 14232 16120 14260
rect 15068 14220 15074 14232
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 17276 14232 17325 14260
rect 17276 14220 17282 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 18064 14260 18092 14359
rect 18138 14356 18144 14408
rect 18196 14405 18202 14408
rect 18196 14399 18245 14405
rect 18196 14365 18199 14399
rect 18233 14365 18245 14399
rect 18196 14359 18245 14365
rect 18196 14356 18202 14359
rect 18322 14356 18328 14408
rect 18380 14356 18386 14408
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14396 18475 14399
rect 18616 14396 18644 14436
rect 19797 14433 19809 14467
rect 19843 14464 19855 14467
rect 20180 14464 20208 14504
rect 19843 14436 20208 14464
rect 19843 14433 19855 14436
rect 19797 14427 19855 14433
rect 20420 14408 20448 14504
rect 20530 14424 20536 14476
rect 20588 14464 20594 14476
rect 21358 14464 21364 14476
rect 20588 14436 21364 14464
rect 20588 14424 20594 14436
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 23106 14464 23112 14476
rect 22787 14436 23112 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 23106 14424 23112 14436
rect 23164 14424 23170 14476
rect 26050 14424 26056 14476
rect 26108 14464 26114 14476
rect 26881 14467 26939 14473
rect 26108 14436 26832 14464
rect 26108 14424 26114 14436
rect 18463 14368 18644 14396
rect 18693 14399 18751 14405
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 18782 14396 18788 14408
rect 18739 14368 18788 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 18966 14356 18972 14408
rect 19024 14396 19030 14408
rect 19024 14368 20116 14396
rect 19024 14356 19030 14368
rect 18340 14328 18368 14356
rect 19794 14328 19800 14340
rect 18340 14300 19800 14328
rect 19794 14288 19800 14300
rect 19852 14288 19858 14340
rect 20088 14328 20116 14368
rect 20254 14356 20260 14408
rect 20312 14356 20318 14408
rect 20420 14368 20444 14408
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20956 14368 21097 14396
rect 20956 14356 20962 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22002 14396 22008 14408
rect 21867 14368 22008 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 22189 14399 22247 14405
rect 22189 14365 22201 14399
rect 22235 14396 22247 14399
rect 22278 14396 22284 14408
rect 22235 14368 22284 14396
rect 22235 14365 22247 14368
rect 22189 14359 22247 14365
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 22462 14356 22468 14408
rect 22520 14396 22526 14408
rect 22649 14399 22707 14405
rect 22649 14396 22661 14399
rect 22520 14368 22661 14396
rect 22520 14356 22526 14368
rect 22649 14365 22661 14368
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14365 22891 14399
rect 22833 14359 22891 14365
rect 22925 14399 22983 14405
rect 22925 14365 22937 14399
rect 22971 14396 22983 14399
rect 23198 14396 23204 14408
rect 22971 14368 23204 14396
rect 22971 14365 22983 14368
rect 22925 14359 22983 14365
rect 22848 14328 22876 14359
rect 23198 14356 23204 14368
rect 23256 14396 23262 14408
rect 23474 14396 23480 14408
rect 23256 14368 23480 14396
rect 23256 14356 23262 14368
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 24854 14356 24860 14408
rect 24912 14356 24918 14408
rect 24946 14356 24952 14408
rect 25004 14396 25010 14408
rect 25225 14399 25283 14405
rect 25225 14396 25237 14399
rect 25004 14368 25237 14396
rect 25004 14356 25010 14368
rect 25225 14365 25237 14368
rect 25271 14365 25283 14399
rect 25225 14359 25283 14365
rect 25590 14356 25596 14408
rect 25648 14356 25654 14408
rect 25682 14356 25688 14408
rect 25740 14396 25746 14408
rect 26804 14405 26832 14436
rect 26881 14433 26893 14467
rect 26927 14464 26939 14467
rect 27264 14464 27292 14572
rect 27430 14492 27436 14544
rect 27488 14492 27494 14544
rect 26927 14436 27292 14464
rect 26927 14433 26939 14436
rect 26881 14427 26939 14433
rect 25869 14399 25927 14405
rect 25869 14396 25881 14399
rect 25740 14368 25881 14396
rect 25740 14356 25746 14368
rect 25869 14365 25881 14368
rect 25915 14365 25927 14399
rect 25869 14359 25927 14365
rect 26421 14399 26479 14405
rect 26421 14365 26433 14399
rect 26467 14365 26479 14399
rect 26421 14359 26479 14365
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14365 26847 14399
rect 26789 14359 26847 14365
rect 23934 14328 23940 14340
rect 20088 14300 22692 14328
rect 22848 14300 23940 14328
rect 18322 14260 18328 14272
rect 18064 14232 18328 14260
rect 17313 14223 17371 14229
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 18782 14260 18788 14272
rect 18564 14232 18788 14260
rect 18564 14220 18570 14232
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19150 14220 19156 14272
rect 19208 14260 19214 14272
rect 20165 14263 20223 14269
rect 20165 14260 20177 14263
rect 19208 14232 20177 14260
rect 19208 14220 19214 14232
rect 20165 14229 20177 14232
rect 20211 14229 20223 14263
rect 20165 14223 20223 14229
rect 21174 14220 21180 14272
rect 21232 14220 21238 14272
rect 21358 14220 21364 14272
rect 21416 14260 21422 14272
rect 22005 14263 22063 14269
rect 22005 14260 22017 14263
rect 21416 14232 22017 14260
rect 21416 14220 21422 14232
rect 22005 14229 22017 14232
rect 22051 14260 22063 14263
rect 22554 14260 22560 14272
rect 22051 14232 22560 14260
rect 22051 14229 22063 14232
rect 22005 14223 22063 14229
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 22664 14260 22692 14300
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 24673 14263 24731 14269
rect 24673 14260 24685 14263
rect 22664 14232 24685 14260
rect 24673 14229 24685 14232
rect 24719 14229 24731 14263
rect 24673 14223 24731 14229
rect 26050 14220 26056 14272
rect 26108 14260 26114 14272
rect 26436 14260 26464 14359
rect 27338 14356 27344 14408
rect 27396 14356 27402 14408
rect 27448 14405 27476 14492
rect 27540 14464 27568 14572
rect 27614 14560 27620 14572
rect 27672 14560 27678 14612
rect 28353 14603 28411 14609
rect 28353 14569 28365 14603
rect 28399 14600 28411 14603
rect 29454 14600 29460 14612
rect 28399 14572 29460 14600
rect 28399 14569 28411 14572
rect 28353 14563 28411 14569
rect 29454 14560 29460 14572
rect 29512 14560 29518 14612
rect 29730 14560 29736 14612
rect 29788 14600 29794 14612
rect 32490 14600 32496 14612
rect 29788 14572 32496 14600
rect 29788 14560 29794 14572
rect 32490 14560 32496 14572
rect 32548 14560 32554 14612
rect 28166 14492 28172 14544
rect 28224 14532 28230 14544
rect 28626 14532 28632 14544
rect 28224 14504 28632 14532
rect 28224 14492 28230 14504
rect 28626 14492 28632 14504
rect 28684 14492 28690 14544
rect 28718 14492 28724 14544
rect 28776 14532 28782 14544
rect 29822 14532 29828 14544
rect 28776 14504 29828 14532
rect 28776 14492 28782 14504
rect 29822 14492 29828 14504
rect 29880 14532 29886 14544
rect 31570 14532 31576 14544
rect 29880 14504 31576 14532
rect 29880 14492 29886 14504
rect 31570 14492 31576 14504
rect 31628 14492 31634 14544
rect 31938 14492 31944 14544
rect 31996 14532 32002 14544
rect 34514 14532 34520 14544
rect 31996 14504 34520 14532
rect 31996 14492 32002 14504
rect 34514 14492 34520 14504
rect 34572 14492 34578 14544
rect 29270 14464 29276 14476
rect 27540 14436 29276 14464
rect 29270 14424 29276 14436
rect 29328 14424 29334 14476
rect 29454 14424 29460 14476
rect 29512 14464 29518 14476
rect 31110 14464 31116 14476
rect 29512 14436 30512 14464
rect 29512 14424 29518 14436
rect 27433 14399 27491 14405
rect 27433 14365 27445 14399
rect 27479 14365 27491 14399
rect 27433 14359 27491 14365
rect 27617 14399 27675 14405
rect 27617 14365 27629 14399
rect 27663 14365 27675 14399
rect 27617 14359 27675 14365
rect 26970 14288 26976 14340
rect 27028 14328 27034 14340
rect 27525 14331 27583 14337
rect 27525 14328 27537 14331
rect 27028 14300 27537 14328
rect 27028 14288 27034 14300
rect 27525 14297 27537 14300
rect 27571 14297 27583 14331
rect 27525 14291 27583 14297
rect 27632 14328 27660 14359
rect 27798 14356 27804 14408
rect 27856 14356 27862 14408
rect 27982 14356 27988 14408
rect 28040 14356 28046 14408
rect 28166 14356 28172 14408
rect 28224 14356 28230 14408
rect 29733 14399 29791 14405
rect 29733 14365 29745 14399
rect 29779 14396 29791 14399
rect 30282 14396 30288 14408
rect 29779 14368 30288 14396
rect 29779 14365 29791 14368
rect 29733 14359 29791 14365
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 30484 14405 30512 14436
rect 30760 14436 31116 14464
rect 30469 14399 30527 14405
rect 30469 14365 30481 14399
rect 30515 14365 30527 14399
rect 30469 14359 30527 14365
rect 30558 14356 30564 14408
rect 30616 14396 30622 14408
rect 30760 14405 30788 14436
rect 31110 14424 31116 14436
rect 31168 14424 31174 14476
rect 31018 14405 31024 14408
rect 30745 14399 30803 14405
rect 30616 14368 30661 14396
rect 30616 14356 30622 14368
rect 30745 14365 30757 14399
rect 30791 14365 30803 14399
rect 30745 14359 30803 14365
rect 30975 14399 31024 14405
rect 30975 14365 30987 14399
rect 31021 14365 31024 14399
rect 30975 14359 31024 14365
rect 31018 14356 31024 14359
rect 31076 14396 31082 14408
rect 31478 14396 31484 14408
rect 31076 14368 31484 14396
rect 31076 14356 31082 14368
rect 31478 14356 31484 14368
rect 31536 14356 31542 14408
rect 27890 14328 27896 14340
rect 27632 14300 27896 14328
rect 27632 14260 27660 14300
rect 27890 14288 27896 14300
rect 27948 14288 27954 14340
rect 28077 14331 28135 14337
rect 28077 14297 28089 14331
rect 28123 14297 28135 14331
rect 28077 14291 28135 14297
rect 26108 14232 27660 14260
rect 26108 14220 26114 14232
rect 27706 14220 27712 14272
rect 27764 14260 27770 14272
rect 28092 14260 28120 14291
rect 29454 14288 29460 14340
rect 29512 14328 29518 14340
rect 29638 14328 29644 14340
rect 29512 14300 29644 14328
rect 29512 14288 29518 14300
rect 29638 14288 29644 14300
rect 29696 14288 29702 14340
rect 30837 14331 30895 14337
rect 30837 14297 30849 14331
rect 30883 14297 30895 14331
rect 30837 14291 30895 14297
rect 27764 14232 28120 14260
rect 27764 14220 27770 14232
rect 28902 14220 28908 14272
rect 28960 14260 28966 14272
rect 29549 14263 29607 14269
rect 29549 14260 29561 14263
rect 28960 14232 29561 14260
rect 28960 14220 28966 14232
rect 29549 14229 29561 14232
rect 29595 14260 29607 14263
rect 30098 14260 30104 14272
rect 29595 14232 30104 14260
rect 29595 14229 29607 14232
rect 29549 14223 29607 14229
rect 30098 14220 30104 14232
rect 30156 14220 30162 14272
rect 30558 14220 30564 14272
rect 30616 14260 30622 14272
rect 30852 14260 30880 14291
rect 30616 14232 30880 14260
rect 31113 14263 31171 14269
rect 30616 14220 30622 14232
rect 31113 14229 31125 14263
rect 31159 14260 31171 14263
rect 32122 14260 32128 14272
rect 31159 14232 32128 14260
rect 31159 14229 31171 14232
rect 31113 14223 31171 14229
rect 32122 14220 32128 14232
rect 32180 14220 32186 14272
rect 1104 14170 36524 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 36524 14170
rect 1104 14096 36524 14118
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14025 4399 14059
rect 4341 14019 4399 14025
rect 5169 14059 5227 14065
rect 5169 14025 5181 14059
rect 5215 14056 5227 14059
rect 5258 14056 5264 14068
rect 5215 14028 5264 14056
rect 5215 14025 5227 14028
rect 5169 14019 5227 14025
rect 4356 13988 4384 14019
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 5718 14016 5724 14068
rect 5776 14056 5782 14068
rect 5911 14059 5969 14065
rect 5911 14056 5923 14059
rect 5776 14028 5923 14056
rect 5776 14016 5782 14028
rect 5911 14025 5923 14028
rect 5957 14025 5969 14059
rect 5911 14019 5969 14025
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 8386 14056 8392 14068
rect 6420 14028 8392 14056
rect 6420 14016 6426 14028
rect 4798 13988 4804 14000
rect 4356 13960 4804 13988
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 5353 13991 5411 13997
rect 5353 13988 5365 13991
rect 5092 13960 5365 13988
rect 2590 13880 2596 13932
rect 2648 13880 2654 13932
rect 3970 13880 3976 13932
rect 4028 13880 4034 13932
rect 4614 13880 4620 13932
rect 4672 13880 4678 13932
rect 5092 13929 5120 13960
rect 5353 13957 5365 13960
rect 5399 13988 5411 13991
rect 5997 13991 6055 13997
rect 5997 13988 6009 13991
rect 5399 13960 6009 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 5997 13957 6009 13960
rect 6043 13957 6055 13991
rect 5997 13951 6055 13957
rect 7852 13951 7880 14028
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 8665 14059 8723 14065
rect 8665 14025 8677 14059
rect 8711 14056 8723 14059
rect 9766 14056 9772 14068
rect 8711 14028 9772 14056
rect 8711 14025 8723 14028
rect 8665 14019 8723 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10137 14059 10195 14065
rect 10137 14025 10149 14059
rect 10183 14056 10195 14059
rect 11330 14056 11336 14068
rect 10183 14028 11336 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12710 14016 12716 14068
rect 12768 14016 12774 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 14700 14028 15240 14056
rect 14700 14016 14706 14028
rect 7832 13945 7890 13951
rect 8018 13948 8024 14000
rect 8076 13948 8082 14000
rect 8205 13991 8263 13997
rect 8205 13957 8217 13991
rect 8251 13988 8263 13991
rect 9033 13991 9091 13997
rect 9033 13988 9045 13991
rect 8251 13960 9045 13988
rect 8251 13957 8263 13960
rect 8205 13951 8263 13957
rect 9033 13957 9045 13960
rect 9079 13957 9091 13991
rect 10686 13988 10692 14000
rect 9033 13951 9091 13957
rect 9140 13960 10180 13988
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5261 13923 5319 13929
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 5442 13920 5448 13932
rect 5307 13892 5448 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 4706 13812 4712 13864
rect 4764 13852 4770 13864
rect 4908 13852 4936 13883
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 4764 13824 4936 13852
rect 4764 13812 4770 13824
rect 5552 13796 5580 13883
rect 5718 13880 5724 13932
rect 5776 13880 5782 13932
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 5828 13852 5856 13883
rect 6086 13880 6092 13932
rect 6144 13880 6150 13932
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13920 7343 13923
rect 7374 13920 7380 13932
rect 7331 13892 7380 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7650 13920 7656 13932
rect 7607 13892 7656 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 7832 13911 7844 13945
rect 7878 13911 7890 13945
rect 7832 13905 7890 13911
rect 7926 13880 7932 13932
rect 7984 13920 7990 13932
rect 7984 13892 8432 13920
rect 7984 13880 7990 13892
rect 5644 13824 5856 13852
rect 4433 13787 4491 13793
rect 4433 13784 4445 13787
rect 3896 13756 4445 13784
rect 2856 13719 2914 13725
rect 2856 13685 2868 13719
rect 2902 13716 2914 13719
rect 3896 13716 3924 13756
rect 4433 13753 4445 13756
rect 4479 13753 4491 13787
rect 4433 13747 4491 13753
rect 5534 13744 5540 13796
rect 5592 13744 5598 13796
rect 2902 13688 3924 13716
rect 2902 13685 2914 13688
rect 2856 13679 2914 13685
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5644 13716 5672 13824
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 5960 13824 7113 13852
rect 5960 13812 5966 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7484 13852 7512 13880
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 7484 13824 8309 13852
rect 7101 13815 7159 13821
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8404 13852 8432 13892
rect 8478 13880 8484 13932
rect 8536 13880 8542 13932
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 8846 13920 8852 13932
rect 8803 13892 8852 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9140 13852 9168 13960
rect 10152 13932 10180 13960
rect 10244 13960 10692 13988
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9398 13920 9404 13932
rect 9263 13892 9404 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9490 13880 9496 13932
rect 9548 13880 9554 13932
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9766 13920 9772 13932
rect 9723 13892 9772 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 10134 13880 10140 13932
rect 10192 13880 10198 13932
rect 10244 13929 10272 13960
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 11054 13988 11060 14000
rect 10796 13960 11060 13988
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10505 13923 10563 13929
rect 10505 13922 10517 13923
rect 10321 13883 10379 13889
rect 10428 13894 10517 13922
rect 8404 13824 9168 13852
rect 9309 13855 9367 13861
rect 8297 13815 8355 13821
rect 9309 13821 9321 13855
rect 9355 13852 9367 13855
rect 9582 13852 9588 13864
rect 9355 13824 9588 13852
rect 9355 13821 9367 13824
rect 9309 13815 9367 13821
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 9784 13852 9812 13880
rect 10336 13852 10364 13883
rect 9784 13824 10364 13852
rect 8202 13744 8208 13796
rect 8260 13744 8266 13796
rect 9401 13787 9459 13793
rect 9401 13753 9413 13787
rect 9447 13784 9459 13787
rect 9447 13756 9674 13784
rect 9447 13753 9459 13756
rect 9401 13747 9459 13753
rect 5408 13688 5672 13716
rect 9646 13716 9674 13756
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10428 13784 10456 13894
rect 10505 13889 10517 13894
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 10796 13920 10824 13960
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 13906 13988 13912 14000
rect 12360 13960 13912 13988
rect 10643 13892 10824 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10870 13880 10876 13932
rect 10928 13880 10934 13932
rect 12360 13929 12388 13960
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 15102 13948 15108 14000
rect 15160 13948 15166 14000
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 12618 13920 12624 13932
rect 12575 13892 12624 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10376 13756 10456 13784
rect 10674 13821 10701 13852
rect 10735 13821 10747 13855
rect 10674 13815 10747 13821
rect 10674 13784 10702 13815
rect 11882 13784 11888 13796
rect 10674 13756 11888 13784
rect 10376 13744 10382 13756
rect 10674 13716 10702 13756
rect 11882 13744 11888 13756
rect 11940 13784 11946 13796
rect 12360 13784 12388 13883
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 13170 13880 13176 13932
rect 13228 13880 13234 13932
rect 13446 13920 13452 13932
rect 13280 13892 13452 13920
rect 12989 13855 13047 13861
rect 12989 13821 13001 13855
rect 13035 13852 13047 13855
rect 13280 13852 13308 13892
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13920 13599 13923
rect 13814 13920 13820 13932
rect 13587 13892 13820 13920
rect 13587 13889 13599 13892
rect 13541 13883 13599 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 13035 13824 13308 13852
rect 13357 13855 13415 13861
rect 13035 13821 13047 13824
rect 12989 13815 13047 13821
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13630 13852 13636 13864
rect 13403 13824 13636 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13630 13812 13636 13824
rect 13688 13852 13694 13864
rect 14292 13852 14320 13883
rect 14458 13880 14464 13932
rect 14516 13920 14522 13932
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 14516 13892 14657 13920
rect 14516 13880 14522 13892
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14826 13880 14832 13932
rect 14884 13920 14890 13932
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14884 13892 15025 13920
rect 14884 13880 14890 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15212 13920 15240 14028
rect 15470 14016 15476 14068
rect 15528 14016 15534 14068
rect 15930 14016 15936 14068
rect 15988 14016 15994 14068
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 17770 14056 17776 14068
rect 17267 14028 17776 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 18322 14016 18328 14068
rect 18380 14056 18386 14068
rect 19150 14056 19156 14068
rect 18380 14028 19156 14056
rect 18380 14016 18386 14028
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20254 14056 20260 14068
rect 20119 14028 20260 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20254 14016 20260 14028
rect 20312 14056 20318 14068
rect 20438 14056 20444 14068
rect 20312 14028 20444 14056
rect 20312 14016 20318 14028
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 21174 14016 21180 14068
rect 21232 14056 21238 14068
rect 23382 14056 23388 14068
rect 21232 14028 23388 14056
rect 21232 14016 21238 14028
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 26602 14016 26608 14068
rect 26660 14016 26666 14068
rect 26970 14016 26976 14068
rect 27028 14056 27034 14068
rect 27065 14059 27123 14065
rect 27065 14056 27077 14059
rect 27028 14028 27077 14056
rect 27028 14016 27034 14028
rect 27065 14025 27077 14028
rect 27111 14025 27123 14059
rect 27065 14019 27123 14025
rect 27709 14059 27767 14065
rect 27709 14025 27721 14059
rect 27755 14056 27767 14059
rect 27982 14056 27988 14068
rect 27755 14028 27988 14056
rect 27755 14025 27767 14028
rect 27709 14019 27767 14025
rect 27982 14016 27988 14028
rect 28040 14056 28046 14068
rect 29914 14056 29920 14068
rect 28040 14028 29040 14056
rect 28040 14016 28046 14028
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 17589 13991 17647 13997
rect 16632 13960 17540 13988
rect 16632 13948 16638 13960
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15212 13892 15301 13920
rect 15013 13883 15071 13889
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15436 13892 15577 13920
rect 15436 13880 15442 13892
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 15749 13923 15807 13929
rect 15749 13889 15761 13923
rect 15795 13920 15807 13923
rect 16390 13920 16396 13932
rect 15795 13892 16396 13920
rect 15795 13889 15807 13892
rect 15749 13883 15807 13889
rect 16390 13880 16396 13892
rect 16448 13920 16454 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 16448 13892 17417 13920
rect 16448 13880 16454 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17512 13920 17540 13960
rect 17589 13957 17601 13991
rect 17635 13988 17647 13991
rect 17678 13988 17684 14000
rect 17635 13960 17684 13988
rect 17635 13957 17647 13960
rect 17589 13951 17647 13957
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 17862 13948 17868 14000
rect 17920 13988 17926 14000
rect 18874 13988 18880 14000
rect 17920 13960 18880 13988
rect 17920 13948 17926 13960
rect 18874 13948 18880 13960
rect 18932 13988 18938 14000
rect 19426 13988 19432 14000
rect 18932 13960 19432 13988
rect 18932 13948 18938 13960
rect 19426 13948 19432 13960
rect 19484 13988 19490 14000
rect 19702 13988 19708 14000
rect 19484 13960 19708 13988
rect 19484 13948 19490 13960
rect 19702 13948 19708 13960
rect 19760 13948 19766 14000
rect 19886 13948 19892 14000
rect 19944 13997 19950 14000
rect 19944 13991 19973 13997
rect 19961 13957 19973 13991
rect 27430 13988 27436 14000
rect 19944 13951 19973 13957
rect 26712 13960 27436 13988
rect 19944 13948 19950 13951
rect 19794 13920 19800 13932
rect 17512 13892 19800 13920
rect 17405 13883 17463 13889
rect 19794 13880 19800 13892
rect 19852 13880 19858 13932
rect 25041 13923 25099 13929
rect 25041 13920 25053 13923
rect 23400 13892 25053 13920
rect 13688 13824 14320 13852
rect 13688 13812 13694 13824
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 18966 13852 18972 13864
rect 15528 13824 18972 13852
rect 15528 13812 15534 13824
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19702 13812 19708 13864
rect 19760 13852 19766 13864
rect 20530 13852 20536 13864
rect 19760 13824 20536 13852
rect 19760 13812 19766 13824
rect 20530 13812 20536 13824
rect 20588 13852 20594 13864
rect 20714 13852 20720 13864
rect 20588 13824 20720 13852
rect 20588 13812 20594 13824
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 13449 13787 13507 13793
rect 13449 13784 13461 13787
rect 11940 13756 12388 13784
rect 13004 13756 13461 13784
rect 11940 13744 11946 13756
rect 13004 13728 13032 13756
rect 13449 13753 13461 13756
rect 13495 13753 13507 13787
rect 13449 13747 13507 13753
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 15620 13756 15700 13784
rect 15620 13744 15626 13756
rect 9646 13688 10702 13716
rect 5408 13676 5414 13688
rect 11054 13676 11060 13728
rect 11112 13676 11118 13728
rect 12526 13676 12532 13728
rect 12584 13676 12590 13728
rect 12986 13676 12992 13728
rect 13044 13676 13050 13728
rect 15672 13725 15700 13756
rect 16758 13744 16764 13796
rect 16816 13784 16822 13796
rect 17862 13784 17868 13796
rect 16816 13756 17868 13784
rect 16816 13744 16822 13756
rect 17862 13744 17868 13756
rect 17920 13784 17926 13796
rect 23198 13784 23204 13796
rect 17920 13756 23204 13784
rect 17920 13744 17926 13756
rect 23198 13744 23204 13756
rect 23256 13784 23262 13796
rect 23400 13784 23428 13892
rect 25041 13889 25053 13892
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13889 25375 13923
rect 25317 13883 25375 13889
rect 25501 13923 25559 13929
rect 25501 13889 25513 13923
rect 25547 13920 25559 13923
rect 25682 13920 25688 13932
rect 25547 13892 25688 13920
rect 25547 13889 25559 13892
rect 25501 13883 25559 13889
rect 24946 13812 24952 13864
rect 25004 13812 25010 13864
rect 25332 13852 25360 13883
rect 25682 13880 25688 13892
rect 25740 13880 25746 13932
rect 26712 13929 26740 13960
rect 27430 13948 27436 13960
rect 27488 13948 27494 14000
rect 29012 13997 29040 14028
rect 29380 14028 29920 14056
rect 28997 13991 29055 13997
rect 28184 13960 28923 13988
rect 28184 13932 28212 13960
rect 28895 13932 28923 13960
rect 28997 13957 29009 13991
rect 29043 13957 29055 13991
rect 29380 13988 29408 14028
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 32585 14059 32643 14065
rect 32585 14025 32597 14059
rect 32631 14056 32643 14059
rect 32950 14056 32956 14068
rect 32631 14028 32956 14056
rect 32631 14025 32643 14028
rect 32585 14019 32643 14025
rect 32950 14016 32956 14028
rect 33008 14016 33014 14068
rect 29733 13991 29791 13997
rect 28997 13951 29055 13957
rect 29288 13960 29593 13988
rect 26513 13923 26571 13929
rect 26513 13889 26525 13923
rect 26559 13889 26571 13923
rect 26513 13883 26571 13889
rect 26697 13923 26755 13929
rect 26697 13889 26709 13923
rect 26743 13889 26755 13923
rect 26697 13883 26755 13889
rect 26973 13923 27031 13929
rect 26973 13889 26985 13923
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27525 13923 27583 13929
rect 27525 13889 27537 13923
rect 27571 13920 27583 13923
rect 27614 13920 27620 13932
rect 27571 13892 27620 13920
rect 27571 13889 27583 13892
rect 27525 13883 27583 13889
rect 25590 13852 25596 13864
rect 25332 13824 25596 13852
rect 25590 13812 25596 13824
rect 25648 13852 25654 13864
rect 26528 13852 26556 13883
rect 25648 13824 26556 13852
rect 25648 13812 25654 13824
rect 23256 13756 23428 13784
rect 26528 13784 26556 13824
rect 26602 13812 26608 13864
rect 26660 13852 26666 13864
rect 26988 13852 27016 13883
rect 26660 13824 27016 13852
rect 26660 13812 26666 13824
rect 26970 13784 26976 13796
rect 26528 13756 26976 13784
rect 23256 13744 23262 13756
rect 26970 13744 26976 13756
rect 27028 13784 27034 13796
rect 27172 13784 27200 13883
rect 27614 13880 27620 13892
rect 27672 13880 27678 13932
rect 28166 13880 28172 13932
rect 28224 13880 28230 13932
rect 28258 13880 28264 13932
rect 28316 13880 28322 13932
rect 28350 13880 28356 13932
rect 28408 13880 28414 13932
rect 28491 13923 28549 13929
rect 28491 13889 28503 13923
rect 28537 13920 28549 13923
rect 28718 13920 28724 13932
rect 28537 13892 28724 13920
rect 28537 13889 28549 13892
rect 28491 13883 28549 13889
rect 28718 13880 28724 13892
rect 28776 13880 28782 13932
rect 28895 13890 28908 13932
rect 28900 13883 28908 13890
rect 28902 13880 28908 13883
rect 28960 13880 28966 13932
rect 29086 13880 29092 13932
rect 29144 13880 29150 13932
rect 29288 13929 29316 13960
rect 29565 13929 29593 13960
rect 29733 13957 29745 13991
rect 29779 13957 29791 13991
rect 29733 13951 29791 13957
rect 29272 13923 29330 13929
rect 29272 13889 29284 13923
rect 29318 13889 29330 13923
rect 29376 13923 29434 13929
rect 29376 13922 29388 13923
rect 29272 13883 29330 13889
rect 29362 13870 29368 13922
rect 29422 13889 29434 13923
rect 29420 13883 29434 13889
rect 29464 13923 29522 13929
rect 29464 13889 29476 13923
rect 29510 13889 29522 13923
rect 29464 13883 29522 13889
rect 29550 13923 29608 13929
rect 29550 13889 29562 13923
rect 29596 13889 29608 13923
rect 29550 13883 29608 13889
rect 29420 13870 29426 13883
rect 27341 13855 27399 13861
rect 27341 13852 27353 13855
rect 27028 13756 27200 13784
rect 27264 13824 27353 13852
rect 27028 13744 27034 13756
rect 15657 13719 15715 13725
rect 15657 13685 15669 13719
rect 15703 13685 15715 13719
rect 15657 13679 15715 13685
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 19334 13716 19340 13728
rect 17368 13688 19340 13716
rect 17368 13676 17374 13688
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 19877 13676 19883 13728
rect 19935 13676 19941 13728
rect 21634 13676 21640 13728
rect 21692 13716 21698 13728
rect 23934 13716 23940 13728
rect 21692 13688 23940 13716
rect 21692 13676 21698 13688
rect 23934 13676 23940 13688
rect 23992 13676 23998 13728
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 27154 13716 27160 13728
rect 26292 13688 27160 13716
rect 26292 13676 26298 13688
rect 27154 13676 27160 13688
rect 27212 13716 27218 13728
rect 27264 13716 27292 13824
rect 27341 13821 27353 13824
rect 27387 13821 27399 13855
rect 27341 13815 27399 13821
rect 27982 13812 27988 13864
rect 28040 13812 28046 13864
rect 28626 13812 28632 13864
rect 28684 13812 28690 13864
rect 29493 13852 29521 13883
rect 29748 13852 29776 13951
rect 32122 13948 32128 14000
rect 32180 13948 32186 14000
rect 29825 13923 29883 13929
rect 29825 13889 29837 13923
rect 29871 13889 29883 13923
rect 29825 13883 29883 13889
rect 29963 13923 30021 13929
rect 29963 13889 29975 13923
rect 30009 13920 30021 13923
rect 30098 13920 30104 13932
rect 30009 13892 30104 13920
rect 30009 13889 30021 13892
rect 29963 13883 30021 13889
rect 29472 13824 29521 13852
rect 29564 13824 29776 13852
rect 27212 13688 27292 13716
rect 27212 13676 27218 13688
rect 27982 13676 27988 13728
rect 28040 13716 28046 13728
rect 28258 13716 28264 13728
rect 28040 13688 28264 13716
rect 28040 13676 28046 13688
rect 28258 13676 28264 13688
rect 28316 13676 28322 13728
rect 28644 13716 28672 13812
rect 29472 13796 29500 13824
rect 28721 13787 28779 13793
rect 28721 13753 28733 13787
rect 28767 13784 28779 13787
rect 28810 13784 28816 13796
rect 28767 13756 28816 13784
rect 28767 13753 28779 13756
rect 28721 13747 28779 13753
rect 28810 13744 28816 13756
rect 28868 13744 28874 13796
rect 28902 13744 28908 13796
rect 28960 13784 28966 13796
rect 29454 13784 29460 13796
rect 28960 13756 29460 13784
rect 28960 13744 28966 13756
rect 29454 13744 29460 13756
rect 29512 13744 29518 13796
rect 29564 13716 29592 13824
rect 29840 13784 29868 13883
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 30650 13880 30656 13932
rect 30708 13880 30714 13932
rect 32401 13923 32459 13929
rect 32401 13889 32413 13923
rect 32447 13920 32459 13923
rect 33594 13920 33600 13932
rect 32447 13892 33600 13920
rect 32447 13889 32459 13892
rect 32401 13883 32459 13889
rect 33594 13880 33600 13892
rect 33652 13880 33658 13932
rect 30190 13852 30196 13864
rect 30116 13824 30196 13852
rect 29914 13784 29920 13796
rect 29840 13756 29920 13784
rect 29914 13744 29920 13756
rect 29972 13744 29978 13796
rect 30116 13793 30144 13824
rect 30190 13812 30196 13824
rect 30248 13812 30254 13864
rect 30745 13855 30803 13861
rect 30745 13821 30757 13855
rect 30791 13852 30803 13855
rect 31938 13852 31944 13864
rect 30791 13824 31944 13852
rect 30791 13821 30803 13824
rect 30745 13815 30803 13821
rect 31938 13812 31944 13824
rect 31996 13852 32002 13864
rect 32217 13855 32275 13861
rect 32217 13852 32229 13855
rect 31996 13824 32229 13852
rect 31996 13812 32002 13824
rect 32217 13821 32229 13824
rect 32263 13821 32275 13855
rect 32217 13815 32275 13821
rect 30101 13787 30159 13793
rect 30101 13753 30113 13787
rect 30147 13753 30159 13787
rect 30101 13747 30159 13753
rect 28644 13688 29592 13716
rect 31754 13676 31760 13728
rect 31812 13716 31818 13728
rect 32125 13719 32183 13725
rect 32125 13716 32137 13719
rect 31812 13688 32137 13716
rect 31812 13676 31818 13688
rect 32125 13685 32137 13688
rect 32171 13685 32183 13719
rect 32125 13679 32183 13685
rect 1104 13626 36524 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 36524 13626
rect 1104 13552 36524 13574
rect 4614 13472 4620 13524
rect 4672 13512 4678 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4672 13484 4905 13512
rect 4672 13472 4678 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 4893 13475 4951 13481
rect 5353 13515 5411 13521
rect 5353 13481 5365 13515
rect 5399 13512 5411 13515
rect 6086 13512 6092 13524
rect 5399 13484 6092 13512
rect 5399 13481 5411 13484
rect 5353 13475 5411 13481
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 9401 13515 9459 13521
rect 9401 13481 9413 13515
rect 9447 13512 9459 13515
rect 9490 13512 9496 13524
rect 9447 13484 9496 13512
rect 9447 13481 9459 13484
rect 9401 13475 9459 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 15289 13515 15347 13521
rect 10192 13484 10824 13512
rect 10192 13472 10198 13484
rect 4264 13416 5580 13444
rect 4264 13317 4292 13416
rect 5552 13388 5580 13416
rect 6730 13404 6736 13456
rect 6788 13444 6794 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 6788 13416 10425 13444
rect 6788 13404 6794 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 10796 13444 10824 13484
rect 15289 13481 15301 13515
rect 15335 13512 15347 13515
rect 15654 13512 15660 13524
rect 15335 13484 15660 13512
rect 15335 13481 15347 13484
rect 15289 13475 15347 13481
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15804 13484 16037 13512
rect 15804 13472 15810 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 16025 13475 16083 13481
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17552 13484 17877 13512
rect 17552 13472 17558 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 18046 13472 18052 13524
rect 18104 13472 18110 13524
rect 18690 13472 18696 13524
rect 18748 13472 18754 13524
rect 18877 13515 18935 13521
rect 18877 13481 18889 13515
rect 18923 13512 18935 13515
rect 19334 13512 19340 13524
rect 18923 13484 19340 13512
rect 18923 13481 18935 13484
rect 18877 13475 18935 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 20346 13512 20352 13524
rect 19725 13484 20352 13512
rect 13354 13444 13360 13456
rect 10796 13416 13360 13444
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13376 4399 13379
rect 5350 13376 5356 13388
rect 4387 13348 5356 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 10796 13376 10824 13416
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 17586 13444 17592 13456
rect 16132 13416 17592 13444
rect 5592 13348 9674 13376
rect 5592 13336 5598 13348
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13277 4307 13311
rect 4801 13311 4859 13317
rect 4801 13308 4813 13311
rect 4249 13271 4307 13277
rect 4632 13280 4813 13308
rect 4632 13181 4660 13280
rect 4801 13277 4813 13280
rect 4847 13277 4859 13311
rect 4801 13271 4859 13277
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13277 5043 13311
rect 4985 13271 5043 13277
rect 5261 13311 5319 13317
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5445 13311 5503 13317
rect 5445 13277 5457 13311
rect 5491 13308 5503 13311
rect 5718 13308 5724 13320
rect 5491 13280 5724 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 4706 13200 4712 13252
rect 4764 13240 4770 13252
rect 5000 13240 5028 13271
rect 4764 13212 5028 13240
rect 5276 13240 5304 13271
rect 5718 13268 5724 13280
rect 5776 13308 5782 13320
rect 6086 13308 6092 13320
rect 5776 13280 6092 13308
rect 5776 13268 5782 13280
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6362 13268 6368 13320
rect 6420 13268 6426 13320
rect 6564 13317 6592 13348
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9398 13308 9404 13320
rect 9355 13280 9404 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 9646 13308 9674 13348
rect 10704 13348 10824 13376
rect 10704 13317 10732 13348
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12124 13348 12633 13376
rect 12124 13336 12130 13348
rect 12621 13345 12633 13348
rect 12667 13345 12679 13379
rect 13722 13376 13728 13388
rect 12621 13339 12679 13345
rect 12820 13348 13728 13376
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 9646 13280 10609 13308
rect 10597 13277 10609 13280
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 5534 13240 5540 13252
rect 5276 13212 5540 13240
rect 4764 13200 4770 13212
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 10226 13240 10232 13252
rect 9732 13212 10232 13240
rect 9732 13200 9738 13212
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 10612 13240 10640 13271
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13308 11023 13311
rect 11054 13308 11060 13320
rect 11011 13280 11060 13308
rect 11011 13277 11023 13280
rect 10965 13271 11023 13277
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 12820 13317 12848 13348
rect 13722 13336 13728 13348
rect 13780 13376 13786 13388
rect 14090 13376 14096 13388
rect 13780 13348 14096 13376
rect 13780 13336 13786 13348
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 16132 13385 16160 13416
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 19725 13444 19753 13484
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 21082 13472 21088 13524
rect 21140 13512 21146 13524
rect 22094 13512 22100 13524
rect 21140 13484 22100 13512
rect 21140 13472 21146 13484
rect 17788 13416 19753 13444
rect 19812 13416 21312 13444
rect 16117 13379 16175 13385
rect 16117 13376 16129 13379
rect 15488 13348 16129 13376
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12805 13271 12863 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13170 13308 13176 13320
rect 13035 13280 13176 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 11238 13240 11244 13252
rect 10612 13212 11244 13240
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13141 4675 13175
rect 4617 13135 4675 13141
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6914 13172 6920 13184
rect 6503 13144 6920 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 8938 13132 8944 13184
rect 8996 13172 9002 13184
rect 12820 13172 12848 13271
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 15488 13317 15516 13348
rect 16117 13345 16129 13348
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13308 15807 13311
rect 16022 13308 16028 13320
rect 15795 13280 16028 13308
rect 15795 13277 15807 13280
rect 15749 13271 15807 13277
rect 15010 13200 15016 13252
rect 15068 13240 15074 13252
rect 15580 13240 15608 13271
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16206 13268 16212 13320
rect 16264 13268 16270 13320
rect 17788 13317 17816 13416
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 18104 13348 19257 13376
rect 18104 13336 18110 13348
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17862 13268 17868 13320
rect 17920 13308 17926 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17920 13280 17969 13308
rect 17920 13268 17926 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13308 18291 13311
rect 18322 13308 18328 13320
rect 18279 13280 18328 13308
rect 18279 13277 18291 13280
rect 18233 13271 18291 13277
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 19521 13311 19579 13317
rect 19521 13277 19533 13311
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 18138 13240 18144 13252
rect 15068 13212 15976 13240
rect 15068 13200 15074 13212
rect 8996 13144 12848 13172
rect 8996 13132 9002 13144
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 15841 13175 15899 13181
rect 15841 13172 15853 13175
rect 15712 13144 15853 13172
rect 15712 13132 15718 13144
rect 15841 13141 15853 13144
rect 15887 13141 15899 13175
rect 15948 13172 15976 13212
rect 16315 13212 18144 13240
rect 16315 13172 16343 13212
rect 18138 13200 18144 13212
rect 18196 13200 18202 13252
rect 19061 13243 19119 13249
rect 19061 13209 19073 13243
rect 19107 13240 19119 13243
rect 19150 13240 19156 13252
rect 19107 13212 19156 13240
rect 19107 13209 19119 13212
rect 19061 13203 19119 13209
rect 19150 13200 19156 13212
rect 19208 13200 19214 13252
rect 19536 13240 19564 13271
rect 19702 13268 19708 13320
rect 19760 13268 19766 13320
rect 19812 13317 19840 13416
rect 20162 13336 20168 13388
rect 20220 13376 20226 13388
rect 20438 13376 20444 13388
rect 20220 13348 20444 13376
rect 20220 13336 20226 13348
rect 20438 13336 20444 13348
rect 20496 13336 20502 13388
rect 21284 13320 21312 13416
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 20254 13268 20260 13320
rect 20312 13268 20318 13320
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 20404 13280 20449 13308
rect 20404 13268 20410 13280
rect 20622 13268 20628 13320
rect 20680 13268 20686 13320
rect 20763 13311 20821 13317
rect 20763 13277 20775 13311
rect 20809 13308 20821 13311
rect 20809 13280 21037 13308
rect 20809 13277 20821 13280
rect 20763 13271 20821 13277
rect 20070 13240 20076 13252
rect 19536 13212 20076 13240
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 20162 13200 20168 13252
rect 20220 13240 20226 13252
rect 20533 13243 20591 13249
rect 20533 13240 20545 13243
rect 20220 13212 20545 13240
rect 20220 13200 20226 13212
rect 20533 13209 20545 13212
rect 20579 13209 20591 13243
rect 20533 13203 20591 13209
rect 15948 13144 16343 13172
rect 15841 13135 15899 13141
rect 17494 13132 17500 13184
rect 17552 13132 17558 13184
rect 17586 13132 17592 13184
rect 17644 13172 17650 13184
rect 18414 13172 18420 13184
rect 17644 13144 18420 13172
rect 17644 13132 17650 13144
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 18861 13175 18919 13181
rect 18861 13141 18873 13175
rect 18907 13172 18919 13175
rect 19518 13172 19524 13184
rect 18907 13144 19524 13172
rect 18907 13141 18919 13144
rect 18861 13135 18919 13141
rect 19518 13132 19524 13144
rect 19576 13132 19582 13184
rect 20254 13132 20260 13184
rect 20312 13172 20318 13184
rect 20901 13175 20959 13181
rect 20901 13172 20913 13175
rect 20312 13144 20913 13172
rect 20312 13132 20318 13144
rect 20901 13141 20913 13144
rect 20947 13141 20959 13175
rect 21009 13172 21037 13280
rect 21266 13268 21272 13320
rect 21324 13268 21330 13320
rect 21468 13317 21496 13484
rect 22094 13472 22100 13484
rect 22152 13512 22158 13524
rect 26237 13515 26295 13521
rect 22152 13484 23152 13512
rect 22152 13472 22158 13484
rect 23124 13456 23152 13484
rect 26237 13481 26249 13515
rect 26283 13512 26295 13515
rect 26418 13512 26424 13524
rect 26283 13484 26424 13512
rect 26283 13481 26295 13484
rect 26237 13475 26295 13481
rect 26418 13472 26424 13484
rect 26476 13472 26482 13524
rect 26694 13472 26700 13524
rect 26752 13512 26758 13524
rect 26789 13515 26847 13521
rect 26789 13512 26801 13515
rect 26752 13484 26801 13512
rect 26752 13472 26758 13484
rect 26789 13481 26801 13484
rect 26835 13481 26847 13515
rect 26789 13475 26847 13481
rect 28166 13472 28172 13524
rect 28224 13512 28230 13524
rect 28718 13512 28724 13524
rect 28224 13484 28724 13512
rect 28224 13472 28230 13484
rect 28718 13472 28724 13484
rect 28776 13472 28782 13524
rect 28902 13472 28908 13524
rect 28960 13512 28966 13524
rect 31570 13512 31576 13524
rect 28960 13484 31576 13512
rect 28960 13472 28966 13484
rect 31570 13472 31576 13484
rect 31628 13472 31634 13524
rect 31665 13515 31723 13521
rect 31665 13481 31677 13515
rect 31711 13481 31723 13515
rect 31665 13475 31723 13481
rect 21542 13404 21548 13456
rect 21600 13444 21606 13456
rect 21600 13416 21956 13444
rect 21600 13404 21606 13416
rect 21928 13320 21956 13416
rect 23106 13404 23112 13456
rect 23164 13444 23170 13456
rect 27338 13444 27344 13456
rect 23164 13416 27344 13444
rect 23164 13404 23170 13416
rect 27338 13404 27344 13416
rect 27396 13404 27402 13456
rect 31680 13444 31708 13475
rect 31754 13472 31760 13524
rect 31812 13512 31818 13524
rect 33321 13515 33379 13521
rect 33321 13512 33333 13515
rect 31812 13484 33333 13512
rect 31812 13472 31818 13484
rect 33321 13481 33333 13484
rect 33367 13512 33379 13515
rect 34149 13515 34207 13521
rect 34149 13512 34161 13515
rect 33367 13484 34161 13512
rect 33367 13481 33379 13484
rect 33321 13475 33379 13481
rect 34149 13481 34161 13484
rect 34195 13481 34207 13515
rect 34149 13475 34207 13481
rect 34790 13472 34796 13524
rect 34848 13512 34854 13524
rect 34977 13515 35035 13521
rect 34977 13512 34989 13515
rect 34848 13484 34989 13512
rect 34848 13472 34854 13484
rect 34977 13481 34989 13484
rect 35023 13481 35035 13515
rect 34977 13475 35035 13481
rect 33042 13444 33048 13456
rect 31680 13416 33048 13444
rect 33042 13404 33048 13416
rect 33100 13404 33106 13456
rect 33134 13404 33140 13456
rect 33192 13404 33198 13456
rect 25682 13336 25688 13388
rect 25740 13336 25746 13388
rect 25777 13379 25835 13385
rect 25777 13345 25789 13379
rect 25823 13376 25835 13379
rect 25823 13348 26832 13376
rect 25823 13345 25835 13348
rect 25777 13339 25835 13345
rect 21453 13311 21511 13317
rect 21453 13277 21465 13311
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 21634 13268 21640 13320
rect 21692 13268 21698 13320
rect 21821 13311 21879 13317
rect 21821 13277 21833 13311
rect 21867 13277 21879 13311
rect 21821 13271 21879 13277
rect 21082 13200 21088 13252
rect 21140 13240 21146 13252
rect 21836 13240 21864 13271
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22189 13311 22247 13317
rect 22189 13308 22201 13311
rect 21968 13280 22201 13308
rect 21968 13268 21974 13280
rect 22189 13277 22201 13280
rect 22235 13277 22247 13311
rect 22189 13271 22247 13277
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 25501 13311 25559 13317
rect 25501 13308 25513 13311
rect 24820 13280 25513 13308
rect 24820 13268 24826 13280
rect 25501 13277 25513 13280
rect 25547 13277 25559 13311
rect 25501 13271 25559 13277
rect 21140 13212 21864 13240
rect 22097 13243 22155 13249
rect 21140 13200 21146 13212
rect 22097 13209 22109 13243
rect 22143 13240 22155 13243
rect 23658 13240 23664 13252
rect 22143 13212 23664 13240
rect 22143 13209 22155 13212
rect 22097 13203 22155 13209
rect 23658 13200 23664 13212
rect 23716 13200 23722 13252
rect 25516 13240 25544 13271
rect 25590 13268 25596 13320
rect 25648 13308 25654 13320
rect 26050 13308 26056 13320
rect 25648 13280 26056 13308
rect 25648 13268 25654 13280
rect 26050 13268 26056 13280
rect 26108 13268 26114 13320
rect 26237 13311 26295 13317
rect 26237 13277 26249 13311
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13308 26479 13311
rect 26602 13308 26608 13320
rect 26467 13280 26608 13308
rect 26467 13277 26479 13280
rect 26421 13271 26479 13277
rect 26252 13240 26280 13271
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 26804 13317 26832 13348
rect 28074 13336 28080 13388
rect 28132 13376 28138 13388
rect 28994 13376 29000 13388
rect 28132 13348 29000 13376
rect 28132 13336 28138 13348
rect 28994 13336 29000 13348
rect 29052 13336 29058 13388
rect 31846 13336 31852 13388
rect 31904 13336 31910 13388
rect 33505 13379 33563 13385
rect 33505 13345 33517 13379
rect 33551 13376 33563 13379
rect 34808 13376 34836 13472
rect 35434 13404 35440 13456
rect 35492 13404 35498 13456
rect 33551 13348 34836 13376
rect 35161 13379 35219 13385
rect 33551 13345 33563 13348
rect 33505 13339 33563 13345
rect 35161 13345 35173 13379
rect 35207 13376 35219 13379
rect 35342 13376 35348 13388
rect 35207 13348 35348 13376
rect 35207 13345 35219 13348
rect 35161 13339 35219 13345
rect 35342 13336 35348 13348
rect 35400 13336 35406 13388
rect 26789 13311 26847 13317
rect 26789 13277 26801 13311
rect 26835 13308 26847 13311
rect 26878 13308 26884 13320
rect 26835 13280 26884 13308
rect 26835 13277 26847 13280
rect 26789 13271 26847 13277
rect 26878 13268 26884 13280
rect 26936 13268 26942 13320
rect 26970 13268 26976 13320
rect 27028 13268 27034 13320
rect 28442 13268 28448 13320
rect 28500 13308 28506 13320
rect 28626 13308 28632 13320
rect 28500 13280 28632 13308
rect 28500 13268 28506 13280
rect 28626 13268 28632 13280
rect 28684 13268 28690 13320
rect 29270 13268 29276 13320
rect 29328 13308 29334 13320
rect 29914 13308 29920 13320
rect 29328 13280 29920 13308
rect 29328 13268 29334 13280
rect 29914 13268 29920 13280
rect 29972 13268 29978 13320
rect 31938 13268 31944 13320
rect 31996 13268 32002 13320
rect 32490 13268 32496 13320
rect 32548 13308 32554 13320
rect 33321 13311 33379 13317
rect 33321 13308 33333 13311
rect 32548 13280 33333 13308
rect 32548 13268 32554 13280
rect 33321 13277 33333 13280
rect 33367 13277 33379 13311
rect 33321 13271 33379 13277
rect 33870 13268 33876 13320
rect 33928 13308 33934 13320
rect 34149 13311 34207 13317
rect 34149 13308 34161 13311
rect 33928 13280 34161 13308
rect 33928 13268 33934 13280
rect 34149 13277 34161 13280
rect 34195 13277 34207 13311
rect 34149 13271 34207 13277
rect 34330 13268 34336 13320
rect 34388 13268 34394 13320
rect 35452 13317 35480 13404
rect 34977 13311 35035 13317
rect 34977 13308 34989 13311
rect 34532 13280 34989 13308
rect 25516 13212 26280 13240
rect 27154 13200 27160 13252
rect 27212 13240 27218 13252
rect 28994 13240 29000 13252
rect 27212 13212 29000 13240
rect 27212 13200 27218 13212
rect 28994 13200 29000 13212
rect 29052 13200 29058 13252
rect 31662 13200 31668 13252
rect 31720 13200 31726 13252
rect 33042 13200 33048 13252
rect 33100 13240 33106 13252
rect 33597 13243 33655 13249
rect 33597 13240 33609 13243
rect 33100 13212 33609 13240
rect 33100 13200 33106 13212
rect 33597 13209 33609 13212
rect 33643 13209 33655 13243
rect 33597 13203 33655 13209
rect 34532 13184 34560 13280
rect 34977 13277 34989 13280
rect 35023 13277 35035 13311
rect 34977 13271 35035 13277
rect 35437 13311 35495 13317
rect 35437 13277 35449 13311
rect 35483 13277 35495 13311
rect 35437 13271 35495 13277
rect 22278 13172 22284 13184
rect 21009 13144 22284 13172
rect 20901 13135 20959 13141
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 23566 13132 23572 13184
rect 23624 13172 23630 13184
rect 25317 13175 25375 13181
rect 25317 13172 25329 13175
rect 23624 13144 25329 13172
rect 23624 13132 23630 13144
rect 25317 13141 25329 13144
rect 25363 13141 25375 13175
rect 25317 13135 25375 13141
rect 26786 13132 26792 13184
rect 26844 13172 26850 13184
rect 27614 13172 27620 13184
rect 26844 13144 27620 13172
rect 26844 13132 26850 13144
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 32122 13132 32128 13184
rect 32180 13132 32186 13184
rect 34514 13132 34520 13184
rect 34572 13132 34578 13184
rect 34790 13132 34796 13184
rect 34848 13132 34854 13184
rect 1104 13082 36524 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 36524 13082
rect 1104 13008 36524 13030
rect 5350 12928 5356 12980
rect 5408 12928 5414 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 9030 12968 9036 12980
rect 8536 12940 9036 12968
rect 8536 12928 8542 12940
rect 9030 12928 9036 12940
rect 9088 12968 9094 12980
rect 9088 12940 9168 12968
rect 9088 12928 9094 12940
rect 5718 12860 5724 12912
rect 5776 12900 5782 12912
rect 6457 12903 6515 12909
rect 6457 12900 6469 12903
rect 5776 12872 6469 12900
rect 5776 12860 5782 12872
rect 6457 12869 6469 12872
rect 6503 12869 6515 12903
rect 7190 12900 7196 12912
rect 6457 12863 6515 12869
rect 6564 12872 7196 12900
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 5902 12832 5908 12844
rect 5583 12804 5908 12832
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6564 12841 6592 12872
rect 7190 12860 7196 12872
rect 7248 12900 7254 12912
rect 7650 12900 7656 12912
rect 7248 12872 7656 12900
rect 7248 12860 7254 12872
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 9140 12909 9168 12940
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10962 12968 10968 12980
rect 10468 12940 10968 12968
rect 10468 12928 10474 12940
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 15286 12928 15292 12980
rect 15344 12928 15350 12980
rect 15746 12928 15752 12980
rect 15804 12928 15810 12980
rect 17221 12971 17279 12977
rect 17221 12937 17233 12971
rect 17267 12968 17279 12971
rect 17310 12968 17316 12980
rect 17267 12940 17316 12968
rect 17267 12937 17279 12940
rect 17221 12931 17279 12937
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 18417 12971 18475 12977
rect 18417 12937 18429 12971
rect 18463 12968 18475 12971
rect 18598 12968 18604 12980
rect 18463 12940 18604 12968
rect 18463 12937 18475 12940
rect 18417 12931 18475 12937
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 19702 12928 19708 12980
rect 19760 12968 19766 12980
rect 19797 12971 19855 12977
rect 19797 12968 19809 12971
rect 19760 12940 19809 12968
rect 19760 12928 19766 12940
rect 19797 12937 19809 12940
rect 19843 12937 19855 12971
rect 19797 12931 19855 12937
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20517 12971 20575 12977
rect 20517 12968 20529 12971
rect 20036 12940 20529 12968
rect 20036 12928 20042 12940
rect 20517 12937 20529 12940
rect 20563 12968 20575 12971
rect 21174 12968 21180 12980
rect 20563 12940 21180 12968
rect 20563 12937 20575 12940
rect 20517 12931 20575 12937
rect 8205 12903 8263 12909
rect 8205 12900 8217 12903
rect 7944 12872 8217 12900
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6380 12764 6408 12795
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 6914 12764 6920 12776
rect 6380 12736 6920 12764
rect 6914 12724 6920 12736
rect 6972 12764 6978 12776
rect 7466 12764 7472 12776
rect 6972 12736 7472 12764
rect 6972 12724 6978 12736
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7558 12724 7564 12776
rect 7616 12724 7622 12776
rect 7944 12705 7972 12872
rect 8205 12869 8217 12872
rect 8251 12900 8263 12903
rect 9125 12903 9183 12909
rect 8251 12872 8892 12900
rect 8251 12869 8263 12872
rect 8205 12863 8263 12869
rect 8110 12792 8116 12844
rect 8168 12792 8174 12844
rect 8294 12792 8300 12844
rect 8352 12792 8358 12844
rect 8568 12835 8626 12841
rect 8568 12801 8580 12835
rect 8614 12801 8626 12835
rect 8568 12795 8626 12801
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8202 12764 8208 12776
rect 8067 12736 8208 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8588 12764 8616 12795
rect 8662 12792 8668 12844
rect 8720 12792 8726 12844
rect 8754 12792 8760 12844
rect 8812 12792 8818 12844
rect 8864 12841 8892 12872
rect 9125 12869 9137 12903
rect 9171 12869 9183 12903
rect 9125 12863 9183 12869
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 12066 12900 12072 12912
rect 9732 12872 12072 12900
rect 9732 12860 9738 12872
rect 8864 12835 8943 12841
rect 8864 12804 8897 12835
rect 8885 12801 8897 12804
rect 8931 12801 8943 12835
rect 8885 12795 8943 12801
rect 9030 12792 9036 12844
rect 9088 12792 9094 12844
rect 9214 12792 9220 12844
rect 9272 12832 9278 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 9272 12804 9321 12832
rect 9272 12792 9278 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 10520 12841 10548 12872
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 14182 12860 14188 12912
rect 14240 12900 14246 12912
rect 17405 12903 17463 12909
rect 17405 12900 17417 12903
rect 14240 12872 17417 12900
rect 14240 12860 14246 12872
rect 17405 12869 17417 12872
rect 17451 12869 17463 12903
rect 17405 12863 17463 12869
rect 17604 12872 19840 12900
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 10192 12804 10241 12832
rect 10192 12792 10198 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 10318 12764 10324 12776
rect 8588 12736 10324 12764
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12764 10471 12767
rect 10594 12764 10600 12776
rect 10459 12736 10600 12764
rect 10459 12733 10471 12736
rect 10413 12727 10471 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 7929 12699 7987 12705
rect 7929 12665 7941 12699
rect 7975 12665 7987 12699
rect 7929 12659 7987 12665
rect 8662 12656 8668 12708
rect 8720 12696 8726 12708
rect 9214 12696 9220 12708
rect 8720 12668 9220 12696
rect 8720 12656 8726 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 9306 12656 9312 12708
rect 9364 12696 9370 12708
rect 9582 12696 9588 12708
rect 9364 12668 9588 12696
rect 9364 12656 9370 12668
rect 9582 12656 9588 12668
rect 9640 12696 9646 12708
rect 10796 12696 10824 12795
rect 10962 12792 10968 12844
rect 11020 12792 11026 12844
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11388 12804 11529 12832
rect 11388 12792 11394 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 11790 12832 11796 12844
rect 11747 12804 11796 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 15010 12792 15016 12844
rect 15068 12792 15074 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15470 12832 15476 12844
rect 15243 12804 15476 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 15562 12792 15568 12844
rect 15620 12792 15626 12844
rect 15654 12792 15660 12844
rect 15712 12792 15718 12844
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12832 15991 12835
rect 16022 12832 16028 12844
rect 15979 12804 16028 12832
rect 15979 12801 15991 12804
rect 15933 12795 15991 12801
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16114 12792 16120 12844
rect 16172 12792 16178 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 16132 12764 16160 12792
rect 14608 12736 16160 12764
rect 17052 12764 17080 12795
rect 17310 12792 17316 12844
rect 17368 12792 17374 12844
rect 17604 12841 17632 12872
rect 19812 12844 19840 12872
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12832 17739 12835
rect 17770 12832 17776 12844
rect 17727 12804 17776 12832
rect 17727 12801 17739 12804
rect 17681 12795 17739 12801
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 17862 12792 17868 12844
rect 17920 12792 17926 12844
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 17957 12795 18015 12801
rect 17880 12764 17908 12792
rect 17052 12736 17908 12764
rect 17972 12764 18000 12795
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12832 18291 12835
rect 19242 12832 19248 12844
rect 18279 12804 19248 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 18248 12764 18276 12795
rect 19242 12792 19248 12804
rect 19300 12792 19306 12844
rect 19794 12792 19800 12844
rect 19852 12792 19858 12844
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19944 12804 19993 12832
rect 19944 12792 19950 12804
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12832 20223 12835
rect 20532 12832 20560 12931
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 26234 12968 26240 12980
rect 25280 12940 26240 12968
rect 25280 12928 25286 12940
rect 26234 12928 26240 12940
rect 26292 12928 26298 12980
rect 26694 12928 26700 12980
rect 26752 12968 26758 12980
rect 31205 12971 31263 12977
rect 26752 12940 28396 12968
rect 26752 12928 26758 12940
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 20717 12903 20775 12909
rect 20717 12900 20729 12903
rect 20680 12872 20729 12900
rect 20680 12860 20686 12872
rect 20717 12869 20729 12872
rect 20763 12869 20775 12903
rect 20717 12863 20775 12869
rect 20990 12860 20996 12912
rect 21048 12900 21054 12912
rect 21726 12900 21732 12912
rect 21048 12872 21732 12900
rect 21048 12860 21054 12872
rect 21726 12860 21732 12872
rect 21784 12860 21790 12912
rect 24578 12860 24584 12912
rect 24636 12900 24642 12912
rect 25866 12900 25872 12912
rect 24636 12872 25872 12900
rect 24636 12860 24642 12872
rect 25866 12860 25872 12872
rect 25924 12900 25930 12912
rect 26602 12900 26608 12912
rect 25924 12872 26188 12900
rect 25924 12860 25930 12872
rect 20211 12804 20560 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 21358 12792 21364 12844
rect 21416 12832 21422 12844
rect 22094 12832 22100 12844
rect 21416 12804 22100 12832
rect 21416 12792 21422 12804
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22554 12792 22560 12844
rect 22612 12792 22618 12844
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 23658 12792 23664 12844
rect 23716 12792 23722 12844
rect 24210 12792 24216 12844
rect 24268 12792 24274 12844
rect 25409 12835 25467 12841
rect 25409 12801 25421 12835
rect 25455 12832 25467 12835
rect 25590 12832 25596 12844
rect 25455 12804 25596 12832
rect 25455 12801 25467 12804
rect 25409 12795 25467 12801
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 26160 12841 26188 12872
rect 26344 12872 26608 12900
rect 26344 12841 26372 12872
rect 26602 12860 26608 12872
rect 26660 12860 26666 12912
rect 27246 12900 27252 12912
rect 26712 12872 27252 12900
rect 26712 12844 26740 12872
rect 27246 12860 27252 12872
rect 27304 12860 27310 12912
rect 27338 12860 27344 12912
rect 27396 12900 27402 12912
rect 27709 12903 27767 12909
rect 27709 12900 27721 12903
rect 27396 12872 27721 12900
rect 27396 12860 27402 12872
rect 27709 12869 27721 12872
rect 27755 12869 27767 12903
rect 27709 12863 27767 12869
rect 28166 12860 28172 12912
rect 28224 12900 28230 12912
rect 28261 12903 28319 12909
rect 28261 12900 28273 12903
rect 28224 12872 28273 12900
rect 28224 12860 28230 12872
rect 28261 12869 28273 12872
rect 28307 12869 28319 12903
rect 28261 12863 28319 12869
rect 26145 12835 26203 12841
rect 26145 12801 26157 12835
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 26513 12835 26571 12841
rect 26513 12801 26525 12835
rect 26559 12801 26571 12835
rect 26513 12795 26571 12801
rect 17972 12736 18276 12764
rect 14608 12724 14614 12736
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 19576 12736 20269 12764
rect 19576 12724 19582 12736
rect 20257 12733 20269 12736
rect 20303 12764 20315 12767
rect 23014 12764 23020 12776
rect 20303 12736 23020 12764
rect 20303 12733 20315 12736
rect 20257 12727 20315 12733
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 24394 12724 24400 12776
rect 24452 12724 24458 12776
rect 24762 12764 24768 12776
rect 24596 12736 24768 12764
rect 9640 12668 10824 12696
rect 9640 12656 9646 12668
rect 11422 12656 11428 12708
rect 11480 12696 11486 12708
rect 12526 12696 12532 12708
rect 11480 12668 12532 12696
rect 11480 12656 11486 12668
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 13170 12656 13176 12708
rect 13228 12696 13234 12708
rect 13354 12696 13360 12708
rect 13228 12668 13360 12696
rect 13228 12656 13234 12668
rect 13354 12656 13360 12668
rect 13412 12656 13418 12708
rect 15194 12656 15200 12708
rect 15252 12696 15258 12708
rect 15746 12696 15752 12708
rect 15252 12668 15752 12696
rect 15252 12656 15258 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 17310 12656 17316 12708
rect 17368 12696 17374 12708
rect 17368 12668 18092 12696
rect 17368 12656 17374 12668
rect 8386 12588 8392 12640
rect 8444 12588 8450 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 8754 12628 8760 12640
rect 8628 12600 8760 12628
rect 8628 12588 8634 12600
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 9490 12588 9496 12640
rect 9548 12588 9554 12640
rect 10042 12588 10048 12640
rect 10100 12588 10106 12640
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10376 12600 10609 12628
rect 10376 12588 10382 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 10597 12591 10655 12597
rect 10962 12588 10968 12640
rect 11020 12588 11026 12640
rect 11701 12631 11759 12637
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 12066 12628 12072 12640
rect 11747 12600 12072 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 13078 12588 13084 12640
rect 13136 12628 13142 12640
rect 15013 12631 15071 12637
rect 15013 12628 15025 12631
rect 13136 12600 15025 12628
rect 13136 12588 13142 12600
rect 15013 12597 15025 12600
rect 15059 12597 15071 12631
rect 15013 12591 15071 12597
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 16298 12628 16304 12640
rect 15712 12600 16304 12628
rect 15712 12588 15718 12600
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 16942 12628 16948 12640
rect 16899 12600 16948 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 18064 12637 18092 12668
rect 18138 12656 18144 12708
rect 18196 12696 18202 12708
rect 18196 12668 20024 12696
rect 18196 12656 18202 12668
rect 18049 12631 18107 12637
rect 18049 12597 18061 12631
rect 18095 12597 18107 12631
rect 19996 12628 20024 12668
rect 24210 12656 24216 12708
rect 24268 12696 24274 12708
rect 24596 12696 24624 12736
rect 24762 12724 24768 12736
rect 24820 12764 24826 12776
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24820 12736 25145 12764
rect 24820 12724 24826 12736
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 25498 12724 25504 12776
rect 25556 12764 25562 12776
rect 25682 12764 25688 12776
rect 25556 12736 25688 12764
rect 25556 12724 25562 12736
rect 25682 12724 25688 12736
rect 25740 12724 25746 12776
rect 25961 12767 26019 12773
rect 25961 12733 25973 12767
rect 26007 12733 26019 12767
rect 26528 12764 26556 12795
rect 26694 12792 26700 12844
rect 26752 12792 26758 12844
rect 27062 12792 27068 12844
rect 27120 12792 27126 12844
rect 27430 12792 27436 12844
rect 27488 12792 27494 12844
rect 27801 12835 27859 12841
rect 27801 12832 27813 12835
rect 27540 12804 27813 12832
rect 26786 12764 26792 12776
rect 26528 12736 26792 12764
rect 25961 12727 26019 12733
rect 24268 12668 24624 12696
rect 24268 12656 24274 12668
rect 24670 12656 24676 12708
rect 24728 12696 24734 12708
rect 24946 12696 24952 12708
rect 24728 12668 24952 12696
rect 24728 12656 24734 12668
rect 24946 12656 24952 12668
rect 25004 12656 25010 12708
rect 25866 12656 25872 12708
rect 25924 12656 25930 12708
rect 25976 12696 26004 12727
rect 26786 12724 26792 12736
rect 26844 12724 26850 12776
rect 27154 12724 27160 12776
rect 27212 12764 27218 12776
rect 27540 12764 27568 12804
rect 27801 12801 27813 12804
rect 27847 12801 27859 12835
rect 27801 12795 27859 12801
rect 27890 12792 27896 12844
rect 27948 12832 27954 12844
rect 27985 12835 28043 12841
rect 27985 12832 27997 12835
rect 27948 12804 27997 12832
rect 27948 12792 27954 12804
rect 27985 12801 27997 12804
rect 28031 12801 28043 12835
rect 27985 12795 28043 12801
rect 28074 12792 28080 12844
rect 28132 12792 28138 12844
rect 28368 12841 28396 12940
rect 29937 12940 30972 12968
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12801 28411 12835
rect 28353 12795 28411 12801
rect 28445 12835 28503 12841
rect 28445 12801 28457 12835
rect 28491 12832 28503 12835
rect 28718 12832 28724 12844
rect 28491 12804 28724 12832
rect 28491 12801 28503 12804
rect 28445 12795 28503 12801
rect 28718 12792 28724 12804
rect 28776 12792 28782 12844
rect 28994 12792 29000 12844
rect 29052 12832 29058 12844
rect 29454 12832 29460 12844
rect 29052 12804 29460 12832
rect 29052 12792 29058 12804
rect 29454 12792 29460 12804
rect 29512 12792 29518 12844
rect 27212 12736 27568 12764
rect 27212 12724 27218 12736
rect 27614 12724 27620 12776
rect 27672 12764 27678 12776
rect 29937 12764 29965 12940
rect 30466 12792 30472 12844
rect 30524 12832 30530 12844
rect 30742 12841 30748 12844
rect 30561 12835 30619 12841
rect 30561 12832 30573 12835
rect 30524 12804 30573 12832
rect 30524 12792 30530 12804
rect 30561 12801 30573 12804
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 30709 12835 30748 12841
rect 30709 12801 30721 12835
rect 30709 12795 30748 12801
rect 30742 12792 30748 12795
rect 30800 12792 30806 12844
rect 30944 12841 30972 12940
rect 31205 12937 31217 12971
rect 31251 12968 31263 12971
rect 32306 12968 32312 12980
rect 31251 12940 32312 12968
rect 31251 12937 31263 12940
rect 31205 12931 31263 12937
rect 32306 12928 32312 12940
rect 32364 12968 32370 12980
rect 32490 12968 32496 12980
rect 32364 12940 32496 12968
rect 32364 12928 32370 12940
rect 32490 12928 32496 12940
rect 32548 12928 32554 12980
rect 33410 12928 33416 12980
rect 33468 12968 33474 12980
rect 33686 12968 33692 12980
rect 33468 12940 33692 12968
rect 33468 12928 33474 12940
rect 33686 12928 33692 12940
rect 33744 12928 33750 12980
rect 30837 12835 30895 12841
rect 30837 12801 30849 12835
rect 30883 12801 30895 12835
rect 30837 12795 30895 12801
rect 30929 12835 30987 12841
rect 30929 12801 30941 12835
rect 30975 12801 30987 12835
rect 30929 12795 30987 12801
rect 27672 12736 29965 12764
rect 30852 12764 30880 12795
rect 31018 12792 31024 12844
rect 31076 12841 31082 12844
rect 31076 12832 31084 12841
rect 31754 12832 31760 12844
rect 31076 12804 31760 12832
rect 31076 12795 31084 12804
rect 31076 12792 31082 12795
rect 31754 12792 31760 12804
rect 31812 12792 31818 12844
rect 30852 12736 30972 12764
rect 27672 12724 27678 12736
rect 30944 12708 30972 12736
rect 26697 12699 26755 12705
rect 26697 12696 26709 12699
rect 25976 12668 26709 12696
rect 26697 12665 26709 12668
rect 26743 12696 26755 12699
rect 26878 12696 26884 12708
rect 26743 12668 26884 12696
rect 26743 12665 26755 12668
rect 26697 12659 26755 12665
rect 26878 12656 26884 12668
rect 26936 12656 26942 12708
rect 28074 12656 28080 12708
rect 28132 12696 28138 12708
rect 28629 12699 28687 12705
rect 28132 12668 28396 12696
rect 28132 12656 28138 12668
rect 20349 12631 20407 12637
rect 20349 12628 20361 12631
rect 19996 12600 20361 12628
rect 18049 12591 18107 12597
rect 20349 12597 20361 12600
rect 20395 12597 20407 12631
rect 20349 12591 20407 12597
rect 20530 12588 20536 12640
rect 20588 12588 20594 12640
rect 22738 12588 22744 12640
rect 22796 12628 22802 12640
rect 26145 12631 26203 12637
rect 26145 12628 26157 12631
rect 22796 12600 26157 12628
rect 22796 12588 22802 12600
rect 26145 12597 26157 12600
rect 26191 12597 26203 12631
rect 26145 12591 26203 12597
rect 27985 12631 28043 12637
rect 27985 12597 27997 12631
rect 28031 12628 28043 12631
rect 28258 12628 28264 12640
rect 28031 12600 28264 12628
rect 28031 12597 28043 12600
rect 27985 12591 28043 12597
rect 28258 12588 28264 12600
rect 28316 12588 28322 12640
rect 28368 12628 28396 12668
rect 28629 12665 28641 12699
rect 28675 12696 28687 12699
rect 30742 12696 30748 12708
rect 28675 12668 30748 12696
rect 28675 12665 28687 12668
rect 28629 12659 28687 12665
rect 30742 12656 30748 12668
rect 30800 12656 30806 12708
rect 30926 12656 30932 12708
rect 30984 12656 30990 12708
rect 28718 12628 28724 12640
rect 28368 12600 28724 12628
rect 28718 12588 28724 12600
rect 28776 12588 28782 12640
rect 28810 12588 28816 12640
rect 28868 12588 28874 12640
rect 29086 12588 29092 12640
rect 29144 12628 29150 12640
rect 32858 12628 32864 12640
rect 29144 12600 32864 12628
rect 29144 12588 29150 12600
rect 32858 12588 32864 12600
rect 32916 12588 32922 12640
rect 1104 12538 36524 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 36524 12538
rect 1104 12464 36524 12486
rect 3970 12384 3976 12436
rect 4028 12384 4034 12436
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5442 12424 5448 12436
rect 4764 12396 5448 12424
rect 4764 12384 4770 12396
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 8757 12427 8815 12433
rect 8260 12396 8524 12424
rect 8260 12384 8266 12396
rect 5534 12316 5540 12368
rect 5592 12356 5598 12368
rect 8386 12356 8392 12368
rect 5592 12328 8392 12356
rect 5592 12316 5598 12328
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 5445 12291 5503 12297
rect 2464 12260 4568 12288
rect 2464 12248 2470 12260
rect 4540 12232 4568 12260
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 5718 12288 5724 12300
rect 5491 12260 5724 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12288 6883 12291
rect 7006 12288 7012 12300
rect 6871 12260 7012 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7558 12248 7564 12300
rect 7616 12248 7622 12300
rect 8294 12288 8300 12300
rect 7852 12260 8300 12288
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4396 12192 4445 12220
rect 4396 12180 4402 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4522 12180 4528 12232
rect 4580 12180 4586 12232
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12220 4859 12223
rect 5258 12220 5264 12232
rect 4847 12192 5264 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 7576 12220 7604 12248
rect 7852 12229 7880 12260
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 7837 12223 7895 12229
rect 6411 12192 7696 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 4065 12155 4123 12161
rect 4065 12121 4077 12155
rect 4111 12152 4123 12155
rect 4617 12155 4675 12161
rect 4111 12124 4476 12152
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 4448 12096 4476 12124
rect 4617 12121 4629 12155
rect 4663 12152 4675 12155
rect 4706 12152 4712 12164
rect 4663 12124 4712 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 6181 12155 6239 12161
rect 6181 12152 6193 12155
rect 5276 12124 6193 12152
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 4212 12056 4261 12084
rect 4212 12044 4218 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 4430 12044 4436 12096
rect 4488 12044 4494 12096
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 5276 12093 5304 12124
rect 6181 12121 6193 12124
rect 6227 12152 6239 12155
rect 6914 12152 6920 12164
rect 6227 12124 6920 12152
rect 6227 12121 6239 12124
rect 6181 12115 6239 12121
rect 6914 12112 6920 12124
rect 6972 12112 6978 12164
rect 7558 12112 7564 12164
rect 7616 12112 7622 12164
rect 7668 12152 7696 12192
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 7929 12155 7987 12161
rect 7929 12152 7941 12155
rect 7668 12124 7941 12152
rect 7929 12121 7941 12124
rect 7975 12152 7987 12155
rect 8128 12152 8156 12183
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8496 12229 8524 12396
rect 8757 12393 8769 12427
rect 8803 12424 8815 12427
rect 9030 12424 9036 12436
rect 8803 12396 9036 12424
rect 8803 12393 8815 12396
rect 8757 12387 8815 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9456 12396 9536 12424
rect 9456 12384 9462 12396
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9508 12356 9536 12396
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 9916 12396 11008 12424
rect 9916 12384 9922 12396
rect 10980 12368 11008 12396
rect 11164 12396 13093 12424
rect 11164 12368 11192 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12393 13783 12427
rect 13725 12387 13783 12393
rect 14185 12427 14243 12433
rect 14185 12393 14197 12427
rect 14231 12424 14243 12427
rect 14642 12424 14648 12436
rect 14231 12396 14648 12424
rect 14231 12393 14243 12396
rect 14185 12387 14243 12393
rect 9766 12356 9772 12368
rect 8996 12328 9444 12356
rect 9508 12328 9772 12356
rect 8996 12316 9002 12328
rect 9416 12300 9444 12328
rect 9766 12316 9772 12328
rect 9824 12356 9830 12368
rect 10226 12356 10232 12368
rect 9824 12328 10232 12356
rect 9824 12316 9830 12328
rect 10226 12316 10232 12328
rect 10284 12316 10290 12368
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12356 10563 12359
rect 10870 12356 10876 12368
rect 10551 12328 10876 12356
rect 10551 12325 10563 12328
rect 10505 12319 10563 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 10962 12316 10968 12368
rect 11020 12316 11026 12368
rect 11146 12316 11152 12368
rect 11204 12316 11210 12368
rect 12894 12356 12900 12368
rect 11440 12328 12900 12356
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9306 12288 9312 12300
rect 9180 12260 9312 12288
rect 9180 12248 9186 12260
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9456 12260 9597 12288
rect 9456 12248 9462 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12288 9919 12291
rect 10594 12288 10600 12300
rect 9907 12260 10600 12288
rect 9907 12257 9919 12260
rect 9861 12251 9919 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 11330 12288 11336 12300
rect 10704 12260 11336 12288
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8570 12180 8576 12232
rect 8628 12180 8634 12232
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12220 9275 12223
rect 9674 12220 9680 12232
rect 9263 12192 9680 12220
rect 9263 12189 9275 12192
rect 9217 12183 9275 12189
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9950 12180 9956 12232
rect 10008 12180 10014 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10324 12223 10382 12229
rect 10324 12220 10336 12223
rect 10100 12192 10336 12220
rect 10100 12180 10106 12192
rect 10324 12189 10336 12192
rect 10370 12220 10382 12223
rect 10704 12220 10732 12260
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 10370 12192 10732 12220
rect 10781 12223 10839 12229
rect 10370 12189 10382 12192
rect 10324 12183 10382 12189
rect 10781 12189 10793 12223
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 10919 12192 11100 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 7975 12124 8156 12152
rect 8271 12155 8329 12161
rect 7975 12121 7987 12124
rect 7929 12115 7987 12121
rect 8271 12121 8283 12155
rect 8317 12152 8329 12155
rect 8317 12124 9260 12152
rect 8317 12121 8329 12124
rect 8271 12115 8329 12121
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4856 12056 4905 12084
rect 4856 12044 4862 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12053 5319 12087
rect 5261 12047 5319 12053
rect 5350 12044 5356 12096
rect 5408 12044 5414 12096
rect 6546 12044 6552 12096
rect 6604 12044 6610 12096
rect 8110 12044 8116 12096
rect 8168 12084 8174 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8168 12056 8953 12084
rect 8168 12044 8174 12056
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 9232 12084 9260 12124
rect 9306 12112 9312 12164
rect 9364 12152 9370 12164
rect 9490 12152 9496 12164
rect 9364 12124 9496 12152
rect 9364 12112 9370 12124
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 10796 12152 10824 12183
rect 10336 12124 10824 12152
rect 10336 12096 10364 12124
rect 10962 12112 10968 12164
rect 11020 12112 11026 12164
rect 11072 12152 11100 12192
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11238 12180 11244 12232
rect 11296 12180 11302 12232
rect 11440 12152 11468 12328
rect 12894 12316 12900 12328
rect 12952 12316 12958 12368
rect 13446 12356 13452 12368
rect 13004 12328 13452 12356
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 12158 12248 12164 12300
rect 12216 12248 12222 12300
rect 13004 12288 13032 12328
rect 13446 12316 13452 12328
rect 13504 12356 13510 12368
rect 13740 12356 13768 12387
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 14734 12384 14740 12436
rect 14792 12384 14798 12436
rect 15194 12384 15200 12436
rect 15252 12384 15258 12436
rect 15654 12384 15660 12436
rect 15712 12384 15718 12436
rect 16853 12427 16911 12433
rect 16853 12424 16865 12427
rect 15764 12396 16865 12424
rect 13504 12328 13768 12356
rect 14553 12359 14611 12365
rect 13504 12316 13510 12328
rect 14553 12325 14565 12359
rect 14599 12356 14611 12359
rect 14829 12359 14887 12365
rect 14829 12356 14841 12359
rect 14599 12328 14841 12356
rect 14599 12325 14611 12328
rect 14553 12319 14611 12325
rect 14829 12325 14841 12328
rect 14875 12356 14887 12359
rect 15764 12356 15792 12396
rect 16853 12393 16865 12396
rect 16899 12393 16911 12427
rect 16853 12387 16911 12393
rect 17310 12384 17316 12436
rect 17368 12384 17374 12436
rect 18046 12384 18052 12436
rect 18104 12384 18110 12436
rect 18509 12427 18567 12433
rect 18509 12393 18521 12427
rect 18555 12424 18567 12427
rect 18690 12424 18696 12436
rect 18555 12396 18696 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 18877 12427 18935 12433
rect 18877 12393 18889 12427
rect 18923 12424 18935 12427
rect 18966 12424 18972 12436
rect 18923 12396 18972 12424
rect 18923 12393 18935 12396
rect 18877 12387 18935 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19242 12384 19248 12436
rect 19300 12384 19306 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 19352 12396 20085 12424
rect 19352 12356 19380 12396
rect 20073 12393 20085 12396
rect 20119 12393 20131 12427
rect 20073 12387 20131 12393
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 20220 12396 20269 12424
rect 20220 12384 20226 12396
rect 20257 12393 20269 12396
rect 20303 12424 20315 12427
rect 20806 12424 20812 12436
rect 20303 12396 20812 12424
rect 20303 12393 20315 12396
rect 20257 12387 20315 12393
rect 20806 12384 20812 12396
rect 20864 12384 20870 12436
rect 21358 12384 21364 12436
rect 21416 12384 21422 12436
rect 22462 12384 22468 12436
rect 22520 12384 22526 12436
rect 23014 12384 23020 12436
rect 23072 12424 23078 12436
rect 23198 12424 23204 12436
rect 23072 12396 23204 12424
rect 23072 12384 23078 12396
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 23382 12384 23388 12436
rect 23440 12424 23446 12436
rect 23658 12424 23664 12436
rect 23440 12396 23664 12424
rect 23440 12384 23446 12396
rect 23658 12384 23664 12396
rect 23716 12384 23722 12436
rect 23750 12384 23756 12436
rect 23808 12424 23814 12436
rect 24302 12424 24308 12436
rect 23808 12396 24308 12424
rect 23808 12384 23814 12396
rect 24302 12384 24308 12396
rect 24360 12384 24366 12436
rect 24394 12384 24400 12436
rect 24452 12384 24458 12436
rect 26142 12384 26148 12436
rect 26200 12424 26206 12436
rect 27341 12427 27399 12433
rect 27341 12424 27353 12427
rect 26200 12396 27353 12424
rect 26200 12384 26206 12396
rect 27341 12393 27353 12396
rect 27387 12393 27399 12427
rect 27341 12387 27399 12393
rect 28442 12384 28448 12436
rect 28500 12424 28506 12436
rect 28718 12424 28724 12436
rect 28500 12396 28724 12424
rect 28500 12384 28506 12396
rect 28718 12384 28724 12396
rect 28776 12384 28782 12436
rect 32214 12384 32220 12436
rect 32272 12424 32278 12436
rect 32493 12427 32551 12433
rect 32493 12424 32505 12427
rect 32272 12396 32505 12424
rect 32272 12384 32278 12396
rect 32493 12393 32505 12396
rect 32539 12424 32551 12427
rect 32539 12396 33088 12424
rect 32539 12393 32551 12396
rect 32493 12387 32551 12393
rect 14875 12328 15792 12356
rect 16315 12328 19380 12356
rect 19521 12359 19579 12365
rect 14875 12325 14887 12328
rect 14829 12319 14887 12325
rect 15381 12291 15439 12297
rect 12820 12260 13032 12288
rect 13280 12260 14688 12288
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 11698 12220 11704 12232
rect 11563 12192 11704 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 11882 12220 11888 12232
rect 11839 12192 11888 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 11974 12180 11980 12232
rect 12032 12180 12038 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 12434 12220 12440 12232
rect 12391 12192 12440 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 12820 12229 12848 12260
rect 13280 12229 13308 12260
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 12805 12183 12863 12189
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13814 12220 13820 12232
rect 13495 12192 13820 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 11992 12152 12020 12180
rect 12897 12155 12955 12161
rect 12897 12152 12909 12155
rect 11072 12124 11468 12152
rect 11624 12124 12909 12152
rect 9766 12084 9772 12096
rect 9232 12056 9772 12084
rect 8941 12047 8999 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10318 12044 10324 12096
rect 10376 12044 10382 12096
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 10597 12087 10655 12093
rect 10597 12084 10609 12087
rect 10560 12056 10609 12084
rect 10560 12044 10566 12056
rect 10597 12053 10609 12056
rect 10643 12053 10655 12087
rect 10597 12047 10655 12053
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 11624 12084 11652 12124
rect 12897 12121 12909 12124
rect 12943 12121 12955 12155
rect 13004 12152 13032 12183
rect 13814 12180 13820 12192
rect 13872 12180 13878 12232
rect 13998 12180 14004 12232
rect 14056 12220 14062 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 14056 12192 14105 12220
rect 14056 12180 14062 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 14550 12220 14556 12232
rect 14415 12192 14556 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 13909 12155 13967 12161
rect 13004 12124 13860 12152
rect 12897 12115 12955 12121
rect 10744 12056 11652 12084
rect 10744 12044 10750 12056
rect 11698 12044 11704 12096
rect 11756 12044 11762 12096
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12710 12084 12716 12096
rect 12575 12056 12716 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13538 12044 13544 12096
rect 13596 12044 13602 12096
rect 13722 12093 13728 12096
rect 13709 12087 13728 12093
rect 13709 12053 13721 12087
rect 13709 12047 13728 12053
rect 13722 12044 13728 12047
rect 13780 12044 13786 12096
rect 13832 12084 13860 12124
rect 13909 12121 13921 12155
rect 13955 12152 13967 12155
rect 14384 12152 14412 12183
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 14660 12164 14688 12260
rect 15381 12257 15393 12291
rect 15427 12288 15439 12291
rect 15427 12260 15608 12288
rect 15427 12257 15439 12260
rect 15381 12251 15439 12257
rect 14918 12180 14924 12232
rect 14976 12180 14982 12232
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 15580 12220 15608 12260
rect 16114 12220 16120 12232
rect 15580 12192 16120 12220
rect 16114 12180 16120 12192
rect 16172 12180 16178 12232
rect 16206 12180 16212 12232
rect 16264 12180 16270 12232
rect 13955 12124 14412 12152
rect 13955 12121 13967 12124
rect 13909 12115 13967 12121
rect 14642 12112 14648 12164
rect 14700 12112 14706 12164
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 16315 12152 16343 12328
rect 19521 12325 19533 12359
rect 19567 12356 19579 12359
rect 19702 12356 19708 12368
rect 19567 12328 19708 12356
rect 19567 12325 19579 12328
rect 19521 12319 19579 12325
rect 19702 12316 19708 12328
rect 19760 12316 19766 12368
rect 19794 12316 19800 12368
rect 19852 12356 19858 12368
rect 21082 12356 21088 12368
rect 19852 12328 21088 12356
rect 19852 12316 19858 12328
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 22480 12356 22508 12384
rect 26421 12359 26479 12365
rect 26421 12356 26433 12359
rect 22480 12328 26433 12356
rect 16942 12248 16948 12300
rect 17000 12248 17006 12300
rect 18417 12291 18475 12297
rect 18417 12257 18429 12291
rect 18463 12288 18475 12291
rect 18598 12288 18604 12300
rect 18463 12260 18604 12288
rect 18463 12257 18475 12260
rect 18417 12251 18475 12257
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 19334 12288 19340 12300
rect 19024 12260 19340 12288
rect 19024 12248 19030 12260
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 21177 12291 21235 12297
rect 19444 12260 20560 12288
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 16574 12180 16580 12232
rect 16632 12229 16638 12232
rect 16632 12183 16640 12229
rect 17034 12220 17040 12232
rect 16776 12192 17040 12220
rect 16632 12180 16638 12183
rect 15243 12124 16343 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 15212 12084 15240 12115
rect 16390 12112 16396 12164
rect 16448 12152 16454 12164
rect 16776 12152 16804 12192
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 19444 12229 19472 12260
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 18196 12192 18245 12220
rect 18196 12180 18202 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 19429 12223 19487 12229
rect 18233 12183 18291 12189
rect 18340 12192 18828 12220
rect 16448 12124 16804 12152
rect 16853 12155 16911 12161
rect 16448 12112 16454 12124
rect 16853 12121 16865 12155
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 13832 12056 15240 12084
rect 16761 12087 16819 12093
rect 16761 12053 16773 12087
rect 16807 12084 16819 12087
rect 16868 12084 16896 12115
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 18340 12152 18368 12192
rect 17000 12124 18368 12152
rect 17000 12112 17006 12124
rect 18414 12112 18420 12164
rect 18472 12152 18478 12164
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 18472 12124 18521 12152
rect 18472 12112 18478 12124
rect 18509 12121 18521 12124
rect 18555 12121 18567 12155
rect 18509 12115 18567 12121
rect 16807 12056 16896 12084
rect 16807 12053 16819 12056
rect 16761 12047 16819 12053
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 17920 12056 18705 12084
rect 17920 12044 17926 12056
rect 18693 12053 18705 12056
rect 18739 12053 18751 12087
rect 18800 12084 18828 12192
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 20532 12220 20560 12260
rect 21177 12257 21189 12291
rect 21223 12288 21235 12291
rect 21542 12288 21548 12300
rect 21223 12260 21548 12288
rect 21223 12257 21235 12260
rect 21177 12251 21235 12257
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 21266 12220 21272 12232
rect 19751 12192 20484 12220
rect 20532 12192 21272 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 18874 12161 18880 12164
rect 18861 12155 18880 12161
rect 18861 12121 18873 12155
rect 18861 12115 18880 12121
rect 18874 12112 18880 12115
rect 18932 12112 18938 12164
rect 19061 12155 19119 12161
rect 19061 12121 19073 12155
rect 19107 12152 19119 12155
rect 19150 12152 19156 12164
rect 19107 12124 19156 12152
rect 19107 12121 19119 12124
rect 19061 12115 19119 12121
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 19628 12152 19656 12183
rect 19794 12152 19800 12164
rect 19628 12124 19800 12152
rect 19794 12112 19800 12124
rect 19852 12112 19858 12164
rect 19886 12112 19892 12164
rect 19944 12152 19950 12164
rect 20070 12152 20076 12164
rect 19944 12124 20076 12152
rect 19944 12112 19950 12124
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 20456 12161 20484 12192
rect 21266 12180 21272 12192
rect 21324 12220 21330 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21324 12192 21373 12220
rect 21324 12180 21330 12192
rect 21361 12189 21373 12192
rect 21407 12220 21419 12223
rect 22480 12220 22508 12328
rect 26421 12325 26433 12328
rect 26467 12356 26479 12359
rect 29730 12356 29736 12368
rect 26467 12328 29736 12356
rect 26467 12325 26479 12328
rect 26421 12319 26479 12325
rect 29730 12316 29736 12328
rect 29788 12316 29794 12368
rect 22554 12248 22560 12300
rect 22612 12248 22618 12300
rect 26510 12288 26516 12300
rect 23676 12260 26516 12288
rect 23676 12229 23704 12260
rect 26510 12248 26516 12260
rect 26568 12248 26574 12300
rect 26878 12248 26884 12300
rect 26936 12288 26942 12300
rect 27614 12288 27620 12300
rect 26936 12260 27620 12288
rect 26936 12248 26942 12260
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 28258 12248 28264 12300
rect 28316 12288 28322 12300
rect 28442 12288 28448 12300
rect 28316 12260 28448 12288
rect 28316 12248 28322 12260
rect 28442 12248 28448 12260
rect 28500 12248 28506 12300
rect 28810 12248 28816 12300
rect 28868 12288 28874 12300
rect 33060 12297 33088 12396
rect 33134 12384 33140 12436
rect 33192 12384 33198 12436
rect 29089 12291 29147 12297
rect 29089 12288 29101 12291
rect 28868 12260 29101 12288
rect 28868 12248 28874 12260
rect 29089 12257 29101 12260
rect 29135 12257 29147 12291
rect 29089 12251 29147 12257
rect 33045 12291 33103 12297
rect 33045 12257 33057 12291
rect 33091 12257 33103 12291
rect 33045 12251 33103 12257
rect 21407 12192 22508 12220
rect 23661 12223 23719 12229
rect 21407 12189 21419 12192
rect 21361 12183 21419 12189
rect 23661 12189 23673 12223
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 24026 12180 24032 12232
rect 24084 12180 24090 12232
rect 24302 12180 24308 12232
rect 24360 12220 24366 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24360 12192 24593 12220
rect 24360 12180 24366 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24857 12223 24915 12229
rect 24857 12189 24869 12223
rect 24903 12220 24915 12223
rect 25866 12220 25872 12232
rect 24903 12192 25872 12220
rect 24903 12189 24915 12192
rect 24857 12183 24915 12189
rect 20441 12155 20499 12161
rect 20441 12121 20453 12155
rect 20487 12152 20499 12155
rect 20622 12152 20628 12164
rect 20487 12124 20628 12152
rect 20487 12121 20499 12124
rect 20441 12115 20499 12121
rect 20622 12112 20628 12124
rect 20680 12112 20686 12164
rect 21082 12112 21088 12164
rect 21140 12152 21146 12164
rect 21450 12152 21456 12164
rect 21140 12124 21456 12152
rect 21140 12112 21146 12124
rect 21450 12112 21456 12124
rect 21508 12112 21514 12164
rect 21910 12112 21916 12164
rect 21968 12152 21974 12164
rect 22005 12155 22063 12161
rect 22005 12152 22017 12155
rect 21968 12124 22017 12152
rect 21968 12112 21974 12124
rect 22005 12121 22017 12124
rect 22051 12121 22063 12155
rect 22005 12115 22063 12121
rect 22189 12155 22247 12161
rect 22189 12121 22201 12155
rect 22235 12121 22247 12155
rect 22189 12115 22247 12121
rect 22373 12155 22431 12161
rect 22373 12121 22385 12155
rect 22419 12152 22431 12155
rect 22554 12152 22560 12164
rect 22419 12124 22560 12152
rect 22419 12121 22431 12124
rect 22373 12115 22431 12121
rect 19426 12084 19432 12096
rect 18800 12056 19432 12084
rect 18693 12047 18751 12053
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20241 12087 20299 12093
rect 20241 12053 20253 12087
rect 20287 12084 20299 12087
rect 20714 12084 20720 12096
rect 20287 12056 20720 12084
rect 20287 12053 20299 12056
rect 20241 12047 20299 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 21174 12044 21180 12096
rect 21232 12084 21238 12096
rect 21545 12087 21603 12093
rect 21545 12084 21557 12087
rect 21232 12056 21557 12084
rect 21232 12044 21238 12056
rect 21545 12053 21557 12056
rect 21591 12053 21603 12087
rect 22204 12084 22232 12115
rect 22554 12112 22560 12124
rect 22612 12112 22618 12164
rect 23382 12112 23388 12164
rect 23440 12112 23446 12164
rect 23566 12112 23572 12164
rect 23624 12152 23630 12164
rect 23753 12155 23811 12161
rect 23753 12152 23765 12155
rect 23624 12124 23765 12152
rect 23624 12112 23630 12124
rect 23753 12121 23765 12124
rect 23799 12121 23811 12155
rect 23753 12115 23811 12121
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 23934 12152 23940 12164
rect 23891 12124 23940 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 23934 12112 23940 12124
rect 23992 12112 23998 12164
rect 24394 12112 24400 12164
rect 24452 12152 24458 12164
rect 24872 12152 24900 12183
rect 25866 12180 25872 12192
rect 25924 12180 25930 12232
rect 26421 12223 26479 12229
rect 26421 12220 26433 12223
rect 25976 12192 26433 12220
rect 25976 12152 26004 12192
rect 26421 12189 26433 12192
rect 26467 12189 26479 12223
rect 26421 12183 26479 12189
rect 26602 12180 26608 12232
rect 26660 12180 26666 12232
rect 26786 12180 26792 12232
rect 26844 12220 26850 12232
rect 27065 12223 27123 12229
rect 27065 12220 27077 12223
rect 26844 12192 27077 12220
rect 26844 12180 26850 12192
rect 27065 12189 27077 12192
rect 27111 12189 27123 12223
rect 27065 12183 27123 12189
rect 27154 12180 27160 12232
rect 27212 12180 27218 12232
rect 27338 12180 27344 12232
rect 27396 12180 27402 12232
rect 28902 12180 28908 12232
rect 28960 12180 28966 12232
rect 32122 12180 32128 12232
rect 32180 12220 32186 12232
rect 32217 12223 32275 12229
rect 32217 12220 32229 12223
rect 32180 12192 32229 12220
rect 32180 12180 32186 12192
rect 32217 12189 32229 12192
rect 32263 12189 32275 12223
rect 32217 12183 32275 12189
rect 32401 12223 32459 12229
rect 32401 12189 32413 12223
rect 32447 12189 32459 12223
rect 32401 12183 32459 12189
rect 24452 12124 24900 12152
rect 25240 12124 26004 12152
rect 24452 12112 24458 12124
rect 25240 12096 25268 12124
rect 26326 12112 26332 12164
rect 26384 12152 26390 12164
rect 26620 12152 26648 12180
rect 27172 12152 27200 12180
rect 26384 12124 27200 12152
rect 26384 12112 26390 12124
rect 27614 12112 27620 12164
rect 27672 12152 27678 12164
rect 28074 12152 28080 12164
rect 27672 12124 28080 12152
rect 27672 12112 27678 12124
rect 28074 12112 28080 12124
rect 28132 12112 28138 12164
rect 28258 12112 28264 12164
rect 28316 12152 28322 12164
rect 28353 12155 28411 12161
rect 28353 12152 28365 12155
rect 28316 12124 28365 12152
rect 28316 12112 28322 12124
rect 28353 12121 28365 12124
rect 28399 12121 28411 12155
rect 32416 12152 32444 12183
rect 32490 12180 32496 12232
rect 32548 12220 32554 12232
rect 32674 12220 32680 12232
rect 32548 12192 32680 12220
rect 32548 12180 32554 12192
rect 32674 12180 32680 12192
rect 32732 12180 32738 12232
rect 32950 12180 32956 12232
rect 33008 12180 33014 12232
rect 33229 12223 33287 12229
rect 33229 12189 33241 12223
rect 33275 12220 33287 12223
rect 34514 12220 34520 12232
rect 33275 12192 34520 12220
rect 33275 12189 33287 12192
rect 33229 12183 33287 12189
rect 34514 12180 34520 12192
rect 34572 12180 34578 12232
rect 35250 12152 35256 12164
rect 32416 12124 35256 12152
rect 28353 12115 28411 12121
rect 35250 12112 35256 12124
rect 35308 12112 35314 12164
rect 23014 12084 23020 12096
rect 22204 12056 23020 12084
rect 21545 12047 21603 12053
rect 23014 12044 23020 12056
rect 23072 12084 23078 12096
rect 23477 12087 23535 12093
rect 23477 12084 23489 12087
rect 23072 12056 23489 12084
rect 23072 12044 23078 12056
rect 23477 12053 23489 12056
rect 23523 12053 23535 12087
rect 23477 12047 23535 12053
rect 24765 12087 24823 12093
rect 24765 12053 24777 12087
rect 24811 12084 24823 12087
rect 24854 12084 24860 12096
rect 24811 12056 24860 12084
rect 24811 12053 24823 12056
rect 24765 12047 24823 12053
rect 24854 12044 24860 12056
rect 24912 12084 24918 12096
rect 25038 12084 25044 12096
rect 24912 12056 25044 12084
rect 24912 12044 24918 12056
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 25222 12044 25228 12096
rect 25280 12044 25286 12096
rect 26234 12044 26240 12096
rect 26292 12084 26298 12096
rect 26881 12087 26939 12093
rect 26881 12084 26893 12087
rect 26292 12056 26893 12084
rect 26292 12044 26298 12056
rect 26881 12053 26893 12056
rect 26927 12053 26939 12087
rect 26881 12047 26939 12053
rect 27154 12044 27160 12096
rect 27212 12084 27218 12096
rect 27982 12084 27988 12096
rect 27212 12056 27988 12084
rect 27212 12044 27218 12056
rect 27982 12044 27988 12056
rect 28040 12044 28046 12096
rect 28718 12044 28724 12096
rect 28776 12044 28782 12096
rect 31478 12044 31484 12096
rect 31536 12084 31542 12096
rect 32030 12084 32036 12096
rect 31536 12056 32036 12084
rect 31536 12044 31542 12056
rect 32030 12044 32036 12056
rect 32088 12044 32094 12096
rect 32582 12044 32588 12096
rect 32640 12084 32646 12096
rect 32677 12087 32735 12093
rect 32677 12084 32689 12087
rect 32640 12056 32689 12084
rect 32640 12044 32646 12056
rect 32677 12053 32689 12056
rect 32723 12053 32735 12087
rect 32677 12047 32735 12053
rect 32766 12044 32772 12096
rect 32824 12044 32830 12096
rect 1104 11994 36524 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 36524 11994
rect 1104 11920 36524 11942
rect 4154 11880 4160 11892
rect 3160 11852 4160 11880
rect 3160 11821 3188 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 4617 11883 4675 11889
rect 4617 11880 4629 11883
rect 4580 11852 4629 11880
rect 4580 11840 4586 11852
rect 4617 11849 4629 11852
rect 4663 11849 4675 11883
rect 4617 11843 4675 11849
rect 4706 11840 4712 11892
rect 4764 11840 4770 11892
rect 5169 11883 5227 11889
rect 5169 11849 5181 11883
rect 5215 11880 5227 11883
rect 5258 11880 5264 11892
rect 5215 11852 5264 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 6181 11883 6239 11889
rect 6181 11849 6193 11883
rect 6227 11849 6239 11883
rect 6181 11843 6239 11849
rect 3145 11815 3203 11821
rect 3145 11781 3157 11815
rect 3191 11781 3203 11815
rect 3145 11775 3203 11781
rect 3878 11772 3884 11824
rect 3936 11772 3942 11824
rect 6196 11812 6224 11843
rect 7558 11840 7564 11892
rect 7616 11840 7622 11892
rect 7650 11840 7656 11892
rect 7708 11840 7714 11892
rect 7745 11883 7803 11889
rect 7745 11849 7757 11883
rect 7791 11880 7803 11883
rect 7834 11880 7840 11892
rect 7791 11852 7840 11880
rect 7791 11849 7803 11852
rect 7745 11843 7803 11849
rect 7834 11840 7840 11852
rect 7892 11880 7898 11892
rect 8202 11880 8208 11892
rect 7892 11852 8208 11880
rect 7892 11840 7898 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 9490 11880 9496 11892
rect 8444 11852 9496 11880
rect 8444 11840 8450 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 10008 11852 10701 11880
rect 10008 11840 10014 11852
rect 10689 11849 10701 11852
rect 10735 11880 10747 11883
rect 10778 11880 10784 11892
rect 10735 11852 10784 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11296 11852 11529 11880
rect 11296 11840 11302 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12894 11880 12900 11892
rect 12483 11852 12900 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12894 11840 12900 11852
rect 12952 11880 12958 11892
rect 13170 11880 13176 11892
rect 12952 11852 13176 11880
rect 12952 11840 12958 11852
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 14642 11840 14648 11892
rect 14700 11880 14706 11892
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 14700 11852 14841 11880
rect 14700 11840 14706 11852
rect 14829 11849 14841 11852
rect 14875 11849 14887 11883
rect 16114 11880 16120 11892
rect 14829 11843 14887 11849
rect 15028 11852 16120 11880
rect 4724 11784 5120 11812
rect 2866 11636 2872 11688
rect 2924 11636 2930 11688
rect 4724 11685 4752 11784
rect 4798 11704 4804 11756
rect 4856 11744 4862 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4856 11716 4905 11744
rect 4856 11704 4862 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 4798 11608 4804 11620
rect 4396 11580 4804 11608
rect 4396 11568 4402 11580
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 5000 11608 5028 11707
rect 5092 11676 5120 11784
rect 5736 11784 6224 11812
rect 7285 11815 7343 11821
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5736 11753 5764 11784
rect 7285 11781 7297 11815
rect 7331 11812 7343 11815
rect 7576 11812 7604 11840
rect 12802 11812 12808 11824
rect 7331 11784 9444 11812
rect 7331 11781 7343 11784
rect 7285 11775 7343 11781
rect 5721 11747 5779 11753
rect 5408 11716 5672 11744
rect 5408 11704 5414 11716
rect 5442 11676 5448 11688
rect 5092 11648 5448 11676
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5644 11676 5672 11716
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5828 11676 5856 11707
rect 7466 11704 7472 11756
rect 7524 11744 7530 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7524 11716 7573 11744
rect 7524 11704 7530 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 8202 11704 8208 11756
rect 8260 11704 8266 11756
rect 8389 11747 8447 11753
rect 8389 11713 8401 11747
rect 8435 11744 8447 11747
rect 8662 11744 8668 11756
rect 8435 11716 8668 11744
rect 8435 11713 8447 11716
rect 8389 11707 8447 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9272 11716 9321 11744
rect 9272 11704 9278 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9416 11744 9444 11784
rect 9600 11784 12808 11812
rect 9600 11744 9628 11784
rect 12802 11772 12808 11784
rect 12860 11812 12866 11824
rect 13722 11812 13728 11824
rect 12860 11784 13728 11812
rect 12860 11772 12866 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 9416 11716 9628 11744
rect 9309 11707 9367 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 9732 11716 10333 11744
rect 9732 11704 9738 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10468 11716 10517 11744
rect 10468 11704 10474 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 10962 11704 10968 11756
rect 11020 11704 11026 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11296 11716 11529 11744
rect 11296 11704 11302 11716
rect 11517 11713 11529 11716
rect 11563 11744 11575 11747
rect 12066 11744 12072 11756
rect 11563 11716 12072 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 12308 11716 12357 11744
rect 12308 11704 12314 11716
rect 12345 11713 12357 11716
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11744 12955 11747
rect 12986 11744 12992 11756
rect 12943 11716 12992 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13262 11744 13268 11756
rect 13219 11716 13268 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 5644 11648 5856 11676
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 5810 11608 5816 11620
rect 5000 11580 5816 11608
rect 5810 11568 5816 11580
rect 5868 11608 5874 11620
rect 5920 11608 5948 11639
rect 6454 11636 6460 11688
rect 6512 11636 6518 11688
rect 8481 11679 8539 11685
rect 8481 11645 8493 11679
rect 8527 11645 8539 11679
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 8481 11639 8539 11645
rect 8772 11648 9413 11676
rect 5868 11580 5948 11608
rect 7929 11611 7987 11617
rect 5868 11568 5874 11580
rect 7929 11577 7941 11611
rect 7975 11608 7987 11611
rect 8202 11608 8208 11620
rect 7975 11580 8208 11608
rect 7975 11577 7987 11580
rect 7929 11571 7987 11577
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8496 11552 8524 11639
rect 5445 11543 5503 11549
rect 5445 11509 5457 11543
rect 5491 11540 5503 11543
rect 5534 11540 5540 11552
rect 5491 11512 5540 11540
rect 5491 11509 5503 11512
rect 5445 11503 5503 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5902 11500 5908 11552
rect 5960 11500 5966 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 7282 11540 7288 11552
rect 6236 11512 7288 11540
rect 6236 11500 6242 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7377 11543 7435 11549
rect 7377 11509 7389 11543
rect 7423 11540 7435 11543
rect 7742 11540 7748 11552
rect 7423 11512 7748 11540
rect 7423 11509 7435 11512
rect 7377 11503 7435 11509
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 8021 11543 8079 11549
rect 8021 11509 8033 11543
rect 8067 11540 8079 11543
rect 8478 11540 8484 11552
rect 8067 11512 8484 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8478 11500 8484 11512
rect 8536 11500 8542 11552
rect 8570 11500 8576 11552
rect 8628 11540 8634 11552
rect 8772 11540 8800 11648
rect 9401 11645 9413 11648
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 9490 11636 9496 11688
rect 9548 11636 9554 11688
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9766 11676 9772 11688
rect 9631 11648 9772 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10980 11676 11008 11704
rect 9916 11648 11008 11676
rect 9916 11636 9922 11648
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11793 11679 11851 11685
rect 11112 11648 11652 11676
rect 11112 11636 11118 11648
rect 8849 11611 8907 11617
rect 8849 11577 8861 11611
rect 8895 11608 8907 11611
rect 9306 11608 9312 11620
rect 8895 11580 9312 11608
rect 8895 11577 8907 11580
rect 8849 11571 8907 11577
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 9508 11608 9536 11636
rect 11624 11617 11652 11648
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 11882 11676 11888 11688
rect 11839 11648 11888 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 11882 11636 11888 11648
rect 11940 11636 11946 11688
rect 12268 11676 12296 11704
rect 11992 11648 12296 11676
rect 11609 11611 11667 11617
rect 9508 11580 11192 11608
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 8628 11512 8953 11540
rect 8628 11500 8634 11512
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 8941 11503 8999 11509
rect 9122 11500 9128 11552
rect 9180 11500 9186 11552
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10284 11512 11069 11540
rect 10284 11500 10290 11512
rect 11057 11509 11069 11512
rect 11103 11509 11115 11543
rect 11164 11540 11192 11580
rect 11609 11577 11621 11611
rect 11655 11608 11667 11611
rect 11992 11608 12020 11648
rect 13096 11620 13124 11707
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 14660 11744 14688 11840
rect 15028 11821 15056 11852
rect 16114 11840 16120 11852
rect 16172 11880 16178 11892
rect 25130 11880 25136 11892
rect 16172 11852 25136 11880
rect 16172 11840 16178 11852
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 26786 11840 26792 11892
rect 26844 11880 26850 11892
rect 26970 11880 26976 11892
rect 26844 11852 26976 11880
rect 26844 11840 26850 11852
rect 26970 11840 26976 11852
rect 27028 11880 27034 11892
rect 27341 11883 27399 11889
rect 27341 11880 27353 11883
rect 27028 11852 27353 11880
rect 27028 11840 27034 11852
rect 27341 11849 27353 11852
rect 27387 11849 27399 11883
rect 27341 11843 27399 11849
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 28166 11880 28172 11892
rect 28040 11852 28172 11880
rect 28040 11840 28046 11852
rect 28166 11840 28172 11852
rect 28224 11880 28230 11892
rect 31478 11880 31484 11892
rect 28224 11852 28672 11880
rect 28224 11840 28230 11852
rect 15013 11815 15071 11821
rect 15013 11781 15025 11815
rect 15059 11781 15071 11815
rect 15013 11775 15071 11781
rect 15378 11772 15384 11824
rect 15436 11812 15442 11824
rect 15565 11815 15623 11821
rect 15565 11812 15577 11815
rect 15436 11784 15577 11812
rect 15436 11772 15442 11784
rect 15565 11781 15577 11784
rect 15611 11781 15623 11815
rect 16666 11812 16672 11824
rect 15565 11775 15623 11781
rect 15672 11784 16672 11812
rect 13587 11716 14688 11744
rect 15197 11747 15255 11753
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15672 11744 15700 11784
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 18325 11815 18383 11821
rect 18325 11812 18337 11815
rect 17920 11784 18337 11812
rect 17920 11772 17926 11784
rect 18325 11781 18337 11784
rect 18371 11781 18383 11815
rect 18325 11775 18383 11781
rect 18414 11772 18420 11824
rect 18472 11772 18478 11824
rect 19058 11812 19064 11824
rect 18524 11784 19064 11812
rect 15243 11716 15700 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 13372 11676 13400 11707
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 15804 11716 17908 11744
rect 15804 11704 15810 11716
rect 13814 11676 13820 11688
rect 13372 11648 13820 11676
rect 13814 11636 13820 11648
rect 13872 11676 13878 11688
rect 14734 11676 14740 11688
rect 13872 11648 14740 11676
rect 13872 11636 13878 11648
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 14826 11636 14832 11688
rect 14884 11676 14890 11688
rect 16942 11676 16948 11688
rect 14884 11648 16948 11676
rect 14884 11636 14890 11648
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 11655 11580 12020 11608
rect 11655 11577 11667 11580
rect 11609 11571 11667 11577
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12713 11611 12771 11617
rect 12713 11608 12725 11611
rect 12308 11580 12725 11608
rect 12308 11568 12314 11580
rect 12713 11577 12725 11580
rect 12759 11577 12771 11611
rect 12713 11571 12771 11577
rect 13078 11568 13084 11620
rect 13136 11568 13142 11620
rect 14844 11540 14872 11636
rect 17126 11608 17132 11620
rect 15948 11580 17132 11608
rect 11164 11512 14872 11540
rect 11057 11503 11115 11509
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 15948 11549 15976 11580
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 17880 11608 17908 11716
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18524 11744 18552 11784
rect 19058 11772 19064 11784
rect 19116 11812 19122 11824
rect 19116 11784 19748 11812
rect 19116 11772 19122 11784
rect 18196 11716 18552 11744
rect 18601 11747 18659 11753
rect 18196 11704 18202 11716
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11713 18843 11747
rect 18785 11707 18843 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 19426 11744 19432 11756
rect 18923 11716 19432 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 18046 11636 18052 11688
rect 18104 11676 18110 11688
rect 18506 11676 18512 11688
rect 18104 11648 18512 11676
rect 18104 11636 18110 11648
rect 18506 11636 18512 11648
rect 18564 11676 18570 11688
rect 18616 11676 18644 11707
rect 18564 11648 18644 11676
rect 18800 11676 18828 11707
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 19720 11744 19748 11784
rect 20346 11772 20352 11824
rect 20404 11812 20410 11824
rect 20533 11815 20591 11821
rect 20533 11812 20545 11815
rect 20404 11784 20545 11812
rect 20404 11772 20410 11784
rect 20533 11781 20545 11784
rect 20579 11812 20591 11815
rect 20622 11812 20628 11824
rect 20579 11784 20628 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 20714 11772 20720 11824
rect 20772 11821 20778 11824
rect 20772 11815 20807 11821
rect 20795 11781 20807 11815
rect 20772 11775 20807 11781
rect 23017 11815 23075 11821
rect 23017 11781 23029 11815
rect 23063 11812 23075 11815
rect 23382 11812 23388 11824
rect 23063 11784 23388 11812
rect 23063 11781 23075 11784
rect 23017 11775 23075 11781
rect 20772 11772 20778 11775
rect 23382 11772 23388 11784
rect 23440 11772 23446 11824
rect 23658 11772 23664 11824
rect 23716 11812 23722 11824
rect 23716 11784 24072 11812
rect 23716 11772 23722 11784
rect 19720 11716 20944 11744
rect 19610 11676 19616 11688
rect 18800 11648 19616 11676
rect 18564 11636 18570 11648
rect 19610 11636 19616 11648
rect 19668 11636 19674 11688
rect 20916 11676 20944 11716
rect 21174 11704 21180 11756
rect 21232 11704 21238 11756
rect 21358 11704 21364 11756
rect 21416 11744 21422 11756
rect 21453 11747 21511 11753
rect 21453 11744 21465 11747
rect 21416 11716 21465 11744
rect 21416 11704 21422 11716
rect 21453 11713 21465 11716
rect 21499 11713 21511 11747
rect 21453 11707 21511 11713
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22833 11747 22891 11753
rect 22060 11716 22784 11744
rect 22060 11704 22066 11716
rect 22278 11676 22284 11688
rect 20916 11648 22284 11676
rect 20916 11617 20944 11648
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 22756 11676 22784 11716
rect 22833 11713 22845 11747
rect 22879 11744 22891 11747
rect 23290 11744 23296 11756
rect 22879 11716 23296 11744
rect 22879 11713 22891 11716
rect 22833 11707 22891 11713
rect 23290 11704 23296 11716
rect 23348 11744 23354 11756
rect 24044 11753 24072 11784
rect 24854 11772 24860 11824
rect 24912 11812 24918 11824
rect 25406 11812 25412 11824
rect 24912 11784 25412 11812
rect 24912 11772 24918 11784
rect 25406 11772 25412 11784
rect 25464 11772 25470 11824
rect 26510 11772 26516 11824
rect 26568 11812 26574 11824
rect 28534 11821 28540 11824
rect 28511 11815 28540 11821
rect 26568 11784 28396 11812
rect 26568 11772 26574 11784
rect 23753 11747 23811 11753
rect 23753 11744 23765 11747
rect 23348 11716 23765 11744
rect 23348 11704 23354 11716
rect 23753 11713 23765 11716
rect 23799 11713 23811 11747
rect 23753 11707 23811 11713
rect 24029 11747 24087 11753
rect 24029 11713 24041 11747
rect 24075 11744 24087 11747
rect 24762 11744 24768 11756
rect 24075 11716 24768 11744
rect 24075 11713 24087 11716
rect 24029 11707 24087 11713
rect 24762 11704 24768 11716
rect 24820 11704 24826 11756
rect 24949 11747 25007 11753
rect 24949 11713 24961 11747
rect 24995 11744 25007 11747
rect 25038 11744 25044 11756
rect 24995 11716 25044 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25222 11704 25228 11756
rect 25280 11704 25286 11756
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11744 25835 11747
rect 26142 11744 26148 11756
rect 25823 11716 26148 11744
rect 25823 11713 25835 11716
rect 25777 11707 25835 11713
rect 26142 11704 26148 11716
rect 26200 11704 26206 11756
rect 26697 11747 26755 11753
rect 26697 11713 26709 11747
rect 26743 11744 26755 11747
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26743 11716 26985 11744
rect 26743 11713 26755 11716
rect 26697 11707 26755 11713
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 27338 11744 27344 11756
rect 26973 11707 27031 11713
rect 27080 11716 27344 11744
rect 27080 11688 27108 11716
rect 27338 11704 27344 11716
rect 27396 11744 27402 11756
rect 27617 11747 27675 11753
rect 27617 11744 27629 11747
rect 27396 11716 27629 11744
rect 27396 11704 27402 11716
rect 27617 11713 27629 11716
rect 27663 11713 27675 11747
rect 27617 11707 27675 11713
rect 28258 11704 28264 11756
rect 28316 11704 28322 11756
rect 28368 11744 28396 11784
rect 28511 11781 28523 11815
rect 28511 11775 28540 11781
rect 28534 11772 28540 11775
rect 28592 11772 28598 11824
rect 28644 11821 28672 11852
rect 31312 11852 31484 11880
rect 28629 11815 28687 11821
rect 28629 11781 28641 11815
rect 28675 11781 28687 11815
rect 28629 11775 28687 11781
rect 28721 11815 28779 11821
rect 28721 11781 28733 11815
rect 28767 11812 28779 11815
rect 28902 11812 28908 11824
rect 28767 11784 28908 11812
rect 28767 11781 28779 11784
rect 28721 11775 28779 11781
rect 28902 11772 28908 11784
rect 28960 11772 28966 11824
rect 30926 11772 30932 11824
rect 30984 11812 30990 11824
rect 31312 11821 31340 11852
rect 31478 11840 31484 11852
rect 31536 11840 31542 11892
rect 31665 11883 31723 11889
rect 31665 11849 31677 11883
rect 31711 11880 31723 11883
rect 31711 11852 31800 11880
rect 31711 11849 31723 11852
rect 31665 11843 31723 11849
rect 31297 11815 31355 11821
rect 30984 11784 31157 11812
rect 30984 11772 30990 11784
rect 28368 11716 28488 11744
rect 23842 11676 23848 11688
rect 22756 11648 23848 11676
rect 23842 11636 23848 11648
rect 23900 11636 23906 11688
rect 24673 11679 24731 11685
rect 24673 11645 24685 11679
rect 24719 11676 24731 11679
rect 25406 11676 25412 11688
rect 24719 11648 25412 11676
rect 24719 11645 24731 11648
rect 24673 11639 24731 11645
rect 25406 11636 25412 11648
rect 25464 11636 25470 11688
rect 25498 11636 25504 11688
rect 25556 11636 25562 11688
rect 27062 11636 27068 11688
rect 27120 11636 27126 11688
rect 27154 11636 27160 11688
rect 27212 11636 27218 11688
rect 27246 11636 27252 11688
rect 27304 11636 27310 11688
rect 27522 11636 27528 11688
rect 27580 11636 27586 11688
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 28353 11679 28411 11685
rect 28353 11676 28365 11679
rect 27856 11648 28365 11676
rect 27856 11636 27862 11648
rect 28353 11645 28365 11648
rect 28399 11645 28411 11679
rect 28460 11676 28488 11716
rect 28810 11704 28816 11756
rect 28868 11704 28874 11756
rect 28997 11747 29055 11753
rect 28997 11713 29009 11747
rect 29043 11744 29055 11747
rect 29089 11747 29147 11753
rect 29089 11744 29101 11747
rect 29043 11716 29101 11744
rect 29043 11713 29055 11716
rect 28997 11707 29055 11713
rect 29089 11713 29101 11716
rect 29135 11713 29147 11747
rect 29089 11707 29147 11713
rect 29181 11747 29239 11753
rect 29181 11713 29193 11747
rect 29227 11744 29239 11747
rect 30282 11744 30288 11756
rect 29227 11716 30288 11744
rect 29227 11713 29239 11716
rect 29181 11707 29239 11713
rect 30282 11704 30288 11716
rect 30340 11704 30346 11756
rect 30558 11704 30564 11756
rect 30616 11744 30622 11756
rect 31129 11753 31157 11784
rect 31297 11781 31309 11815
rect 31343 11781 31355 11815
rect 31772 11812 31800 11852
rect 32030 11840 32036 11892
rect 32088 11880 32094 11892
rect 33686 11880 33692 11892
rect 32088 11852 33692 11880
rect 32088 11840 32094 11852
rect 33686 11840 33692 11852
rect 33744 11840 33750 11892
rect 35250 11840 35256 11892
rect 35308 11880 35314 11892
rect 35345 11883 35403 11889
rect 35345 11880 35357 11883
rect 35308 11852 35357 11880
rect 35308 11840 35314 11852
rect 35345 11849 35357 11852
rect 35391 11849 35403 11883
rect 35345 11843 35403 11849
rect 32309 11815 32367 11821
rect 32309 11812 32321 11815
rect 31772 11784 32321 11812
rect 31297 11775 31355 11781
rect 32309 11781 32321 11784
rect 32355 11781 32367 11815
rect 34422 11812 34428 11824
rect 32309 11775 32367 11781
rect 33152 11784 34428 11812
rect 31021 11747 31079 11753
rect 31021 11744 31033 11747
rect 30616 11716 31033 11744
rect 30616 11704 30622 11716
rect 31021 11713 31033 11716
rect 31067 11713 31079 11747
rect 31021 11707 31079 11713
rect 31114 11747 31172 11753
rect 31114 11713 31126 11747
rect 31160 11713 31172 11747
rect 31114 11707 31172 11713
rect 31202 11704 31208 11756
rect 31260 11744 31266 11756
rect 31389 11747 31447 11753
rect 31389 11744 31401 11747
rect 31260 11716 31401 11744
rect 31260 11704 31266 11716
rect 31389 11713 31401 11716
rect 31435 11713 31447 11747
rect 31389 11707 31447 11713
rect 31527 11747 31585 11753
rect 31527 11713 31539 11747
rect 31573 11744 31585 11747
rect 31754 11744 31760 11756
rect 31573 11716 31760 11744
rect 31573 11713 31585 11716
rect 31527 11707 31585 11713
rect 31754 11704 31760 11716
rect 31812 11704 31818 11756
rect 33152 11753 33180 11784
rect 34422 11772 34428 11784
rect 34480 11772 34486 11824
rect 34882 11772 34888 11824
rect 34940 11772 34946 11824
rect 33318 11753 33324 11756
rect 32585 11747 32643 11753
rect 32585 11713 32597 11747
rect 32631 11744 32643 11747
rect 33137 11747 33195 11753
rect 32631 11716 33088 11744
rect 32631 11713 32643 11716
rect 32585 11707 32643 11713
rect 29546 11676 29552 11688
rect 28460 11648 29552 11676
rect 28353 11639 28411 11645
rect 29546 11636 29552 11648
rect 29604 11636 29610 11688
rect 32398 11636 32404 11688
rect 32456 11636 32462 11688
rect 33060 11676 33088 11716
rect 33137 11713 33149 11747
rect 33183 11713 33195 11747
rect 33137 11707 33195 11713
rect 33295 11747 33324 11753
rect 33295 11713 33307 11747
rect 33295 11707 33324 11713
rect 33318 11704 33324 11707
rect 33376 11704 33382 11756
rect 33410 11704 33416 11756
rect 33468 11704 33474 11756
rect 33502 11704 33508 11756
rect 33560 11704 33566 11756
rect 33594 11704 33600 11756
rect 33652 11704 33658 11756
rect 33686 11704 33692 11756
rect 33744 11744 33750 11756
rect 33873 11747 33931 11753
rect 33873 11744 33885 11747
rect 33744 11716 33885 11744
rect 33744 11704 33750 11716
rect 33873 11713 33885 11716
rect 33919 11713 33931 11747
rect 33873 11707 33931 11713
rect 33962 11704 33968 11756
rect 34020 11704 34026 11756
rect 34606 11704 34612 11756
rect 34664 11744 34670 11756
rect 35161 11747 35219 11753
rect 35161 11744 35173 11747
rect 34664 11716 35173 11744
rect 34664 11704 34670 11716
rect 35161 11713 35173 11716
rect 35207 11713 35219 11747
rect 35161 11707 35219 11713
rect 33980 11676 34008 11704
rect 33060 11648 34008 11676
rect 34977 11679 35035 11685
rect 34977 11645 34989 11679
rect 35023 11645 35035 11679
rect 34977 11639 35035 11645
rect 20901 11611 20959 11617
rect 17880 11580 20852 11608
rect 15933 11543 15991 11549
rect 15933 11540 15945 11543
rect 15712 11512 15945 11540
rect 15712 11500 15718 11512
rect 15933 11509 15945 11512
rect 15979 11509 15991 11543
rect 15933 11503 15991 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16942 11540 16948 11552
rect 16724 11512 16948 11540
rect 16724 11500 16730 11512
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17957 11543 18015 11549
rect 17957 11509 17969 11543
rect 18003 11540 18015 11543
rect 18506 11540 18512 11552
rect 18003 11512 18512 11540
rect 18003 11509 18015 11512
rect 17957 11503 18015 11509
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 20530 11540 20536 11552
rect 19392 11512 20536 11540
rect 19392 11500 19398 11512
rect 20530 11500 20536 11512
rect 20588 11540 20594 11552
rect 20714 11540 20720 11552
rect 20588 11512 20720 11540
rect 20588 11500 20594 11512
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 20824 11540 20852 11580
rect 20901 11577 20913 11611
rect 20947 11577 20959 11611
rect 24765 11611 24823 11617
rect 24765 11608 24777 11611
rect 20901 11571 20959 11577
rect 21008 11580 24777 11608
rect 21008 11540 21036 11580
rect 24765 11577 24777 11580
rect 24811 11577 24823 11611
rect 24765 11571 24823 11577
rect 25774 11568 25780 11620
rect 25832 11608 25838 11620
rect 26053 11611 26111 11617
rect 26053 11608 26065 11611
rect 25832 11580 26065 11608
rect 25832 11568 25838 11580
rect 26053 11577 26065 11580
rect 26099 11577 26111 11611
rect 26053 11571 26111 11577
rect 27614 11568 27620 11620
rect 27672 11608 27678 11620
rect 29270 11608 29276 11620
rect 27672 11580 29276 11608
rect 27672 11568 27678 11580
rect 29270 11568 29276 11580
rect 29328 11568 29334 11620
rect 29457 11611 29515 11617
rect 29457 11577 29469 11611
rect 29503 11608 29515 11611
rect 34330 11608 34336 11620
rect 29503 11580 34336 11608
rect 29503 11577 29515 11580
rect 29457 11571 29515 11577
rect 34330 11568 34336 11580
rect 34388 11568 34394 11620
rect 34606 11568 34612 11620
rect 34664 11608 34670 11620
rect 34992 11608 35020 11639
rect 34664 11580 35020 11608
rect 34664 11568 34670 11580
rect 20824 11512 21036 11540
rect 21266 11500 21272 11552
rect 21324 11500 21330 11552
rect 21637 11543 21695 11549
rect 21637 11509 21649 11543
rect 21683 11540 21695 11543
rect 22462 11540 22468 11552
rect 21683 11512 22468 11540
rect 21683 11509 21695 11512
rect 21637 11503 21695 11509
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 23842 11500 23848 11552
rect 23900 11540 23906 11552
rect 24213 11543 24271 11549
rect 24213 11540 24225 11543
rect 23900 11512 24225 11540
rect 23900 11500 23906 11512
rect 24213 11509 24225 11512
rect 24259 11540 24271 11543
rect 24486 11540 24492 11552
rect 24259 11512 24492 11540
rect 24259 11509 24271 11512
rect 24213 11503 24271 11509
rect 24486 11500 24492 11512
rect 24544 11500 24550 11552
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 28442 11540 28448 11552
rect 24636 11512 28448 11540
rect 24636 11500 24642 11512
rect 28442 11500 28448 11512
rect 28500 11500 28506 11552
rect 29178 11500 29184 11552
rect 29236 11500 29242 11552
rect 32490 11500 32496 11552
rect 32548 11500 32554 11552
rect 32674 11500 32680 11552
rect 32732 11540 32738 11552
rect 32769 11543 32827 11549
rect 32769 11540 32781 11543
rect 32732 11512 32781 11540
rect 32732 11500 32738 11512
rect 32769 11509 32781 11512
rect 32815 11509 32827 11543
rect 32769 11503 32827 11509
rect 33778 11500 33784 11552
rect 33836 11500 33842 11552
rect 33870 11500 33876 11552
rect 33928 11500 33934 11552
rect 33962 11500 33968 11552
rect 34020 11540 34026 11552
rect 34241 11543 34299 11549
rect 34241 11540 34253 11543
rect 34020 11512 34253 11540
rect 34020 11500 34026 11512
rect 34241 11509 34253 11512
rect 34287 11509 34299 11543
rect 34348 11540 34376 11568
rect 34885 11543 34943 11549
rect 34885 11540 34897 11543
rect 34348 11512 34897 11540
rect 34241 11503 34299 11509
rect 34885 11509 34897 11512
rect 34931 11509 34943 11543
rect 34885 11503 34943 11509
rect 1104 11450 36524 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 36524 11450
rect 1104 11376 36524 11398
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5350 11336 5356 11348
rect 5307 11308 5356 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 5810 11296 5816 11348
rect 5868 11296 5874 11348
rect 6270 11336 6276 11348
rect 5920 11308 6276 11336
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 5920 11268 5948 11308
rect 6270 11296 6276 11308
rect 6328 11336 6334 11348
rect 7469 11339 7527 11345
rect 6328 11308 7420 11336
rect 6328 11296 6334 11308
rect 5500 11240 5948 11268
rect 5500 11228 5506 11240
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 7285 11271 7343 11277
rect 7285 11268 7297 11271
rect 6696 11240 7297 11268
rect 6696 11228 6702 11240
rect 7285 11237 7297 11240
rect 7331 11237 7343 11271
rect 7392 11268 7420 11308
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 7650 11336 7656 11348
rect 7515 11308 7656 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 11146 11336 11152 11348
rect 7760 11308 11152 11336
rect 7760 11268 7788 11308
rect 11146 11296 11152 11308
rect 11204 11336 11210 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 11204 11308 12541 11336
rect 11204 11296 11210 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 12529 11299 12587 11305
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 17954 11336 17960 11348
rect 13504 11308 17960 11336
rect 13504 11296 13510 11308
rect 17954 11296 17960 11308
rect 18012 11296 18018 11348
rect 18138 11296 18144 11348
rect 18196 11296 18202 11348
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 19058 11336 19064 11348
rect 18288 11308 19064 11336
rect 18288 11296 18294 11308
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 19242 11296 19248 11348
rect 19300 11296 19306 11348
rect 19886 11336 19892 11348
rect 19444 11308 19892 11336
rect 9122 11268 9128 11280
rect 7392 11240 7788 11268
rect 8220 11240 9128 11268
rect 7285 11231 7343 11237
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5092 11172 6193 11200
rect 5092 11141 5120 11172
rect 6181 11169 6193 11172
rect 6227 11200 6239 11203
rect 6914 11200 6920 11212
rect 6227 11172 6920 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 6972 11172 7696 11200
rect 6972 11160 6978 11172
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5261 11135 5319 11141
rect 5261 11101 5273 11135
rect 5307 11132 5319 11135
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5307 11104 6009 11132
rect 5307 11101 5319 11104
rect 5261 11095 5319 11101
rect 5997 11101 6009 11104
rect 6043 11132 6055 11135
rect 6086 11132 6092 11144
rect 6043 11104 6092 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6365 11135 6423 11141
rect 6365 11101 6377 11135
rect 6411 11132 6423 11135
rect 6454 11132 6460 11144
rect 6411 11104 6460 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 5626 11064 5632 11076
rect 4120 11036 5632 11064
rect 4120 11024 4126 11036
rect 5626 11024 5632 11036
rect 5684 11064 5690 11076
rect 6380 11064 6408 11095
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 7466 11073 7472 11076
rect 5684 11036 6408 11064
rect 7453 11067 7472 11073
rect 5684 11024 5690 11036
rect 7453 11033 7465 11067
rect 7453 11027 7472 11033
rect 7466 11024 7472 11027
rect 7524 11024 7530 11076
rect 7668 11073 7696 11172
rect 8110 11092 8116 11144
rect 8168 11092 8174 11144
rect 8220 11141 8248 11240
rect 9122 11228 9128 11240
rect 9180 11228 9186 11280
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 13538 11268 13544 11280
rect 9456 11240 13544 11268
rect 9456 11228 9462 11240
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 15470 11228 15476 11280
rect 15528 11268 15534 11280
rect 15838 11268 15844 11280
rect 15528 11240 15844 11268
rect 15528 11228 15534 11240
rect 15838 11228 15844 11240
rect 15896 11268 15902 11280
rect 19444 11268 19472 11308
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20533 11339 20591 11345
rect 20036 11308 20484 11336
rect 20036 11296 20042 11308
rect 15896 11240 19472 11268
rect 19521 11271 19579 11277
rect 15896 11228 15902 11240
rect 19521 11237 19533 11271
rect 19567 11268 19579 11271
rect 19702 11268 19708 11280
rect 19567 11240 19708 11268
rect 19567 11237 19579 11240
rect 19521 11231 19579 11237
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 20162 11228 20168 11280
rect 20220 11268 20226 11280
rect 20346 11268 20352 11280
rect 20220 11240 20352 11268
rect 20220 11228 20226 11240
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 10134 11200 10140 11212
rect 8435 11172 10140 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 13078 11200 13084 11212
rect 12728 11172 13084 11200
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 12250 11132 12256 11144
rect 9364 11104 12256 11132
rect 9364 11092 9370 11104
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12728 11141 12756 11172
rect 13078 11160 13084 11172
rect 13136 11200 13142 11212
rect 13446 11200 13452 11212
rect 13136 11172 13452 11200
rect 13136 11160 13142 11172
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 16850 11200 16856 11212
rect 16408 11172 16856 11200
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 12894 11132 12900 11144
rect 12851 11104 12900 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 7653 11067 7711 11073
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 7834 11064 7840 11076
rect 7699 11036 7840 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 7926 11024 7932 11076
rect 7984 11024 7990 11076
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 12544 11064 12572 11095
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 12986 11092 12992 11144
rect 13044 11092 13050 11144
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16408 11141 16436 11172
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11200 17555 11203
rect 17543 11172 18368 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 18340 11144 18368 11172
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 20456 11209 20484 11308
rect 20533 11305 20545 11339
rect 20579 11336 20591 11339
rect 20714 11336 20720 11348
rect 20579 11308 20720 11336
rect 20579 11305 20591 11308
rect 20533 11299 20591 11305
rect 20714 11296 20720 11308
rect 20772 11336 20778 11348
rect 21266 11336 21272 11348
rect 20772 11308 21272 11336
rect 20772 11296 20778 11308
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 21450 11296 21456 11348
rect 21508 11296 21514 11348
rect 21542 11296 21548 11348
rect 21600 11336 21606 11348
rect 22278 11336 22284 11348
rect 21600 11308 22284 11336
rect 21600 11296 21606 11308
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22465 11339 22523 11345
rect 22465 11305 22477 11339
rect 22511 11305 22523 11339
rect 22465 11299 22523 11305
rect 22649 11339 22707 11345
rect 22649 11305 22661 11339
rect 22695 11336 22707 11339
rect 22830 11336 22836 11348
rect 22695 11308 22836 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 20806 11228 20812 11280
rect 20864 11228 20870 11280
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 22002 11268 22008 11280
rect 21232 11240 22008 11268
rect 21232 11228 21238 11240
rect 22002 11228 22008 11240
rect 22060 11268 22066 11280
rect 22097 11271 22155 11277
rect 22097 11268 22109 11271
rect 22060 11240 22109 11268
rect 22060 11228 22066 11240
rect 22097 11237 22109 11240
rect 22143 11237 22155 11271
rect 22480 11268 22508 11299
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23014 11296 23020 11348
rect 23072 11296 23078 11348
rect 23109 11339 23167 11345
rect 23109 11305 23121 11339
rect 23155 11336 23167 11339
rect 23658 11336 23664 11348
rect 23155 11308 23664 11336
rect 23155 11305 23167 11308
rect 23109 11299 23167 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24210 11296 24216 11348
rect 24268 11336 24274 11348
rect 24765 11339 24823 11345
rect 24765 11336 24777 11339
rect 24268 11308 24777 11336
rect 24268 11296 24274 11308
rect 24765 11305 24777 11308
rect 24811 11336 24823 11339
rect 24854 11336 24860 11348
rect 24811 11308 24860 11336
rect 24811 11305 24823 11308
rect 24765 11299 24823 11305
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25130 11296 25136 11348
rect 25188 11296 25194 11348
rect 25406 11336 25412 11348
rect 25240 11308 25412 11336
rect 23382 11268 23388 11280
rect 22480 11240 23388 11268
rect 22097 11231 22155 11237
rect 23382 11228 23388 11240
rect 23440 11228 23446 11280
rect 25240 11277 25268 11308
rect 25406 11296 25412 11308
rect 25464 11336 25470 11348
rect 27154 11336 27160 11348
rect 25464 11308 27160 11336
rect 25464 11296 25470 11308
rect 27154 11296 27160 11308
rect 27212 11336 27218 11348
rect 27890 11336 27896 11348
rect 27212 11308 27896 11336
rect 27212 11296 27218 11308
rect 27890 11296 27896 11308
rect 27948 11296 27954 11348
rect 28534 11296 28540 11348
rect 28592 11336 28598 11348
rect 28994 11336 29000 11348
rect 28592 11308 29000 11336
rect 28592 11296 28598 11308
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 29178 11296 29184 11348
rect 29236 11336 29242 11348
rect 29236 11308 30328 11336
rect 29236 11296 29242 11308
rect 25225 11271 25283 11277
rect 25225 11237 25237 11271
rect 25271 11237 25283 11271
rect 25866 11268 25872 11280
rect 25225 11231 25283 11237
rect 25700 11240 25872 11268
rect 19613 11203 19671 11209
rect 19392 11172 19564 11200
rect 19392 11160 19398 11172
rect 16300 11135 16358 11141
rect 16300 11132 16312 11135
rect 16264 11104 16312 11132
rect 16264 11092 16270 11104
rect 16300 11101 16312 11104
rect 16346 11101 16358 11135
rect 16300 11095 16358 11101
rect 16393 11135 16451 11141
rect 16393 11101 16405 11135
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16482 11092 16488 11144
rect 16540 11092 16546 11144
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11132 16727 11135
rect 16758 11132 16764 11144
rect 16715 11104 16764 11132
rect 16715 11101 16727 11104
rect 16669 11095 16727 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 17092 11104 17141 11132
rect 17092 11092 17098 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17129 11095 17187 11101
rect 9456 11036 11100 11064
rect 12544 11036 13032 11064
rect 9456 11024 9462 11036
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 9674 10996 9680 11008
rect 5960 10968 9680 10996
rect 5960 10956 5966 10968
rect 9674 10956 9680 10968
rect 9732 10996 9738 11008
rect 10962 10996 10968 11008
rect 9732 10968 10968 10996
rect 9732 10956 9738 10968
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 11072 10996 11100 11036
rect 12618 10996 12624 11008
rect 11072 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 13004 11005 13032 11036
rect 15378 11024 15384 11076
rect 15436 11064 15442 11076
rect 16025 11067 16083 11073
rect 16025 11064 16037 11067
rect 15436 11036 16037 11064
rect 15436 11024 15442 11036
rect 16025 11033 16037 11036
rect 16071 11033 16083 11067
rect 17144 11064 17172 11095
rect 17310 11092 17316 11144
rect 17368 11092 17374 11144
rect 18046 11092 18052 11144
rect 18104 11092 18110 11144
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18156 11064 18184 11095
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 19536 11132 19564 11172
rect 19613 11169 19625 11203
rect 19659 11200 19671 11203
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 19659 11172 19993 11200
rect 19659 11169 19671 11172
rect 19613 11163 19671 11169
rect 19981 11169 19993 11172
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 20441 11203 20499 11209
rect 20441 11169 20453 11203
rect 20487 11200 20499 11203
rect 20530 11200 20536 11212
rect 20487 11172 20536 11200
rect 20487 11169 20499 11172
rect 20441 11163 20499 11169
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19536 11104 19717 11132
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19886 11132 19892 11144
rect 19705 11095 19763 11101
rect 19801 11104 19892 11132
rect 18782 11064 18788 11076
rect 17144 11036 18092 11064
rect 18156 11036 18788 11064
rect 16025 11027 16083 11033
rect 12989 10999 13047 11005
rect 12989 10965 13001 10999
rect 13035 10996 13047 10999
rect 13262 10996 13268 11008
rect 13035 10968 13268 10996
rect 13035 10965 13047 10968
rect 12989 10959 13047 10965
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 14918 10956 14924 11008
rect 14976 10996 14982 11008
rect 17770 10996 17776 11008
rect 14976 10968 17776 10996
rect 14976 10956 14982 10968
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 17862 10956 17868 11008
rect 17920 10956 17926 11008
rect 18064 10996 18092 11036
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 19801 11064 19829 11104
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 20128 11104 20177 11132
rect 20128 11092 20134 11104
rect 20165 11101 20177 11104
rect 20211 11132 20223 11135
rect 20622 11132 20628 11144
rect 20211 11104 20628 11132
rect 20211 11101 20223 11104
rect 20165 11095 20223 11101
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 20824 11141 20852 11228
rect 20898 11160 20904 11212
rect 20956 11160 20962 11212
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 22830 11200 22836 11212
rect 22419 11172 22836 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 23566 11200 23572 11212
rect 23124 11172 23572 11200
rect 20809 11135 20867 11141
rect 20809 11101 20821 11135
rect 20855 11101 20867 11135
rect 20916 11132 20944 11160
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 20916 11104 21189 11132
rect 20809 11095 20867 11101
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11132 21327 11135
rect 21358 11132 21364 11144
rect 21315 11104 21364 11132
rect 21315 11101 21327 11104
rect 21269 11095 21327 11101
rect 19668 11036 19829 11064
rect 19668 11024 19674 11036
rect 20898 11024 20904 11076
rect 20956 11073 20962 11076
rect 20956 11067 21005 11073
rect 20956 11033 20959 11067
rect 20993 11033 21005 11067
rect 20956 11027 21005 11033
rect 21085 11067 21143 11073
rect 21085 11033 21097 11067
rect 21131 11033 21143 11067
rect 21192 11064 21220 11095
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 21542 11092 21548 11144
rect 21600 11092 21606 11144
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 21775 11104 22048 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 21913 11067 21971 11073
rect 21913 11064 21925 11067
rect 21192 11036 21925 11064
rect 21085 11027 21143 11033
rect 21913 11033 21925 11036
rect 21959 11033 21971 11067
rect 22020 11064 22048 11104
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22462 11092 22468 11144
rect 22520 11092 22526 11144
rect 23124 11132 23152 11172
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 25038 11160 25044 11212
rect 25096 11200 25102 11212
rect 25409 11203 25467 11209
rect 25409 11200 25421 11203
rect 25096 11172 25421 11200
rect 25096 11160 25102 11172
rect 25409 11169 25421 11172
rect 25455 11169 25467 11203
rect 25409 11163 25467 11169
rect 25590 11160 25596 11212
rect 25648 11160 25654 11212
rect 22848 11104 23152 11132
rect 23201 11135 23259 11141
rect 22278 11064 22284 11076
rect 22020 11036 22284 11064
rect 21913 11027 21971 11033
rect 20956 11024 20962 11027
rect 19628 10996 19656 11024
rect 18064 10968 19656 10996
rect 21100 10996 21128 11027
rect 21542 10996 21548 11008
rect 21100 10968 21548 10996
rect 21542 10956 21548 10968
rect 21600 10956 21606 11008
rect 21634 10956 21640 11008
rect 21692 10996 21698 11008
rect 21821 10999 21879 11005
rect 21821 10996 21833 10999
rect 21692 10968 21833 10996
rect 21692 10956 21698 10968
rect 21821 10965 21833 10968
rect 21867 10965 21879 10999
rect 21928 10996 21956 11027
rect 22278 11024 22284 11036
rect 22336 11024 22342 11076
rect 22738 11024 22744 11076
rect 22796 11024 22802 11076
rect 22646 10996 22652 11008
rect 21928 10968 22652 10996
rect 21821 10959 21879 10965
rect 22646 10956 22652 10968
rect 22704 10996 22710 11008
rect 22848 10996 22876 11104
rect 23201 11101 23213 11135
rect 23247 11101 23259 11135
rect 23201 11095 23259 11101
rect 23477 11135 23535 11141
rect 23477 11101 23489 11135
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 22922 11024 22928 11076
rect 22980 11064 22986 11076
rect 23216 11064 23244 11095
rect 22980 11036 23244 11064
rect 23492 11064 23520 11095
rect 24486 11092 24492 11144
rect 24544 11132 24550 11144
rect 24949 11135 25007 11141
rect 24949 11132 24961 11135
rect 24544 11104 24961 11132
rect 24544 11092 24550 11104
rect 24949 11101 24961 11104
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11132 25191 11135
rect 25608 11132 25636 11160
rect 25700 11141 25728 11240
rect 25866 11228 25872 11240
rect 25924 11228 25930 11280
rect 28810 11268 28816 11280
rect 28552 11240 28816 11268
rect 25792 11172 28304 11200
rect 25179 11104 25636 11132
rect 25685 11135 25743 11141
rect 25179 11101 25191 11104
rect 25133 11095 25191 11101
rect 25685 11101 25697 11135
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 23566 11064 23572 11076
rect 23492 11036 23572 11064
rect 22980 11024 22986 11036
rect 23124 11008 23152 11036
rect 23566 11024 23572 11036
rect 23624 11064 23630 11076
rect 24578 11064 24584 11076
rect 23624 11036 24584 11064
rect 23624 11024 23630 11036
rect 24578 11024 24584 11036
rect 24636 11024 24642 11076
rect 25590 11024 25596 11076
rect 25648 11064 25654 11076
rect 25792 11073 25820 11172
rect 25869 11135 25927 11141
rect 25869 11101 25881 11135
rect 25915 11101 25927 11135
rect 25869 11095 25927 11101
rect 25777 11067 25835 11073
rect 25777 11064 25789 11067
rect 25648 11036 25789 11064
rect 25648 11024 25654 11036
rect 25777 11033 25789 11036
rect 25823 11033 25835 11067
rect 25777 11027 25835 11033
rect 22704 10968 22876 10996
rect 22704 10956 22710 10968
rect 23106 10956 23112 11008
rect 23164 10956 23170 11008
rect 23385 10999 23443 11005
rect 23385 10965 23397 10999
rect 23431 10996 23443 10999
rect 23842 10996 23848 11008
rect 23431 10968 23848 10996
rect 23431 10965 23443 10968
rect 23385 10959 23443 10965
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 25222 10956 25228 11008
rect 25280 10996 25286 11008
rect 25884 10996 25912 11095
rect 26878 11092 26884 11144
rect 26936 11132 26942 11144
rect 27249 11135 27307 11141
rect 27249 11132 27261 11135
rect 26936 11104 27261 11132
rect 26936 11092 26942 11104
rect 27249 11101 27261 11104
rect 27295 11101 27307 11135
rect 27249 11095 27307 11101
rect 28074 11092 28080 11144
rect 28132 11092 28138 11144
rect 28166 11092 28172 11144
rect 28224 11092 28230 11144
rect 28276 11064 28304 11172
rect 28350 11092 28356 11144
rect 28408 11092 28414 11144
rect 28442 11092 28448 11144
rect 28500 11092 28506 11144
rect 28552 11141 28580 11240
rect 28810 11228 28816 11240
rect 28868 11268 28874 11280
rect 29365 11271 29423 11277
rect 28868 11240 29224 11268
rect 28868 11228 28874 11240
rect 28913 11172 29132 11200
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28626 11092 28632 11144
rect 28684 11132 28690 11144
rect 28813 11135 28871 11141
rect 28813 11132 28825 11135
rect 28684 11104 28825 11132
rect 28684 11092 28690 11104
rect 28813 11101 28825 11104
rect 28859 11101 28871 11135
rect 28813 11095 28871 11101
rect 28913 11064 28941 11172
rect 28994 11092 29000 11144
rect 29052 11092 29058 11144
rect 29104 11141 29132 11172
rect 29196 11144 29224 11240
rect 29365 11237 29377 11271
rect 29411 11237 29423 11271
rect 30300 11268 30328 11308
rect 30374 11296 30380 11348
rect 30432 11296 30438 11348
rect 30561 11339 30619 11345
rect 30561 11305 30573 11339
rect 30607 11305 30619 11339
rect 30561 11299 30619 11305
rect 33505 11339 33563 11345
rect 33505 11305 33517 11339
rect 33551 11336 33563 11339
rect 33686 11336 33692 11348
rect 33551 11308 33692 11336
rect 33551 11305 33563 11308
rect 33505 11299 33563 11305
rect 30576 11268 30604 11299
rect 33686 11296 33692 11308
rect 33744 11296 33750 11348
rect 33778 11296 33784 11348
rect 33836 11296 33842 11348
rect 34330 11268 34336 11280
rect 30300 11240 30604 11268
rect 31726 11240 34336 11268
rect 29365 11231 29423 11237
rect 29089 11135 29147 11141
rect 29089 11101 29101 11135
rect 29135 11101 29147 11135
rect 29089 11095 29147 11101
rect 29178 11092 29184 11144
rect 29236 11092 29242 11144
rect 29380 11132 29408 11231
rect 30374 11160 30380 11212
rect 30432 11200 30438 11212
rect 30653 11203 30711 11209
rect 30653 11200 30665 11203
rect 30432 11172 30665 11200
rect 30432 11160 30438 11172
rect 30653 11169 30665 11172
rect 30699 11169 30711 11203
rect 30653 11163 30711 11169
rect 30558 11132 30564 11144
rect 29380 11104 30564 11132
rect 30558 11092 30564 11104
rect 30616 11092 30622 11144
rect 30837 11135 30895 11141
rect 30837 11101 30849 11135
rect 30883 11132 30895 11135
rect 31726 11132 31754 11240
rect 34330 11228 34336 11240
rect 34388 11228 34394 11280
rect 33873 11203 33931 11209
rect 33873 11169 33885 11203
rect 33919 11200 33931 11203
rect 34606 11200 34612 11212
rect 33919 11172 34612 11200
rect 33919 11169 33931 11172
rect 33873 11163 33931 11169
rect 34606 11160 34612 11172
rect 34664 11160 34670 11212
rect 30883 11104 31754 11132
rect 30883 11101 30895 11104
rect 30837 11095 30895 11101
rect 32674 11092 32680 11144
rect 32732 11092 32738 11144
rect 33686 11092 33692 11144
rect 33744 11092 33750 11144
rect 33965 11135 34023 11141
rect 33965 11101 33977 11135
rect 34011 11132 34023 11135
rect 34790 11132 34796 11144
rect 34011 11104 34796 11132
rect 34011 11101 34023 11104
rect 33965 11095 34023 11101
rect 34790 11092 34796 11104
rect 34848 11092 34854 11144
rect 30650 11064 30656 11076
rect 28276 11036 28941 11064
rect 29104 11036 30656 11064
rect 25280 10968 25912 10996
rect 25280 10956 25286 10968
rect 28442 10956 28448 11008
rect 28500 10996 28506 11008
rect 28626 10996 28632 11008
rect 28500 10968 28632 10996
rect 28500 10956 28506 10968
rect 28626 10956 28632 10968
rect 28684 10956 28690 11008
rect 28721 10999 28779 11005
rect 28721 10965 28733 10999
rect 28767 10996 28779 10999
rect 29104 10996 29132 11036
rect 30650 11024 30656 11036
rect 30708 11064 30714 11076
rect 32309 11067 32367 11073
rect 30708 11036 30880 11064
rect 30708 11024 30714 11036
rect 30852 11008 30880 11036
rect 32309 11033 32321 11067
rect 32355 11064 32367 11067
rect 32398 11064 32404 11076
rect 32355 11036 32404 11064
rect 32355 11033 32367 11036
rect 32309 11027 32367 11033
rect 32398 11024 32404 11036
rect 32456 11024 32462 11076
rect 32493 11067 32551 11073
rect 32493 11033 32505 11067
rect 32539 11064 32551 11067
rect 32950 11064 32956 11076
rect 32539 11036 32956 11064
rect 32539 11033 32551 11036
rect 32493 11027 32551 11033
rect 32950 11024 32956 11036
rect 33008 11024 33014 11076
rect 28767 10968 29132 10996
rect 28767 10965 28779 10968
rect 28721 10959 28779 10965
rect 29178 10956 29184 11008
rect 29236 10996 29242 11008
rect 30098 10996 30104 11008
rect 29236 10968 30104 10996
rect 29236 10956 29242 10968
rect 30098 10956 30104 10968
rect 30156 10956 30162 11008
rect 30834 10956 30840 11008
rect 30892 10956 30898 11008
rect 33226 10956 33232 11008
rect 33284 10996 33290 11008
rect 33502 10996 33508 11008
rect 33284 10968 33508 10996
rect 33284 10956 33290 10968
rect 33502 10956 33508 10968
rect 33560 10956 33566 11008
rect 1104 10906 36524 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 36524 10906
rect 1104 10832 36524 10854
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5994 10792 6000 10804
rect 4856 10764 6000 10792
rect 4856 10752 4862 10764
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6089 10795 6147 10801
rect 6089 10761 6101 10795
rect 6135 10792 6147 10795
rect 7006 10792 7012 10804
rect 6135 10764 7012 10792
rect 6135 10761 6147 10764
rect 6089 10755 6147 10761
rect 5902 10684 5908 10736
rect 5960 10684 5966 10736
rect 6380 10733 6408 10764
rect 7006 10752 7012 10764
rect 7064 10792 7070 10804
rect 7064 10764 7972 10792
rect 7064 10752 7070 10764
rect 6365 10727 6423 10733
rect 6365 10693 6377 10727
rect 6411 10693 6423 10727
rect 7944 10724 7972 10764
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 8260 10764 8401 10792
rect 8260 10752 8266 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 8389 10755 8447 10761
rect 11514 10752 11520 10804
rect 11572 10792 11578 10804
rect 18506 10792 18512 10804
rect 11572 10764 14504 10792
rect 11572 10752 11578 10764
rect 8220 10724 8248 10752
rect 6365 10687 6423 10693
rect 6840 10696 7788 10724
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10656 6239 10659
rect 6546 10656 6552 10668
rect 6227 10628 6552 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6840 10665 6868 10696
rect 7760 10668 7788 10696
rect 7944 10696 8248 10724
rect 10413 10727 10471 10733
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 6748 10588 6776 10619
rect 7006 10616 7012 10668
rect 7064 10616 7070 10668
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 6656 10560 6776 10588
rect 6656 10529 6684 10560
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 7116 10588 7144 10619
rect 7650 10616 7656 10668
rect 7708 10616 7714 10668
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 7944 10665 7972 10696
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 10459 10696 11100 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8297 10659 8355 10665
rect 8297 10656 8309 10659
rect 8076 10628 8309 10656
rect 8076 10616 8082 10628
rect 8297 10625 8309 10628
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8478 10588 8484 10600
rect 6972 10560 7144 10588
rect 6972 10548 6978 10560
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10489 6699 10523
rect 7116 10520 7144 10560
rect 8128 10560 8484 10588
rect 8018 10520 8024 10532
rect 7116 10492 8024 10520
rect 6641 10483 6699 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 5905 10455 5963 10461
rect 5905 10421 5917 10455
rect 5951 10452 5963 10455
rect 7190 10452 7196 10464
rect 5951 10424 7196 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7374 10452 7380 10464
rect 7331 10424 7380 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8128 10452 8156 10560
rect 8478 10548 8484 10560
rect 8536 10588 8542 10600
rect 8588 10588 8616 10619
rect 9674 10616 9680 10668
rect 9732 10616 9738 10668
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 10134 10656 10140 10668
rect 9907 10628 10140 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10226 10616 10232 10668
rect 10284 10616 10290 10668
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 10870 10616 10876 10668
rect 10928 10616 10934 10668
rect 11072 10665 11100 10696
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 14476 10733 14504 10764
rect 15764 10764 18512 10792
rect 14461 10727 14519 10733
rect 11388 10696 13216 10724
rect 11388 10684 11394 10696
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11698 10656 11704 10668
rect 11204 10628 11704 10656
rect 11204 10616 11210 10628
rect 11698 10616 11704 10628
rect 11756 10656 11762 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 11756 10628 12081 10656
rect 11756 10616 11762 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 13188 10665 13216 10696
rect 14461 10693 14473 10727
rect 14507 10693 14519 10727
rect 14461 10687 14519 10693
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 8536 10560 8616 10588
rect 8536 10548 8542 10560
rect 9950 10548 9956 10600
rect 10008 10548 10014 10600
rect 10045 10591 10103 10597
rect 10045 10557 10057 10591
rect 10091 10557 10103 10591
rect 10152 10588 10180 10616
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 10152 10560 11805 10588
rect 10045 10551 10103 10557
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10588 12035 10591
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12023 10560 12541 10588
rect 12023 10557 12035 10560
rect 11977 10551 12035 10557
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 10060 10520 10088 10551
rect 11698 10520 11704 10532
rect 10060 10492 11704 10520
rect 11698 10480 11704 10492
rect 11756 10520 11762 10532
rect 13004 10520 13032 10619
rect 13262 10616 13268 10668
rect 13320 10616 13326 10668
rect 13446 10616 13452 10668
rect 13504 10616 13510 10668
rect 13906 10616 13912 10668
rect 13964 10616 13970 10668
rect 14090 10616 14096 10668
rect 14148 10616 14154 10668
rect 14734 10616 14740 10668
rect 14792 10616 14798 10668
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10656 15163 10659
rect 15565 10659 15623 10665
rect 15151 10628 15516 10656
rect 15151 10625 15163 10628
rect 15105 10619 15163 10625
rect 13464 10588 13492 10616
rect 14001 10591 14059 10597
rect 14001 10588 14013 10591
rect 13464 10560 14013 10588
rect 14001 10557 14013 10560
rect 14047 10557 14059 10591
rect 14001 10551 14059 10557
rect 11756 10492 13032 10520
rect 11756 10480 11762 10492
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 14108 10520 14136 10616
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14752 10588 14780 10616
rect 14240 10560 14780 10588
rect 14240 10548 14246 10560
rect 14642 10520 14648 10532
rect 13412 10492 14648 10520
rect 13412 10480 13418 10492
rect 14642 10480 14648 10492
rect 14700 10480 14706 10532
rect 15488 10520 15516 10628
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15611 10628 15669 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15764 10656 15792 10764
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 19484 10764 21097 10792
rect 19484 10752 19490 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 25590 10792 25596 10804
rect 21085 10755 21143 10761
rect 21192 10764 25596 10792
rect 15841 10727 15899 10733
rect 15841 10693 15853 10727
rect 15887 10724 15899 10727
rect 16574 10724 16580 10736
rect 15887 10696 16580 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 16574 10684 16580 10696
rect 16632 10724 16638 10736
rect 17129 10727 17187 10733
rect 16632 10696 16896 10724
rect 16632 10684 16638 10696
rect 16868 10665 16896 10696
rect 17129 10693 17141 10727
rect 17175 10724 17187 10727
rect 17862 10724 17868 10736
rect 17175 10696 17868 10724
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 17862 10684 17868 10696
rect 17920 10684 17926 10736
rect 17954 10684 17960 10736
rect 18012 10724 18018 10736
rect 21192 10724 21220 10764
rect 25590 10752 25596 10764
rect 25648 10752 25654 10804
rect 27338 10792 27344 10804
rect 25700 10764 27344 10792
rect 18012 10696 21220 10724
rect 21253 10727 21311 10733
rect 18012 10684 18018 10696
rect 21253 10693 21265 10727
rect 21299 10724 21311 10727
rect 21358 10724 21364 10736
rect 21299 10696 21364 10724
rect 21299 10693 21311 10696
rect 21253 10687 21311 10693
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 21453 10727 21511 10733
rect 21453 10693 21465 10727
rect 21499 10724 21511 10727
rect 21542 10724 21548 10736
rect 21499 10696 21548 10724
rect 21499 10693 21511 10696
rect 21453 10687 21511 10693
rect 21542 10684 21548 10696
rect 21600 10684 21606 10736
rect 23842 10684 23848 10736
rect 23900 10684 23906 10736
rect 24305 10727 24363 10733
rect 24305 10693 24317 10727
rect 24351 10724 24363 10727
rect 24486 10724 24492 10736
rect 24351 10696 24492 10724
rect 24351 10693 24363 10696
rect 24305 10687 24363 10693
rect 24486 10684 24492 10696
rect 24544 10684 24550 10736
rect 25700 10724 25728 10764
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 27798 10752 27804 10804
rect 27856 10792 27862 10804
rect 27893 10795 27951 10801
rect 27893 10792 27905 10795
rect 27856 10764 27905 10792
rect 27856 10752 27862 10764
rect 27893 10761 27905 10764
rect 27939 10761 27951 10795
rect 27893 10755 27951 10761
rect 28534 10752 28540 10804
rect 28592 10792 28598 10804
rect 29178 10792 29184 10804
rect 28592 10764 28856 10792
rect 28592 10752 28598 10764
rect 27246 10724 27252 10736
rect 24872 10696 25728 10724
rect 25884 10696 27252 10724
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15764 10628 16037 10656
rect 15657 10619 15715 10625
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17310 10616 17316 10668
rect 17368 10656 17374 10668
rect 19426 10656 19432 10668
rect 17368 10628 19432 10656
rect 17368 10616 17374 10628
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10625 19947 10659
rect 19889 10619 19947 10625
rect 16206 10548 16212 10600
rect 16264 10588 16270 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16264 10560 16957 10588
rect 16264 10548 16270 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 16945 10551 17003 10557
rect 18690 10548 18696 10600
rect 18748 10588 18754 10600
rect 19904 10588 19932 10619
rect 19978 10616 19984 10668
rect 20036 10616 20042 10668
rect 20162 10616 20168 10668
rect 20220 10616 20226 10668
rect 20254 10616 20260 10668
rect 20312 10616 20318 10668
rect 21376 10656 21404 10684
rect 22002 10656 22008 10668
rect 21376 10628 22008 10656
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 23566 10616 23572 10668
rect 23624 10616 23630 10668
rect 23658 10616 23664 10668
rect 23716 10656 23722 10668
rect 23716 10628 23888 10656
rect 23716 10616 23722 10628
rect 22462 10588 22468 10600
rect 18748 10560 22468 10588
rect 18748 10548 18754 10560
rect 22462 10548 22468 10560
rect 22520 10588 22526 10600
rect 22922 10588 22928 10600
rect 22520 10560 22928 10588
rect 22520 10548 22526 10560
rect 22922 10548 22928 10560
rect 22980 10588 22986 10600
rect 23753 10591 23811 10597
rect 23753 10588 23765 10591
rect 22980 10560 23765 10588
rect 22980 10548 22986 10560
rect 23753 10557 23765 10560
rect 23799 10557 23811 10591
rect 23860 10588 23888 10628
rect 24210 10616 24216 10668
rect 24268 10616 24274 10668
rect 24397 10659 24455 10665
rect 24397 10625 24409 10659
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 24762 10656 24768 10668
rect 24627 10628 24768 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 24412 10588 24440 10619
rect 24762 10616 24768 10628
rect 24820 10616 24826 10668
rect 24872 10588 24900 10696
rect 25222 10616 25228 10668
rect 25280 10616 25286 10668
rect 25406 10616 25412 10668
rect 25464 10656 25470 10668
rect 25590 10656 25596 10668
rect 25464 10628 25596 10656
rect 25464 10616 25470 10628
rect 25590 10616 25596 10628
rect 25648 10616 25654 10668
rect 25884 10665 25912 10696
rect 27246 10684 27252 10696
rect 27304 10684 27310 10736
rect 28166 10684 28172 10736
rect 28224 10724 28230 10736
rect 28224 10696 28672 10724
rect 28224 10684 28230 10696
rect 25685 10659 25743 10665
rect 25685 10625 25697 10659
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 25869 10659 25927 10665
rect 25869 10625 25881 10659
rect 25915 10625 25927 10659
rect 25869 10619 25927 10625
rect 25961 10659 26019 10665
rect 25961 10625 25973 10659
rect 26007 10656 26019 10659
rect 26142 10656 26148 10668
rect 26007 10628 26148 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 23860 10560 24900 10588
rect 23753 10551 23811 10557
rect 25314 10548 25320 10600
rect 25372 10588 25378 10600
rect 25501 10591 25559 10597
rect 25501 10588 25513 10591
rect 25372 10560 25513 10588
rect 25372 10548 25378 10560
rect 25501 10557 25513 10560
rect 25547 10557 25559 10591
rect 25700 10588 25728 10619
rect 26142 10616 26148 10628
rect 26200 10616 26206 10668
rect 26234 10616 26240 10668
rect 26292 10616 26298 10668
rect 26329 10659 26387 10665
rect 26329 10625 26341 10659
rect 26375 10656 26387 10659
rect 26418 10656 26424 10668
rect 26375 10628 26424 10656
rect 26375 10625 26387 10628
rect 26329 10619 26387 10625
rect 26418 10616 26424 10628
rect 26476 10616 26482 10668
rect 26694 10616 26700 10668
rect 26752 10616 26758 10668
rect 27062 10616 27068 10668
rect 27120 10656 27126 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 27120 10628 27169 10656
rect 27120 10616 27126 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 27430 10616 27436 10668
rect 27488 10616 27494 10668
rect 27982 10616 27988 10668
rect 28040 10656 28046 10668
rect 28077 10659 28135 10665
rect 28077 10656 28089 10659
rect 28040 10628 28089 10656
rect 28040 10616 28046 10628
rect 28077 10625 28089 10628
rect 28123 10625 28135 10659
rect 28353 10659 28411 10665
rect 28353 10656 28365 10659
rect 28077 10619 28135 10625
rect 28184 10628 28365 10656
rect 27249 10591 27307 10597
rect 25700 10560 26280 10588
rect 25501 10551 25559 10557
rect 26252 10532 26280 10560
rect 27249 10557 27261 10591
rect 27295 10588 27307 10591
rect 27338 10588 27344 10600
rect 27295 10560 27344 10588
rect 27295 10557 27307 10560
rect 27249 10551 27307 10557
rect 27338 10548 27344 10560
rect 27396 10548 27402 10600
rect 27890 10548 27896 10600
rect 27948 10588 27954 10600
rect 28184 10588 28212 10628
rect 28353 10625 28365 10628
rect 28399 10625 28411 10659
rect 28353 10619 28411 10625
rect 28534 10616 28540 10668
rect 28592 10616 28598 10668
rect 28644 10665 28672 10696
rect 28718 10684 28724 10736
rect 28776 10684 28782 10736
rect 28828 10733 28856 10764
rect 29017 10764 29184 10792
rect 28813 10727 28871 10733
rect 28813 10693 28825 10727
rect 28859 10693 28871 10727
rect 28813 10687 28871 10693
rect 28629 10659 28687 10665
rect 28629 10625 28641 10659
rect 28675 10625 28687 10659
rect 28736 10656 28764 10684
rect 29017 10665 29045 10764
rect 29178 10752 29184 10764
rect 29236 10752 29242 10804
rect 29270 10752 29276 10804
rect 29328 10752 29334 10804
rect 32585 10795 32643 10801
rect 32585 10761 32597 10795
rect 32631 10792 32643 10795
rect 33134 10792 33140 10804
rect 32631 10764 33140 10792
rect 32631 10761 32643 10764
rect 32585 10755 32643 10761
rect 33134 10752 33140 10764
rect 33192 10752 33198 10804
rect 34698 10752 34704 10804
rect 34756 10792 34762 10804
rect 35161 10795 35219 10801
rect 35161 10792 35173 10795
rect 34756 10764 35173 10792
rect 34756 10752 34762 10764
rect 35161 10761 35173 10764
rect 35207 10761 35219 10795
rect 35161 10755 35219 10761
rect 31294 10724 31300 10736
rect 30668 10696 31300 10724
rect 28905 10659 28963 10665
rect 28905 10656 28917 10659
rect 28736 10628 28917 10656
rect 28629 10619 28687 10625
rect 28905 10625 28917 10628
rect 28951 10625 28963 10659
rect 29017 10659 29079 10665
rect 29017 10628 29033 10659
rect 28905 10619 28963 10625
rect 29021 10625 29033 10628
rect 29067 10625 29079 10659
rect 29021 10619 29079 10625
rect 29457 10659 29515 10665
rect 29457 10625 29469 10659
rect 29503 10625 29515 10659
rect 29457 10619 29515 10625
rect 29641 10659 29699 10665
rect 29641 10625 29653 10659
rect 29687 10656 29699 10659
rect 29730 10656 29736 10668
rect 29687 10628 29736 10656
rect 29687 10625 29699 10628
rect 29641 10619 29699 10625
rect 27948 10560 28212 10588
rect 28261 10591 28319 10597
rect 27948 10548 27954 10560
rect 28261 10557 28273 10591
rect 28307 10588 28319 10591
rect 28718 10588 28724 10600
rect 28307 10560 28724 10588
rect 28307 10557 28319 10560
rect 28261 10551 28319 10557
rect 28718 10548 28724 10560
rect 28776 10548 28782 10600
rect 29472 10588 29500 10619
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 30668 10656 30696 10696
rect 31294 10684 31300 10696
rect 31352 10684 31358 10736
rect 34330 10684 34336 10736
rect 34388 10684 34394 10736
rect 34517 10727 34575 10733
rect 34517 10693 34529 10727
rect 34563 10724 34575 10727
rect 34790 10724 34796 10736
rect 34563 10696 34796 10724
rect 34563 10693 34575 10696
rect 34517 10687 34575 10693
rect 34790 10684 34796 10696
rect 34848 10724 34854 10736
rect 35621 10727 35679 10733
rect 35621 10724 35633 10727
rect 34848 10696 35633 10724
rect 34848 10684 34854 10696
rect 35621 10693 35633 10696
rect 35667 10693 35679 10727
rect 35621 10687 35679 10693
rect 29972 10628 30696 10656
rect 29972 10616 29978 10628
rect 31018 10616 31024 10668
rect 31076 10656 31082 10668
rect 32125 10659 32183 10665
rect 32125 10656 32137 10659
rect 31076 10628 32137 10656
rect 31076 10616 31082 10628
rect 32125 10625 32137 10628
rect 32171 10625 32183 10659
rect 32125 10619 32183 10625
rect 32401 10659 32459 10665
rect 32401 10625 32413 10659
rect 32447 10656 32459 10659
rect 33686 10656 33692 10668
rect 32447 10628 33692 10656
rect 32447 10625 32459 10628
rect 32401 10619 32459 10625
rect 33686 10616 33692 10628
rect 33744 10616 33750 10668
rect 34606 10616 34612 10668
rect 34664 10656 34670 10668
rect 34701 10659 34759 10665
rect 34701 10656 34713 10659
rect 34664 10628 34713 10656
rect 34664 10616 34670 10628
rect 34701 10625 34713 10628
rect 34747 10625 34759 10659
rect 34701 10619 34759 10625
rect 35345 10659 35403 10665
rect 35345 10625 35357 10659
rect 35391 10625 35403 10659
rect 35345 10619 35403 10625
rect 28920 10560 29500 10588
rect 30024 10560 30328 10588
rect 19705 10523 19763 10529
rect 19705 10520 19717 10523
rect 15488 10492 19717 10520
rect 19705 10489 19717 10492
rect 19751 10489 19763 10523
rect 19705 10483 19763 10489
rect 21450 10480 21456 10532
rect 21508 10520 21514 10532
rect 25225 10523 25283 10529
rect 25225 10520 25237 10523
rect 21508 10492 25237 10520
rect 21508 10480 21514 10492
rect 25225 10489 25237 10492
rect 25271 10520 25283 10523
rect 25406 10520 25412 10532
rect 25271 10492 25412 10520
rect 25271 10489 25283 10492
rect 25225 10483 25283 10489
rect 25406 10480 25412 10492
rect 25464 10480 25470 10532
rect 26234 10480 26240 10532
rect 26292 10480 26298 10532
rect 26421 10523 26479 10529
rect 26421 10489 26433 10523
rect 26467 10520 26479 10523
rect 27798 10520 27804 10532
rect 26467 10492 27804 10520
rect 26467 10489 26479 10492
rect 26421 10483 26479 10489
rect 27798 10480 27804 10492
rect 27856 10480 27862 10532
rect 28074 10480 28080 10532
rect 28132 10520 28138 10532
rect 28132 10492 28304 10520
rect 28132 10480 28138 10492
rect 7708 10424 8156 10452
rect 8205 10455 8263 10461
rect 7708 10412 7714 10424
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 8294 10452 8300 10464
rect 8251 10424 8300 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8573 10455 8631 10461
rect 8573 10421 8585 10455
rect 8619 10452 8631 10455
rect 9674 10452 9680 10464
rect 8619 10424 9680 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 9824 10424 10517 10452
rect 9824 10412 9830 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 12400 10424 12449 10452
rect 12400 10412 12406 10424
rect 12437 10421 12449 10424
rect 12483 10421 12495 10455
rect 12437 10415 12495 10421
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 16669 10455 16727 10461
rect 16669 10421 16681 10455
rect 16715 10452 16727 10455
rect 16758 10452 16764 10464
rect 16715 10424 16764 10452
rect 16715 10421 16727 10424
rect 16669 10415 16727 10421
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 17129 10455 17187 10461
rect 17129 10421 17141 10455
rect 17175 10452 17187 10455
rect 17218 10452 17224 10464
rect 17175 10424 17224 10452
rect 17175 10421 17187 10424
rect 17129 10415 17187 10421
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 22186 10412 22192 10464
rect 22244 10452 22250 10464
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 22244 10424 23397 10452
rect 22244 10412 22250 10424
rect 23385 10421 23397 10424
rect 23431 10421 23443 10455
rect 23385 10415 23443 10421
rect 23845 10455 23903 10461
rect 23845 10421 23857 10455
rect 23891 10452 23903 10455
rect 23934 10452 23940 10464
rect 23891 10424 23940 10452
rect 23891 10421 23903 10424
rect 23845 10415 23903 10421
rect 23934 10412 23940 10424
rect 23992 10412 23998 10464
rect 24029 10455 24087 10461
rect 24029 10421 24041 10455
rect 24075 10452 24087 10455
rect 24394 10452 24400 10464
rect 24075 10424 24400 10452
rect 24075 10421 24087 10424
rect 24029 10415 24087 10421
rect 24394 10412 24400 10424
rect 24452 10412 24458 10464
rect 24578 10412 24584 10464
rect 24636 10452 24642 10464
rect 26513 10455 26571 10461
rect 26513 10452 26525 10455
rect 24636 10424 26525 10452
rect 24636 10412 24642 10424
rect 26513 10421 26525 10424
rect 26559 10452 26571 10455
rect 27154 10452 27160 10464
rect 26559 10424 27160 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 27154 10412 27160 10424
rect 27212 10412 27218 10464
rect 27338 10412 27344 10464
rect 27396 10452 27402 10464
rect 28166 10452 28172 10464
rect 27396 10424 28172 10452
rect 27396 10412 27402 10424
rect 28166 10412 28172 10424
rect 28224 10412 28230 10464
rect 28276 10452 28304 10492
rect 28350 10480 28356 10532
rect 28408 10520 28414 10532
rect 28537 10523 28595 10529
rect 28537 10520 28549 10523
rect 28408 10492 28549 10520
rect 28408 10480 28414 10492
rect 28537 10489 28549 10492
rect 28583 10489 28595 10523
rect 28537 10483 28595 10489
rect 28920 10452 28948 10560
rect 30024 10520 30052 10560
rect 30300 10532 30328 10560
rect 30650 10548 30656 10600
rect 30708 10588 30714 10600
rect 32217 10591 32275 10597
rect 32217 10588 32229 10591
rect 30708 10560 32229 10588
rect 30708 10548 30714 10560
rect 32217 10557 32229 10560
rect 32263 10557 32275 10591
rect 32217 10551 32275 10557
rect 29288 10492 30052 10520
rect 28276 10424 28948 10452
rect 29181 10455 29239 10461
rect 29181 10421 29193 10455
rect 29227 10452 29239 10455
rect 29288 10452 29316 10492
rect 30282 10480 30288 10532
rect 30340 10520 30346 10532
rect 35360 10520 35388 10619
rect 35434 10616 35440 10668
rect 35492 10616 35498 10668
rect 30340 10492 35388 10520
rect 30340 10480 30346 10492
rect 29227 10424 29316 10452
rect 29227 10421 29239 10424
rect 29181 10415 29239 10421
rect 32306 10412 32312 10464
rect 32364 10412 32370 10464
rect 35621 10455 35679 10461
rect 35621 10421 35633 10455
rect 35667 10452 35679 10455
rect 36170 10452 36176 10464
rect 35667 10424 36176 10452
rect 35667 10421 35679 10424
rect 35621 10415 35679 10421
rect 36170 10412 36176 10424
rect 36228 10412 36234 10464
rect 1104 10362 36524 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 36524 10362
rect 1104 10288 36524 10310
rect 6270 10208 6276 10260
rect 6328 10208 6334 10260
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6914 10248 6920 10260
rect 6604 10220 6920 10248
rect 6604 10208 6610 10220
rect 6914 10208 6920 10220
rect 6972 10248 6978 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6972 10220 7021 10248
rect 6972 10208 6978 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 7926 10248 7932 10260
rect 7883 10220 7932 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8754 10248 8760 10260
rect 8619 10220 8760 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 9950 10248 9956 10260
rect 9447 10220 9956 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10686 10248 10692 10260
rect 10091 10220 10692 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11330 10208 11336 10260
rect 11388 10208 11394 10260
rect 16025 10251 16083 10257
rect 16025 10217 16037 10251
rect 16071 10248 16083 10251
rect 16206 10248 16212 10260
rect 16071 10220 16212 10248
rect 16071 10217 16083 10220
rect 16025 10211 16083 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16574 10208 16580 10260
rect 16632 10208 16638 10260
rect 17494 10208 17500 10260
rect 17552 10208 17558 10260
rect 17678 10208 17684 10260
rect 17736 10208 17742 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 17828 10220 19809 10248
rect 17828 10208 17834 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 19797 10211 19855 10217
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20220 10220 20637 10248
rect 20220 10208 20226 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 20809 10251 20867 10257
rect 20809 10248 20821 10251
rect 20772 10220 20821 10248
rect 20772 10208 20778 10220
rect 20809 10217 20821 10220
rect 20855 10217 20867 10251
rect 20809 10211 20867 10217
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22097 10251 22155 10257
rect 22097 10248 22109 10251
rect 21968 10220 22109 10248
rect 21968 10208 21974 10220
rect 22097 10217 22109 10220
rect 22143 10217 22155 10251
rect 22097 10211 22155 10217
rect 22186 10208 22192 10260
rect 22244 10208 22250 10260
rect 22557 10251 22615 10257
rect 22557 10217 22569 10251
rect 22603 10248 22615 10251
rect 22830 10248 22836 10260
rect 22603 10220 22836 10248
rect 22603 10217 22615 10220
rect 22557 10211 22615 10217
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 25406 10208 25412 10260
rect 25464 10248 25470 10260
rect 29089 10251 29147 10257
rect 25464 10220 28856 10248
rect 25464 10208 25470 10220
rect 5537 10183 5595 10189
rect 5537 10149 5549 10183
rect 5583 10180 5595 10183
rect 6086 10180 6092 10192
rect 5583 10152 6092 10180
rect 5583 10149 5595 10152
rect 5537 10143 5595 10149
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 9766 10180 9772 10192
rect 6380 10152 9772 10180
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 2924 10084 3801 10112
rect 2924 10072 2930 10084
rect 3789 10081 3801 10084
rect 3835 10112 3847 10115
rect 4062 10112 4068 10124
rect 3835 10084 4068 10112
rect 3835 10081 3847 10084
rect 3789 10075 3847 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 6380 10121 6408 10152
rect 9766 10140 9772 10152
rect 9824 10140 9830 10192
rect 10318 10180 10324 10192
rect 9876 10152 10324 10180
rect 6365 10115 6423 10121
rect 4672 10084 5212 10112
rect 4672 10072 4678 10084
rect 5184 10044 5212 10084
rect 6365 10081 6377 10115
rect 6411 10081 6423 10115
rect 6365 10075 6423 10081
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7006 10112 7012 10124
rect 6963 10084 7012 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7098 10072 7104 10124
rect 7156 10112 7162 10124
rect 7377 10115 7435 10121
rect 7156 10084 7328 10112
rect 7156 10072 7162 10084
rect 5718 10044 5724 10056
rect 5184 10030 5724 10044
rect 5198 10016 5724 10030
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5902 10044 5908 10056
rect 5863 10016 5908 10044
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7116 10044 7144 10072
rect 6880 10016 7144 10044
rect 6880 10004 6886 10016
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 7300 10044 7328 10084
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7423 10084 7941 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 8662 10072 8668 10124
rect 8720 10072 8726 10124
rect 9398 10112 9404 10124
rect 8956 10084 9404 10112
rect 8956 10056 8984 10084
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9674 10072 9680 10124
rect 9732 10072 9738 10124
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 7300 10016 7665 10044
rect 7653 10013 7665 10016
rect 7699 10044 7711 10047
rect 8202 10047 8260 10053
rect 7699 10016 8156 10044
rect 7699 10013 7711 10016
rect 7653 10007 7711 10013
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9945 4123 9979
rect 8128 9976 8156 10016
rect 8202 10013 8214 10047
rect 8248 10044 8260 10047
rect 8386 10044 8392 10056
rect 8248 10016 8392 10044
rect 8248 10013 8260 10016
rect 8202 10007 8260 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8938 10004 8944 10056
rect 8996 10004 9002 10056
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 9582 10044 9588 10056
rect 9539 10016 9588 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 9122 9976 9128 9988
rect 4065 9939 4123 9945
rect 5460 9948 8064 9976
rect 8128 9948 9128 9976
rect 4080 9908 4108 9939
rect 5460 9908 5488 9948
rect 4080 9880 5488 9908
rect 5718 9868 5724 9920
rect 5776 9868 5782 9920
rect 5905 9911 5963 9917
rect 5905 9877 5917 9911
rect 5951 9908 5963 9911
rect 5994 9908 6000 9920
rect 5951 9880 6000 9908
rect 5951 9877 5963 9880
rect 5905 9871 5963 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 7466 9868 7472 9920
rect 7524 9868 7530 9920
rect 8036 9917 8064 9948
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 9232 9976 9260 10007
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 9876 10044 9904 10152
rect 10318 10140 10324 10152
rect 10376 10180 10382 10192
rect 10376 10152 10824 10180
rect 10376 10140 10382 10152
rect 10226 10072 10232 10124
rect 10284 10112 10290 10124
rect 10284 10084 10732 10112
rect 10284 10072 10290 10084
rect 9815 10016 9904 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10410 10044 10416 10056
rect 10008 10016 10416 10044
rect 10008 10004 10014 10016
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 10704 10053 10732 10084
rect 10796 10053 10824 10152
rect 16390 10140 16396 10192
rect 16448 10180 16454 10192
rect 16448 10152 18644 10180
rect 16448 10140 16454 10152
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 12069 10115 12127 10121
rect 11103 10084 11928 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11900 10056 11928 10084
rect 12069 10081 12081 10115
rect 12115 10112 12127 10115
rect 12989 10115 13047 10121
rect 12989 10112 13001 10115
rect 12115 10084 13001 10112
rect 12115 10081 12127 10084
rect 12069 10075 12127 10081
rect 12989 10081 13001 10084
rect 13035 10081 13047 10115
rect 12989 10075 13047 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13262 10112 13268 10124
rect 13127 10084 13268 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10112 13415 10115
rect 13906 10112 13912 10124
rect 13403 10084 13912 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 13906 10072 13912 10084
rect 13964 10112 13970 10124
rect 13964 10084 14780 10112
rect 13964 10072 13970 10084
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10044 10839 10047
rect 10962 10044 10968 10056
rect 10827 10016 10968 10044
rect 10827 10013 10839 10016
rect 10781 10007 10839 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11146 10004 11152 10056
rect 11204 10004 11210 10056
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 11296 10016 11345 10044
rect 11296 10004 11302 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10044 11483 10047
rect 11514 10044 11520 10056
rect 11471 10016 11520 10044
rect 11471 10013 11483 10016
rect 11425 10007 11483 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 11882 10004 11888 10056
rect 11940 10004 11946 10056
rect 12342 10004 12348 10056
rect 12400 10004 12406 10056
rect 12618 10004 12624 10056
rect 12676 10004 12682 10056
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 14752 10053 14780 10084
rect 16482 10072 16488 10124
rect 16540 10072 16546 10124
rect 16666 10072 16672 10124
rect 16724 10112 16730 10124
rect 16945 10115 17003 10121
rect 16724 10084 16804 10112
rect 16724 10072 16730 10084
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 14826 10044 14832 10056
rect 14783 10016 14832 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10013 14979 10047
rect 14921 10007 14979 10013
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 9232 9948 12173 9976
rect 12161 9945 12173 9948
rect 12207 9945 12219 9979
rect 13538 9976 13544 9988
rect 12161 9939 12219 9945
rect 12406 9948 13544 9976
rect 8021 9911 8079 9917
rect 8021 9877 8033 9911
rect 8067 9877 8079 9911
rect 8021 9871 8079 9877
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 9039 9911 9097 9917
rect 9039 9908 9051 9911
rect 8251 9880 9051 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 9039 9877 9051 9880
rect 9085 9877 9097 9911
rect 9140 9908 9168 9936
rect 12406 9908 12434 9948
rect 13538 9936 13544 9948
rect 13596 9936 13602 9988
rect 14645 9979 14703 9985
rect 14645 9945 14657 9979
rect 14691 9976 14703 9979
rect 14936 9976 14964 10007
rect 16206 10004 16212 10056
rect 16264 10004 16270 10056
rect 16776 10053 16804 10084
rect 16945 10081 16957 10115
rect 16991 10112 17003 10115
rect 17218 10112 17224 10124
rect 16991 10084 17224 10112
rect 16991 10081 17003 10084
rect 16945 10075 17003 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10112 17463 10115
rect 18414 10112 18420 10124
rect 17451 10084 18420 10112
rect 17451 10081 17463 10084
rect 17405 10075 17463 10081
rect 18414 10072 18420 10084
rect 18472 10112 18478 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18472 10084 18521 10112
rect 18472 10072 18478 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18616 10112 18644 10152
rect 18690 10140 18696 10192
rect 18748 10180 18754 10192
rect 18785 10183 18843 10189
rect 18785 10180 18797 10183
rect 18748 10152 18797 10180
rect 18748 10140 18754 10152
rect 18785 10149 18797 10152
rect 18831 10149 18843 10183
rect 18785 10143 18843 10149
rect 18874 10140 18880 10192
rect 18932 10140 18938 10192
rect 19610 10180 19616 10192
rect 19306 10152 19616 10180
rect 19306 10112 19334 10152
rect 19610 10140 19616 10152
rect 19668 10180 19674 10192
rect 25961 10183 26019 10189
rect 25961 10180 25973 10183
rect 19668 10152 25973 10180
rect 19668 10140 19674 10152
rect 25961 10149 25973 10152
rect 26007 10149 26019 10183
rect 25961 10143 26019 10149
rect 26344 10152 26740 10180
rect 18616 10084 19334 10112
rect 18509 10075 18567 10081
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 19760 10084 20177 10112
rect 19760 10072 19766 10084
rect 20165 10081 20177 10084
rect 20211 10112 20223 10115
rect 21085 10115 21143 10121
rect 21085 10112 21097 10115
rect 20211 10084 21097 10112
rect 20211 10081 20223 10084
rect 20165 10075 20223 10081
rect 21085 10081 21097 10084
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 22922 10072 22928 10124
rect 22980 10112 22986 10124
rect 24857 10115 24915 10121
rect 24857 10112 24869 10115
rect 22980 10084 24869 10112
rect 22980 10072 22986 10084
rect 24857 10081 24869 10084
rect 24903 10081 24915 10115
rect 24857 10075 24915 10081
rect 25317 10115 25375 10121
rect 25317 10081 25329 10115
rect 25363 10112 25375 10115
rect 25682 10112 25688 10124
rect 25363 10084 25688 10112
rect 25363 10081 25375 10084
rect 25317 10075 25375 10081
rect 25682 10072 25688 10084
rect 25740 10072 25746 10124
rect 25869 10115 25927 10121
rect 25869 10081 25881 10115
rect 25915 10112 25927 10115
rect 26234 10112 26240 10124
rect 25915 10084 26240 10112
rect 25915 10081 25927 10084
rect 25869 10075 25927 10081
rect 26234 10072 26240 10084
rect 26292 10112 26298 10124
rect 26344 10112 26372 10152
rect 26712 10124 26740 10152
rect 27890 10140 27896 10192
rect 27948 10180 27954 10192
rect 28169 10183 28227 10189
rect 28169 10180 28181 10183
rect 27948 10152 28181 10180
rect 27948 10140 27954 10152
rect 28169 10149 28181 10152
rect 28215 10149 28227 10183
rect 28169 10143 28227 10149
rect 28718 10140 28724 10192
rect 28776 10140 28782 10192
rect 28828 10180 28856 10220
rect 29089 10217 29101 10251
rect 29135 10248 29147 10251
rect 29454 10248 29460 10260
rect 29135 10220 29460 10248
rect 29135 10217 29147 10220
rect 29089 10211 29147 10217
rect 29454 10208 29460 10220
rect 29512 10208 29518 10260
rect 31018 10208 31024 10260
rect 31076 10208 31082 10260
rect 31202 10180 31208 10192
rect 28828 10152 31208 10180
rect 31202 10140 31208 10152
rect 31260 10140 31266 10192
rect 26292 10084 26372 10112
rect 26292 10072 26298 10084
rect 26418 10072 26424 10124
rect 26476 10072 26482 10124
rect 26694 10072 26700 10124
rect 26752 10112 26758 10124
rect 27249 10115 27307 10121
rect 27249 10112 27261 10115
rect 26752 10084 27261 10112
rect 26752 10072 26758 10084
rect 27249 10081 27261 10084
rect 27295 10081 27307 10115
rect 27249 10075 27307 10081
rect 28350 10072 28356 10124
rect 28408 10112 28414 10124
rect 28408 10084 31340 10112
rect 28408 10072 28414 10084
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 18432 10016 18705 10044
rect 18432 10010 18460 10016
rect 17954 9976 17960 9988
rect 14691 9948 17960 9976
rect 14691 9945 14703 9948
rect 14645 9939 14703 9945
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 18138 9936 18144 9988
rect 18196 9976 18202 9988
rect 18340 9982 18460 10010
rect 18693 10013 18705 10016
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 18969 10047 19027 10053
rect 18969 10013 18981 10047
rect 19015 10044 19027 10047
rect 19426 10044 19432 10056
rect 19015 10016 19432 10044
rect 19015 10013 19027 10016
rect 18969 10007 19027 10013
rect 18340 9976 18368 9982
rect 18196 9948 18368 9976
rect 18708 9976 18736 10007
rect 19426 10004 19432 10016
rect 19484 10044 19490 10056
rect 19978 10044 19984 10056
rect 19484 10016 19984 10044
rect 19484 10004 19490 10016
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 19334 9976 19340 9988
rect 18708 9948 19340 9976
rect 18196 9936 18202 9948
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 20088 9976 20116 10007
rect 20254 10004 20260 10056
rect 20312 10004 20318 10056
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20622 10044 20628 10056
rect 20579 10016 20628 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 19944 9948 20116 9976
rect 19944 9936 19950 9948
rect 9140 9880 12434 9908
rect 12529 9911 12587 9917
rect 9039 9871 9097 9877
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12894 9908 12900 9920
rect 12575 9880 12900 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 13354 9908 13360 9920
rect 13311 9880 13360 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 13814 9908 13820 9920
rect 13679 9880 13820 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 14734 9868 14740 9920
rect 14792 9908 14798 9920
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 14792 9880 14841 9908
rect 14792 9868 14798 9880
rect 14829 9877 14841 9880
rect 14875 9877 14887 9911
rect 14829 9871 14887 9877
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 19702 9908 19708 9920
rect 14976 9880 19708 9908
rect 14976 9868 14982 9880
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 20088 9908 20116 9948
rect 20162 9936 20168 9988
rect 20220 9976 20226 9988
rect 20364 9976 20392 10007
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 20732 10016 21036 10044
rect 20220 9948 20392 9976
rect 20220 9936 20226 9948
rect 20732 9908 20760 10016
rect 21008 9985 21036 10016
rect 21450 10004 21456 10056
rect 21508 10004 21514 10056
rect 21821 10047 21879 10053
rect 21821 10013 21833 10047
rect 21867 10013 21879 10047
rect 21821 10007 21879 10013
rect 20993 9979 21051 9985
rect 20993 9945 21005 9979
rect 21039 9945 21051 9979
rect 20993 9939 21051 9945
rect 21266 9936 21272 9988
rect 21324 9936 21330 9988
rect 21836 9976 21864 10007
rect 22002 10004 22008 10056
rect 22060 10004 22066 10056
rect 22281 10047 22339 10053
rect 22281 10013 22293 10047
rect 22327 10044 22339 10047
rect 23934 10044 23940 10056
rect 22327 10016 23940 10044
rect 22327 10013 22339 10016
rect 22281 10007 22339 10013
rect 23934 10004 23940 10016
rect 23992 10004 23998 10056
rect 24765 10047 24823 10053
rect 24765 10013 24777 10047
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 25133 10047 25191 10053
rect 25133 10013 25145 10047
rect 25179 10044 25191 10047
rect 25222 10044 25228 10056
rect 25179 10016 25228 10044
rect 25179 10013 25191 10016
rect 25133 10007 25191 10013
rect 22922 9976 22928 9988
rect 21836 9948 22928 9976
rect 22922 9936 22928 9948
rect 22980 9976 22986 9988
rect 24302 9976 24308 9988
rect 22980 9948 24308 9976
rect 22980 9936 22986 9948
rect 24302 9936 24308 9948
rect 24360 9936 24366 9988
rect 24780 9976 24808 10007
rect 25222 10004 25228 10016
rect 25280 10044 25286 10056
rect 26145 10047 26203 10053
rect 26145 10044 26157 10047
rect 25280 10016 26157 10044
rect 25280 10004 25286 10016
rect 26145 10013 26157 10016
rect 26191 10013 26203 10047
rect 26605 10047 26663 10053
rect 26605 10044 26617 10047
rect 26145 10007 26203 10013
rect 26436 10016 26617 10044
rect 25590 9976 25596 9988
rect 24780 9948 25596 9976
rect 25590 9936 25596 9948
rect 25648 9976 25654 9988
rect 26050 9976 26056 9988
rect 25648 9948 26056 9976
rect 25648 9936 25654 9948
rect 26050 9936 26056 9948
rect 26108 9936 26114 9988
rect 20088 9880 20760 9908
rect 20793 9911 20851 9917
rect 20793 9877 20805 9911
rect 20839 9908 20851 9911
rect 21358 9908 21364 9920
rect 20839 9880 21364 9908
rect 20839 9877 20851 9880
rect 20793 9871 20851 9877
rect 21358 9868 21364 9880
rect 21416 9908 21422 9920
rect 21818 9908 21824 9920
rect 21416 9880 21824 9908
rect 21416 9868 21422 9880
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 26436 9908 26464 10016
rect 26605 10013 26617 10016
rect 26651 10013 26663 10047
rect 26605 10007 26663 10013
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10044 27031 10047
rect 27019 10016 27292 10044
rect 27019 10013 27031 10016
rect 26973 10007 27031 10013
rect 26510 9936 26516 9988
rect 26568 9976 26574 9988
rect 26988 9976 27016 10007
rect 26568 9948 27016 9976
rect 26568 9936 26574 9948
rect 27062 9908 27068 9920
rect 26436 9880 27068 9908
rect 27062 9868 27068 9880
rect 27120 9868 27126 9920
rect 27264 9908 27292 10016
rect 27338 10004 27344 10056
rect 27396 10044 27402 10056
rect 27890 10044 27896 10056
rect 27396 10016 27896 10044
rect 27396 10004 27402 10016
rect 27890 10004 27896 10016
rect 27948 10044 27954 10056
rect 28166 10044 28172 10056
rect 27948 10016 28172 10044
rect 27948 10004 27954 10016
rect 28166 10004 28172 10016
rect 28224 10004 28230 10056
rect 28917 10047 28975 10053
rect 28917 10034 28929 10047
rect 28074 9936 28080 9988
rect 28132 9976 28138 9988
rect 28463 9979 28521 9985
rect 28902 9982 28908 10034
rect 28963 10013 28975 10047
rect 28960 10007 28975 10013
rect 28960 9982 28966 10007
rect 29178 10004 29184 10056
rect 29236 10044 29242 10056
rect 29273 10047 29331 10053
rect 29273 10044 29285 10047
rect 29236 10016 29285 10044
rect 29236 10004 29242 10016
rect 29273 10013 29285 10016
rect 29319 10013 29331 10047
rect 29273 10007 29331 10013
rect 29546 10004 29552 10056
rect 29604 10044 29610 10056
rect 29822 10053 29828 10056
rect 29641 10047 29699 10053
rect 29641 10044 29653 10047
rect 29604 10016 29653 10044
rect 29604 10004 29610 10016
rect 29641 10013 29653 10016
rect 29687 10013 29699 10047
rect 29641 10007 29699 10013
rect 29799 10047 29828 10053
rect 29799 10013 29811 10047
rect 29799 10007 29828 10013
rect 29822 10004 29828 10007
rect 29880 10004 29886 10056
rect 30098 10004 30104 10056
rect 30156 10004 30162 10056
rect 30190 10004 30196 10056
rect 30248 10044 30254 10056
rect 30377 10047 30435 10053
rect 30377 10044 30389 10047
rect 30248 10016 30389 10044
rect 30248 10004 30254 10016
rect 30377 10013 30389 10016
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 30742 10004 30748 10056
rect 30800 10004 30806 10056
rect 31202 10053 31208 10056
rect 31200 10044 31208 10053
rect 30852 10016 31208 10044
rect 28463 9976 28475 9979
rect 28132 9948 28475 9976
rect 28132 9936 28138 9948
rect 28463 9945 28475 9948
rect 28509 9945 28521 9979
rect 28463 9939 28521 9945
rect 29012 9948 29776 9976
rect 29012 9908 29040 9948
rect 29748 9920 29776 9948
rect 29914 9936 29920 9988
rect 29972 9936 29978 9988
rect 30009 9979 30067 9985
rect 30009 9945 30021 9979
rect 30055 9945 30067 9979
rect 30116 9976 30144 10004
rect 30852 9976 30880 10016
rect 31200 10007 31208 10016
rect 31202 10004 31208 10007
rect 31260 10004 31266 10056
rect 31312 10053 31340 10084
rect 31386 10072 31392 10124
rect 31444 10112 31450 10124
rect 31444 10084 31560 10112
rect 31444 10072 31450 10084
rect 31532 10053 31560 10084
rect 31297 10047 31355 10053
rect 31297 10013 31309 10047
rect 31343 10013 31355 10047
rect 31297 10007 31355 10013
rect 31517 10047 31575 10053
rect 31517 10013 31529 10047
rect 31563 10013 31575 10047
rect 31517 10007 31575 10013
rect 31662 10004 31668 10056
rect 31720 10004 31726 10056
rect 30116 9948 30880 9976
rect 30009 9939 30067 9945
rect 27264 9880 29040 9908
rect 29730 9868 29736 9920
rect 29788 9868 29794 9920
rect 29822 9868 29828 9920
rect 29880 9908 29886 9920
rect 30024 9908 30052 9939
rect 30926 9936 30932 9988
rect 30984 9976 30990 9988
rect 31389 9979 31447 9985
rect 31389 9976 31401 9979
rect 30984 9948 31401 9976
rect 30984 9936 30990 9948
rect 31389 9945 31401 9948
rect 31435 9976 31447 9979
rect 34330 9976 34336 9988
rect 31435 9948 34336 9976
rect 31435 9945 31447 9948
rect 31389 9939 31447 9945
rect 34330 9936 34336 9948
rect 34388 9936 34394 9988
rect 30190 9908 30196 9920
rect 29880 9880 30196 9908
rect 29880 9868 29886 9880
rect 30190 9868 30196 9880
rect 30248 9868 30254 9920
rect 30285 9911 30343 9917
rect 30285 9877 30297 9911
rect 30331 9908 30343 9911
rect 30374 9908 30380 9920
rect 30331 9880 30380 9908
rect 30331 9877 30343 9880
rect 30285 9871 30343 9877
rect 30374 9868 30380 9880
rect 30432 9868 30438 9920
rect 31110 9868 31116 9920
rect 31168 9908 31174 9920
rect 31478 9908 31484 9920
rect 31168 9880 31484 9908
rect 31168 9868 31174 9880
rect 31478 9868 31484 9880
rect 31536 9908 31542 9920
rect 36262 9908 36268 9920
rect 31536 9880 36268 9908
rect 31536 9868 31542 9880
rect 36262 9868 36268 9880
rect 36320 9868 36326 9920
rect 1104 9818 36524 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 36524 9818
rect 1104 9744 36524 9766
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10781 9707 10839 9713
rect 10781 9704 10793 9707
rect 10652 9676 10793 9704
rect 10652 9664 10658 9676
rect 10781 9673 10793 9676
rect 10827 9673 10839 9707
rect 10781 9667 10839 9673
rect 13446 9664 13452 9716
rect 13504 9664 13510 9716
rect 14369 9707 14427 9713
rect 14369 9704 14381 9707
rect 13740 9676 14381 9704
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6236 9608 6837 9636
rect 6236 9596 6242 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 11054 9636 11060 9648
rect 6825 9599 6883 9605
rect 10152 9608 11060 9636
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 6728 9571 6786 9577
rect 6728 9568 6740 9571
rect 6052 9540 6740 9568
rect 6052 9528 6058 9540
rect 6728 9537 6740 9540
rect 6774 9568 6786 9571
rect 6774 9540 6868 9568
rect 6774 9537 6786 9540
rect 6728 9531 6786 9537
rect 4062 9460 4068 9512
rect 4120 9500 4126 9512
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 4120 9472 4445 9500
rect 4120 9460 4126 9472
rect 4433 9469 4445 9472
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 6840 9500 6868 9540
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7098 9568 7104 9580
rect 7059 9540 7104 9568
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 7466 9568 7472 9580
rect 7239 9540 7472 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 10152 9577 10180 9608
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 13740 9645 13768 9676
rect 14369 9673 14381 9676
rect 14415 9704 14427 9707
rect 14415 9676 15516 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 13725 9639 13783 9645
rect 13725 9605 13737 9639
rect 13771 9605 13783 9639
rect 13725 9599 13783 9605
rect 13817 9639 13875 9645
rect 13817 9605 13829 9639
rect 13863 9636 13875 9639
rect 14182 9636 14188 9648
rect 13863 9608 14188 9636
rect 13863 9605 13875 9608
rect 13817 9599 13875 9605
rect 14182 9596 14188 9608
rect 14240 9636 14246 9648
rect 14918 9636 14924 9648
rect 14240 9608 14924 9636
rect 14240 9596 14246 9608
rect 10137 9571 10195 9577
rect 10137 9537 10149 9571
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10520 9540 10885 9568
rect 8938 9500 8944 9512
rect 4755 9472 6592 9500
rect 6840 9472 8944 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 6178 9392 6184 9444
rect 6236 9392 6242 9444
rect 6564 9441 6592 9472
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 10318 9460 10324 9512
rect 10376 9500 10382 9512
rect 10520 9500 10548 9540
rect 10873 9537 10885 9540
rect 10919 9568 10931 9571
rect 11146 9568 11152 9580
rect 10919 9540 11152 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 11698 9568 11704 9580
rect 11256 9540 11704 9568
rect 10376 9472 10548 9500
rect 10597 9503 10655 9509
rect 10376 9460 10382 9472
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 11256 9500 11284 9540
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 13630 9568 13636 9580
rect 12584 9540 13636 9568
rect 12584 9528 12590 9540
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 14292 9577 14320 9608
rect 14918 9596 14924 9608
rect 14976 9636 14982 9648
rect 15488 9636 15516 9676
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 17954 9704 17960 9716
rect 16080 9676 17960 9704
rect 16080 9664 16086 9676
rect 17954 9664 17960 9676
rect 18012 9704 18018 9716
rect 18138 9704 18144 9716
rect 18012 9676 18144 9704
rect 18012 9664 18018 9676
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 18230 9664 18236 9716
rect 18288 9704 18294 9716
rect 18690 9704 18696 9716
rect 18288 9676 18696 9704
rect 18288 9664 18294 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 17310 9636 17316 9648
rect 14976 9608 15424 9636
rect 15488 9608 17316 9636
rect 14976 9596 14982 9608
rect 13955 9571 14013 9577
rect 13955 9537 13967 9571
rect 14001 9568 14013 9571
rect 14292 9571 14368 9577
rect 14001 9540 14228 9568
rect 14292 9540 14322 9571
rect 14001 9537 14013 9540
rect 13955 9531 14013 9537
rect 10643 9472 11284 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 11330 9460 11336 9512
rect 11388 9500 11394 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11388 9472 11621 9500
rect 11388 9460 11394 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 14090 9460 14096 9512
rect 14148 9460 14154 9512
rect 6549 9435 6607 9441
rect 6549 9401 6561 9435
rect 6595 9401 6607 9435
rect 6549 9395 6607 9401
rect 12069 9435 12127 9441
rect 12069 9401 12081 9435
rect 12115 9432 12127 9435
rect 12618 9432 12624 9444
rect 12115 9404 12624 9432
rect 12115 9401 12127 9404
rect 12069 9395 12127 9401
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 14200 9441 14228 9540
rect 14310 9537 14322 9540
rect 14356 9537 14368 9571
rect 14310 9531 14368 9537
rect 14734 9528 14740 9580
rect 14792 9528 14798 9580
rect 15396 9577 15424 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 18800 9642 19012 9670
rect 24578 9664 24584 9716
rect 24636 9664 24642 9716
rect 28534 9704 28540 9716
rect 28184 9676 28540 9704
rect 18800 9636 18828 9642
rect 17926 9608 18257 9636
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 15562 9528 15568 9580
rect 15620 9568 15626 9580
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 15620 9540 15761 9568
rect 15620 9528 15626 9540
rect 15749 9537 15761 9540
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 15930 9528 15936 9580
rect 15988 9528 15994 9580
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16390 9568 16396 9580
rect 16255 9540 16396 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 15102 9500 15108 9512
rect 14875 9472 15108 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 15654 9460 15660 9512
rect 15712 9460 15718 9512
rect 15948 9500 15976 9528
rect 17034 9500 17040 9512
rect 15948 9472 17040 9500
rect 17034 9460 17040 9472
rect 17092 9500 17098 9512
rect 17926 9500 17954 9608
rect 18229 9577 18257 9608
rect 18340 9608 18828 9636
rect 18984 9636 19012 9642
rect 19245 9639 19303 9645
rect 19245 9636 19257 9639
rect 18984 9608 19257 9636
rect 18340 9580 18368 9608
rect 19245 9605 19257 9608
rect 19291 9605 19303 9639
rect 20441 9639 20499 9645
rect 20441 9636 20453 9639
rect 19245 9599 19303 9605
rect 19720 9608 20453 9636
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9558 18107 9571
rect 18214 9571 18272 9577
rect 18095 9537 18184 9558
rect 18049 9531 18184 9537
rect 18214 9537 18226 9571
rect 18260 9537 18272 9571
rect 18214 9531 18272 9537
rect 18064 9530 18184 9531
rect 17092 9472 17954 9500
rect 18156 9500 18184 9530
rect 18322 9528 18328 9580
rect 18380 9528 18386 9580
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 18506 9568 18512 9580
rect 18463 9540 18512 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18690 9528 18696 9580
rect 18748 9574 18754 9580
rect 18877 9577 18935 9583
rect 18785 9574 18843 9577
rect 18748 9571 18843 9574
rect 18748 9546 18797 9571
rect 18748 9528 18754 9546
rect 18785 9537 18797 9546
rect 18831 9537 18843 9571
rect 18877 9543 18889 9577
rect 18923 9574 18935 9577
rect 18966 9574 18972 9580
rect 18923 9546 18972 9574
rect 18923 9543 18935 9546
rect 18877 9537 18935 9543
rect 18785 9531 18843 9537
rect 18966 9528 18972 9546
rect 19024 9528 19030 9580
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19521 9571 19579 9577
rect 19521 9568 19533 9571
rect 19484 9540 19533 9568
rect 19484 9528 19490 9540
rect 19521 9537 19533 9540
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19610 9528 19616 9580
rect 19668 9528 19674 9580
rect 19720 9577 19748 9608
rect 20441 9605 20453 9608
rect 20487 9636 20499 9639
rect 21266 9636 21272 9648
rect 20487 9608 21272 9636
rect 20487 9605 20499 9608
rect 20441 9599 20499 9605
rect 21266 9596 21272 9608
rect 21324 9636 21330 9648
rect 21324 9608 23428 9636
rect 21324 9596 21330 9608
rect 19705 9571 19763 9577
rect 19705 9537 19717 9571
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 19981 9571 20039 9577
rect 19981 9537 19993 9571
rect 20027 9568 20039 9571
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 20027 9540 20269 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 20257 9537 20269 9540
rect 20303 9568 20315 9571
rect 20622 9568 20628 9580
rect 20303 9540 20628 9568
rect 20303 9537 20315 9540
rect 20257 9531 20315 9537
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9537 22523 9571
rect 22465 9531 22523 9537
rect 19794 9500 19800 9512
rect 18156 9472 19800 9500
rect 17092 9460 17098 9472
rect 19794 9460 19800 9472
rect 19852 9460 19858 9512
rect 22480 9500 22508 9531
rect 22554 9528 22560 9580
rect 22612 9528 22618 9580
rect 22922 9528 22928 9580
rect 22980 9528 22986 9580
rect 23198 9528 23204 9580
rect 23256 9568 23262 9580
rect 23400 9577 23428 9608
rect 23842 9596 23848 9648
rect 23900 9636 23906 9648
rect 24596 9636 24624 9664
rect 23900 9608 24624 9636
rect 25792 9608 26372 9636
rect 23900 9596 23906 9608
rect 23293 9571 23351 9577
rect 23293 9568 23305 9571
rect 23256 9540 23305 9568
rect 23256 9528 23262 9540
rect 23293 9537 23305 9540
rect 23339 9537 23351 9571
rect 23293 9531 23351 9537
rect 23385 9571 23443 9577
rect 23385 9537 23397 9571
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23569 9571 23627 9577
rect 23569 9537 23581 9571
rect 23615 9568 23627 9571
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 23615 9540 24317 9568
rect 23615 9537 23627 9540
rect 23569 9531 23627 9537
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 23216 9500 23244 9528
rect 22480 9472 23244 9500
rect 23400 9500 23428 9531
rect 24320 9500 24348 9531
rect 24394 9528 24400 9580
rect 24452 9528 24458 9580
rect 24578 9528 24584 9580
rect 24636 9528 24642 9580
rect 25498 9528 25504 9580
rect 25556 9568 25562 9580
rect 25792 9577 25820 9608
rect 25777 9571 25835 9577
rect 25777 9568 25789 9571
rect 25556 9540 25789 9568
rect 25556 9528 25562 9540
rect 25777 9537 25789 9540
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 26050 9528 26056 9580
rect 26108 9528 26114 9580
rect 26344 9577 26372 9608
rect 26970 9596 26976 9648
rect 27028 9636 27034 9648
rect 28077 9639 28135 9645
rect 28077 9636 28089 9639
rect 27028 9608 28089 9636
rect 27028 9596 27034 9608
rect 28077 9605 28089 9608
rect 28123 9605 28135 9639
rect 28077 9599 28135 9605
rect 26329 9571 26387 9577
rect 26329 9537 26341 9571
rect 26375 9537 26387 9571
rect 26329 9531 26387 9537
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9568 26663 9571
rect 26694 9568 26700 9580
rect 26651 9540 26700 9568
rect 26651 9537 26663 9540
rect 26605 9531 26663 9537
rect 26694 9528 26700 9540
rect 26752 9528 26758 9580
rect 27154 9528 27160 9580
rect 27212 9528 27218 9580
rect 27709 9571 27767 9577
rect 27709 9537 27721 9571
rect 27755 9537 27767 9571
rect 27709 9531 27767 9537
rect 27985 9571 28043 9577
rect 27985 9537 27997 9571
rect 28031 9568 28043 9571
rect 28184 9568 28212 9676
rect 28534 9664 28540 9676
rect 28592 9664 28598 9716
rect 32030 9704 32036 9716
rect 30300 9676 32036 9704
rect 28718 9636 28724 9648
rect 28552 9608 28724 9636
rect 28552 9577 28580 9608
rect 28718 9596 28724 9608
rect 28776 9596 28782 9648
rect 29454 9636 29460 9648
rect 29104 9608 29460 9636
rect 28031 9540 28212 9568
rect 28537 9571 28595 9577
rect 28031 9537 28043 9540
rect 27985 9531 28043 9537
rect 28537 9537 28549 9571
rect 28583 9537 28595 9571
rect 28537 9531 28595 9537
rect 28629 9571 28687 9577
rect 28629 9537 28641 9571
rect 28675 9568 28687 9571
rect 29104 9568 29132 9608
rect 29454 9596 29460 9608
rect 29512 9596 29518 9648
rect 29546 9596 29552 9648
rect 29604 9636 29610 9648
rect 30300 9636 30328 9676
rect 32030 9664 32036 9676
rect 32088 9664 32094 9716
rect 33505 9707 33563 9713
rect 33505 9673 33517 9707
rect 33551 9704 33563 9707
rect 33686 9704 33692 9716
rect 33551 9676 33692 9704
rect 33551 9673 33563 9676
rect 33505 9667 33563 9673
rect 33686 9664 33692 9676
rect 33744 9664 33750 9716
rect 34330 9664 34336 9716
rect 34388 9664 34394 9716
rect 34790 9664 34796 9716
rect 34848 9704 34854 9716
rect 34885 9707 34943 9713
rect 34885 9704 34897 9707
rect 34848 9676 34897 9704
rect 34848 9664 34854 9676
rect 34885 9673 34897 9676
rect 34931 9673 34943 9707
rect 34885 9667 34943 9673
rect 29604 9608 30328 9636
rect 29604 9596 29610 9608
rect 30374 9596 30380 9648
rect 30432 9636 30438 9648
rect 34348 9636 34376 9664
rect 34517 9639 34575 9645
rect 34517 9636 34529 9639
rect 30432 9608 34284 9636
rect 34348 9608 34529 9636
rect 30432 9596 30438 9608
rect 28675 9540 29132 9568
rect 29181 9571 29239 9577
rect 28675 9537 28687 9540
rect 28629 9531 28687 9537
rect 29181 9537 29193 9571
rect 29227 9568 29239 9571
rect 29270 9568 29276 9580
rect 29227 9540 29276 9568
rect 29227 9537 29239 9540
rect 29181 9531 29239 9537
rect 25038 9500 25044 9512
rect 23400 9472 23704 9500
rect 24320 9472 25044 9500
rect 14185 9435 14243 9441
rect 14185 9401 14197 9435
rect 14231 9401 14243 9435
rect 14185 9395 14243 9401
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9432 16175 9435
rect 16758 9432 16764 9444
rect 16163 9404 16764 9432
rect 16163 9401 16175 9404
rect 16117 9395 16175 9401
rect 16758 9392 16764 9404
rect 16816 9392 16822 9444
rect 18874 9392 18880 9444
rect 18932 9432 18938 9444
rect 20073 9435 20131 9441
rect 20073 9432 20085 9435
rect 18932 9404 20085 9432
rect 18932 9392 18938 9404
rect 20073 9401 20085 9404
rect 20119 9401 20131 9435
rect 22554 9432 22560 9444
rect 20073 9395 20131 9401
rect 20180 9404 22560 9432
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15286 9364 15292 9376
rect 15243 9336 15292 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 17865 9367 17923 9373
rect 17865 9364 17877 9367
rect 17552 9336 17877 9364
rect 17552 9324 17558 9336
rect 17865 9333 17877 9336
rect 17911 9333 17923 9367
rect 17865 9327 17923 9333
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 18196 9336 18521 9364
rect 18196 9324 18202 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 18598 9324 18604 9376
rect 18656 9364 18662 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 18656 9336 18705 9364
rect 18656 9324 18662 9336
rect 18693 9333 18705 9336
rect 18739 9333 18751 9367
rect 18693 9327 18751 9333
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 19116 9336 19809 9364
rect 19116 9324 19122 9336
rect 19797 9333 19809 9336
rect 19843 9364 19855 9367
rect 20180 9364 20208 9404
rect 22554 9392 22560 9404
rect 22612 9392 22618 9444
rect 22649 9435 22707 9441
rect 22649 9401 22661 9435
rect 22695 9432 22707 9435
rect 23014 9432 23020 9444
rect 22695 9404 23020 9432
rect 22695 9401 22707 9404
rect 22649 9395 22707 9401
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 23566 9392 23572 9444
rect 23624 9392 23630 9444
rect 23676 9432 23704 9472
rect 25038 9460 25044 9472
rect 25096 9460 25102 9512
rect 25130 9460 25136 9512
rect 25188 9500 25194 9512
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 25188 9472 25697 9500
rect 25188 9460 25194 9472
rect 25685 9469 25697 9472
rect 25731 9500 25743 9503
rect 25958 9500 25964 9512
rect 25731 9472 25964 9500
rect 25731 9469 25743 9472
rect 25685 9463 25743 9469
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 27341 9503 27399 9509
rect 27341 9500 27353 9503
rect 26252 9472 27353 9500
rect 23676 9404 25544 9432
rect 19843 9336 20208 9364
rect 22189 9367 22247 9373
rect 19843 9333 19855 9336
rect 19797 9327 19855 9333
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 22462 9364 22468 9376
rect 22235 9336 22468 9364
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 22741 9367 22799 9373
rect 22741 9333 22753 9367
rect 22787 9364 22799 9367
rect 22830 9364 22836 9376
rect 22787 9336 22836 9364
rect 22787 9333 22799 9336
rect 22741 9327 22799 9333
rect 22830 9324 22836 9336
rect 22888 9324 22894 9376
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 24121 9367 24179 9373
rect 24121 9364 24133 9367
rect 23440 9336 24133 9364
rect 23440 9324 23446 9336
rect 24121 9333 24133 9336
rect 24167 9333 24179 9367
rect 24121 9327 24179 9333
rect 24581 9367 24639 9373
rect 24581 9333 24593 9367
rect 24627 9364 24639 9367
rect 25406 9364 25412 9376
rect 24627 9336 25412 9364
rect 24627 9333 24639 9336
rect 24581 9327 24639 9333
rect 25406 9324 25412 9336
rect 25464 9324 25470 9376
rect 25516 9364 25544 9404
rect 25866 9392 25872 9444
rect 25924 9432 25930 9444
rect 26252 9432 26280 9472
rect 27341 9469 27353 9472
rect 27387 9500 27399 9503
rect 27430 9500 27436 9512
rect 27387 9472 27436 9500
rect 27387 9469 27399 9472
rect 27341 9463 27399 9469
rect 27430 9460 27436 9472
rect 27488 9500 27494 9512
rect 27724 9500 27752 9531
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29641 9571 29699 9577
rect 29641 9537 29653 9571
rect 29687 9568 29699 9571
rect 29822 9568 29828 9580
rect 29687 9540 29828 9568
rect 29687 9537 29699 9540
rect 29641 9531 29699 9537
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 30006 9528 30012 9580
rect 30064 9568 30070 9580
rect 30101 9571 30159 9577
rect 30101 9568 30113 9571
rect 30064 9540 30113 9568
rect 30064 9528 30070 9540
rect 30101 9537 30113 9540
rect 30147 9537 30159 9571
rect 30101 9531 30159 9537
rect 32858 9528 32864 9580
rect 32916 9528 32922 9580
rect 33042 9577 33048 9580
rect 33019 9571 33048 9577
rect 33019 9537 33031 9571
rect 33019 9531 33048 9537
rect 33042 9528 33048 9531
rect 33100 9528 33106 9580
rect 33134 9528 33140 9580
rect 33192 9528 33198 9580
rect 33226 9528 33232 9580
rect 33284 9528 33290 9580
rect 33318 9528 33324 9580
rect 33376 9568 33382 9580
rect 33502 9568 33508 9580
rect 33376 9540 33508 9568
rect 33376 9528 33382 9540
rect 33502 9528 33508 9540
rect 33560 9528 33566 9580
rect 33594 9528 33600 9580
rect 33652 9528 33658 9580
rect 34256 9577 34284 9608
rect 34517 9605 34529 9608
rect 34563 9605 34575 9639
rect 34517 9599 34575 9605
rect 34241 9571 34299 9577
rect 34241 9537 34253 9571
rect 34287 9537 34299 9571
rect 34241 9531 34299 9537
rect 34330 9528 34336 9580
rect 34388 9568 34394 9580
rect 34609 9571 34667 9577
rect 34388 9540 34433 9568
rect 34388 9528 34394 9540
rect 34609 9537 34621 9571
rect 34655 9537 34667 9571
rect 34609 9531 34667 9537
rect 34706 9571 34764 9577
rect 34706 9537 34718 9571
rect 34752 9537 34764 9571
rect 34706 9531 34764 9537
rect 27488 9472 27752 9500
rect 27488 9460 27494 9472
rect 27798 9460 27804 9512
rect 27856 9500 27862 9512
rect 28442 9500 28448 9512
rect 27856 9472 28448 9500
rect 27856 9460 27862 9472
rect 28442 9460 28448 9472
rect 28500 9500 28506 9512
rect 28902 9500 28908 9512
rect 28500 9472 28908 9500
rect 28500 9460 28506 9472
rect 28902 9460 28908 9472
rect 28960 9500 28966 9512
rect 28997 9503 29055 9509
rect 28997 9500 29009 9503
rect 28960 9472 29009 9500
rect 28960 9460 28966 9472
rect 28997 9469 29009 9472
rect 29043 9469 29055 9503
rect 34624 9500 34652 9531
rect 28997 9463 29055 9469
rect 32968 9472 34652 9500
rect 25924 9404 26280 9432
rect 25924 9392 25930 9404
rect 26326 9392 26332 9444
rect 26384 9432 26390 9444
rect 27706 9432 27712 9444
rect 26384 9404 27712 9432
rect 26384 9392 26390 9404
rect 27706 9392 27712 9404
rect 27764 9392 27770 9444
rect 29365 9435 29423 9441
rect 29365 9432 29377 9435
rect 27816 9404 29377 9432
rect 27816 9364 27844 9404
rect 29365 9401 29377 9404
rect 29411 9432 29423 9435
rect 32968 9432 32996 9472
rect 29411 9404 32996 9432
rect 29411 9401 29423 9404
rect 29365 9395 29423 9401
rect 33226 9392 33232 9444
rect 33284 9432 33290 9444
rect 33781 9435 33839 9441
rect 33781 9432 33793 9435
rect 33284 9404 33793 9432
rect 33284 9392 33290 9404
rect 33781 9401 33793 9404
rect 33827 9401 33839 9435
rect 33781 9395 33839 9401
rect 25516 9336 27844 9364
rect 28718 9324 28724 9376
rect 28776 9364 28782 9376
rect 28813 9367 28871 9373
rect 28813 9364 28825 9367
rect 28776 9336 28825 9364
rect 28776 9324 28782 9336
rect 28813 9333 28825 9336
rect 28859 9333 28871 9367
rect 28813 9327 28871 9333
rect 28902 9324 28908 9376
rect 28960 9364 28966 9376
rect 29549 9367 29607 9373
rect 29549 9364 29561 9367
rect 28960 9336 29561 9364
rect 28960 9324 28966 9336
rect 29549 9333 29561 9336
rect 29595 9333 29607 9367
rect 29549 9327 29607 9333
rect 29914 9324 29920 9376
rect 29972 9364 29978 9376
rect 30098 9364 30104 9376
rect 29972 9336 30104 9364
rect 29972 9324 29978 9336
rect 30098 9324 30104 9336
rect 30156 9364 30162 9376
rect 30285 9367 30343 9373
rect 30285 9364 30297 9367
rect 30156 9336 30297 9364
rect 30156 9324 30162 9336
rect 30285 9333 30297 9336
rect 30331 9333 30343 9367
rect 30285 9327 30343 9333
rect 33318 9324 33324 9376
rect 33376 9364 33382 9376
rect 34716 9364 34744 9531
rect 33376 9336 34744 9364
rect 33376 9324 33382 9336
rect 1104 9274 36524 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 36524 9274
rect 1104 9200 36524 9222
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 5960 9132 6285 9160
rect 5960 9120 5966 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 6914 9160 6920 9172
rect 6871 9132 6920 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7156 9132 7297 9160
rect 7156 9120 7162 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 15194 9160 15200 9172
rect 7285 9123 7343 9129
rect 7392 9132 15200 9160
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 7392 9024 7420 9132
rect 15194 9120 15200 9132
rect 15252 9160 15258 9172
rect 16114 9160 16120 9172
rect 15252 9132 16120 9160
rect 15252 9120 15258 9132
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 17402 9120 17408 9172
rect 17460 9160 17466 9172
rect 18141 9163 18199 9169
rect 18141 9160 18153 9163
rect 17460 9132 18153 9160
rect 17460 9120 17466 9132
rect 18141 9129 18153 9132
rect 18187 9129 18199 9163
rect 18141 9123 18199 9129
rect 18598 9120 18604 9172
rect 18656 9120 18662 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 21085 9163 21143 9169
rect 21085 9160 21097 9163
rect 19392 9132 21097 9160
rect 19392 9120 19398 9132
rect 21085 9129 21097 9132
rect 21131 9160 21143 9163
rect 21358 9160 21364 9172
rect 21131 9132 21364 9160
rect 21131 9129 21143 9132
rect 21085 9123 21143 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 21450 9120 21456 9172
rect 21508 9160 21514 9172
rect 21545 9163 21603 9169
rect 21545 9160 21557 9163
rect 21508 9132 21557 9160
rect 21508 9120 21514 9132
rect 21545 9129 21557 9132
rect 21591 9129 21603 9163
rect 21545 9123 21603 9129
rect 21913 9163 21971 9169
rect 21913 9129 21925 9163
rect 21959 9160 21971 9163
rect 22002 9160 22008 9172
rect 21959 9132 22008 9160
rect 21959 9129 21971 9132
rect 21913 9123 21971 9129
rect 22002 9120 22008 9132
rect 22060 9120 22066 9172
rect 22646 9120 22652 9172
rect 22704 9120 22710 9172
rect 22738 9120 22744 9172
rect 22796 9160 22802 9172
rect 22833 9163 22891 9169
rect 22833 9160 22845 9163
rect 22796 9132 22845 9160
rect 22796 9120 22802 9132
rect 22833 9129 22845 9132
rect 22879 9129 22891 9163
rect 22833 9123 22891 9129
rect 24394 9120 24400 9172
rect 24452 9120 24458 9172
rect 25038 9120 25044 9172
rect 25096 9120 25102 9172
rect 25409 9163 25467 9169
rect 25409 9129 25421 9163
rect 25455 9160 25467 9163
rect 25958 9160 25964 9172
rect 25455 9132 25964 9160
rect 25455 9129 25467 9132
rect 25409 9123 25467 9129
rect 25958 9120 25964 9132
rect 26016 9160 26022 9172
rect 27709 9163 27767 9169
rect 27709 9160 27721 9163
rect 26016 9132 27721 9160
rect 26016 9120 26022 9132
rect 27709 9129 27721 9132
rect 27755 9129 27767 9163
rect 31389 9163 31447 9169
rect 27709 9123 27767 9129
rect 28552 9132 30696 9160
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 8352 9064 9720 9092
rect 8352 9052 8358 9064
rect 5868 8996 7420 9024
rect 5868 8984 5874 8996
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4525 8959 4583 8965
rect 4525 8956 4537 8959
rect 4120 8928 4537 8956
rect 4120 8916 4126 8928
rect 4525 8925 4537 8928
rect 4571 8925 4583 8959
rect 5920 8942 5948 8996
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 4525 8919 4583 8925
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 6880 8928 7144 8956
rect 6880 8916 6886 8928
rect 4798 8848 4804 8900
rect 4856 8848 4862 8900
rect 7009 8891 7067 8897
rect 7009 8888 7021 8891
rect 6932 8860 7021 8888
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 6932 8820 6960 8860
rect 7009 8857 7021 8860
rect 7055 8857 7067 8891
rect 7116 8888 7144 8928
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7248 8928 7573 8956
rect 7248 8916 7254 8928
rect 7561 8925 7573 8928
rect 7607 8956 7619 8959
rect 8202 8956 8208 8968
rect 7607 8928 8208 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8956 8355 8959
rect 9030 8956 9036 8968
rect 8343 8928 9036 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9692 8965 9720 9064
rect 17494 9052 17500 9104
rect 17552 9052 17558 9104
rect 17589 9095 17647 9101
rect 17589 9061 17601 9095
rect 17635 9092 17647 9095
rect 17862 9092 17868 9104
rect 17635 9064 17868 9092
rect 17635 9061 17647 9064
rect 17589 9055 17647 9061
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 20530 9052 20536 9104
rect 20588 9092 20594 9104
rect 22554 9092 22560 9104
rect 20588 9064 22560 9092
rect 20588 9052 20594 9064
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 24765 9095 24823 9101
rect 24765 9061 24777 9095
rect 24811 9092 24823 9095
rect 25590 9092 25596 9104
rect 24811 9064 25596 9092
rect 24811 9061 24823 9064
rect 24765 9055 24823 9061
rect 25590 9052 25596 9064
rect 25648 9052 25654 9104
rect 25869 9095 25927 9101
rect 25869 9061 25881 9095
rect 25915 9092 25927 9095
rect 26234 9092 26240 9104
rect 25915 9064 26240 9092
rect 25915 9061 25927 9064
rect 25869 9055 25927 9061
rect 26234 9052 26240 9064
rect 26292 9052 26298 9104
rect 26786 9052 26792 9104
rect 26844 9052 26850 9104
rect 26970 9052 26976 9104
rect 27028 9052 27034 9104
rect 27065 9095 27123 9101
rect 27065 9061 27077 9095
rect 27111 9061 27123 9095
rect 27065 9055 27123 9061
rect 10042 8984 10048 9036
rect 10100 9024 10106 9036
rect 12710 9024 12716 9036
rect 10100 8996 12716 9024
rect 10100 8984 10106 8996
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 9024 14795 9027
rect 17221 9027 17279 9033
rect 17221 9024 17233 9027
rect 14783 8996 17233 9024
rect 14783 8993 14795 8996
rect 14737 8987 14795 8993
rect 17221 8993 17233 8996
rect 17267 8993 17279 9027
rect 18233 9027 18291 9033
rect 18233 9024 18245 9027
rect 17221 8987 17279 8993
rect 17604 8996 18245 9024
rect 17604 8968 17632 8996
rect 18233 8993 18245 8996
rect 18279 9024 18291 9027
rect 18693 9027 18751 9033
rect 18693 9024 18705 9027
rect 18279 8996 18705 9024
rect 18279 8993 18291 8996
rect 18233 8987 18291 8993
rect 18693 8993 18705 8996
rect 18739 9024 18751 9027
rect 18966 9024 18972 9036
rect 18739 8996 18972 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 18966 8984 18972 8996
rect 19024 8984 19030 9036
rect 20622 8984 20628 9036
rect 20680 9024 20686 9036
rect 21637 9027 21695 9033
rect 21637 9024 21649 9027
rect 20680 8996 21649 9024
rect 20680 8984 20686 8996
rect 21637 8993 21649 8996
rect 21683 8993 21695 9027
rect 21637 8987 21695 8993
rect 25682 8984 25688 9036
rect 25740 8984 25746 9036
rect 26694 8984 26700 9036
rect 26752 9024 26758 9036
rect 26881 9027 26939 9033
rect 26881 9024 26893 9027
rect 26752 8996 26893 9024
rect 26752 8984 26758 8996
rect 26881 8993 26893 8996
rect 26927 8993 26939 9027
rect 26881 8987 26939 8993
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9916 8928 9965 8956
rect 9916 8916 9922 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 11054 8956 11060 8968
rect 10459 8928 11060 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11514 8956 11520 8968
rect 11195 8928 11520 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 7285 8891 7343 8897
rect 7285 8888 7297 8891
rect 7116 8860 7297 8888
rect 7009 8851 7067 8857
rect 7285 8857 7297 8860
rect 7331 8857 7343 8891
rect 7285 8851 7343 8857
rect 7374 8848 7380 8900
rect 7432 8888 7438 8900
rect 7469 8891 7527 8897
rect 7469 8888 7481 8891
rect 7432 8860 7481 8888
rect 7432 8848 7438 8860
rect 7469 8857 7481 8860
rect 7515 8888 7527 8891
rect 8110 8888 8116 8900
rect 7515 8860 8116 8888
rect 7515 8857 7527 8860
rect 7469 8851 7527 8857
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 8386 8848 8392 8900
rect 8444 8888 8450 8900
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 8444 8860 8493 8888
rect 8444 8848 8450 8860
rect 8481 8857 8493 8860
rect 8527 8857 8539 8891
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 8481 8851 8539 8857
rect 9784 8860 10333 8888
rect 7392 8820 7420 8848
rect 6696 8792 7420 8820
rect 6696 8780 6702 8792
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9784 8829 9812 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 11716 8888 11744 8919
rect 12802 8916 12808 8968
rect 12860 8916 12866 8968
rect 14918 8916 14924 8968
rect 14976 8916 14982 8968
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 15930 8956 15936 8968
rect 15151 8928 15936 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 18141 8959 18199 8965
rect 18141 8925 18153 8959
rect 18187 8956 18199 8959
rect 18322 8956 18328 8968
rect 18187 8928 18328 8956
rect 18187 8925 18199 8928
rect 18141 8919 18199 8925
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 18414 8916 18420 8968
rect 18472 8916 18478 8968
rect 18598 8916 18604 8968
rect 18656 8956 18662 8968
rect 19426 8956 19432 8968
rect 18656 8928 19432 8956
rect 18656 8916 18662 8928
rect 19426 8916 19432 8928
rect 19484 8956 19490 8968
rect 19978 8956 19984 8968
rect 19484 8928 19984 8956
rect 19484 8916 19490 8928
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 20254 8916 20260 8968
rect 20312 8956 20318 8968
rect 20916 8965 21036 8966
rect 20916 8959 21051 8965
rect 20916 8956 21005 8959
rect 20312 8938 21005 8956
rect 20312 8928 20944 8938
rect 20312 8916 20318 8928
rect 20993 8925 21005 8938
rect 21039 8925 21051 8959
rect 20993 8919 21051 8925
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8956 21327 8959
rect 21450 8956 21456 8968
rect 21315 8928 21456 8956
rect 21315 8925 21327 8928
rect 21269 8919 21327 8925
rect 21450 8916 21456 8928
rect 21508 8916 21514 8968
rect 21542 8916 21548 8968
rect 21600 8916 21606 8968
rect 23106 8916 23112 8968
rect 23164 8956 23170 8968
rect 24581 8959 24639 8965
rect 24581 8956 24593 8959
rect 23164 8928 24593 8956
rect 23164 8916 23170 8928
rect 24581 8925 24593 8928
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 24670 8916 24676 8968
rect 24728 8916 24734 8968
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 25225 8959 25283 8965
rect 25225 8956 25237 8959
rect 24903 8928 25237 8956
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 25225 8925 25237 8928
rect 25271 8925 25283 8959
rect 25225 8919 25283 8925
rect 25501 8959 25559 8965
rect 25501 8925 25513 8959
rect 25547 8956 25559 8959
rect 25547 8928 26096 8956
rect 25547 8925 25559 8928
rect 25501 8919 25559 8925
rect 12066 8888 12072 8900
rect 11716 8860 12072 8888
rect 10321 8851 10379 8857
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 14461 8891 14519 8897
rect 14461 8857 14473 8891
rect 14507 8888 14519 8891
rect 14826 8888 14832 8900
rect 14507 8860 14832 8888
rect 14507 8857 14519 8860
rect 14461 8851 14519 8857
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 16264 8860 17264 8888
rect 16264 8848 16270 8860
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 8720 8792 9781 8820
rect 8720 8780 8726 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 10137 8823 10195 8829
rect 10137 8789 10149 8823
rect 10183 8820 10195 8823
rect 10410 8820 10416 8832
rect 10183 8792 10416 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 10410 8780 10416 8792
rect 10468 8820 10474 8832
rect 10870 8820 10876 8832
rect 10468 8792 10876 8820
rect 10468 8780 10474 8792
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13412 8792 14105 8820
rect 13412 8780 13418 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 14550 8780 14556 8832
rect 14608 8780 14614 8832
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 17034 8820 17040 8832
rect 15160 8792 17040 8820
rect 15160 8780 15166 8792
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17236 8820 17264 8860
rect 17310 8848 17316 8900
rect 17368 8888 17374 8900
rect 18506 8888 18512 8900
rect 17368 8860 18512 8888
rect 17368 8848 17374 8860
rect 18506 8848 18512 8860
rect 18564 8848 18570 8900
rect 18782 8848 18788 8900
rect 18840 8888 18846 8900
rect 18877 8891 18935 8897
rect 18877 8888 18889 8891
rect 18840 8860 18889 8888
rect 18840 8848 18846 8860
rect 18877 8857 18889 8860
rect 18923 8857 18935 8891
rect 18877 8851 18935 8857
rect 19058 8848 19064 8900
rect 19116 8848 19122 8900
rect 22830 8897 22836 8900
rect 22817 8891 22836 8897
rect 22817 8857 22829 8891
rect 22817 8851 22836 8857
rect 22830 8848 22836 8851
rect 22888 8848 22894 8900
rect 23017 8891 23075 8897
rect 23017 8857 23029 8891
rect 23063 8857 23075 8891
rect 23017 8851 23075 8857
rect 21266 8820 21272 8832
rect 17236 8792 21272 8820
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 22832 8820 22860 8848
rect 21968 8792 22860 8820
rect 21968 8780 21974 8792
rect 22922 8780 22928 8832
rect 22980 8820 22986 8832
rect 23032 8820 23060 8851
rect 23934 8848 23940 8900
rect 23992 8888 23998 8900
rect 24872 8888 24900 8919
rect 23992 8860 24900 8888
rect 23992 8848 23998 8860
rect 22980 8792 23060 8820
rect 22980 8780 22986 8792
rect 24578 8780 24584 8832
rect 24636 8820 24642 8832
rect 26068 8820 26096 8928
rect 26234 8916 26240 8968
rect 26292 8956 26298 8968
rect 27080 8956 27108 9055
rect 27982 8984 27988 9036
rect 28040 8984 28046 9036
rect 28552 9024 28580 9132
rect 28629 9095 28687 9101
rect 28629 9061 28641 9095
rect 28675 9092 28687 9095
rect 29362 9092 29368 9104
rect 28675 9064 29368 9092
rect 28675 9061 28687 9064
rect 28629 9055 28687 9061
rect 28276 8996 28764 9024
rect 26292 8928 27108 8956
rect 27433 8959 27491 8965
rect 26292 8916 26298 8928
rect 27433 8925 27445 8959
rect 27479 8925 27491 8959
rect 27433 8919 27491 8925
rect 26145 8891 26203 8897
rect 26145 8857 26157 8891
rect 26191 8888 26203 8891
rect 26510 8888 26516 8900
rect 26191 8860 26516 8888
rect 26191 8857 26203 8860
rect 26145 8851 26203 8857
rect 26510 8848 26516 8860
rect 26568 8888 26574 8900
rect 27448 8888 27476 8919
rect 27890 8916 27896 8968
rect 27948 8916 27954 8968
rect 28000 8956 28028 8984
rect 28166 8956 28172 8968
rect 28000 8928 28172 8956
rect 28166 8916 28172 8928
rect 28224 8956 28230 8968
rect 28276 8965 28304 8996
rect 28261 8959 28319 8965
rect 28261 8956 28273 8959
rect 28224 8928 28273 8956
rect 28224 8916 28230 8928
rect 28261 8925 28273 8928
rect 28307 8925 28319 8959
rect 28261 8919 28319 8925
rect 28350 8916 28356 8968
rect 28408 8956 28414 8968
rect 28445 8959 28503 8965
rect 28445 8956 28457 8959
rect 28408 8928 28457 8956
rect 28408 8916 28414 8928
rect 28445 8925 28457 8928
rect 28491 8925 28503 8959
rect 28736 8956 28764 8996
rect 29012 8965 29040 9064
rect 29362 9052 29368 9064
rect 29420 9052 29426 9104
rect 29730 9052 29736 9104
rect 29788 9092 29794 9104
rect 30469 9095 30527 9101
rect 30469 9092 30481 9095
rect 29788 9064 30481 9092
rect 29788 9052 29794 9064
rect 30469 9061 30481 9064
rect 30515 9061 30527 9095
rect 30469 9055 30527 9061
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 29236 8996 30604 9024
rect 29236 8984 29242 8996
rect 28997 8959 29055 8965
rect 28736 8928 28948 8956
rect 28445 8919 28503 8925
rect 26568 8860 27476 8888
rect 26568 8848 26574 8860
rect 27798 8848 27804 8900
rect 27856 8888 27862 8900
rect 27985 8891 28043 8897
rect 27985 8888 27997 8891
rect 27856 8860 27997 8888
rect 27856 8848 27862 8860
rect 27985 8857 27997 8860
rect 28031 8857 28043 8891
rect 27985 8851 28043 8857
rect 28077 8891 28135 8897
rect 28077 8857 28089 8891
rect 28123 8888 28135 8891
rect 28810 8888 28816 8900
rect 28123 8860 28816 8888
rect 28123 8857 28135 8860
rect 28077 8851 28135 8857
rect 28810 8848 28816 8860
rect 28868 8848 28874 8900
rect 28920 8888 28948 8928
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 29546 8916 29552 8968
rect 29604 8916 29610 8968
rect 29638 8916 29644 8968
rect 29696 8956 29702 8968
rect 30285 8959 30343 8965
rect 30285 8956 30297 8959
rect 29696 8928 30297 8956
rect 29696 8916 29702 8928
rect 30285 8925 30297 8928
rect 30331 8925 30343 8959
rect 30285 8919 30343 8925
rect 30101 8891 30159 8897
rect 28920 8860 29776 8888
rect 28626 8820 28632 8832
rect 24636 8792 28632 8820
rect 24636 8780 24642 8792
rect 28626 8780 28632 8792
rect 28684 8780 28690 8832
rect 28905 8823 28963 8829
rect 28905 8789 28917 8823
rect 28951 8820 28963 8823
rect 28994 8820 29000 8832
rect 28951 8792 29000 8820
rect 28951 8789 28963 8792
rect 28905 8783 28963 8789
rect 28994 8780 29000 8792
rect 29052 8780 29058 8832
rect 29748 8829 29776 8860
rect 30101 8857 30113 8891
rect 30147 8888 30159 8891
rect 30190 8888 30196 8900
rect 30147 8860 30196 8888
rect 30147 8857 30159 8860
rect 30101 8851 30159 8857
rect 30190 8848 30196 8860
rect 30248 8848 30254 8900
rect 29733 8823 29791 8829
rect 29733 8789 29745 8823
rect 29779 8789 29791 8823
rect 29733 8783 29791 8789
rect 29914 8780 29920 8832
rect 29972 8820 29978 8832
rect 30009 8823 30067 8829
rect 30009 8820 30021 8823
rect 29972 8792 30021 8820
rect 29972 8780 29978 8792
rect 30009 8789 30021 8792
rect 30055 8789 30067 8823
rect 30576 8820 30604 8996
rect 30668 8888 30696 9132
rect 31389 9129 31401 9163
rect 31435 9160 31447 9163
rect 31570 9160 31576 9172
rect 31435 9132 31576 9160
rect 31435 9129 31447 9132
rect 31389 9123 31447 9129
rect 31570 9120 31576 9132
rect 31628 9120 31634 9172
rect 32674 9120 32680 9172
rect 32732 9160 32738 9172
rect 32769 9163 32827 9169
rect 32769 9160 32781 9163
rect 32732 9132 32781 9160
rect 32732 9120 32738 9132
rect 32769 9129 32781 9132
rect 32815 9160 32827 9163
rect 33594 9160 33600 9172
rect 32815 9132 33600 9160
rect 32815 9129 32827 9132
rect 32769 9123 32827 9129
rect 33594 9120 33600 9132
rect 33652 9120 33658 9172
rect 33505 9095 33563 9101
rect 32876 9064 33272 9092
rect 31386 8984 31392 9036
rect 31444 9024 31450 9036
rect 32033 9027 32091 9033
rect 32033 9024 32045 9027
rect 31444 8996 32045 9024
rect 31444 8984 31450 8996
rect 32033 8993 32045 8996
rect 32079 8993 32091 9027
rect 32033 8987 32091 8993
rect 32490 8984 32496 9036
rect 32548 9024 32554 9036
rect 32876 9024 32904 9064
rect 32548 8996 32904 9024
rect 32548 8984 32554 8996
rect 31202 8916 31208 8968
rect 31260 8956 31266 8968
rect 31573 8959 31631 8965
rect 31573 8956 31585 8959
rect 31260 8928 31585 8956
rect 31260 8916 31266 8928
rect 31573 8925 31585 8928
rect 31619 8925 31631 8959
rect 31573 8919 31631 8925
rect 31662 8916 31668 8968
rect 31720 8916 31726 8968
rect 31757 8959 31815 8965
rect 31757 8925 31769 8959
rect 31803 8956 31815 8959
rect 33134 8956 33140 8968
rect 31803 8928 33140 8956
rect 31803 8925 31815 8928
rect 31757 8919 31815 8925
rect 31772 8888 31800 8919
rect 33134 8916 33140 8928
rect 33192 8916 33198 8968
rect 33244 8956 33272 9064
rect 33505 9061 33517 9095
rect 33551 9092 33563 9095
rect 33870 9092 33876 9104
rect 33551 9064 33876 9092
rect 33551 9061 33563 9064
rect 33505 9055 33563 9061
rect 33870 9052 33876 9064
rect 33928 9052 33934 9104
rect 35986 8956 35992 8968
rect 33244 8928 35992 8956
rect 35986 8916 35992 8928
rect 36044 8916 36050 8968
rect 30668 8860 31800 8888
rect 31895 8891 31953 8897
rect 31895 8857 31907 8891
rect 31941 8888 31953 8891
rect 32858 8888 32864 8900
rect 31941 8860 32864 8888
rect 31941 8857 31953 8860
rect 31895 8851 31953 8857
rect 32858 8848 32864 8860
rect 32916 8848 32922 8900
rect 32968 8860 33364 8888
rect 32490 8820 32496 8832
rect 30576 8792 32496 8820
rect 30009 8783 30067 8789
rect 32490 8780 32496 8792
rect 32548 8780 32554 8832
rect 32674 8780 32680 8832
rect 32732 8820 32738 8832
rect 32968 8829 32996 8860
rect 32953 8823 33011 8829
rect 32953 8820 32965 8823
rect 32732 8792 32965 8820
rect 32732 8780 32738 8792
rect 32953 8789 32965 8792
rect 32999 8789 33011 8823
rect 32953 8783 33011 8789
rect 33042 8780 33048 8832
rect 33100 8780 33106 8832
rect 33336 8820 33364 8860
rect 33502 8848 33508 8900
rect 33560 8848 33566 8900
rect 34974 8820 34980 8832
rect 33336 8792 34980 8820
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 1104 8730 36524 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 36524 8730
rect 1104 8656 36524 8678
rect 4798 8576 4804 8628
rect 4856 8616 4862 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 4856 8588 5549 8616
rect 4856 8576 4862 8588
rect 5537 8585 5549 8588
rect 5583 8585 5595 8619
rect 5537 8579 5595 8585
rect 9030 8576 9036 8628
rect 9088 8576 9094 8628
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 15194 8616 15200 8628
rect 12124 8588 15200 8616
rect 12124 8576 12130 8588
rect 9122 8508 9128 8560
rect 9180 8548 9186 8560
rect 10502 8548 10508 8560
rect 9180 8520 9536 8548
rect 9180 8508 9186 8520
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 6730 8480 6736 8492
rect 5307 8452 6736 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7098 8480 7104 8492
rect 6871 8452 7104 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 8294 8440 8300 8492
rect 8352 8440 8358 8492
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 9398 8440 9404 8492
rect 9456 8440 9462 8492
rect 9508 8480 9536 8520
rect 10060 8520 10508 8548
rect 10060 8489 10088 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 12802 8548 12808 8560
rect 12483 8520 12808 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 12802 8508 12808 8520
rect 12860 8508 12866 8560
rect 10045 8483 10103 8489
rect 9508 8452 9996 8480
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5718 8412 5724 8424
rect 5583 8384 5724 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 6914 8372 6920 8424
rect 6972 8372 6978 8424
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7190 8412 7196 8424
rect 7055 8384 7196 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 7837 8415 7895 8421
rect 7837 8381 7849 8415
rect 7883 8381 7895 8415
rect 7837 8375 7895 8381
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 5399 8316 6469 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 6457 8313 6469 8316
rect 6503 8313 6515 8347
rect 6932 8344 6960 8372
rect 7852 8344 7880 8375
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9968 8412 9996 8452
rect 10045 8449 10057 8483
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10336 8412 10364 8443
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11330 8480 11336 8492
rect 11020 8452 11336 8480
rect 11020 8440 11026 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 13096 8489 13124 8588
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 17678 8616 17684 8628
rect 16776 8588 17684 8616
rect 13354 8508 13360 8560
rect 13412 8508 13418 8560
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 13081 8443 13139 8449
rect 14458 8440 14464 8492
rect 14516 8440 14522 8492
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 16025 8483 16083 8489
rect 16025 8480 16037 8483
rect 14700 8452 16037 8480
rect 14700 8440 14706 8452
rect 16025 8449 16037 8452
rect 16071 8449 16083 8483
rect 16025 8443 16083 8449
rect 16206 8440 16212 8492
rect 16264 8440 16270 8492
rect 16776 8489 16804 8588
rect 16945 8493 17003 8499
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16945 8459 16957 8493
rect 16991 8459 17003 8493
rect 17328 8489 17356 8588
rect 17678 8576 17684 8588
rect 17736 8616 17742 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 17736 8588 17969 8616
rect 17736 8576 17742 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 18690 8576 18696 8628
rect 18748 8576 18754 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 21174 8616 21180 8628
rect 19484 8588 21180 8616
rect 19484 8576 19490 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 21692 8588 22232 8616
rect 21692 8576 21698 8588
rect 18414 8548 18420 8560
rect 17788 8520 18420 8548
rect 16945 8453 17003 8459
rect 17313 8483 17371 8489
rect 16761 8443 16819 8449
rect 9968 8384 10364 8412
rect 9585 8375 9643 8381
rect 9306 8344 9312 8356
rect 6932 8316 7880 8344
rect 8220 8316 9312 8344
rect 6457 8307 6515 8313
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 8220 8276 8248 8316
rect 9306 8304 9312 8316
rect 9364 8344 9370 8356
rect 9600 8344 9628 8375
rect 10870 8372 10876 8424
rect 10928 8372 10934 8424
rect 11514 8372 11520 8424
rect 11572 8412 11578 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11572 8384 11621 8412
rect 11572 8372 11578 8384
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 14734 8412 14740 8424
rect 11609 8375 11667 8381
rect 12406 8384 14740 8412
rect 9364 8316 9628 8344
rect 9364 8304 9370 8316
rect 10134 8304 10140 8356
rect 10192 8304 10198 8356
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 10505 8347 10563 8353
rect 10505 8313 10517 8347
rect 10551 8344 10563 8347
rect 12406 8344 12434 8384
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 14826 8372 14832 8424
rect 14884 8372 14890 8424
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 16776 8412 16804 8443
rect 14976 8384 16804 8412
rect 16960 8412 16988 8453
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17494 8480 17500 8492
rect 17451 8452 17500 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17788 8489 17816 8520
rect 18414 8508 18420 8520
rect 18472 8508 18478 8560
rect 19150 8508 19156 8560
rect 19208 8548 19214 8560
rect 19208 8520 19472 8548
rect 19208 8508 19214 8520
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 18104 8452 18153 8480
rect 18104 8440 18110 8452
rect 18141 8449 18153 8452
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18322 8440 18328 8492
rect 18380 8440 18386 8492
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 16960 8384 17724 8412
rect 14976 8372 14982 8384
rect 17696 8356 17724 8384
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18233 8415 18291 8421
rect 18233 8412 18245 8415
rect 18012 8384 18245 8412
rect 18012 8372 18018 8384
rect 18233 8381 18245 8384
rect 18279 8381 18291 8415
rect 18233 8375 18291 8381
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 10551 8316 12434 8344
rect 14384 8316 17049 8344
rect 10551 8313 10563 8316
rect 10505 8307 10563 8313
rect 7340 8248 8248 8276
rect 7340 8236 7346 8248
rect 10686 8236 10692 8288
rect 10744 8236 10750 8288
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14384 8276 14412 8316
rect 17037 8313 17049 8316
rect 17083 8313 17095 8347
rect 17037 8307 17095 8313
rect 17402 8304 17408 8356
rect 17460 8304 17466 8356
rect 17494 8304 17500 8356
rect 17552 8304 17558 8356
rect 17589 8347 17647 8353
rect 17589 8313 17601 8347
rect 17635 8313 17647 8347
rect 17589 8307 17647 8313
rect 13964 8248 14412 8276
rect 13964 8236 13970 8248
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 15102 8276 15108 8288
rect 14792 8248 15108 8276
rect 14792 8236 14798 8248
rect 15102 8236 15108 8248
rect 15160 8236 15166 8288
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 16080 8248 16129 8276
rect 16080 8236 16086 8248
rect 16117 8245 16129 8248
rect 16163 8245 16175 8279
rect 16117 8239 16175 8245
rect 16850 8236 16856 8288
rect 16908 8236 16914 8288
rect 17420 8276 17448 8304
rect 17604 8276 17632 8307
rect 17678 8304 17684 8356
rect 17736 8344 17742 8356
rect 18969 8347 19027 8353
rect 18969 8344 18981 8347
rect 17736 8316 18981 8344
rect 17736 8304 17742 8316
rect 18969 8313 18981 8316
rect 19015 8313 19027 8347
rect 18969 8307 19027 8313
rect 17420 8248 17632 8276
rect 19260 8294 19288 8443
rect 19334 8440 19340 8492
rect 19392 8440 19398 8492
rect 19444 8489 19472 8520
rect 19518 8508 19524 8560
rect 19576 8548 19582 8560
rect 20714 8548 20720 8560
rect 19576 8520 20116 8548
rect 19576 8508 19582 8520
rect 20088 8489 20116 8520
rect 20548 8520 20720 8548
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8480 20131 8483
rect 20438 8480 20444 8492
rect 20119 8452 20444 8480
rect 20119 8449 20131 8452
rect 20073 8443 20131 8449
rect 19628 8412 19656 8443
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20548 8489 20576 8520
rect 20714 8508 20720 8520
rect 20772 8548 20778 8560
rect 21450 8548 21456 8560
rect 20772 8520 21456 8548
rect 20772 8508 20778 8520
rect 21450 8508 21456 8520
rect 21508 8548 21514 8560
rect 22204 8557 22232 8588
rect 22554 8576 22560 8628
rect 22612 8576 22618 8628
rect 22738 8576 22744 8628
rect 22796 8576 22802 8628
rect 24394 8616 24400 8628
rect 24044 8588 24400 8616
rect 22189 8551 22247 8557
rect 21508 8520 22032 8548
rect 21508 8508 21514 8520
rect 21959 8517 22032 8520
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8449 20591 8483
rect 20533 8443 20591 8449
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20680 8452 20821 8480
rect 20680 8440 20686 8452
rect 20809 8449 20821 8452
rect 20855 8480 20867 8483
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20855 8452 20913 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 20901 8449 20913 8452
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 21959 8483 21971 8517
rect 22005 8483 22032 8517
rect 22189 8517 22201 8551
rect 22235 8517 22247 8551
rect 22572 8548 22600 8576
rect 23842 8548 23848 8560
rect 22572 8520 23848 8548
rect 22189 8511 22247 8517
rect 23842 8508 23848 8520
rect 23900 8508 23906 8560
rect 21959 8480 22032 8483
rect 21407 8452 21680 8480
rect 21959 8477 22140 8480
rect 22004 8452 22140 8477
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 20714 8412 20720 8424
rect 19628 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 21177 8415 21235 8421
rect 21177 8381 21189 8415
rect 21223 8412 21235 8415
rect 21542 8412 21548 8424
rect 21223 8384 21548 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 21652 8412 21680 8452
rect 22002 8412 22008 8424
rect 21652 8384 22008 8412
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 22112 8412 22140 8452
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 22462 8440 22468 8492
rect 22520 8440 22526 8492
rect 22557 8483 22615 8489
rect 22557 8449 22569 8483
rect 22603 8480 22615 8483
rect 23753 8483 23811 8489
rect 23753 8480 23765 8483
rect 22603 8452 23765 8480
rect 22603 8449 22615 8452
rect 22557 8443 22615 8449
rect 23753 8449 23765 8452
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 24044 8412 24072 8588
rect 24394 8576 24400 8588
rect 24452 8576 24458 8628
rect 24670 8576 24676 8628
rect 24728 8616 24734 8628
rect 24765 8619 24823 8625
rect 24765 8616 24777 8619
rect 24728 8588 24777 8616
rect 24728 8576 24734 8588
rect 24765 8585 24777 8588
rect 24811 8585 24823 8619
rect 24765 8579 24823 8585
rect 27065 8619 27123 8625
rect 27065 8585 27077 8619
rect 27111 8616 27123 8619
rect 27246 8616 27252 8628
rect 27111 8588 27252 8616
rect 27111 8585 27123 8588
rect 27065 8579 27123 8585
rect 27246 8576 27252 8588
rect 27304 8576 27310 8628
rect 28169 8619 28227 8625
rect 28169 8585 28181 8619
rect 28215 8616 28227 8619
rect 28534 8616 28540 8628
rect 28215 8588 28540 8616
rect 28215 8585 28227 8588
rect 28169 8579 28227 8585
rect 28534 8576 28540 8588
rect 28592 8576 28598 8628
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 29089 8619 29147 8625
rect 29089 8616 29101 8619
rect 28684 8588 29101 8616
rect 28684 8576 28690 8588
rect 29089 8585 29101 8588
rect 29135 8585 29147 8619
rect 30466 8616 30472 8628
rect 29089 8579 29147 8585
rect 29748 8588 30472 8616
rect 24688 8548 24716 8576
rect 24228 8520 24716 8548
rect 24228 8489 24256 8520
rect 25498 8508 25504 8560
rect 25556 8548 25562 8560
rect 29748 8557 29776 8588
rect 30466 8576 30472 8588
rect 30524 8576 30530 8628
rect 31202 8576 31208 8628
rect 31260 8616 31266 8628
rect 31754 8616 31760 8628
rect 31260 8588 31760 8616
rect 31260 8576 31266 8588
rect 31754 8576 31760 8588
rect 31812 8616 31818 8628
rect 31812 8588 32720 8616
rect 31812 8576 31818 8588
rect 25777 8551 25835 8557
rect 25777 8548 25789 8551
rect 25556 8520 25789 8548
rect 25556 8508 25562 8520
rect 25777 8517 25789 8520
rect 25823 8517 25835 8551
rect 29733 8551 29791 8557
rect 25777 8511 25835 8517
rect 25976 8520 29684 8548
rect 24209 8483 24267 8489
rect 24209 8449 24221 8483
rect 24255 8449 24267 8483
rect 24209 8443 24267 8449
rect 24394 8440 24400 8492
rect 24452 8440 24458 8492
rect 24578 8440 24584 8492
rect 24636 8440 24642 8492
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 24820 8452 24869 8480
rect 24820 8440 24826 8452
rect 24857 8449 24869 8452
rect 24903 8480 24915 8483
rect 25866 8480 25872 8492
rect 24903 8452 25872 8480
rect 24903 8449 24915 8452
rect 24857 8443 24915 8449
rect 25866 8440 25872 8452
rect 25924 8440 25930 8492
rect 22112 8384 24072 8412
rect 24118 8372 24124 8424
rect 24176 8412 24182 8424
rect 24176 8404 24256 8412
rect 24305 8407 24363 8413
rect 24305 8404 24317 8407
rect 24176 8384 24317 8404
rect 24176 8372 24182 8384
rect 24228 8376 24317 8384
rect 24305 8373 24317 8376
rect 24351 8373 24363 8407
rect 24412 8412 24440 8440
rect 25976 8412 26004 8520
rect 26605 8483 26663 8489
rect 26605 8449 26617 8483
rect 26651 8480 26663 8483
rect 26786 8480 26792 8492
rect 26651 8452 26792 8480
rect 26651 8449 26663 8452
rect 26605 8443 26663 8449
rect 26786 8440 26792 8452
rect 26844 8480 26850 8492
rect 26970 8480 26976 8492
rect 26844 8452 26976 8480
rect 26844 8440 26850 8452
rect 26970 8440 26976 8452
rect 27028 8480 27034 8492
rect 27801 8483 27859 8489
rect 27801 8480 27813 8483
rect 27028 8452 27813 8480
rect 27028 8440 27034 8452
rect 27801 8449 27813 8452
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 28626 8480 28632 8492
rect 27939 8452 28632 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 24412 8384 26004 8412
rect 26145 8415 26203 8421
rect 26145 8381 26157 8415
rect 26191 8412 26203 8415
rect 26234 8412 26240 8424
rect 26191 8384 26240 8412
rect 26191 8381 26203 8384
rect 26145 8375 26203 8381
rect 24305 8367 24363 8373
rect 26234 8372 26240 8384
rect 26292 8372 26298 8424
rect 26694 8372 26700 8424
rect 26752 8372 26758 8424
rect 27356 8421 27476 8423
rect 27341 8415 27476 8421
rect 27341 8381 27353 8415
rect 27387 8412 27476 8415
rect 27816 8412 27844 8443
rect 28626 8440 28632 8452
rect 28684 8440 28690 8492
rect 28810 8440 28816 8492
rect 28868 8480 28874 8492
rect 29273 8483 29331 8489
rect 29273 8480 29285 8483
rect 28868 8452 29285 8480
rect 28868 8440 28874 8452
rect 29273 8449 29285 8452
rect 29319 8449 29331 8483
rect 29656 8480 29684 8520
rect 29733 8517 29745 8551
rect 29779 8517 29791 8551
rect 29733 8511 29791 8517
rect 29822 8508 29828 8560
rect 29880 8548 29886 8560
rect 30282 8548 30288 8560
rect 29880 8520 30288 8548
rect 29880 8508 29886 8520
rect 30282 8508 30288 8520
rect 30340 8508 30346 8560
rect 30377 8551 30435 8557
rect 30377 8517 30389 8551
rect 30423 8548 30435 8551
rect 30423 8520 31064 8548
rect 30423 8517 30435 8520
rect 30377 8511 30435 8517
rect 30098 8480 30104 8492
rect 29656 8452 30104 8480
rect 29273 8443 29331 8449
rect 30098 8440 30104 8452
rect 30156 8440 30162 8492
rect 30190 8440 30196 8492
rect 30248 8480 30254 8492
rect 30926 8480 30932 8492
rect 30248 8452 30932 8480
rect 30248 8440 30254 8452
rect 30926 8440 30932 8452
rect 30984 8440 30990 8492
rect 31036 8489 31064 8520
rect 32692 8492 32720 8588
rect 33410 8576 33416 8628
rect 33468 8616 33474 8628
rect 33597 8619 33655 8625
rect 33597 8616 33609 8619
rect 33468 8588 33609 8616
rect 33468 8576 33474 8588
rect 33597 8585 33609 8588
rect 33643 8585 33655 8619
rect 33597 8579 33655 8585
rect 33870 8576 33876 8628
rect 33928 8616 33934 8628
rect 34333 8619 34391 8625
rect 34333 8616 34345 8619
rect 33928 8588 34345 8616
rect 33928 8576 33934 8588
rect 34333 8585 34345 8588
rect 34379 8585 34391 8619
rect 34333 8579 34391 8585
rect 34974 8576 34980 8628
rect 35032 8576 35038 8628
rect 34514 8508 34520 8560
rect 34572 8548 34578 8560
rect 35069 8551 35127 8557
rect 35069 8548 35081 8551
rect 34572 8520 35081 8548
rect 34572 8508 34578 8520
rect 35069 8517 35081 8520
rect 35115 8517 35127 8551
rect 35069 8511 35127 8517
rect 31021 8483 31079 8489
rect 31021 8449 31033 8483
rect 31067 8449 31079 8483
rect 31021 8443 31079 8449
rect 31113 8483 31171 8489
rect 31113 8449 31125 8483
rect 31159 8480 31171 8483
rect 31386 8480 31392 8492
rect 31159 8452 31392 8480
rect 31159 8449 31171 8452
rect 31113 8443 31171 8449
rect 28445 8415 28503 8421
rect 28445 8412 28457 8415
rect 27387 8395 27752 8412
rect 27387 8381 27399 8395
rect 27448 8384 27752 8395
rect 27816 8384 28457 8412
rect 27341 8375 27399 8381
rect 27724 8356 27752 8384
rect 28445 8381 28457 8384
rect 28491 8381 28503 8415
rect 28445 8375 28503 8381
rect 28534 8372 28540 8424
rect 28592 8412 28598 8424
rect 28902 8412 28908 8424
rect 28592 8384 28908 8412
rect 28592 8372 28598 8384
rect 28902 8372 28908 8384
rect 28960 8372 28966 8424
rect 29086 8372 29092 8424
rect 29144 8412 29150 8424
rect 29457 8415 29515 8421
rect 29457 8412 29469 8415
rect 29144 8384 29469 8412
rect 29144 8372 29150 8384
rect 29457 8381 29469 8384
rect 29503 8381 29515 8415
rect 29457 8375 29515 8381
rect 29822 8372 29828 8424
rect 29880 8372 29886 8424
rect 31036 8412 31064 8443
rect 31386 8440 31392 8452
rect 31444 8480 31450 8492
rect 31444 8452 31800 8480
rect 31444 8440 31450 8452
rect 31036 8384 31340 8412
rect 19518 8304 19524 8356
rect 19576 8344 19582 8356
rect 20257 8347 20315 8353
rect 20257 8344 20269 8347
rect 19576 8316 20269 8344
rect 19576 8304 19582 8316
rect 20257 8313 20269 8316
rect 20303 8313 20315 8347
rect 20257 8307 20315 8313
rect 20349 8347 20407 8353
rect 20349 8313 20361 8347
rect 20395 8344 20407 8347
rect 20530 8344 20536 8356
rect 20395 8316 20536 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 20530 8304 20536 8316
rect 20588 8304 20594 8356
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 20956 8316 21281 8344
rect 20956 8304 20962 8316
rect 21269 8313 21281 8316
rect 21315 8344 21327 8347
rect 21637 8347 21695 8353
rect 21315 8316 21588 8344
rect 21315 8313 21327 8316
rect 21269 8307 21327 8313
rect 19260 8276 19334 8294
rect 19610 8276 19616 8288
rect 19260 8266 19616 8276
rect 19306 8248 19616 8266
rect 19610 8236 19616 8248
rect 19668 8276 19674 8288
rect 20070 8276 20076 8288
rect 19668 8248 20076 8276
rect 19668 8236 19674 8248
rect 20070 8236 20076 8248
rect 20128 8276 20134 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 20128 8248 20453 8276
rect 20128 8236 20134 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 21560 8276 21588 8316
rect 21637 8313 21649 8347
rect 21683 8344 21695 8347
rect 21683 8316 22324 8344
rect 21683 8313 21695 8316
rect 21637 8307 21695 8313
rect 21821 8279 21879 8285
rect 21821 8276 21833 8279
rect 21560 8248 21833 8276
rect 20441 8239 20499 8245
rect 21821 8245 21833 8248
rect 21867 8245 21879 8279
rect 21821 8239 21879 8245
rect 22002 8236 22008 8288
rect 22060 8236 22066 8288
rect 22296 8285 22324 8316
rect 24394 8304 24400 8356
rect 24452 8304 24458 8356
rect 24489 8347 24547 8353
rect 24489 8313 24501 8347
rect 24535 8344 24547 8347
rect 25498 8344 25504 8356
rect 24535 8316 25504 8344
rect 24535 8313 24547 8316
rect 24489 8307 24547 8313
rect 22281 8279 22339 8285
rect 22281 8245 22293 8279
rect 22327 8245 22339 8279
rect 22281 8239 22339 8245
rect 24121 8279 24179 8285
rect 24121 8245 24133 8279
rect 24167 8276 24179 8279
rect 24504 8276 24532 8307
rect 25498 8304 25504 8316
rect 25556 8304 25562 8356
rect 27706 8304 27712 8356
rect 27764 8344 27770 8356
rect 28997 8347 29055 8353
rect 28997 8344 29009 8347
rect 27764 8316 29009 8344
rect 27764 8304 27770 8316
rect 28997 8313 29009 8316
rect 29043 8344 29055 8347
rect 31202 8344 31208 8356
rect 29043 8316 31208 8344
rect 29043 8313 29055 8316
rect 28997 8307 29055 8313
rect 31202 8304 31208 8316
rect 31260 8304 31266 8356
rect 31312 8344 31340 8384
rect 31478 8372 31484 8424
rect 31536 8372 31542 8424
rect 31665 8415 31723 8421
rect 31665 8381 31677 8415
rect 31711 8381 31723 8415
rect 31772 8412 31800 8452
rect 32674 8440 32680 8492
rect 32732 8440 32738 8492
rect 33045 8483 33103 8489
rect 33045 8480 33057 8483
rect 32876 8452 33057 8480
rect 32876 8412 32904 8452
rect 33045 8449 33057 8452
rect 33091 8449 33103 8483
rect 33045 8443 33103 8449
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8449 33471 8483
rect 33413 8443 33471 8449
rect 31772 8384 32904 8412
rect 33428 8412 33456 8443
rect 33502 8440 33508 8492
rect 33560 8480 33566 8492
rect 33597 8483 33655 8489
rect 33597 8480 33609 8483
rect 33560 8452 33609 8480
rect 33560 8440 33566 8452
rect 33597 8449 33609 8452
rect 33643 8449 33655 8483
rect 33597 8443 33655 8449
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 34790 8440 34796 8492
rect 34848 8440 34854 8492
rect 34164 8412 34192 8440
rect 33428 8384 34192 8412
rect 31665 8375 31723 8381
rect 31570 8344 31576 8356
rect 31312 8316 31576 8344
rect 31570 8304 31576 8316
rect 31628 8304 31634 8356
rect 24167 8248 24532 8276
rect 26237 8279 26295 8285
rect 24167 8245 24179 8248
rect 24121 8239 24179 8245
rect 26237 8245 26249 8279
rect 26283 8276 26295 8279
rect 26510 8276 26516 8288
rect 26283 8248 26516 8276
rect 26283 8245 26295 8248
rect 26237 8239 26295 8245
rect 26510 8236 26516 8248
rect 26568 8236 26574 8288
rect 27433 8279 27491 8285
rect 27433 8245 27445 8279
rect 27479 8276 27491 8279
rect 27982 8276 27988 8288
rect 27479 8248 27988 8276
rect 27479 8245 27491 8248
rect 27433 8239 27491 8245
rect 27982 8236 27988 8248
rect 28040 8236 28046 8288
rect 28534 8236 28540 8288
rect 28592 8236 28598 8288
rect 28626 8236 28632 8288
rect 28684 8236 28690 8288
rect 31018 8236 31024 8288
rect 31076 8276 31082 8288
rect 31680 8276 31708 8375
rect 32876 8356 32904 8384
rect 32858 8304 32864 8356
rect 32916 8304 32922 8356
rect 33042 8304 33048 8356
rect 33100 8344 33106 8356
rect 34057 8347 34115 8353
rect 34057 8344 34069 8347
rect 33100 8316 34069 8344
rect 33100 8304 33106 8316
rect 34057 8313 34069 8316
rect 34103 8344 34115 8347
rect 34238 8344 34244 8356
rect 34103 8316 34244 8344
rect 34103 8313 34115 8316
rect 34057 8307 34115 8313
rect 34238 8304 34244 8316
rect 34296 8344 34302 8356
rect 34609 8347 34667 8353
rect 34609 8344 34621 8347
rect 34296 8316 34621 8344
rect 34296 8304 34302 8316
rect 34609 8313 34621 8316
rect 34655 8313 34667 8347
rect 34609 8307 34667 8313
rect 33502 8276 33508 8288
rect 31076 8248 33508 8276
rect 31076 8236 31082 8248
rect 33502 8236 33508 8248
rect 33560 8236 33566 8288
rect 1104 8186 36524 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 36524 8186
rect 1104 8112 36524 8134
rect 7098 8032 7104 8084
rect 7156 8032 7162 8084
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 8536 8044 9229 8072
rect 8536 8032 8542 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9548 8044 9689 8072
rect 9548 8032 9554 8044
rect 8113 8007 8171 8013
rect 8113 7973 8125 8007
rect 8159 8004 8171 8007
rect 9398 8004 9404 8016
rect 8159 7976 9404 8004
rect 8159 7973 8171 7976
rect 8113 7967 8171 7973
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 9600 8004 9628 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9677 8035 9735 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 9916 8044 9965 8072
rect 9916 8032 9922 8044
rect 9953 8041 9965 8044
rect 9999 8072 10011 8075
rect 10134 8072 10140 8084
rect 9999 8044 10140 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 10284 8044 10517 8072
rect 10284 8032 10290 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 11440 8044 13400 8072
rect 9600 7976 10548 8004
rect 6638 7896 6644 7948
rect 6696 7896 6702 7948
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 6963 7908 7297 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 8205 7939 8263 7945
rect 8205 7936 8217 7939
rect 7285 7899 7343 7905
rect 7944 7908 8217 7936
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6564 7800 6592 7831
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 7944 7877 7972 7908
rect 8205 7905 8217 7908
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 9600 7936 9628 7976
rect 8619 7908 9628 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 6914 7800 6920 7812
rect 6564 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7800 6978 7812
rect 7944 7800 7972 7831
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8168 7840 8401 7868
rect 8168 7828 8174 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9033 7871 9091 7877
rect 9033 7837 9045 7871
rect 9079 7868 9091 7871
rect 9122 7868 9128 7880
rect 9079 7840 9128 7868
rect 9079 7837 9091 7840
rect 9033 7831 9091 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9263 7840 9781 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 6972 7772 7972 7800
rect 9784 7800 9812 7831
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 10318 7868 10324 7880
rect 10183 7840 10324 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 10520 7877 10548 7976
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 11146 7828 11152 7880
rect 11204 7828 11210 7880
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11440 7877 11468 8044
rect 13372 8004 13400 8044
rect 13446 8032 13452 8084
rect 13504 8032 13510 8084
rect 13630 8032 13636 8084
rect 13688 8072 13694 8084
rect 14734 8072 14740 8084
rect 13688 8044 14740 8072
rect 13688 8032 13694 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 16850 8072 16856 8084
rect 16623 8044 16856 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 17310 8032 17316 8084
rect 17368 8032 17374 8084
rect 18877 8075 18935 8081
rect 18877 8041 18889 8075
rect 18923 8041 18935 8075
rect 18877 8035 18935 8041
rect 13648 8004 13676 8032
rect 15381 8007 15439 8013
rect 15381 8004 15393 8007
rect 13372 7976 13676 8004
rect 14660 7976 15393 8004
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 14660 7877 14688 7976
rect 15381 7973 15393 7976
rect 15427 7973 15439 8007
rect 18892 8004 18920 8035
rect 19058 8032 19064 8084
rect 19116 8072 19122 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 19116 8044 19257 8072
rect 19116 8032 19122 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19426 8072 19432 8084
rect 19245 8035 19303 8041
rect 19352 8044 19432 8072
rect 19352 8004 19380 8044
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 20990 8032 20996 8084
rect 21048 8032 21054 8084
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 21542 8072 21548 8084
rect 21407 8044 21548 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 24026 8072 24032 8084
rect 21652 8044 24032 8072
rect 18892 7976 19380 8004
rect 15381 7967 15439 7973
rect 16022 7896 16028 7948
rect 16080 7896 16086 7948
rect 19334 7936 19340 7948
rect 19076 7908 19340 7936
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11572 7840 11713 7868
rect 11572 7828 11578 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 14738 7871 14796 7877
rect 14738 7837 14750 7871
rect 14784 7837 14796 7871
rect 14738 7831 14796 7837
rect 10704 7800 10732 7828
rect 9784 7772 10732 7800
rect 11348 7800 11376 7828
rect 11348 7772 11836 7800
rect 6972 7760 6978 7772
rect 11808 7744 11836 7772
rect 11974 7760 11980 7812
rect 12032 7760 12038 7812
rect 14458 7800 14464 7812
rect 13202 7772 14464 7800
rect 14458 7760 14464 7772
rect 14516 7760 14522 7812
rect 14752 7800 14780 7831
rect 15102 7828 15108 7880
rect 15160 7877 15166 7880
rect 15160 7868 15168 7877
rect 15160 7840 15205 7868
rect 15160 7831 15168 7840
rect 15160 7828 15166 7831
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 15344 7840 16221 7868
rect 15344 7828 15350 7840
rect 16209 7837 16221 7840
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 17126 7868 17132 7880
rect 16632 7840 17132 7868
rect 16632 7828 16638 7840
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17678 7828 17684 7880
rect 17736 7828 17742 7880
rect 14826 7800 14832 7812
rect 14752 7772 14832 7800
rect 14826 7760 14832 7772
rect 14884 7760 14890 7812
rect 14918 7760 14924 7812
rect 14976 7760 14982 7812
rect 15013 7803 15071 7809
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 15304 7800 15332 7828
rect 15059 7772 15332 7800
rect 15841 7803 15899 7809
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15841 7769 15853 7803
rect 15887 7800 15899 7803
rect 15887 7772 16804 7800
rect 15887 7769 15899 7772
rect 15841 7763 15899 7769
rect 8202 7692 8208 7744
rect 8260 7732 8266 7744
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 8260 7704 9505 7732
rect 8260 7692 8266 7704
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 9493 7695 9551 7701
rect 10321 7735 10379 7741
rect 10321 7701 10333 7735
rect 10367 7732 10379 7735
rect 10962 7732 10968 7744
rect 10367 7704 10968 7732
rect 10367 7701 10379 7704
rect 10321 7695 10379 7701
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11514 7692 11520 7744
rect 11572 7732 11578 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11572 7704 11621 7732
rect 11572 7692 11578 7704
rect 11609 7701 11621 7704
rect 11655 7701 11667 7735
rect 11609 7695 11667 7701
rect 11790 7692 11796 7744
rect 11848 7692 11854 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 14550 7732 14556 7744
rect 11940 7704 14556 7732
rect 11940 7692 11946 7704
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 15286 7692 15292 7744
rect 15344 7692 15350 7744
rect 15746 7692 15752 7744
rect 15804 7692 15810 7744
rect 16574 7692 16580 7744
rect 16632 7692 16638 7744
rect 16776 7741 16804 7772
rect 16942 7760 16948 7812
rect 17000 7800 17006 7812
rect 19076 7809 19104 7908
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 21652 7936 21680 8044
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 26786 8032 26792 8084
rect 26844 8032 26850 8084
rect 27062 8032 27068 8084
rect 27120 8072 27126 8084
rect 27157 8075 27215 8081
rect 27157 8072 27169 8075
rect 27120 8044 27169 8072
rect 27120 8032 27126 8044
rect 27157 8041 27169 8044
rect 27203 8041 27215 8075
rect 27157 8035 27215 8041
rect 28537 8075 28595 8081
rect 28537 8041 28549 8075
rect 28583 8072 28595 8075
rect 28810 8072 28816 8084
rect 28583 8044 28816 8072
rect 28583 8041 28595 8044
rect 28537 8035 28595 8041
rect 28810 8032 28816 8044
rect 28868 8032 28874 8084
rect 28905 8075 28963 8081
rect 28905 8041 28917 8075
rect 28951 8072 28963 8075
rect 29178 8072 29184 8084
rect 28951 8044 29184 8072
rect 28951 8041 28963 8044
rect 28905 8035 28963 8041
rect 29178 8032 29184 8044
rect 29236 8032 29242 8084
rect 29270 8032 29276 8084
rect 29328 8072 29334 8084
rect 36538 8072 36544 8084
rect 29328 8044 36544 8072
rect 29328 8032 29334 8044
rect 36538 8032 36544 8044
rect 36596 8032 36602 8084
rect 21726 7964 21732 8016
rect 21784 7964 21790 8016
rect 22094 7964 22100 8016
rect 22152 8004 22158 8016
rect 25041 8007 25099 8013
rect 25041 8004 25053 8007
rect 22152 7976 25053 8004
rect 22152 7964 22158 7976
rect 25041 7973 25053 7976
rect 25087 8004 25099 8007
rect 25498 8004 25504 8016
rect 25087 7976 25504 8004
rect 25087 7973 25099 7976
rect 25041 7967 25099 7973
rect 25498 7964 25504 7976
rect 25556 7964 25562 8016
rect 26234 7964 26240 8016
rect 26292 8004 26298 8016
rect 26329 8007 26387 8013
rect 26329 8004 26341 8007
rect 26292 7976 26341 8004
rect 26292 7964 26298 7976
rect 26329 7973 26341 7976
rect 26375 7973 26387 8007
rect 26329 7967 26387 7973
rect 26510 7964 26516 8016
rect 26568 8004 26574 8016
rect 26697 8007 26755 8013
rect 26697 8004 26709 8007
rect 26568 7976 26709 8004
rect 26568 7964 26574 7976
rect 26697 7973 26709 7976
rect 26743 7973 26755 8007
rect 27798 8004 27804 8016
rect 26697 7967 26755 7973
rect 26804 7976 27804 8004
rect 20824 7908 21680 7936
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7868 19947 7871
rect 19978 7868 19984 7880
rect 19935 7840 19984 7868
rect 19935 7837 19947 7840
rect 19889 7831 19947 7837
rect 19978 7828 19984 7840
rect 20036 7868 20042 7880
rect 20824 7868 20852 7908
rect 20036 7840 20852 7868
rect 20901 7871 20959 7877
rect 20036 7828 20042 7840
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 21082 7868 21088 7880
rect 20947 7840 21088 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 21082 7828 21088 7840
rect 21140 7828 21146 7880
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 21450 7868 21456 7880
rect 21223 7840 21456 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 21737 7877 21765 7964
rect 24118 7896 24124 7948
rect 24176 7936 24182 7948
rect 26804 7936 26832 7976
rect 27798 7964 27804 7976
rect 27856 7964 27862 8016
rect 29089 8007 29147 8013
rect 29089 7973 29101 8007
rect 29135 8004 29147 8007
rect 29362 8004 29368 8016
rect 29135 7976 29368 8004
rect 29135 7973 29147 7976
rect 29089 7967 29147 7973
rect 29362 7964 29368 7976
rect 29420 8004 29426 8016
rect 29730 8004 29736 8016
rect 29420 7976 29736 8004
rect 29420 7964 29426 7976
rect 29730 7964 29736 7976
rect 29788 7964 29794 8016
rect 30374 7964 30380 8016
rect 30432 8004 30438 8016
rect 30926 8004 30932 8016
rect 30432 7976 30932 8004
rect 30432 7964 30438 7976
rect 30926 7964 30932 7976
rect 30984 8004 30990 8016
rect 31938 8004 31944 8016
rect 30984 7976 31944 8004
rect 30984 7964 30990 7976
rect 31938 7964 31944 7976
rect 31996 8004 32002 8016
rect 33042 8004 33048 8016
rect 31996 7976 33048 8004
rect 31996 7964 32002 7976
rect 33042 7964 33048 7976
rect 33100 7964 33106 8016
rect 34238 8004 34244 8016
rect 34072 7976 34244 8004
rect 24176 7908 26832 7936
rect 26881 7939 26939 7945
rect 24176 7896 24182 7908
rect 26881 7905 26893 7939
rect 26927 7905 26939 7939
rect 26881 7899 26939 7905
rect 28261 7939 28319 7945
rect 28261 7905 28273 7939
rect 28307 7936 28319 7939
rect 28626 7936 28632 7948
rect 28307 7908 28632 7936
rect 28307 7905 28319 7908
rect 28261 7899 28319 7905
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 24578 7868 24584 7880
rect 23808 7840 24584 7868
rect 23808 7828 23814 7840
rect 24578 7828 24584 7840
rect 24636 7828 24642 7880
rect 24854 7828 24860 7880
rect 24912 7868 24918 7880
rect 25682 7868 25688 7880
rect 24912 7840 25688 7868
rect 24912 7828 24918 7840
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 26896 7868 26924 7899
rect 28626 7896 28632 7908
rect 28684 7936 28690 7948
rect 29914 7936 29920 7948
rect 28684 7908 29920 7936
rect 28684 7896 28690 7908
rect 27617 7871 27675 7877
rect 27617 7868 27629 7871
rect 26896 7840 27629 7868
rect 27617 7837 27629 7840
rect 27663 7868 27675 7871
rect 27706 7868 27712 7880
rect 27663 7840 27712 7868
rect 27663 7837 27675 7840
rect 27617 7831 27675 7837
rect 27706 7828 27712 7840
rect 27764 7828 27770 7880
rect 27890 7828 27896 7880
rect 27948 7828 27954 7880
rect 27982 7828 27988 7880
rect 28040 7868 28046 7880
rect 28169 7871 28227 7877
rect 28169 7868 28181 7871
rect 28040 7840 28181 7868
rect 28040 7828 28046 7840
rect 28169 7837 28181 7840
rect 28215 7868 28227 7871
rect 28902 7868 28908 7880
rect 28215 7840 28908 7868
rect 28215 7837 28227 7840
rect 28169 7831 28227 7837
rect 28902 7828 28908 7840
rect 28960 7868 28966 7880
rect 29748 7877 29776 7908
rect 29914 7896 29920 7908
rect 29972 7896 29978 7948
rect 30466 7936 30472 7948
rect 30392 7908 30472 7936
rect 30392 7877 30420 7908
rect 30466 7896 30472 7908
rect 30524 7936 30530 7948
rect 31386 7936 31392 7948
rect 30524 7908 31392 7936
rect 30524 7896 30530 7908
rect 31386 7896 31392 7908
rect 31444 7896 31450 7948
rect 32674 7896 32680 7948
rect 32732 7936 32738 7948
rect 33870 7936 33876 7948
rect 32732 7908 33088 7936
rect 32732 7896 32738 7908
rect 29733 7871 29791 7877
rect 28960 7840 29684 7868
rect 28960 7828 28966 7840
rect 17497 7803 17555 7809
rect 17497 7800 17509 7803
rect 17000 7772 17509 7800
rect 17000 7760 17006 7772
rect 17497 7769 17509 7772
rect 17543 7800 17555 7803
rect 19061 7803 19119 7809
rect 17543 7772 18736 7800
rect 17543 7769 17555 7772
rect 17497 7763 17555 7769
rect 18708 7741 18736 7772
rect 19061 7769 19073 7803
rect 19107 7769 19119 7803
rect 19061 7763 19119 7769
rect 19150 7760 19156 7812
rect 19208 7800 19214 7812
rect 19208 7772 19472 7800
rect 19208 7760 19214 7772
rect 16761 7735 16819 7741
rect 16761 7701 16773 7735
rect 16807 7701 16819 7735
rect 16761 7695 16819 7701
rect 18693 7735 18751 7741
rect 18693 7701 18705 7735
rect 18739 7701 18751 7735
rect 18693 7695 18751 7701
rect 18861 7735 18919 7741
rect 18861 7701 18873 7735
rect 18907 7732 18919 7735
rect 19334 7732 19340 7744
rect 18907 7704 19340 7732
rect 18907 7701 18919 7704
rect 18861 7695 18919 7701
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 19444 7732 19472 7772
rect 24670 7760 24676 7812
rect 24728 7800 24734 7812
rect 25590 7800 25596 7812
rect 24728 7772 25596 7800
rect 24728 7760 24734 7772
rect 25590 7760 25596 7772
rect 25648 7800 25654 7812
rect 28378 7803 28436 7809
rect 25648 7772 27568 7800
rect 25648 7760 25654 7772
rect 19610 7732 19616 7744
rect 19444 7704 19616 7732
rect 19610 7692 19616 7704
rect 19668 7692 19674 7744
rect 21545 7735 21603 7741
rect 21545 7701 21557 7735
rect 21591 7732 21603 7735
rect 21910 7732 21916 7744
rect 21591 7704 21916 7732
rect 21591 7701 21603 7704
rect 21545 7695 21603 7701
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 26050 7732 26056 7744
rect 22980 7704 26056 7732
rect 22980 7692 22986 7704
rect 26050 7692 26056 7704
rect 26108 7692 26114 7744
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 27430 7732 27436 7744
rect 26752 7704 27436 7732
rect 26752 7692 26758 7704
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 27540 7732 27568 7772
rect 28378 7769 28390 7803
rect 28424 7800 28436 7803
rect 28810 7800 28816 7812
rect 28424 7772 28816 7800
rect 28424 7769 28436 7772
rect 28378 7763 28436 7769
rect 28810 7760 28816 7772
rect 28868 7760 28874 7812
rect 29178 7760 29184 7812
rect 29236 7800 29242 7812
rect 29365 7803 29423 7809
rect 29365 7800 29377 7803
rect 29236 7772 29377 7800
rect 29236 7760 29242 7772
rect 29365 7769 29377 7772
rect 29411 7769 29423 7803
rect 29365 7763 29423 7769
rect 29454 7760 29460 7812
rect 29512 7800 29518 7812
rect 29549 7803 29607 7809
rect 29549 7800 29561 7803
rect 29512 7772 29561 7800
rect 29512 7760 29518 7772
rect 29549 7769 29561 7772
rect 29595 7769 29607 7803
rect 29656 7800 29684 7840
rect 29733 7837 29745 7871
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 29825 7871 29883 7877
rect 29825 7837 29837 7871
rect 29871 7837 29883 7871
rect 29825 7831 29883 7837
rect 30101 7871 30159 7877
rect 30101 7837 30113 7871
rect 30147 7837 30159 7871
rect 30101 7831 30159 7837
rect 30377 7871 30435 7877
rect 30377 7837 30389 7871
rect 30423 7837 30435 7871
rect 30561 7871 30619 7877
rect 30561 7868 30573 7871
rect 30377 7831 30435 7837
rect 30484 7840 30573 7868
rect 29840 7800 29868 7831
rect 29656 7772 29868 7800
rect 29549 7763 29607 7769
rect 30116 7744 30144 7831
rect 30190 7760 30196 7812
rect 30248 7800 30254 7812
rect 30484 7800 30512 7840
rect 30561 7837 30573 7840
rect 30607 7837 30619 7871
rect 30561 7831 30619 7837
rect 31018 7828 31024 7880
rect 31076 7828 31082 7880
rect 31849 7871 31907 7877
rect 31849 7837 31861 7871
rect 31895 7868 31907 7871
rect 31938 7868 31944 7880
rect 31895 7840 31944 7868
rect 31895 7837 31907 7840
rect 31849 7831 31907 7837
rect 31938 7828 31944 7840
rect 31996 7828 32002 7880
rect 32033 7871 32091 7877
rect 32033 7837 32045 7871
rect 32079 7837 32091 7871
rect 32033 7831 32091 7837
rect 32585 7871 32643 7877
rect 32585 7837 32597 7871
rect 32631 7868 32643 7871
rect 32858 7868 32864 7880
rect 32631 7840 32864 7868
rect 32631 7837 32643 7840
rect 32585 7831 32643 7837
rect 30834 7800 30840 7812
rect 30248 7772 30512 7800
rect 30576 7772 30840 7800
rect 30248 7760 30254 7772
rect 29270 7732 29276 7744
rect 27540 7704 29276 7732
rect 29270 7692 29276 7704
rect 29328 7692 29334 7744
rect 30098 7692 30104 7744
rect 30156 7732 30162 7744
rect 30576 7732 30604 7772
rect 30834 7760 30840 7772
rect 30892 7800 30898 7812
rect 32048 7800 32076 7831
rect 32858 7828 32864 7840
rect 32916 7828 32922 7880
rect 33060 7877 33088 7908
rect 33428 7908 33876 7936
rect 33045 7871 33103 7877
rect 33045 7837 33057 7871
rect 33091 7837 33103 7871
rect 33045 7831 33103 7837
rect 33428 7800 33456 7908
rect 33502 7828 33508 7880
rect 33560 7828 33566 7880
rect 33612 7877 33640 7908
rect 33870 7896 33876 7908
rect 33928 7896 33934 7948
rect 34072 7945 34100 7976
rect 34238 7964 34244 7976
rect 34296 7964 34302 8016
rect 34057 7939 34115 7945
rect 34057 7905 34069 7939
rect 34103 7905 34115 7939
rect 34057 7899 34115 7905
rect 33597 7871 33655 7877
rect 33597 7837 33609 7871
rect 33643 7837 33655 7871
rect 34241 7871 34299 7877
rect 34241 7868 34253 7871
rect 33597 7831 33655 7837
rect 33704 7840 34253 7868
rect 30892 7772 33456 7800
rect 33520 7800 33548 7828
rect 33704 7800 33732 7840
rect 34241 7837 34253 7840
rect 34287 7837 34299 7871
rect 34241 7831 34299 7837
rect 34330 7828 34336 7880
rect 34388 7868 34394 7880
rect 34793 7871 34851 7877
rect 34793 7868 34805 7871
rect 34388 7840 34805 7868
rect 34388 7828 34394 7840
rect 34793 7837 34805 7840
rect 34839 7837 34851 7871
rect 34793 7831 34851 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7868 35035 7871
rect 36078 7868 36084 7880
rect 35023 7840 36084 7868
rect 35023 7837 35035 7840
rect 34977 7831 35035 7837
rect 36078 7828 36084 7840
rect 36136 7828 36142 7880
rect 33520 7772 33732 7800
rect 33965 7803 34023 7809
rect 30892 7760 30898 7772
rect 33965 7769 33977 7803
rect 34011 7800 34023 7803
rect 34054 7800 34060 7812
rect 34011 7772 34060 7800
rect 34011 7769 34023 7772
rect 33965 7763 34023 7769
rect 34054 7760 34060 7772
rect 34112 7760 34118 7812
rect 34422 7760 34428 7812
rect 34480 7760 34486 7812
rect 30156 7704 30604 7732
rect 30156 7692 30162 7704
rect 30650 7692 30656 7744
rect 30708 7692 30714 7744
rect 31481 7735 31539 7741
rect 31481 7701 31493 7735
rect 31527 7732 31539 7735
rect 31662 7732 31668 7744
rect 31527 7704 31668 7732
rect 31527 7701 31539 7704
rect 31481 7695 31539 7701
rect 31662 7692 31668 7704
rect 31720 7692 31726 7744
rect 1104 7642 36524 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 36524 7642
rect 1104 7568 36524 7590
rect 11606 7488 11612 7540
rect 11664 7488 11670 7540
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 12066 7488 12072 7540
rect 12124 7488 12130 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 11514 7420 11520 7472
rect 11572 7420 11578 7472
rect 11882 7420 11888 7472
rect 11940 7420 11946 7472
rect 12084 7460 12112 7488
rect 13280 7460 13308 7491
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14918 7528 14924 7540
rect 14056 7500 14924 7528
rect 14056 7488 14062 7500
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 15013 7531 15071 7537
rect 15013 7497 15025 7531
rect 15059 7528 15071 7531
rect 15746 7528 15752 7540
rect 15059 7500 15752 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 21910 7528 21916 7540
rect 16868 7500 21916 7528
rect 12084 7432 12296 7460
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12268 7401 12296 7432
rect 12452 7432 13308 7460
rect 13449 7463 13507 7469
rect 12452 7401 12480 7432
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 13495 7432 14136 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 12161 7395 12219 7401
rect 12161 7392 12173 7395
rect 12124 7364 12173 7392
rect 12124 7352 12130 7364
rect 12161 7361 12173 7364
rect 12207 7361 12219 7395
rect 12161 7355 12219 7361
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 12422 7395 12480 7401
rect 12422 7361 12434 7395
rect 12468 7361 12480 7395
rect 12422 7355 12480 7361
rect 12268 7324 12296 7355
rect 12526 7352 12532 7404
rect 12584 7352 12590 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12805 7395 12863 7401
rect 12805 7392 12817 7395
rect 12768 7364 12817 7392
rect 12768 7352 12774 7364
rect 12805 7361 12817 7364
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7392 13231 7395
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13219 7364 13829 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13817 7361 13829 7364
rect 13863 7392 13875 7395
rect 13906 7392 13912 7404
rect 13863 7364 13912 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14108 7401 14136 7432
rect 15102 7420 15108 7472
rect 15160 7420 15166 7472
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 14139 7364 14381 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14369 7361 14381 7364
rect 14415 7392 14427 7395
rect 15120 7392 15148 7420
rect 16868 7401 16896 7500
rect 21910 7488 21916 7500
rect 21968 7488 21974 7540
rect 22186 7488 22192 7540
rect 22244 7488 22250 7540
rect 23658 7488 23664 7540
rect 23716 7528 23722 7540
rect 23716 7500 24440 7528
rect 23716 7488 23722 7500
rect 18782 7420 18788 7472
rect 18840 7460 18846 7472
rect 18969 7463 19027 7469
rect 18969 7460 18981 7463
rect 18840 7432 18981 7460
rect 18840 7420 18846 7432
rect 18969 7429 18981 7432
rect 19015 7429 19027 7463
rect 19518 7460 19524 7472
rect 18969 7423 19027 7429
rect 19168 7432 19524 7460
rect 16853 7395 16911 7401
rect 14415 7364 15056 7392
rect 15120 7364 15240 7392
rect 14415 7361 14427 7364
rect 14369 7355 14427 7361
rect 12268 7296 12756 7324
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 11747 7228 12204 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 11790 7148 11796 7200
rect 11848 7148 11854 7200
rect 12176 7188 12204 7228
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 12176 7160 12633 7188
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 12728 7188 12756 7296
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 13320 7296 13952 7324
rect 13320 7284 13326 7296
rect 13924 7256 13952 7296
rect 14182 7284 14188 7336
rect 14240 7284 14246 7336
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7324 14611 7327
rect 14599 7296 14872 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 14645 7259 14703 7265
rect 14645 7256 14657 7259
rect 13924 7228 14657 7256
rect 14645 7225 14657 7228
rect 14691 7225 14703 7259
rect 14844 7256 14872 7296
rect 15028 7256 15056 7364
rect 15102 7284 15108 7336
rect 15160 7284 15166 7336
rect 15212 7333 15240 7364
rect 16853 7361 16865 7395
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 17000 7364 17141 7392
rect 17000 7352 17006 7364
rect 17129 7361 17141 7364
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17310 7352 17316 7404
rect 17368 7352 17374 7404
rect 17770 7352 17776 7404
rect 17828 7392 17834 7404
rect 19168 7392 19196 7432
rect 19518 7420 19524 7432
rect 19576 7460 19582 7472
rect 20717 7463 20775 7469
rect 19576 7432 20024 7460
rect 19576 7420 19582 7432
rect 17828 7364 19196 7392
rect 17828 7352 17834 7364
rect 19242 7352 19248 7404
rect 19300 7352 19306 7404
rect 19334 7352 19340 7404
rect 19392 7352 19398 7404
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19794 7392 19800 7404
rect 19659 7364 19800 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 19996 7401 20024 7432
rect 20487 7429 20545 7435
rect 19981 7395 20039 7401
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 20487 7395 20499 7429
rect 20533 7426 20545 7429
rect 20717 7429 20729 7463
rect 20763 7460 20775 7463
rect 20898 7460 20904 7472
rect 20763 7432 20904 7460
rect 20763 7429 20775 7432
rect 20533 7395 20560 7426
rect 20717 7423 20775 7429
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 21453 7463 21511 7469
rect 21453 7429 21465 7463
rect 21499 7460 21511 7463
rect 21634 7460 21640 7472
rect 21499 7432 21640 7460
rect 21499 7429 21511 7432
rect 21453 7423 21511 7429
rect 21634 7420 21640 7432
rect 21692 7460 21698 7472
rect 21821 7463 21879 7469
rect 21821 7460 21833 7463
rect 21692 7432 21833 7460
rect 21692 7420 21698 7432
rect 21821 7429 21833 7432
rect 21867 7429 21879 7463
rect 21821 7423 21879 7429
rect 22002 7420 22008 7472
rect 22060 7420 22066 7472
rect 22094 7420 22100 7472
rect 22152 7460 22158 7472
rect 22646 7460 22652 7472
rect 22152 7432 22652 7460
rect 22152 7420 22158 7432
rect 22646 7420 22652 7432
rect 22704 7460 22710 7472
rect 23201 7463 23259 7469
rect 23201 7460 23213 7463
rect 22704 7432 23213 7460
rect 22704 7420 22710 7432
rect 23201 7429 23213 7432
rect 23247 7460 23259 7463
rect 23382 7460 23388 7472
rect 23247 7432 23388 7460
rect 23247 7429 23259 7432
rect 23201 7423 23259 7429
rect 23382 7420 23388 7432
rect 23440 7420 23446 7472
rect 23934 7420 23940 7472
rect 23992 7460 23998 7472
rect 23992 7432 24348 7460
rect 23992 7420 23998 7432
rect 20487 7392 20560 7395
rect 21266 7392 21272 7404
rect 20487 7389 21272 7392
rect 20532 7364 21272 7389
rect 19981 7355 20039 7361
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21542 7392 21548 7404
rect 21407 7364 21548 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21542 7352 21548 7364
rect 21600 7392 21606 7404
rect 22922 7392 22928 7404
rect 21600 7364 22928 7392
rect 21600 7352 21606 7364
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7392 23075 7395
rect 24118 7392 24124 7404
rect 23063 7364 24124 7392
rect 23063 7361 23075 7364
rect 23017 7355 23075 7361
rect 15197 7327 15255 7333
rect 15197 7293 15209 7327
rect 15243 7293 15255 7327
rect 15197 7287 15255 7293
rect 15746 7284 15752 7336
rect 15804 7324 15810 7336
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 15804 7296 19717 7324
rect 15804 7284 15810 7296
rect 19705 7293 19717 7296
rect 19751 7293 19763 7327
rect 19705 7287 19763 7293
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7293 19947 7327
rect 19889 7287 19947 7293
rect 16850 7256 16856 7268
rect 14844 7228 14964 7256
rect 15028 7228 16856 7256
rect 14645 7219 14703 7225
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12728 7160 12817 7188
rect 12621 7151 12679 7157
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 13446 7148 13452 7200
rect 13504 7148 13510 7200
rect 14936 7188 14964 7228
rect 16850 7216 16856 7228
rect 16908 7216 16914 7268
rect 16945 7259 17003 7265
rect 16945 7225 16957 7259
rect 16991 7225 17003 7259
rect 16945 7219 17003 7225
rect 15102 7188 15108 7200
rect 14936 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 16666 7148 16672 7200
rect 16724 7148 16730 7200
rect 16960 7188 16988 7219
rect 17034 7216 17040 7268
rect 17092 7216 17098 7268
rect 19610 7216 19616 7268
rect 19668 7256 19674 7268
rect 19904 7256 19932 7287
rect 20070 7284 20076 7336
rect 20128 7284 20134 7336
rect 20162 7284 20168 7336
rect 20220 7284 20226 7336
rect 20346 7256 20352 7268
rect 19668 7228 20352 7256
rect 19668 7216 19674 7228
rect 20346 7216 20352 7228
rect 20404 7216 20410 7268
rect 20898 7216 20904 7268
rect 20956 7256 20962 7268
rect 21818 7256 21824 7268
rect 20956 7228 21824 7256
rect 20956 7216 20962 7228
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 23032 7256 23060 7355
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 24320 7401 24348 7432
rect 24412 7404 24440 7500
rect 24486 7488 24492 7540
rect 24544 7528 24550 7540
rect 24544 7500 25360 7528
rect 24544 7488 24550 7500
rect 24765 7463 24823 7469
rect 24765 7429 24777 7463
rect 24811 7460 24823 7463
rect 25332 7460 25360 7500
rect 25406 7488 25412 7540
rect 25464 7488 25470 7540
rect 25590 7488 25596 7540
rect 25648 7488 25654 7540
rect 25869 7531 25927 7537
rect 25869 7497 25881 7531
rect 25915 7528 25927 7531
rect 26418 7528 26424 7540
rect 25915 7500 26424 7528
rect 25915 7497 25927 7500
rect 25869 7491 25927 7497
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 27065 7531 27123 7537
rect 27065 7497 27077 7531
rect 27111 7497 27123 7531
rect 28077 7531 28135 7537
rect 28077 7528 28089 7531
rect 27065 7491 27123 7497
rect 27264 7500 28089 7528
rect 27080 7460 27108 7491
rect 24811 7432 24900 7460
rect 25332 7432 27108 7460
rect 24811 7429 24823 7432
rect 24765 7423 24823 7429
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24394 7352 24400 7404
rect 24452 7352 24458 7404
rect 24872 7401 24900 7432
rect 24489 7395 24547 7401
rect 24489 7361 24501 7395
rect 24535 7361 24547 7395
rect 24489 7355 24547 7361
rect 24857 7395 24915 7401
rect 24857 7361 24869 7395
rect 24903 7361 24915 7395
rect 24857 7355 24915 7361
rect 24949 7395 25007 7401
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 25225 7395 25283 7401
rect 25225 7361 25237 7395
rect 25271 7392 25283 7395
rect 25314 7392 25320 7404
rect 25271 7364 25320 7392
rect 25271 7361 25283 7364
rect 25225 7355 25283 7361
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 24504 7324 24532 7355
rect 23900 7296 24532 7324
rect 23900 7284 23906 7296
rect 24762 7284 24768 7336
rect 24820 7324 24826 7336
rect 24964 7324 24992 7355
rect 24820 7296 24992 7324
rect 25148 7324 25176 7355
rect 25314 7352 25320 7364
rect 25372 7352 25378 7404
rect 25498 7352 25504 7404
rect 25556 7352 25562 7404
rect 26510 7352 26516 7404
rect 26568 7392 26574 7404
rect 26605 7395 26663 7401
rect 26605 7392 26617 7395
rect 26568 7364 26617 7392
rect 26568 7352 26574 7364
rect 26605 7361 26617 7364
rect 26651 7392 26663 7395
rect 26786 7392 26792 7404
rect 26651 7364 26792 7392
rect 26651 7361 26663 7364
rect 26605 7355 26663 7361
rect 26786 7352 26792 7364
rect 26844 7392 26850 7404
rect 27264 7401 27292 7500
rect 28077 7497 28089 7500
rect 28123 7497 28135 7531
rect 28077 7491 28135 7497
rect 28994 7488 29000 7540
rect 29052 7488 29058 7540
rect 30101 7531 30159 7537
rect 30101 7497 30113 7531
rect 30147 7528 30159 7531
rect 30374 7528 30380 7540
rect 30147 7500 30380 7528
rect 30147 7497 30159 7500
rect 30101 7491 30159 7497
rect 30374 7488 30380 7500
rect 30432 7488 30438 7540
rect 30561 7531 30619 7537
rect 30561 7497 30573 7531
rect 30607 7528 30619 7531
rect 30742 7528 30748 7540
rect 30607 7500 30748 7528
rect 30607 7497 30619 7500
rect 30561 7491 30619 7497
rect 30742 7488 30748 7500
rect 30800 7488 30806 7540
rect 34146 7528 34152 7540
rect 32968 7500 34152 7528
rect 27890 7420 27896 7472
rect 27948 7460 27954 7472
rect 27985 7463 28043 7469
rect 27985 7460 27997 7463
rect 27948 7432 27997 7460
rect 27948 7420 27954 7432
rect 27985 7429 27997 7432
rect 28031 7460 28043 7463
rect 28031 7432 28764 7460
rect 28031 7429 28043 7432
rect 27985 7423 28043 7429
rect 28736 7404 28764 7432
rect 28810 7420 28816 7472
rect 28868 7460 28874 7472
rect 29181 7463 29239 7469
rect 29181 7460 29193 7463
rect 28868 7432 29193 7460
rect 28868 7420 28874 7432
rect 29181 7429 29193 7432
rect 29227 7460 29239 7463
rect 29227 7432 30788 7460
rect 29227 7429 29239 7432
rect 29181 7423 29239 7429
rect 27249 7395 27307 7401
rect 27249 7392 27261 7395
rect 26844 7364 27261 7392
rect 26844 7352 26850 7364
rect 27249 7361 27261 7364
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 27430 7352 27436 7404
rect 27488 7392 27494 7404
rect 27617 7395 27675 7401
rect 27617 7392 27629 7395
rect 27488 7364 27629 7392
rect 27488 7352 27494 7364
rect 27617 7361 27629 7364
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 28074 7352 28080 7404
rect 28132 7392 28138 7404
rect 28629 7395 28687 7401
rect 28629 7392 28641 7395
rect 28132 7364 28641 7392
rect 28132 7352 28138 7364
rect 28629 7361 28641 7364
rect 28675 7361 28687 7395
rect 28629 7355 28687 7361
rect 28718 7352 28724 7404
rect 28776 7392 28782 7404
rect 29273 7395 29331 7401
rect 29273 7392 29285 7395
rect 28776 7364 29285 7392
rect 28776 7352 28782 7364
rect 29273 7361 29285 7364
rect 29319 7392 29331 7395
rect 29641 7395 29699 7401
rect 29319 7364 29592 7392
rect 29319 7361 29331 7364
rect 29273 7355 29331 7361
rect 25774 7324 25780 7336
rect 25148 7296 25780 7324
rect 24820 7284 24826 7296
rect 25148 7256 25176 7296
rect 25774 7284 25780 7296
rect 25832 7284 25838 7336
rect 26050 7284 26056 7336
rect 26108 7324 26114 7336
rect 26145 7327 26203 7333
rect 26145 7324 26157 7327
rect 26108 7296 26157 7324
rect 26108 7284 26114 7296
rect 26145 7293 26157 7296
rect 26191 7293 26203 7327
rect 26145 7287 26203 7293
rect 22296 7228 23060 7256
rect 23860 7228 25176 7256
rect 26160 7256 26188 7287
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 26697 7327 26755 7333
rect 26697 7324 26709 7327
rect 26292 7296 26709 7324
rect 26292 7284 26298 7296
rect 26697 7293 26709 7296
rect 26743 7324 26755 7327
rect 27709 7327 27767 7333
rect 27709 7324 27721 7327
rect 26743 7296 27721 7324
rect 26743 7293 26755 7296
rect 26697 7287 26755 7293
rect 27709 7293 27721 7296
rect 27755 7293 27767 7327
rect 27709 7287 27767 7293
rect 28166 7284 28172 7336
rect 28224 7324 28230 7336
rect 28813 7327 28871 7333
rect 28813 7324 28825 7327
rect 28224 7296 28825 7324
rect 28224 7284 28230 7296
rect 28813 7293 28825 7296
rect 28859 7293 28871 7327
rect 28813 7287 28871 7293
rect 28902 7284 28908 7336
rect 28960 7324 28966 7336
rect 29365 7327 29423 7333
rect 29365 7324 29377 7327
rect 28960 7296 29377 7324
rect 28960 7284 28966 7296
rect 29365 7293 29377 7296
rect 29411 7293 29423 7327
rect 29564 7324 29592 7364
rect 29641 7361 29653 7395
rect 29687 7392 29699 7395
rect 29914 7392 29920 7404
rect 29687 7364 29920 7392
rect 29687 7361 29699 7364
rect 29641 7355 29699 7361
rect 29914 7352 29920 7364
rect 29972 7352 29978 7404
rect 30009 7395 30067 7401
rect 30009 7361 30021 7395
rect 30055 7392 30067 7395
rect 30098 7392 30104 7404
rect 30055 7364 30104 7392
rect 30055 7361 30067 7364
rect 30009 7355 30067 7361
rect 30024 7324 30052 7355
rect 30098 7352 30104 7364
rect 30156 7352 30162 7404
rect 30193 7395 30251 7401
rect 30193 7361 30205 7395
rect 30239 7392 30251 7395
rect 30282 7392 30288 7404
rect 30239 7364 30288 7392
rect 30239 7361 30251 7364
rect 30193 7355 30251 7361
rect 30282 7352 30288 7364
rect 30340 7352 30346 7404
rect 30760 7401 30788 7432
rect 30926 7420 30932 7472
rect 30984 7420 30990 7472
rect 31021 7463 31079 7469
rect 31021 7429 31033 7463
rect 31067 7460 31079 7463
rect 31294 7460 31300 7472
rect 31067 7432 31300 7460
rect 31067 7429 31079 7432
rect 31021 7423 31079 7429
rect 31294 7420 31300 7432
rect 31352 7420 31358 7472
rect 30745 7395 30803 7401
rect 30745 7361 30757 7395
rect 30791 7392 30803 7395
rect 31386 7392 31392 7404
rect 30791 7364 31392 7392
rect 30791 7361 30803 7364
rect 30745 7355 30803 7361
rect 31386 7352 31392 7364
rect 31444 7352 31450 7404
rect 31481 7395 31539 7401
rect 31481 7361 31493 7395
rect 31527 7361 31539 7395
rect 31481 7355 31539 7361
rect 29564 7296 30052 7324
rect 30300 7324 30328 7352
rect 31018 7324 31024 7336
rect 30300 7296 31024 7324
rect 29365 7287 29423 7293
rect 31018 7284 31024 7296
rect 31076 7324 31082 7336
rect 31294 7324 31300 7336
rect 31076 7296 31300 7324
rect 31076 7284 31082 7296
rect 31294 7284 31300 7296
rect 31352 7324 31358 7336
rect 31496 7324 31524 7355
rect 31570 7352 31576 7404
rect 31628 7392 31634 7404
rect 31941 7395 31999 7401
rect 31941 7392 31953 7395
rect 31628 7364 31953 7392
rect 31628 7352 31634 7364
rect 31941 7361 31953 7364
rect 31987 7392 31999 7395
rect 32968 7392 32996 7500
rect 34146 7488 34152 7500
rect 34204 7488 34210 7540
rect 34790 7488 34796 7540
rect 34848 7528 34854 7540
rect 35345 7531 35403 7537
rect 35345 7528 35357 7531
rect 34848 7500 35357 7528
rect 34848 7488 34854 7500
rect 35345 7497 35357 7500
rect 35391 7497 35403 7531
rect 35345 7491 35403 7497
rect 33873 7463 33931 7469
rect 33873 7429 33885 7463
rect 33919 7460 33931 7463
rect 33962 7460 33968 7472
rect 33919 7432 33968 7460
rect 33919 7429 33931 7432
rect 33873 7423 33931 7429
rect 33962 7420 33968 7432
rect 34020 7420 34026 7472
rect 34330 7420 34336 7472
rect 34388 7420 34394 7472
rect 31987 7364 32996 7392
rect 31987 7361 31999 7364
rect 31941 7355 31999 7361
rect 31352 7296 31524 7324
rect 31352 7284 31358 7296
rect 33134 7284 33140 7336
rect 33192 7324 33198 7336
rect 33597 7327 33655 7333
rect 33597 7324 33609 7327
rect 33192 7296 33609 7324
rect 33192 7284 33198 7296
rect 33597 7293 33609 7296
rect 33643 7293 33655 7327
rect 33597 7287 33655 7293
rect 26786 7256 26792 7268
rect 26160 7228 26792 7256
rect 19150 7188 19156 7200
rect 16960 7160 19156 7188
rect 19150 7148 19156 7160
rect 19208 7148 19214 7200
rect 20438 7148 20444 7200
rect 20496 7188 20502 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 20496 7160 20545 7188
rect 20496 7148 20502 7160
rect 20533 7157 20545 7160
rect 20579 7157 20591 7191
rect 20533 7151 20591 7157
rect 20806 7148 20812 7200
rect 20864 7188 20870 7200
rect 22296 7188 22324 7228
rect 23860 7200 23888 7228
rect 26786 7216 26792 7228
rect 26844 7216 26850 7268
rect 27614 7216 27620 7268
rect 27672 7256 27678 7268
rect 28445 7259 28503 7265
rect 28445 7256 28457 7259
rect 27672 7228 28457 7256
rect 27672 7216 27678 7228
rect 28445 7225 28457 7228
rect 28491 7225 28503 7259
rect 28445 7219 28503 7225
rect 28534 7216 28540 7268
rect 28592 7256 28598 7268
rect 28920 7256 28948 7284
rect 28592 7228 28948 7256
rect 28592 7216 28598 7228
rect 20864 7160 22324 7188
rect 22373 7191 22431 7197
rect 20864 7148 20870 7160
rect 22373 7157 22385 7191
rect 22419 7188 22431 7191
rect 22646 7188 22652 7200
rect 22419 7160 22652 7188
rect 22419 7157 22431 7160
rect 22373 7151 22431 7157
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 23842 7148 23848 7200
rect 23900 7148 23906 7200
rect 26237 7191 26295 7197
rect 26237 7157 26249 7191
rect 26283 7188 26295 7191
rect 26418 7188 26424 7200
rect 26283 7160 26424 7188
rect 26283 7157 26295 7160
rect 26237 7151 26295 7157
rect 26418 7148 26424 7160
rect 26476 7188 26482 7200
rect 26602 7188 26608 7200
rect 26476 7160 26608 7188
rect 26476 7148 26482 7160
rect 26602 7148 26608 7160
rect 26660 7188 26666 7200
rect 27249 7191 27307 7197
rect 27249 7188 27261 7191
rect 26660 7160 27261 7188
rect 26660 7148 26666 7160
rect 27249 7157 27261 7160
rect 27295 7188 27307 7191
rect 27430 7188 27436 7200
rect 27295 7160 27436 7188
rect 27295 7157 27307 7160
rect 27249 7151 27307 7157
rect 27430 7148 27436 7160
rect 27488 7148 27494 7200
rect 1104 7098 36524 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 36524 7098
rect 1104 7024 36524 7046
rect 15286 6944 15292 6996
rect 15344 6984 15350 6996
rect 15454 6987 15512 6993
rect 15454 6984 15466 6987
rect 15344 6956 15466 6984
rect 15344 6944 15350 6956
rect 15454 6953 15466 6956
rect 15500 6953 15512 6987
rect 15454 6947 15512 6953
rect 21174 6944 21180 6996
rect 21232 6944 21238 6996
rect 21361 6987 21419 6993
rect 21361 6953 21373 6987
rect 21407 6984 21419 6987
rect 22002 6984 22008 6996
rect 21407 6956 22008 6984
rect 21407 6953 21419 6956
rect 21361 6947 21419 6953
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22373 6987 22431 6993
rect 22373 6984 22385 6987
rect 22336 6956 22385 6984
rect 22336 6944 22342 6956
rect 22373 6953 22385 6956
rect 22419 6953 22431 6987
rect 22373 6947 22431 6953
rect 22646 6944 22652 6996
rect 22704 6944 22710 6996
rect 23382 6944 23388 6996
rect 23440 6944 23446 6996
rect 25866 6984 25872 6996
rect 24596 6956 25872 6984
rect 14182 6916 14188 6928
rect 13188 6888 14188 6916
rect 12986 6808 12992 6860
rect 13044 6848 13050 6860
rect 13188 6857 13216 6888
rect 14182 6876 14188 6888
rect 14240 6876 14246 6928
rect 15120 6888 15332 6916
rect 13173 6851 13231 6857
rect 13173 6848 13185 6851
rect 13044 6820 13185 6848
rect 13044 6808 13050 6820
rect 13173 6817 13185 6820
rect 13219 6817 13231 6851
rect 13173 6811 13231 6817
rect 13814 6808 13820 6860
rect 13872 6808 13878 6860
rect 11422 6740 11428 6792
rect 11480 6740 11486 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 11698 6672 11704 6724
rect 11756 6672 11762 6724
rect 13556 6712 13584 6743
rect 13630 6740 13636 6792
rect 13688 6740 13694 6792
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 15120 6712 15148 6888
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15304 6848 15332 6888
rect 20162 6876 20168 6928
rect 20220 6916 20226 6928
rect 24596 6916 24624 6956
rect 25866 6944 25872 6956
rect 25924 6944 25930 6996
rect 26145 6987 26203 6993
rect 26145 6984 26157 6987
rect 25976 6956 26157 6984
rect 24762 6916 24768 6928
rect 20220 6888 24624 6916
rect 24688 6888 24768 6916
rect 20220 6876 20226 6888
rect 15304 6820 16712 6848
rect 16684 6780 16712 6820
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 17184 6820 17233 6848
rect 17184 6808 17190 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 22741 6851 22799 6857
rect 22741 6817 22753 6851
rect 22787 6848 22799 6851
rect 24688 6848 24716 6888
rect 24762 6876 24768 6888
rect 24820 6916 24826 6928
rect 24857 6919 24915 6925
rect 24857 6916 24869 6919
rect 24820 6888 24869 6916
rect 24820 6876 24826 6888
rect 24857 6885 24869 6888
rect 24903 6885 24915 6919
rect 24857 6879 24915 6885
rect 25317 6919 25375 6925
rect 25317 6885 25329 6919
rect 25363 6885 25375 6919
rect 25317 6879 25375 6885
rect 22787 6820 24716 6848
rect 22787 6817 22799 6820
rect 22741 6811 22799 6817
rect 16758 6780 16764 6792
rect 16684 6752 16764 6780
rect 16758 6740 16764 6752
rect 16816 6780 16822 6792
rect 17589 6783 17647 6789
rect 16816 6752 17172 6780
rect 16816 6740 16822 6752
rect 17034 6712 17040 6724
rect 12926 6684 13492 6712
rect 13556 6684 15148 6712
rect 16698 6684 17040 6712
rect 13354 6604 13360 6656
rect 13412 6604 13418 6656
rect 13464 6644 13492 6684
rect 13998 6644 14004 6656
rect 13464 6616 14004 6644
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 16776 6644 16804 6684
rect 17034 6672 17040 6684
rect 17092 6672 17098 6724
rect 17144 6712 17172 6752
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17678 6780 17684 6792
rect 17635 6752 17684 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 17770 6740 17776 6792
rect 17828 6740 17834 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19518 6780 19524 6792
rect 19475 6752 19524 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 22094 6780 22100 6792
rect 21376 6752 22100 6780
rect 19245 6715 19303 6721
rect 17144 6684 17816 6712
rect 14516 6616 16804 6644
rect 14516 6604 14522 6616
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17644 6616 17693 6644
rect 17644 6604 17650 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17788 6644 17816 6684
rect 19245 6681 19257 6715
rect 19291 6712 19303 6715
rect 19334 6712 19340 6724
rect 19291 6684 19340 6712
rect 19291 6681 19303 6684
rect 19245 6675 19303 6681
rect 19334 6672 19340 6684
rect 19392 6712 19398 6724
rect 20070 6712 20076 6724
rect 19392 6684 20076 6712
rect 19392 6672 19398 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 21376 6721 21404 6752
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6749 22891 6783
rect 22833 6743 22891 6749
rect 22925 6783 22983 6789
rect 22925 6749 22937 6783
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 21329 6715 21404 6721
rect 21329 6712 21341 6715
rect 20772 6684 21341 6712
rect 20772 6672 20778 6684
rect 21329 6681 21341 6684
rect 21375 6684 21404 6715
rect 21375 6681 21387 6684
rect 21329 6675 21387 6681
rect 21542 6672 21548 6724
rect 21600 6672 21606 6724
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 17788 6616 19533 6644
rect 17681 6607 17739 6613
rect 19521 6613 19533 6616
rect 19567 6613 19579 6647
rect 19521 6607 19579 6613
rect 19702 6604 19708 6656
rect 19760 6644 19766 6656
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 19760 6616 19809 6644
rect 19760 6604 19766 6616
rect 19797 6613 19809 6616
rect 19843 6613 19855 6647
rect 22848 6644 22876 6743
rect 22940 6712 22968 6743
rect 23106 6740 23112 6792
rect 23164 6740 23170 6792
rect 23474 6740 23480 6792
rect 23532 6780 23538 6792
rect 24029 6783 24087 6789
rect 24029 6780 24041 6783
rect 23532 6752 24041 6780
rect 23532 6740 23538 6752
rect 24029 6749 24041 6752
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6780 24639 6783
rect 24670 6780 24676 6792
rect 24627 6752 24676 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 24762 6740 24768 6792
rect 24820 6740 24826 6792
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6749 24915 6783
rect 25332 6780 25360 6879
rect 25593 6851 25651 6857
rect 25593 6817 25605 6851
rect 25639 6848 25651 6851
rect 25976 6848 26004 6956
rect 26145 6953 26157 6956
rect 26191 6984 26203 6987
rect 26326 6984 26332 6996
rect 26191 6956 26332 6984
rect 26191 6953 26203 6956
rect 26145 6947 26203 6953
rect 26326 6944 26332 6956
rect 26384 6944 26390 6996
rect 27157 6987 27215 6993
rect 27157 6953 27169 6987
rect 27203 6984 27215 6987
rect 27522 6984 27528 6996
rect 27203 6956 27528 6984
rect 27203 6953 27215 6956
rect 27157 6947 27215 6953
rect 27522 6944 27528 6956
rect 27580 6944 27586 6996
rect 29178 6984 29184 6996
rect 27632 6956 29184 6984
rect 26237 6919 26295 6925
rect 26237 6885 26249 6919
rect 26283 6885 26295 6919
rect 26237 6879 26295 6885
rect 25639 6820 26004 6848
rect 25639 6817 25651 6820
rect 25593 6811 25651 6817
rect 26050 6808 26056 6860
rect 26108 6808 26114 6860
rect 26252 6780 26280 6879
rect 27246 6876 27252 6928
rect 27304 6916 27310 6928
rect 27632 6916 27660 6956
rect 27304 6888 27660 6916
rect 28721 6919 28779 6925
rect 27304 6876 27310 6888
rect 28721 6885 28733 6919
rect 28767 6916 28779 6919
rect 28810 6916 28816 6928
rect 28767 6888 28816 6916
rect 28767 6885 28779 6888
rect 28721 6879 28779 6885
rect 28810 6876 28816 6888
rect 28868 6876 28874 6928
rect 29012 6925 29040 6956
rect 29178 6944 29184 6956
rect 29236 6984 29242 6996
rect 30650 6984 30656 6996
rect 29236 6956 30656 6984
rect 29236 6944 29242 6956
rect 28997 6919 29055 6925
rect 28997 6885 29009 6919
rect 29043 6885 29055 6919
rect 28997 6879 29055 6885
rect 26326 6808 26332 6860
rect 26384 6848 26390 6860
rect 29273 6851 29331 6857
rect 26384 6820 27384 6848
rect 26384 6808 26390 6820
rect 27356 6792 27384 6820
rect 29273 6817 29285 6851
rect 29319 6848 29331 6851
rect 29362 6848 29368 6860
rect 29319 6820 29368 6848
rect 29319 6817 29331 6820
rect 29273 6811 29331 6817
rect 29362 6808 29368 6820
rect 29420 6808 29426 6860
rect 29641 6851 29699 6857
rect 29641 6817 29653 6851
rect 29687 6848 29699 6851
rect 29914 6848 29920 6860
rect 29687 6820 29920 6848
rect 29687 6817 29699 6820
rect 29641 6811 29699 6817
rect 29914 6808 29920 6820
rect 29972 6808 29978 6860
rect 30024 6857 30052 6956
rect 30009 6851 30067 6857
rect 30009 6817 30021 6851
rect 30055 6817 30067 6851
rect 30009 6811 30067 6817
rect 26418 6780 26424 6792
rect 25332 6752 26424 6780
rect 24857 6743 24915 6749
rect 23492 6712 23520 6740
rect 22940 6684 23520 6712
rect 23569 6715 23627 6721
rect 23569 6681 23581 6715
rect 23615 6681 23627 6715
rect 23569 6675 23627 6681
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 22848 6616 23213 6644
rect 19797 6607 19855 6613
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 23369 6647 23427 6653
rect 23369 6613 23381 6647
rect 23415 6644 23427 6647
rect 23474 6644 23480 6656
rect 23415 6616 23480 6644
rect 23415 6613 23427 6616
rect 23369 6607 23427 6613
rect 23474 6604 23480 6616
rect 23532 6604 23538 6656
rect 23584 6644 23612 6675
rect 23658 6672 23664 6724
rect 23716 6672 23722 6724
rect 23842 6672 23848 6724
rect 23900 6672 23906 6724
rect 24872 6712 24900 6743
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 26510 6740 26516 6792
rect 26568 6780 26574 6792
rect 26605 6783 26663 6789
rect 26605 6780 26617 6783
rect 26568 6752 26617 6780
rect 26568 6740 26574 6752
rect 26605 6749 26617 6752
rect 26651 6749 26663 6783
rect 26605 6743 26663 6749
rect 26697 6783 26755 6789
rect 26697 6749 26709 6783
rect 26743 6780 26755 6783
rect 26786 6780 26792 6792
rect 26743 6752 26792 6780
rect 26743 6749 26755 6752
rect 26697 6743 26755 6749
rect 25222 6712 25228 6724
rect 24872 6684 25228 6712
rect 25222 6672 25228 6684
rect 25280 6712 25286 6724
rect 25685 6715 25743 6721
rect 25685 6712 25697 6715
rect 25280 6684 25697 6712
rect 25280 6672 25286 6684
rect 25685 6681 25697 6684
rect 25731 6681 25743 6715
rect 26620 6712 26648 6743
rect 26786 6740 26792 6752
rect 26844 6740 26850 6792
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6749 27123 6783
rect 27065 6743 27123 6749
rect 27080 6712 27108 6743
rect 27338 6740 27344 6792
rect 27396 6740 27402 6792
rect 27522 6740 27528 6792
rect 27580 6780 27586 6792
rect 27617 6783 27675 6789
rect 27617 6780 27629 6783
rect 27580 6752 27629 6780
rect 27580 6740 27586 6752
rect 27617 6749 27629 6752
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 28353 6783 28411 6789
rect 28353 6749 28365 6783
rect 28399 6780 28411 6783
rect 28626 6780 28632 6792
rect 28399 6752 28632 6780
rect 28399 6749 28411 6752
rect 28353 6743 28411 6749
rect 28626 6740 28632 6752
rect 28684 6740 28690 6792
rect 29380 6780 29408 6808
rect 29825 6783 29883 6789
rect 29825 6780 29837 6783
rect 29380 6752 29837 6780
rect 29825 6749 29837 6752
rect 29871 6780 29883 6783
rect 30193 6783 30251 6789
rect 30193 6780 30205 6783
rect 29871 6752 30205 6780
rect 29871 6749 29883 6752
rect 29825 6743 29883 6749
rect 30193 6749 30205 6752
rect 30239 6749 30251 6783
rect 30300 6780 30328 6956
rect 30650 6944 30656 6956
rect 30708 6944 30714 6996
rect 32480 6987 32538 6993
rect 32480 6953 32492 6987
rect 32526 6984 32538 6987
rect 32582 6984 32588 6996
rect 32526 6956 32588 6984
rect 32526 6953 32538 6956
rect 32480 6947 32538 6953
rect 32582 6944 32588 6956
rect 32640 6944 32646 6996
rect 33965 6987 34023 6993
rect 33965 6953 33977 6987
rect 34011 6984 34023 6987
rect 34422 6984 34428 6996
rect 34011 6956 34428 6984
rect 34011 6953 34023 6956
rect 33965 6947 34023 6953
rect 34422 6944 34428 6956
rect 34480 6944 34486 6996
rect 30834 6857 30840 6860
rect 30812 6851 30840 6857
rect 30812 6817 30824 6851
rect 30812 6811 30840 6817
rect 30834 6808 30840 6811
rect 30892 6808 30898 6860
rect 30926 6808 30932 6860
rect 30984 6848 30990 6860
rect 31021 6851 31079 6857
rect 31021 6848 31033 6851
rect 30984 6820 31033 6848
rect 30984 6808 30990 6820
rect 31021 6817 31033 6820
rect 31067 6817 31079 6851
rect 31021 6811 31079 6817
rect 31294 6808 31300 6860
rect 31352 6808 31358 6860
rect 32217 6851 32275 6857
rect 32217 6817 32229 6851
rect 32263 6848 32275 6851
rect 33134 6848 33140 6860
rect 32263 6820 33140 6848
rect 32263 6817 32275 6820
rect 32217 6811 32275 6817
rect 33134 6808 33140 6820
rect 33192 6808 33198 6860
rect 30377 6783 30435 6789
rect 30377 6780 30389 6783
rect 30300 6752 30389 6780
rect 30193 6743 30251 6749
rect 30377 6749 30389 6752
rect 30423 6749 30435 6783
rect 30377 6743 30435 6749
rect 26620 6684 27108 6712
rect 25685 6675 25743 6681
rect 28442 6672 28448 6724
rect 28500 6672 28506 6724
rect 28537 6715 28595 6721
rect 28537 6681 28549 6715
rect 28583 6712 28595 6715
rect 28718 6712 28724 6724
rect 28583 6684 28724 6712
rect 28583 6681 28595 6684
rect 28537 6675 28595 6681
rect 28718 6672 28724 6684
rect 28776 6672 28782 6724
rect 29546 6672 29552 6724
rect 29604 6712 29610 6724
rect 30101 6715 30159 6721
rect 30101 6712 30113 6715
rect 29604 6684 30113 6712
rect 29604 6672 29610 6684
rect 30101 6681 30113 6684
rect 30147 6681 30159 6715
rect 33778 6712 33784 6724
rect 33718 6684 33784 6712
rect 30101 6675 30159 6681
rect 33778 6672 33784 6684
rect 33836 6712 33842 6724
rect 34330 6712 34336 6724
rect 33836 6684 34336 6712
rect 33836 6672 33842 6684
rect 34330 6672 34336 6684
rect 34388 6672 34394 6724
rect 23934 6644 23940 6656
rect 23584 6616 23940 6644
rect 23934 6604 23940 6616
rect 23992 6604 23998 6656
rect 25130 6604 25136 6656
rect 25188 6604 25194 6656
rect 26602 6604 26608 6656
rect 26660 6644 26666 6656
rect 28074 6644 28080 6656
rect 26660 6616 28080 6644
rect 26660 6604 26666 6616
rect 28074 6604 28080 6616
rect 28132 6644 28138 6656
rect 28169 6647 28227 6653
rect 28169 6644 28181 6647
rect 28132 6616 28181 6644
rect 28132 6604 28138 6616
rect 28169 6613 28181 6616
rect 28215 6613 28227 6647
rect 28169 6607 28227 6613
rect 28350 6604 28356 6656
rect 28408 6644 28414 6656
rect 28813 6647 28871 6653
rect 28813 6644 28825 6647
rect 28408 6616 28825 6644
rect 28408 6604 28414 6616
rect 28813 6613 28825 6616
rect 28859 6613 28871 6647
rect 28813 6607 28871 6613
rect 30558 6604 30564 6656
rect 30616 6644 30622 6656
rect 30653 6647 30711 6653
rect 30653 6644 30665 6647
rect 30616 6616 30665 6644
rect 30616 6604 30622 6616
rect 30653 6613 30665 6616
rect 30699 6613 30711 6647
rect 30653 6607 30711 6613
rect 30929 6647 30987 6653
rect 30929 6613 30941 6647
rect 30975 6644 30987 6647
rect 31754 6644 31760 6656
rect 30975 6616 31760 6644
rect 30975 6613 30987 6616
rect 30929 6607 30987 6613
rect 31754 6604 31760 6616
rect 31812 6604 31818 6656
rect 32122 6604 32128 6656
rect 32180 6644 32186 6656
rect 36354 6644 36360 6656
rect 32180 6616 36360 6644
rect 32180 6604 32186 6616
rect 36354 6604 36360 6616
rect 36412 6604 36418 6656
rect 1104 6554 36524 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 36524 6554
rect 1104 6480 36524 6502
rect 11609 6443 11667 6449
rect 11609 6409 11621 6443
rect 11655 6440 11667 6443
rect 11698 6440 11704 6452
rect 11655 6412 11704 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 17678 6440 17684 6452
rect 16132 6412 17684 6440
rect 13262 6372 13268 6384
rect 11808 6344 13268 6372
rect 11808 6313 11836 6344
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13354 6332 13360 6384
rect 13412 6332 13418 6384
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15105 6375 15163 6381
rect 15105 6372 15117 6375
rect 15068 6344 15117 6372
rect 15068 6332 15074 6344
rect 15105 6341 15117 6344
rect 15151 6341 15163 6375
rect 16132 6372 16160 6412
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 23106 6400 23112 6452
rect 23164 6440 23170 6452
rect 25038 6440 25044 6452
rect 23164 6412 25044 6440
rect 23164 6400 23170 6412
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 26602 6440 26608 6452
rect 25332 6412 26608 6440
rect 15105 6335 15163 6341
rect 16040 6344 16160 6372
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11974 6264 11980 6316
rect 12032 6264 12038 6316
rect 12066 6264 12072 6316
rect 12124 6264 12130 6316
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11940 6208 12173 6236
rect 11940 6196 11946 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 13078 6196 13084 6248
rect 13136 6196 13142 6248
rect 13998 6196 14004 6248
rect 14056 6236 14062 6248
rect 14476 6236 14504 6290
rect 14918 6264 14924 6316
rect 14976 6304 14982 6316
rect 15749 6307 15807 6313
rect 15749 6304 15761 6307
rect 14976 6276 15761 6304
rect 14976 6264 14982 6276
rect 15749 6273 15761 6276
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16040 6313 16068 6344
rect 17586 6332 17592 6384
rect 17644 6332 17650 6384
rect 18874 6372 18880 6384
rect 18814 6344 18880 6372
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 20073 6375 20131 6381
rect 20073 6341 20085 6375
rect 20119 6372 20131 6375
rect 20438 6372 20444 6384
rect 20119 6344 20444 6372
rect 20119 6341 20131 6344
rect 20073 6335 20131 6341
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 20530 6332 20536 6384
rect 20588 6332 20594 6384
rect 24394 6332 24400 6384
rect 24452 6372 24458 6384
rect 25332 6372 25360 6412
rect 26602 6400 26608 6412
rect 26660 6400 26666 6452
rect 27522 6440 27528 6452
rect 26804 6412 27528 6440
rect 24452 6344 25360 6372
rect 25409 6375 25467 6381
rect 24452 6332 24458 6344
rect 25409 6341 25421 6375
rect 25455 6372 25467 6375
rect 26694 6372 26700 6384
rect 25455 6344 26700 6372
rect 25455 6341 25467 6344
rect 25409 6335 25467 6341
rect 26694 6332 26700 6344
rect 26752 6332 26758 6384
rect 26804 6381 26832 6412
rect 27522 6400 27528 6412
rect 27580 6400 27586 6452
rect 28442 6440 28448 6452
rect 27816 6412 28448 6440
rect 26789 6375 26847 6381
rect 26789 6341 26801 6375
rect 26835 6341 26847 6375
rect 26789 6335 26847 6341
rect 27338 6332 27344 6384
rect 27396 6372 27402 6384
rect 27816 6381 27844 6412
rect 28442 6400 28448 6412
rect 28500 6400 28506 6452
rect 30190 6400 30196 6452
rect 30248 6400 30254 6452
rect 33134 6440 33140 6452
rect 32140 6412 33140 6440
rect 27617 6375 27675 6381
rect 27617 6372 27629 6375
rect 27396 6344 27629 6372
rect 27396 6332 27402 6344
rect 27617 6341 27629 6344
rect 27663 6341 27675 6375
rect 27617 6335 27675 6341
rect 27801 6375 27859 6381
rect 27801 6341 27813 6375
rect 27847 6341 27859 6375
rect 27801 6335 27859 6341
rect 28169 6375 28227 6381
rect 28169 6341 28181 6375
rect 28215 6372 28227 6375
rect 28626 6372 28632 6384
rect 28215 6344 28632 6372
rect 28215 6341 28227 6344
rect 28169 6335 28227 6341
rect 28626 6332 28632 6344
rect 28684 6332 28690 6384
rect 28718 6332 28724 6384
rect 28776 6332 28782 6384
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16666 6304 16672 6316
rect 16163 6276 16672 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16666 6264 16672 6276
rect 16724 6264 16730 6316
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 17313 6307 17371 6313
rect 17313 6304 17325 6307
rect 17276 6276 17325 6304
rect 17276 6264 17282 6276
rect 17313 6273 17325 6276
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19024 6276 19625 6304
rect 19024 6264 19030 6276
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6273 20407 6307
rect 20349 6267 20407 6273
rect 17052 6236 17080 6264
rect 19150 6236 19156 6248
rect 14056 6208 16804 6236
rect 17052 6208 19156 6236
rect 14056 6196 14062 6208
rect 16776 6112 16804 6208
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19334 6196 19340 6248
rect 19392 6196 19398 6248
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 19705 6239 19763 6245
rect 19705 6236 19717 6239
rect 19576 6208 19717 6236
rect 19576 6196 19582 6208
rect 19705 6205 19717 6208
rect 19751 6236 19763 6239
rect 20180 6236 20208 6267
rect 19751 6208 20208 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 19352 6168 19380 6196
rect 19352 6140 19656 6168
rect 19628 6112 19656 6140
rect 19794 6128 19800 6180
rect 19852 6168 19858 6180
rect 20364 6168 20392 6267
rect 21634 6264 21640 6316
rect 21692 6304 21698 6316
rect 21910 6304 21916 6316
rect 21692 6276 21916 6304
rect 21692 6264 21698 6276
rect 21910 6264 21916 6276
rect 21968 6304 21974 6316
rect 23658 6304 23664 6316
rect 21968 6276 23664 6304
rect 21968 6264 21974 6276
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 25225 6307 25283 6313
rect 25225 6273 25237 6307
rect 25271 6304 25283 6307
rect 25774 6304 25780 6316
rect 25271 6276 25780 6304
rect 25271 6273 25283 6276
rect 25225 6267 25283 6273
rect 25774 6264 25780 6276
rect 25832 6264 25838 6316
rect 25866 6264 25872 6316
rect 25924 6304 25930 6316
rect 27246 6304 27252 6316
rect 25924 6276 27252 6304
rect 25924 6264 25930 6276
rect 27246 6264 27252 6276
rect 27304 6304 27310 6316
rect 27433 6307 27491 6313
rect 27433 6304 27445 6307
rect 27304 6276 27445 6304
rect 27304 6264 27310 6276
rect 27433 6273 27445 6276
rect 27479 6273 27491 6307
rect 27433 6267 27491 6273
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 27985 6307 28043 6313
rect 27985 6304 27997 6307
rect 27580 6276 27997 6304
rect 27580 6264 27586 6276
rect 27985 6273 27997 6276
rect 28031 6273 28043 6307
rect 27985 6267 28043 6273
rect 28258 6264 28264 6316
rect 28316 6304 28322 6316
rect 32140 6313 32168 6412
rect 33134 6400 33140 6412
rect 33192 6400 33198 6452
rect 33873 6443 33931 6449
rect 33873 6409 33885 6443
rect 33919 6440 33931 6443
rect 34514 6440 34520 6452
rect 33919 6412 34520 6440
rect 33919 6409 33931 6412
rect 33873 6403 33931 6409
rect 34514 6400 34520 6412
rect 34572 6400 34578 6452
rect 33778 6372 33784 6384
rect 33626 6344 33784 6372
rect 33778 6332 33784 6344
rect 33836 6332 33842 6384
rect 28445 6307 28503 6313
rect 28445 6304 28457 6307
rect 28316 6276 28457 6304
rect 28316 6264 28322 6276
rect 28445 6273 28457 6276
rect 28491 6273 28503 6307
rect 32125 6307 32183 6313
rect 28445 6267 28503 6273
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 26053 6239 26111 6245
rect 26053 6236 26065 6239
rect 24636 6208 26065 6236
rect 24636 6196 24642 6208
rect 26053 6205 26065 6208
rect 26099 6205 26111 6239
rect 26053 6199 26111 6205
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6236 26479 6239
rect 26786 6236 26792 6248
rect 26467 6208 26792 6236
rect 26467 6205 26479 6208
rect 26421 6199 26479 6205
rect 26786 6196 26792 6208
rect 26844 6196 26850 6248
rect 27062 6196 27068 6248
rect 27120 6196 27126 6248
rect 27157 6239 27215 6245
rect 27157 6205 27169 6239
rect 27203 6236 27215 6239
rect 29362 6236 29368 6248
rect 27203 6208 29368 6236
rect 27203 6205 27215 6208
rect 27157 6199 27215 6205
rect 29362 6196 29368 6208
rect 29420 6196 29426 6248
rect 29840 6236 29868 6290
rect 32125 6273 32137 6307
rect 32171 6273 32183 6307
rect 32125 6267 32183 6273
rect 29914 6236 29920 6248
rect 29840 6208 29920 6236
rect 29914 6196 29920 6208
rect 29972 6236 29978 6248
rect 32401 6239 32459 6245
rect 29972 6208 31754 6236
rect 29972 6196 29978 6208
rect 19852 6140 20392 6168
rect 19852 6128 19858 6140
rect 23014 6128 23020 6180
rect 23072 6168 23078 6180
rect 23934 6168 23940 6180
rect 23072 6140 23940 6168
rect 23072 6128 23078 6140
rect 23934 6128 23940 6140
rect 23992 6128 23998 6180
rect 24762 6128 24768 6180
rect 24820 6168 24826 6180
rect 31726 6168 31754 6208
rect 32401 6205 32413 6239
rect 32447 6236 32459 6239
rect 32766 6236 32772 6248
rect 32447 6208 32772 6236
rect 32447 6205 32459 6208
rect 32401 6199 32459 6205
rect 32766 6196 32772 6208
rect 32824 6196 32830 6248
rect 24820 6140 28212 6168
rect 31726 6140 32260 6168
rect 24820 6128 24826 6140
rect 12802 6060 12808 6112
rect 12860 6060 12866 6112
rect 15470 6060 15476 6112
rect 15528 6100 15534 6112
rect 15565 6103 15623 6109
rect 15565 6100 15577 6103
rect 15528 6072 15577 6100
rect 15528 6060 15534 6072
rect 15565 6069 15577 6072
rect 15611 6069 15623 6103
rect 15565 6063 15623 6069
rect 16758 6060 16764 6112
rect 16816 6060 16822 6112
rect 17218 6060 17224 6112
rect 17276 6100 17282 6112
rect 17770 6100 17776 6112
rect 17276 6072 17776 6100
rect 17276 6060 17282 6072
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 19426 6060 19432 6112
rect 19484 6060 19490 6112
rect 19610 6060 19616 6112
rect 19668 6060 19674 6112
rect 22002 6060 22008 6112
rect 22060 6100 22066 6112
rect 25130 6100 25136 6112
rect 22060 6072 25136 6100
rect 22060 6060 22066 6072
rect 25130 6060 25136 6072
rect 25188 6060 25194 6112
rect 25682 6060 25688 6112
rect 25740 6060 25746 6112
rect 26510 6060 26516 6112
rect 26568 6060 26574 6112
rect 26651 6103 26709 6109
rect 26651 6069 26663 6103
rect 26697 6100 26709 6103
rect 27338 6100 27344 6112
rect 26697 6072 27344 6100
rect 26697 6069 26709 6072
rect 26651 6063 26709 6069
rect 27338 6060 27344 6072
rect 27396 6060 27402 6112
rect 28184 6100 28212 6140
rect 32122 6100 32128 6112
rect 28184 6072 32128 6100
rect 32122 6060 32128 6072
rect 32180 6060 32186 6112
rect 32232 6100 32260 6140
rect 33778 6100 33784 6112
rect 32232 6072 33784 6100
rect 33778 6060 33784 6072
rect 33836 6060 33842 6112
rect 1104 6010 36524 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 36524 6010
rect 1104 5936 36524 5958
rect 10400 5899 10458 5905
rect 10400 5865 10412 5899
rect 10446 5896 10458 5899
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 10446 5868 11989 5896
rect 10446 5865 10458 5868
rect 10400 5859 10458 5865
rect 11977 5865 11989 5868
rect 12023 5865 12035 5899
rect 11977 5859 12035 5865
rect 13081 5899 13139 5905
rect 13081 5865 13093 5899
rect 13127 5896 13139 5899
rect 13722 5896 13728 5908
rect 13127 5868 13728 5896
rect 13127 5865 13139 5868
rect 13081 5859 13139 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 14274 5856 14280 5908
rect 14332 5896 14338 5908
rect 16945 5899 17003 5905
rect 14332 5868 16896 5896
rect 14332 5856 14338 5868
rect 12618 5828 12624 5840
rect 12452 5800 12624 5828
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5760 10195 5763
rect 11422 5760 11428 5772
rect 10183 5732 11428 5760
rect 10183 5729 10195 5732
rect 10137 5723 10195 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 12452 5769 12480 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 16868 5828 16896 5868
rect 16945 5865 16957 5899
rect 16991 5896 17003 5899
rect 17310 5896 17316 5908
rect 16991 5868 17316 5896
rect 16991 5865 17003 5868
rect 16945 5859 17003 5865
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 18874 5856 18880 5908
rect 18932 5896 18938 5908
rect 19058 5896 19064 5908
rect 18932 5868 19064 5896
rect 18932 5856 18938 5868
rect 19058 5856 19064 5868
rect 19116 5896 19122 5908
rect 19429 5899 19487 5905
rect 19429 5896 19441 5899
rect 19116 5868 19441 5896
rect 19116 5856 19122 5868
rect 19429 5865 19441 5868
rect 19475 5865 19487 5899
rect 23753 5899 23811 5905
rect 23753 5896 23765 5899
rect 19429 5859 19487 5865
rect 21744 5868 23765 5896
rect 21744 5840 21772 5868
rect 19610 5828 19616 5840
rect 16868 5800 19616 5828
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 12529 5763 12587 5769
rect 12529 5729 12541 5763
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5760 13323 5763
rect 13630 5760 13636 5772
rect 13311 5732 13636 5760
rect 13311 5729 13323 5732
rect 13265 5723 13323 5729
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 12544 5692 12572 5723
rect 13630 5720 13636 5732
rect 13688 5760 13694 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 13688 5732 14565 5760
rect 13688 5720 13694 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 12308 5664 12572 5692
rect 13173 5695 13231 5701
rect 12308 5652 12314 5664
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 12345 5627 12403 5633
rect 11638 5596 12296 5624
rect 11882 5516 11888 5568
rect 11940 5516 11946 5568
rect 12268 5556 12296 5596
rect 12345 5593 12357 5627
rect 12391 5624 12403 5627
rect 12802 5624 12808 5636
rect 12391 5596 12808 5624
rect 12391 5593 12403 5596
rect 12345 5587 12403 5593
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 13188 5624 13216 5655
rect 13814 5652 13820 5704
rect 13872 5652 13878 5704
rect 14752 5624 14780 5723
rect 15470 5720 15476 5772
rect 15528 5720 15534 5772
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 18414 5652 18420 5704
rect 18472 5692 18478 5704
rect 18892 5701 18920 5800
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 21726 5828 21732 5840
rect 20680 5800 21732 5828
rect 20680 5788 20686 5800
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 21818 5788 21824 5840
rect 21876 5828 21882 5840
rect 21876 5800 22600 5828
rect 21876 5788 21882 5800
rect 21082 5760 21088 5772
rect 20916 5732 21088 5760
rect 18693 5695 18751 5701
rect 18693 5692 18705 5695
rect 18472 5664 18705 5692
rect 18472 5652 18478 5664
rect 18693 5661 18705 5664
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 18966 5652 18972 5704
rect 19024 5652 19030 5704
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 19208 5664 19257 5692
rect 19208 5652 19214 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 20916 5701 20944 5732
rect 21082 5720 21088 5732
rect 21140 5720 21146 5772
rect 21284 5732 22140 5760
rect 21284 5704 21312 5732
rect 22112 5704 22140 5732
rect 19889 5695 19947 5701
rect 19889 5692 19901 5695
rect 19576 5664 19901 5692
rect 19576 5652 19582 5664
rect 19889 5661 19901 5664
rect 19935 5661 19947 5695
rect 19889 5655 19947 5661
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 20625 5695 20683 5701
rect 20625 5692 20637 5695
rect 20579 5664 20637 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 20625 5661 20637 5664
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 21048 5664 21189 5692
rect 21048 5652 21054 5664
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 21266 5652 21272 5704
rect 21324 5652 21330 5704
rect 21726 5652 21732 5704
rect 21784 5652 21790 5704
rect 22002 5652 22008 5704
rect 22060 5652 22066 5704
rect 22094 5652 22100 5704
rect 22152 5652 22158 5704
rect 16758 5624 16764 5636
rect 13188 5596 14504 5624
rect 14752 5596 15884 5624
rect 16698 5596 16764 5624
rect 13998 5556 14004 5568
rect 12268 5528 14004 5556
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 14476 5565 14504 5596
rect 14461 5559 14519 5565
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 14826 5556 14832 5568
rect 14507 5528 14832 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 15856 5556 15884 5596
rect 16758 5584 16764 5596
rect 16816 5584 16822 5636
rect 17310 5584 17316 5636
rect 17368 5624 17374 5636
rect 18984 5624 19012 5652
rect 17368 5596 19012 5624
rect 17368 5584 17374 5596
rect 20806 5584 20812 5636
rect 20864 5624 20870 5636
rect 21085 5627 21143 5633
rect 21085 5624 21097 5627
rect 20864 5596 21097 5624
rect 20864 5584 20870 5596
rect 21085 5593 21097 5596
rect 21131 5624 21143 5627
rect 21818 5624 21824 5636
rect 21131 5596 21824 5624
rect 21131 5593 21143 5596
rect 21085 5587 21143 5593
rect 21818 5584 21824 5596
rect 21876 5624 21882 5636
rect 21913 5627 21971 5633
rect 21913 5624 21925 5627
rect 21876 5596 21925 5624
rect 21876 5584 21882 5596
rect 21913 5593 21925 5596
rect 21959 5593 21971 5627
rect 22020 5624 22048 5652
rect 22572 5624 22600 5800
rect 22649 5695 22707 5701
rect 22649 5661 22661 5695
rect 22695 5692 22707 5695
rect 22922 5692 22928 5704
rect 22695 5664 22928 5692
rect 22695 5661 22707 5664
rect 22649 5655 22707 5661
rect 22922 5652 22928 5664
rect 22980 5652 22986 5704
rect 23014 5652 23020 5704
rect 23072 5652 23078 5704
rect 23124 5692 23152 5868
rect 23753 5865 23765 5868
rect 23799 5896 23811 5899
rect 23842 5896 23848 5908
rect 23799 5868 23848 5896
rect 23799 5865 23811 5868
rect 23753 5859 23811 5865
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 29549 5899 29607 5905
rect 29549 5865 29561 5899
rect 29595 5896 29607 5899
rect 29638 5896 29644 5908
rect 29595 5868 29644 5896
rect 29595 5865 29607 5868
rect 29549 5859 29607 5865
rect 29638 5856 29644 5868
rect 29696 5856 29702 5908
rect 33873 5899 33931 5905
rect 33873 5865 33885 5899
rect 33919 5896 33931 5899
rect 34146 5896 34152 5908
rect 33919 5868 34152 5896
rect 33919 5865 33931 5868
rect 33873 5859 33931 5865
rect 34146 5856 34152 5868
rect 34204 5856 34210 5908
rect 23934 5788 23940 5840
rect 23992 5828 23998 5840
rect 25317 5831 25375 5837
rect 25317 5828 25329 5831
rect 23992 5800 25329 5828
rect 23992 5788 23998 5800
rect 24486 5760 24492 5772
rect 23400 5732 24492 5760
rect 23400 5704 23428 5732
rect 24486 5720 24492 5732
rect 24544 5720 24550 5772
rect 23293 5695 23351 5701
rect 23293 5692 23305 5695
rect 23124 5664 23305 5692
rect 23293 5661 23305 5664
rect 23339 5661 23351 5695
rect 23293 5655 23351 5661
rect 23382 5652 23388 5704
rect 23440 5652 23446 5704
rect 23934 5652 23940 5704
rect 23992 5652 23998 5704
rect 24670 5652 24676 5704
rect 24728 5652 24734 5704
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 24964 5701 24992 5800
rect 25317 5797 25329 5800
rect 25363 5797 25375 5831
rect 25317 5791 25375 5797
rect 28258 5720 28264 5772
rect 28316 5760 28322 5772
rect 31297 5763 31355 5769
rect 31297 5760 31309 5763
rect 28316 5732 31309 5760
rect 28316 5720 28322 5732
rect 31297 5729 31309 5732
rect 31343 5760 31355 5763
rect 32125 5763 32183 5769
rect 32125 5760 32137 5763
rect 31343 5732 32137 5760
rect 31343 5729 31355 5732
rect 31297 5723 31355 5729
rect 32125 5729 32137 5732
rect 32171 5760 32183 5763
rect 33134 5760 33140 5772
rect 32171 5732 33140 5760
rect 32171 5729 32183 5732
rect 32125 5723 32183 5729
rect 33134 5720 33140 5732
rect 33192 5720 33198 5772
rect 24857 5695 24915 5701
rect 24857 5692 24869 5695
rect 24820 5664 24869 5692
rect 24820 5652 24826 5664
rect 24857 5661 24869 5664
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 25041 5695 25099 5701
rect 25041 5661 25053 5695
rect 25087 5661 25099 5695
rect 25041 5655 25099 5661
rect 25501 5695 25559 5701
rect 25501 5661 25513 5695
rect 25547 5692 25559 5695
rect 25682 5692 25688 5704
rect 25547 5664 25688 5692
rect 25547 5661 25559 5664
rect 25501 5655 25559 5661
rect 23201 5627 23259 5633
rect 23201 5624 23213 5627
rect 22020 5596 22508 5624
rect 22572 5596 23213 5624
rect 21913 5587 21971 5593
rect 16850 5556 16856 5568
rect 15856 5528 16856 5556
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17494 5516 17500 5568
rect 17552 5556 17558 5568
rect 17773 5559 17831 5565
rect 17773 5556 17785 5559
rect 17552 5528 17785 5556
rect 17552 5516 17558 5528
rect 17773 5525 17785 5528
rect 17819 5525 17831 5559
rect 17773 5519 17831 5525
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18509 5559 18567 5565
rect 18509 5556 18521 5559
rect 18012 5528 18521 5556
rect 18012 5516 18018 5528
rect 18509 5525 18521 5528
rect 18555 5525 18567 5559
rect 18509 5519 18567 5525
rect 20714 5516 20720 5568
rect 20772 5516 20778 5568
rect 21453 5559 21511 5565
rect 21453 5525 21465 5559
rect 21499 5556 21511 5559
rect 22094 5556 22100 5568
rect 21499 5528 22100 5556
rect 21499 5525 21511 5528
rect 21453 5519 21511 5525
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 22278 5516 22284 5568
rect 22336 5516 22342 5568
rect 22480 5565 22508 5596
rect 23201 5593 23213 5596
rect 23247 5593 23259 5627
rect 24780 5624 24808 5652
rect 25056 5624 25084 5655
rect 25682 5652 25688 5664
rect 25740 5652 25746 5704
rect 29914 5652 29920 5704
rect 29972 5652 29978 5704
rect 23201 5587 23259 5593
rect 23400 5596 24808 5624
rect 24964 5596 25084 5624
rect 22465 5559 22523 5565
rect 22465 5525 22477 5559
rect 22511 5525 22523 5559
rect 23216 5556 23244 5587
rect 23400 5556 23428 5596
rect 23216 5528 23428 5556
rect 22465 5519 22523 5525
rect 23566 5516 23572 5568
rect 23624 5516 23630 5568
rect 24486 5516 24492 5568
rect 24544 5556 24550 5568
rect 24964 5556 24992 5596
rect 31018 5584 31024 5636
rect 31076 5584 31082 5636
rect 32398 5584 32404 5636
rect 32456 5584 32462 5636
rect 33778 5624 33784 5636
rect 33626 5596 33784 5624
rect 33778 5584 33784 5596
rect 33836 5584 33842 5636
rect 24544 5528 24992 5556
rect 25225 5559 25283 5565
rect 24544 5516 24550 5528
rect 25225 5525 25237 5559
rect 25271 5556 25283 5559
rect 25314 5556 25320 5568
rect 25271 5528 25320 5556
rect 25271 5525 25283 5528
rect 25225 5519 25283 5525
rect 25314 5516 25320 5528
rect 25372 5516 25378 5568
rect 1104 5466 36524 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 36524 5466
rect 1104 5392 36524 5414
rect 12158 5312 12164 5364
rect 12216 5352 12222 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 12216 5324 12265 5352
rect 12216 5312 12222 5324
rect 12253 5321 12265 5324
rect 12299 5321 12311 5355
rect 12253 5315 12311 5321
rect 12621 5355 12679 5361
rect 12621 5321 12633 5355
rect 12667 5352 12679 5355
rect 13814 5352 13820 5364
rect 12667 5324 13820 5352
rect 12667 5321 12679 5324
rect 12621 5315 12679 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 17586 5352 17592 5364
rect 17236 5324 17592 5352
rect 13998 5284 14004 5296
rect 13662 5256 14004 5284
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 14090 5244 14096 5296
rect 14148 5244 14154 5296
rect 15286 5284 15292 5296
rect 14384 5256 15292 5284
rect 12158 5176 12164 5228
rect 12216 5176 12222 5228
rect 14384 5225 14412 5256
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 17236 5225 17264 5324
rect 17586 5312 17592 5324
rect 17644 5352 17650 5364
rect 17862 5352 17868 5364
rect 17644 5324 17868 5352
rect 17644 5312 17650 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 19518 5312 19524 5364
rect 19576 5312 19582 5364
rect 19610 5312 19616 5364
rect 19668 5352 19674 5364
rect 26418 5352 26424 5364
rect 19668 5324 21864 5352
rect 19668 5312 19674 5324
rect 17954 5284 17960 5296
rect 17420 5256 17960 5284
rect 17420 5225 17448 5256
rect 17954 5244 17960 5256
rect 18012 5244 18018 5296
rect 19334 5284 19340 5296
rect 19274 5256 19340 5284
rect 19334 5244 19340 5256
rect 19392 5284 19398 5296
rect 20346 5284 20352 5296
rect 19392 5256 20352 5284
rect 19392 5244 19398 5256
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 21836 5284 21864 5324
rect 24872 5324 26424 5352
rect 22370 5284 22376 5296
rect 21836 5256 22376 5284
rect 14369 5219 14427 5225
rect 14369 5185 14381 5219
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15749 5219 15807 5225
rect 15749 5216 15761 5219
rect 15243 5188 15761 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 15749 5185 15761 5188
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 17221 5219 17279 5225
rect 17221 5185 17233 5219
rect 17267 5185 17279 5219
rect 17221 5179 17279 5185
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 17678 5176 17684 5228
rect 17736 5176 17742 5228
rect 19610 5176 19616 5228
rect 19668 5176 19674 5228
rect 21836 5225 21864 5256
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 22554 5244 22560 5296
rect 22612 5244 22618 5296
rect 24305 5287 24363 5293
rect 24305 5253 24317 5287
rect 24351 5284 24363 5287
rect 24762 5284 24768 5296
rect 24351 5256 24768 5284
rect 24351 5253 24363 5256
rect 24305 5247 24363 5253
rect 24762 5244 24768 5256
rect 24820 5244 24826 5296
rect 24872 5228 24900 5324
rect 26418 5312 26424 5324
rect 26476 5352 26482 5364
rect 26878 5352 26884 5364
rect 26476 5324 26884 5352
rect 26476 5312 26482 5324
rect 26878 5312 26884 5324
rect 26936 5312 26942 5364
rect 25130 5244 25136 5296
rect 25188 5284 25194 5296
rect 25188 5256 25622 5284
rect 25188 5244 25194 5256
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 24121 5219 24179 5225
rect 24121 5185 24133 5219
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 12345 5151 12403 5157
rect 12345 5148 12357 5151
rect 12308 5120 12357 5148
rect 12308 5108 12314 5120
rect 12345 5117 12357 5120
rect 12391 5117 12403 5151
rect 12345 5111 12403 5117
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 14976 5120 15301 5148
rect 14976 5108 14982 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 15378 5108 15384 5160
rect 15436 5108 15442 5160
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 16301 5151 16359 5157
rect 16301 5148 16313 5151
rect 16264 5120 16313 5148
rect 16264 5108 16270 5120
rect 16301 5117 16313 5120
rect 16347 5117 16359 5151
rect 16301 5111 16359 5117
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 16908 5120 17325 5148
rect 16908 5108 16914 5120
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 17770 5108 17776 5160
rect 17828 5108 17834 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 19242 5148 19248 5160
rect 18095 5120 19248 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 19242 5108 19248 5120
rect 19300 5108 19306 5160
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5148 19947 5151
rect 20346 5148 20352 5160
rect 19935 5120 20352 5148
rect 19935 5117 19947 5120
rect 19889 5111 19947 5117
rect 20346 5108 20352 5120
rect 20404 5108 20410 5160
rect 21637 5151 21695 5157
rect 21637 5117 21649 5151
rect 21683 5117 21695 5151
rect 21637 5111 21695 5117
rect 21082 5080 21088 5092
rect 16316 5052 17908 5080
rect 16316 5024 16344 5052
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 11572 4984 11805 5012
rect 11572 4972 11578 4984
rect 11793 4981 11805 4984
rect 11839 4981 11851 5015
rect 11793 4975 11851 4981
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 14829 5015 14887 5021
rect 14829 5012 14841 5015
rect 14700 4984 14841 5012
rect 14700 4972 14706 4984
rect 14829 4981 14841 4984
rect 14875 4981 14887 5015
rect 14829 4975 14887 4981
rect 16298 4972 16304 5024
rect 16356 4972 16362 5024
rect 16482 4972 16488 5024
rect 16540 5012 16546 5024
rect 17037 5015 17095 5021
rect 17037 5012 17049 5015
rect 16540 4984 17049 5012
rect 16540 4972 16546 4984
rect 17037 4981 17049 4984
rect 17083 4981 17095 5015
rect 17880 5012 17908 5052
rect 20916 5052 21088 5080
rect 20916 5012 20944 5052
rect 21082 5040 21088 5052
rect 21140 5080 21146 5092
rect 21652 5080 21680 5111
rect 22094 5108 22100 5160
rect 22152 5108 22158 5160
rect 23845 5151 23903 5157
rect 23845 5117 23857 5151
rect 23891 5148 23903 5151
rect 24136 5148 24164 5179
rect 24394 5176 24400 5228
rect 24452 5176 24458 5228
rect 24486 5176 24492 5228
rect 24544 5176 24550 5228
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 25133 5151 25191 5157
rect 25133 5148 25145 5151
rect 23891 5120 24164 5148
rect 24688 5120 25145 5148
rect 23891 5117 23903 5120
rect 23845 5111 23903 5117
rect 21140 5052 21680 5080
rect 21140 5040 21146 5052
rect 17880 4984 20944 5012
rect 17037 4975 17095 4981
rect 20990 4972 20996 5024
rect 21048 5012 21054 5024
rect 23860 5012 23888 5111
rect 24688 5089 24716 5120
rect 25133 5117 25145 5120
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 24673 5083 24731 5089
rect 24673 5049 24685 5083
rect 24719 5049 24731 5083
rect 24673 5043 24731 5049
rect 21048 4984 23888 5012
rect 21048 4972 21054 4984
rect 24394 4972 24400 5024
rect 24452 5012 24458 5024
rect 26605 5015 26663 5021
rect 26605 5012 26617 5015
rect 24452 4984 26617 5012
rect 24452 4972 24458 4984
rect 26605 4981 26617 4984
rect 26651 4981 26663 5015
rect 26605 4975 26663 4981
rect 1104 4922 36524 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 36524 4922
rect 1104 4848 36524 4870
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 19610 4808 19616 4820
rect 16172 4780 19616 4808
rect 16172 4768 16178 4780
rect 19610 4768 19616 4780
rect 19668 4808 19674 4820
rect 20073 4811 20131 4817
rect 20073 4808 20085 4811
rect 19668 4780 20085 4808
rect 19668 4768 19674 4780
rect 20073 4777 20085 4780
rect 20119 4777 20131 4811
rect 20073 4771 20131 4777
rect 20346 4768 20352 4820
rect 20404 4768 20410 4820
rect 22922 4768 22928 4820
rect 22980 4808 22986 4820
rect 23845 4811 23903 4817
rect 23845 4808 23857 4811
rect 22980 4780 23857 4808
rect 22980 4768 22986 4780
rect 23845 4777 23857 4780
rect 23891 4777 23903 4811
rect 23845 4771 23903 4777
rect 26694 4768 26700 4820
rect 26752 4808 26758 4820
rect 26789 4811 26847 4817
rect 26789 4808 26801 4811
rect 26752 4780 26801 4808
rect 26752 4768 26758 4780
rect 26789 4777 26801 4780
rect 26835 4777 26847 4811
rect 26789 4771 26847 4777
rect 17957 4743 18015 4749
rect 17957 4709 17969 4743
rect 18003 4740 18015 4743
rect 18414 4740 18420 4752
rect 18003 4712 18420 4740
rect 18003 4709 18015 4712
rect 17957 4703 18015 4709
rect 18414 4700 18420 4712
rect 18472 4740 18478 4752
rect 20254 4740 20260 4752
rect 18472 4712 20260 4740
rect 18472 4700 18478 4712
rect 20254 4700 20260 4712
rect 20312 4700 20318 4752
rect 13078 4672 13084 4684
rect 11256 4644 13084 4672
rect 11256 4613 11284 4644
rect 13078 4632 13084 4644
rect 13136 4672 13142 4684
rect 14369 4675 14427 4681
rect 14369 4672 14381 4675
rect 13136 4644 14381 4672
rect 13136 4632 13142 4644
rect 14369 4641 14381 4644
rect 14415 4672 14427 4675
rect 15194 4672 15200 4684
rect 14415 4644 15200 4672
rect 14415 4641 14427 4644
rect 14369 4635 14427 4641
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15344 4644 16221 4672
rect 15344 4632 15350 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16209 4635 16267 4641
rect 16482 4632 16488 4684
rect 16540 4632 16546 4684
rect 16850 4632 16856 4684
rect 16908 4672 16914 4684
rect 21266 4672 21272 4684
rect 16908 4644 21272 4672
rect 16908 4632 16914 4644
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 13814 4604 13820 4616
rect 13403 4576 13820 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 11256 4536 11284 4567
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 18690 4564 18696 4616
rect 18748 4564 18754 4616
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19886 4564 19892 4616
rect 19944 4564 19950 4616
rect 20548 4613 20576 4644
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 22094 4632 22100 4684
rect 22152 4672 22158 4684
rect 23106 4672 23112 4684
rect 22152 4644 23112 4672
rect 22152 4632 22158 4644
rect 23106 4632 23112 4644
rect 23164 4632 23170 4684
rect 24854 4632 24860 4684
rect 24912 4672 24918 4684
rect 25041 4675 25099 4681
rect 25041 4672 25053 4675
rect 24912 4644 25053 4672
rect 24912 4632 24918 4644
rect 25041 4641 25053 4644
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 25314 4632 25320 4684
rect 25372 4632 25378 4684
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20533 4607 20591 4613
rect 20533 4573 20545 4607
rect 20579 4573 20591 4607
rect 20533 4567 20591 4573
rect 20717 4607 20775 4613
rect 20717 4573 20729 4607
rect 20763 4604 20775 4607
rect 20806 4604 20812 4616
rect 20763 4576 20812 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 11422 4536 11428 4548
rect 11256 4508 11428 4536
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 11514 4496 11520 4548
rect 11572 4496 11578 4548
rect 13170 4536 13176 4548
rect 12742 4508 13176 4536
rect 13170 4496 13176 4508
rect 13228 4536 13234 4548
rect 13998 4536 14004 4548
rect 13228 4508 14004 4536
rect 13228 4496 13234 4508
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 14642 4496 14648 4548
rect 14700 4496 14706 4548
rect 18230 4536 18236 4548
rect 15870 4508 16896 4536
rect 17710 4508 18236 4536
rect 12986 4428 12992 4480
rect 13044 4428 13050 4480
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14918 4468 14924 4480
rect 13955 4440 14924 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 16117 4471 16175 4477
rect 16117 4437 16129 4471
rect 16163 4468 16175 4471
rect 16206 4468 16212 4480
rect 16163 4440 16212 4468
rect 16163 4437 16175 4440
rect 16117 4431 16175 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 16868 4468 16896 4508
rect 17788 4468 17816 4508
rect 18230 4496 18236 4508
rect 18288 4536 18294 4548
rect 19058 4536 19064 4548
rect 18288 4508 19064 4536
rect 18288 4496 18294 4508
rect 19058 4496 19064 4508
rect 19116 4496 19122 4548
rect 16868 4440 17816 4468
rect 18138 4428 18144 4480
rect 18196 4428 18202 4480
rect 20272 4468 20300 4567
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21910 4604 21916 4616
rect 20947 4576 21916 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 20625 4539 20683 4545
rect 20625 4505 20637 4539
rect 20671 4536 20683 4539
rect 21082 4536 21088 4548
rect 20671 4508 21088 4536
rect 20671 4505 20683 4508
rect 20625 4499 20683 4505
rect 21082 4496 21088 4508
rect 21140 4496 21146 4548
rect 22278 4496 22284 4548
rect 22336 4536 22342 4548
rect 22373 4539 22431 4545
rect 22373 4536 22385 4539
rect 22336 4508 22385 4536
rect 22336 4496 22342 4508
rect 22373 4505 22385 4508
rect 22419 4505 22431 4539
rect 22373 4499 22431 4505
rect 22646 4496 22652 4548
rect 22704 4536 22710 4548
rect 22704 4508 22862 4536
rect 22704 4496 22710 4508
rect 25222 4496 25228 4548
rect 25280 4536 25286 4548
rect 25280 4508 25806 4536
rect 25280 4496 25286 4508
rect 27338 4468 27344 4480
rect 20272 4440 27344 4468
rect 27338 4428 27344 4440
rect 27396 4428 27402 4480
rect 1104 4378 36524 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 36524 4378
rect 1104 4304 36524 4326
rect 11977 4267 12035 4273
rect 11977 4233 11989 4267
rect 12023 4264 12035 4267
rect 12158 4264 12164 4276
rect 12023 4236 12164 4264
rect 12023 4233 12035 4236
rect 11977 4227 12035 4233
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 14918 4224 14924 4276
rect 14976 4224 14982 4276
rect 17678 4264 17684 4276
rect 17420 4236 17684 4264
rect 13170 4156 13176 4208
rect 13228 4156 13234 4208
rect 15286 4196 15292 4208
rect 14476 4168 15292 4196
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 4062 4128 4068 4140
rect 2087 4100 4068 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 14476 4137 14504 4168
rect 15286 4156 15292 4168
rect 15344 4156 15350 4208
rect 16025 4199 16083 4205
rect 16025 4165 16037 4199
rect 16071 4196 16083 4199
rect 16669 4199 16727 4205
rect 16669 4196 16681 4199
rect 16071 4168 16681 4196
rect 16071 4165 16083 4168
rect 16025 4159 16083 4165
rect 16669 4165 16681 4168
rect 16715 4165 16727 4199
rect 16669 4159 16727 4165
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14792 4100 15025 4128
rect 14792 4088 14798 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 15838 4088 15844 4140
rect 15896 4128 15902 4140
rect 17420 4137 17448 4236
rect 17678 4224 17684 4236
rect 17736 4264 17742 4276
rect 17736 4236 19380 4264
rect 17736 4224 17742 4236
rect 17497 4199 17555 4205
rect 17497 4165 17509 4199
rect 17543 4196 17555 4199
rect 17586 4196 17592 4208
rect 17543 4168 17592 4196
rect 17543 4165 17555 4168
rect 17497 4159 17555 4165
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 18049 4199 18107 4205
rect 18049 4165 18061 4199
rect 18095 4196 18107 4199
rect 18138 4196 18144 4208
rect 18095 4168 18144 4196
rect 18095 4165 18107 4168
rect 18049 4159 18107 4165
rect 18138 4156 18144 4168
rect 18196 4156 18202 4208
rect 19058 4156 19064 4208
rect 19116 4156 19122 4208
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15896 4100 16129 4128
rect 15896 4088 15902 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 17678 4088 17684 4140
rect 17736 4088 17742 4140
rect 11330 4020 11336 4072
rect 11388 4020 11394 4072
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4060 12679 4063
rect 12986 4060 12992 4072
rect 12667 4032 12992 4060
rect 12667 4029 12679 4032
rect 12621 4023 12679 4029
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 15197 4063 15255 4069
rect 14231 4032 14596 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 934 3952 940 4004
rect 992 3992 998 4004
rect 14568 4001 14596 4032
rect 15197 4029 15209 4063
rect 15243 4060 15255 4063
rect 15378 4060 15384 4072
rect 15243 4032 15384 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 15378 4020 15384 4032
rect 15436 4060 15442 4072
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 15436 4032 16221 4060
rect 15436 4020 15442 4032
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 1857 3995 1915 4001
rect 1857 3992 1869 3995
rect 992 3964 1869 3992
rect 992 3952 998 3964
rect 1857 3961 1869 3964
rect 1903 3961 1915 3995
rect 1857 3955 1915 3961
rect 14553 3995 14611 4001
rect 14553 3961 14565 3995
rect 14599 3961 14611 3995
rect 14553 3955 14611 3961
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 17328 3992 17356 4023
rect 17770 4020 17776 4072
rect 17828 4020 17834 4072
rect 18506 4060 18512 4072
rect 17880 4032 18512 4060
rect 17880 3992 17908 4032
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 17000 3964 17908 3992
rect 19352 3992 19380 4236
rect 19886 4224 19892 4276
rect 19944 4224 19950 4276
rect 25608 4236 27200 4264
rect 22646 4156 22652 4208
rect 22704 4196 22710 4208
rect 24026 4196 24032 4208
rect 22704 4168 24032 4196
rect 22704 4156 22710 4168
rect 24026 4156 24032 4168
rect 24084 4156 24090 4208
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 20165 4131 20223 4137
rect 19484 4100 19932 4128
rect 19484 4088 19490 4100
rect 19518 4020 19524 4072
rect 19576 4060 19582 4072
rect 19794 4060 19800 4072
rect 19576 4032 19800 4060
rect 19576 4020 19582 4032
rect 19794 4020 19800 4032
rect 19852 4020 19858 4072
rect 19904 4069 19932 4100
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4029 19947 4063
rect 20180 4060 20208 4091
rect 20254 4088 20260 4140
rect 20312 4088 20318 4140
rect 23290 4088 23296 4140
rect 23348 4088 23354 4140
rect 24854 4088 24860 4140
rect 24912 4128 24918 4140
rect 25133 4131 25191 4137
rect 25133 4128 25145 4131
rect 24912 4100 25145 4128
rect 24912 4088 24918 4100
rect 25133 4097 25145 4100
rect 25179 4128 25191 4131
rect 25608 4128 25636 4236
rect 27172 4205 27200 4236
rect 26973 4199 27031 4205
rect 26973 4196 26985 4199
rect 25179 4100 25636 4128
rect 26436 4168 26985 4196
rect 25179 4097 25191 4100
rect 25133 4091 25191 4097
rect 20714 4060 20720 4072
rect 20180 4032 20720 4060
rect 19889 4023 19947 4029
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 23566 4020 23572 4072
rect 23624 4020 23630 4072
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 23992 4032 25053 4060
rect 23992 4020 23998 4032
rect 25041 4029 25053 4032
rect 25087 4029 25099 4063
rect 25041 4023 25099 4029
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26436 4069 26464 4168
rect 26973 4165 26985 4168
rect 27019 4165 27031 4199
rect 26973 4159 27031 4165
rect 27157 4199 27215 4205
rect 27157 4165 27169 4199
rect 27203 4165 27215 4199
rect 27157 4159 27215 4165
rect 26789 4131 26847 4137
rect 26789 4097 26801 4131
rect 26835 4097 26847 4131
rect 26789 4091 26847 4097
rect 27341 4131 27399 4137
rect 27341 4097 27353 4131
rect 27387 4128 27399 4131
rect 36446 4128 36452 4140
rect 27387 4100 36452 4128
rect 27387 4097 27399 4100
rect 27341 4091 27399 4097
rect 26421 4063 26479 4069
rect 26421 4060 26433 4063
rect 26384 4032 26433 4060
rect 26384 4020 26390 4032
rect 26421 4029 26433 4032
rect 26467 4029 26479 4063
rect 26804 4060 26832 4091
rect 27356 4060 27384 4091
rect 36446 4088 36452 4100
rect 36504 4088 36510 4140
rect 26804 4032 27384 4060
rect 26421 4023 26479 4029
rect 19702 3992 19708 4004
rect 19352 3964 19708 3992
rect 17000 3952 17006 3964
rect 19702 3952 19708 3964
rect 19760 3992 19766 4004
rect 20073 3995 20131 4001
rect 20073 3992 20085 3995
rect 19760 3964 20085 3992
rect 19760 3952 19766 3964
rect 20073 3961 20085 3964
rect 20119 3961 20131 3995
rect 20073 3955 20131 3961
rect 25501 3995 25559 4001
rect 25501 3961 25513 3995
rect 25547 3992 25559 3995
rect 25869 3995 25927 4001
rect 25869 3992 25881 3995
rect 25547 3964 25881 3992
rect 25547 3961 25559 3964
rect 25501 3955 25559 3961
rect 25869 3961 25881 3964
rect 25915 3961 25927 3995
rect 25869 3955 25927 3961
rect 10689 3927 10747 3933
rect 10689 3893 10701 3927
rect 10735 3924 10747 3927
rect 10962 3924 10968 3936
rect 10735 3896 10968 3924
rect 10735 3893 10747 3896
rect 10689 3887 10747 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3924 12771 3927
rect 13814 3924 13820 3936
rect 12759 3896 13820 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15620 3896 15669 3924
rect 15620 3884 15626 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 17681 3927 17739 3933
rect 17681 3893 17693 3927
rect 17727 3924 17739 3927
rect 18690 3924 18696 3936
rect 17727 3896 18696 3924
rect 17727 3893 17739 3896
rect 17681 3887 17739 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 20346 3884 20352 3936
rect 20404 3884 20410 3936
rect 25593 3927 25651 3933
rect 25593 3893 25605 3927
rect 25639 3924 25651 3927
rect 26602 3924 26608 3936
rect 25639 3896 26608 3924
rect 25639 3893 25651 3896
rect 25593 3887 25651 3893
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 26694 3884 26700 3936
rect 26752 3924 26758 3936
rect 36722 3924 36728 3936
rect 26752 3896 36728 3924
rect 26752 3884 26758 3896
rect 36722 3884 36728 3896
rect 36780 3884 36786 3936
rect 1104 3834 36524 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 36524 3834
rect 1104 3760 36524 3782
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12308 3692 14780 3720
rect 12308 3680 12314 3692
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 12250 3584 12256 3596
rect 11195 3556 12256 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 13173 3587 13231 3593
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 13630 3584 13636 3596
rect 13219 3556 13636 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 13630 3544 13636 3556
rect 13688 3584 13694 3596
rect 13817 3587 13875 3593
rect 13817 3584 13829 3587
rect 13688 3556 13829 3584
rect 13688 3544 13694 3556
rect 13817 3553 13829 3556
rect 13863 3553 13875 3587
rect 13817 3547 13875 3553
rect 14550 3544 14556 3596
rect 14608 3544 14614 3596
rect 14752 3593 14780 3692
rect 16942 3680 16948 3732
rect 17000 3680 17006 3732
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 17773 3723 17831 3729
rect 17773 3720 17785 3723
rect 17736 3692 17785 3720
rect 17736 3680 17742 3692
rect 17773 3689 17785 3692
rect 17819 3689 17831 3723
rect 17773 3683 17831 3689
rect 26145 3723 26203 3729
rect 26145 3689 26157 3723
rect 26191 3720 26203 3723
rect 26326 3720 26332 3732
rect 26191 3692 26332 3720
rect 26191 3689 26203 3692
rect 26145 3683 26203 3689
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 27338 3680 27344 3732
rect 27396 3720 27402 3732
rect 35989 3723 36047 3729
rect 35989 3720 36001 3723
rect 27396 3692 36001 3720
rect 27396 3680 27402 3692
rect 35989 3689 36001 3692
rect 36035 3720 36047 3723
rect 36078 3720 36084 3732
rect 36035 3692 36084 3720
rect 36035 3689 36047 3692
rect 35989 3683 36047 3689
rect 36078 3680 36084 3692
rect 36136 3680 36142 3732
rect 17586 3612 17592 3664
rect 17644 3652 17650 3664
rect 20346 3652 20352 3664
rect 17644 3624 17816 3652
rect 17644 3612 17650 3624
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3516 11115 3519
rect 11238 3516 11244 3528
rect 11103 3488 11244 3516
rect 11103 3485 11115 3488
rect 11057 3479 11115 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 12802 3476 12808 3528
rect 12860 3516 12866 3528
rect 13078 3516 13084 3528
rect 12860 3488 13084 3516
rect 12860 3476 12866 3488
rect 13078 3476 13084 3488
rect 13136 3516 13142 3528
rect 13722 3516 13728 3528
rect 13136 3488 13728 3516
rect 13136 3476 13142 3488
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 11698 3408 11704 3460
rect 11756 3408 11762 3460
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 13004 3420 13277 3448
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10597 3383 10655 3389
rect 10597 3380 10609 3383
rect 9916 3352 10609 3380
rect 9916 3340 9922 3352
rect 10597 3349 10609 3352
rect 10643 3349 10655 3383
rect 10597 3343 10655 3349
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 13004 3380 13032 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 13265 3411 13323 3417
rect 14461 3451 14519 3457
rect 14461 3417 14473 3451
rect 14507 3448 14519 3451
rect 14642 3448 14648 3460
rect 14507 3420 14648 3448
rect 14507 3417 14519 3420
rect 14461 3411 14519 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 14752 3448 14780 3547
rect 15194 3544 15200 3596
rect 15252 3584 15258 3596
rect 15470 3584 15476 3596
rect 15252 3556 15476 3584
rect 15252 3544 15258 3556
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17589 3519 17647 3525
rect 17589 3516 17601 3519
rect 16816 3488 17601 3516
rect 16816 3476 16822 3488
rect 17589 3485 17601 3488
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 15378 3448 15384 3460
rect 14752 3420 15384 3448
rect 15378 3408 15384 3420
rect 15436 3408 15442 3460
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 15562 3448 15568 3460
rect 15519 3420 15568 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 15562 3408 15568 3420
rect 15620 3408 15626 3460
rect 16114 3408 16120 3460
rect 16172 3408 16178 3460
rect 17788 3457 17816 3624
rect 17972 3624 20352 3652
rect 17972 3525 18000 3624
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 23934 3612 23940 3664
rect 23992 3652 23998 3664
rect 26694 3652 26700 3664
rect 23992 3624 24532 3652
rect 23992 3612 23998 3624
rect 18598 3544 18604 3596
rect 18656 3584 18662 3596
rect 18656 3556 19656 3584
rect 18656 3544 18662 3556
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3485 18015 3519
rect 17957 3479 18015 3485
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3516 18107 3519
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 18095 3488 18153 3516
rect 18095 3485 18107 3488
rect 18049 3479 18107 3485
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18693 3519 18751 3525
rect 18693 3516 18705 3519
rect 18472 3488 18705 3516
rect 18472 3476 18478 3488
rect 18693 3485 18705 3488
rect 18739 3485 18751 3519
rect 18693 3479 18751 3485
rect 18782 3476 18788 3528
rect 18840 3516 18846 3528
rect 18877 3519 18935 3525
rect 18877 3516 18889 3519
rect 18840 3488 18889 3516
rect 18840 3476 18846 3488
rect 18877 3485 18889 3488
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 19150 3476 19156 3528
rect 19208 3516 19214 3528
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 19208 3488 19257 3516
rect 19208 3476 19214 3488
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3516 19487 3519
rect 19518 3516 19524 3528
rect 19475 3488 19524 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 19628 3525 19656 3556
rect 23290 3544 23296 3596
rect 23348 3584 23354 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 23348 3556 24409 3584
rect 23348 3544 23354 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 24504 3584 24532 3624
rect 25700 3624 26700 3652
rect 24673 3587 24731 3593
rect 24673 3584 24685 3587
rect 24504 3556 24685 3584
rect 24397 3547 24455 3553
rect 24673 3553 24685 3556
rect 24719 3584 24731 3587
rect 25700 3584 25728 3624
rect 26694 3612 26700 3624
rect 26752 3612 26758 3664
rect 24719 3556 25728 3584
rect 24719 3553 24731 3556
rect 24673 3547 24731 3553
rect 26602 3544 26608 3596
rect 26660 3584 26666 3596
rect 26789 3587 26847 3593
rect 26789 3584 26801 3587
rect 26660 3556 26801 3584
rect 26660 3544 26666 3556
rect 26789 3553 26801 3556
rect 26835 3553 26847 3587
rect 26789 3547 26847 3553
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 27338 3476 27344 3528
rect 27396 3476 27402 3528
rect 17773 3451 17831 3457
rect 17773 3417 17785 3451
rect 17819 3417 17831 3451
rect 18969 3451 19027 3457
rect 18969 3448 18981 3451
rect 17773 3411 17831 3417
rect 17880 3420 18981 3448
rect 12768 3352 13032 3380
rect 12768 3340 12774 3352
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13504 3352 14105 3380
rect 13504 3340 13510 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 17034 3340 17040 3392
rect 17092 3340 17098 3392
rect 17126 3340 17132 3392
rect 17184 3380 17190 3392
rect 17880 3380 17908 3420
rect 18969 3417 18981 3420
rect 19015 3417 19027 3451
rect 18969 3411 19027 3417
rect 24026 3408 24032 3460
rect 24084 3448 24090 3460
rect 25130 3448 25136 3460
rect 24084 3420 25136 3448
rect 24084 3408 24090 3420
rect 17184 3352 17908 3380
rect 17184 3340 17190 3352
rect 18138 3340 18144 3392
rect 18196 3380 18202 3392
rect 19705 3383 19763 3389
rect 19705 3380 19717 3383
rect 18196 3352 19717 3380
rect 18196 3340 18202 3352
rect 19705 3349 19717 3352
rect 19751 3349 19763 3383
rect 25056 3380 25084 3420
rect 25130 3408 25136 3420
rect 25188 3408 25194 3460
rect 26973 3451 27031 3457
rect 26973 3448 26985 3451
rect 25976 3420 26985 3448
rect 25976 3380 26004 3420
rect 26973 3417 26985 3420
rect 27019 3417 27031 3451
rect 26973 3411 27031 3417
rect 36078 3408 36084 3460
rect 36136 3408 36142 3460
rect 25056 3352 26004 3380
rect 19705 3343 19763 3349
rect 26234 3340 26240 3392
rect 26292 3340 26298 3392
rect 1104 3290 36524 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 36524 3290
rect 1104 3216 36524 3238
rect 11422 3176 11428 3188
rect 9600 3148 11428 3176
rect 9600 3049 9628 3148
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11756 3148 11897 3176
rect 11756 3136 11762 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12710 3176 12716 3188
rect 12299 3148 12716 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 12912 3148 14780 3176
rect 9858 3068 9864 3120
rect 9916 3068 9922 3120
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 10980 2904 11008 3026
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12912 3049 12940 3148
rect 13173 3111 13231 3117
rect 13173 3077 13185 3111
rect 13219 3108 13231 3111
rect 13446 3108 13452 3120
rect 13219 3080 13452 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 13722 3068 13728 3120
rect 13780 3068 13786 3120
rect 14752 3108 14780 3148
rect 15304 3148 16896 3176
rect 15304 3120 15332 3148
rect 15286 3108 15292 3120
rect 14752 3080 15292 3108
rect 14752 3049 14780 3080
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 12032 3012 12357 3040
rect 12032 3000 12038 3012
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 16114 3000 16120 3052
rect 16172 3000 16178 3052
rect 16868 3049 16896 3148
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 22094 3176 22100 3188
rect 17828 3148 22100 3176
rect 17828 3136 17834 3148
rect 17126 3068 17132 3120
rect 17184 3068 17190 3120
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 18230 3000 18236 3052
rect 18288 3000 18294 3052
rect 18708 3049 18736 3148
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 24397 3179 24455 3185
rect 24084 3148 24164 3176
rect 24084 3136 24090 3148
rect 19426 3068 19432 3120
rect 19484 3068 19490 3120
rect 23290 3068 23296 3120
rect 23348 3108 23354 3120
rect 24136 3108 24164 3148
rect 24397 3145 24409 3179
rect 24443 3176 24455 3179
rect 24854 3176 24860 3188
rect 24443 3148 24860 3176
rect 24443 3145 24455 3148
rect 24397 3139 24455 3145
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 25869 3111 25927 3117
rect 23348 3080 24072 3108
rect 24136 3080 24702 3108
rect 23348 3068 23354 3080
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 23934 3000 23940 3052
rect 23992 3000 23998 3052
rect 24044 3049 24072 3080
rect 25869 3077 25881 3111
rect 25915 3108 25927 3111
rect 26234 3108 26240 3120
rect 25915 3080 26240 3108
rect 25915 3077 25927 3080
rect 25869 3071 25927 3077
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 26418 3040 26424 3052
rect 26191 3012 26424 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 26418 3000 26424 3012
rect 26476 3000 26482 3052
rect 11330 2932 11336 2984
rect 11388 2932 11394 2984
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12308 2944 12449 2972
rect 12308 2932 12314 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2972 15071 2975
rect 15059 2944 16068 2972
rect 15059 2941 15071 2944
rect 15013 2935 15071 2941
rect 12802 2904 12808 2916
rect 10980 2876 12808 2904
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 14645 2839 14703 2845
rect 14645 2805 14657 2839
rect 14691 2836 14703 2839
rect 15194 2836 15200 2848
rect 14691 2808 15200 2836
rect 14691 2805 14703 2808
rect 14645 2799 14703 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 16040 2836 16068 2944
rect 16132 2904 16160 3000
rect 16485 2975 16543 2981
rect 16485 2941 16497 2975
rect 16531 2972 16543 2975
rect 16758 2972 16764 2984
rect 16531 2944 16764 2972
rect 16531 2941 16543 2944
rect 16485 2935 16543 2941
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 18248 2972 18276 3000
rect 16868 2944 18276 2972
rect 16868 2904 16896 2944
rect 18966 2932 18972 2984
rect 19024 2932 19030 2984
rect 20438 2932 20444 2984
rect 20496 2932 20502 2984
rect 16132 2876 16896 2904
rect 18138 2836 18144 2848
rect 16040 2808 18144 2836
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 18601 2839 18659 2845
rect 18601 2805 18613 2839
rect 18647 2836 18659 2839
rect 19702 2836 19708 2848
rect 18647 2808 19708 2836
rect 18647 2805 18659 2808
rect 18601 2799 18659 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 23753 2839 23811 2845
rect 23753 2805 23765 2839
rect 23799 2836 23811 2839
rect 23842 2836 23848 2848
rect 23799 2808 23848 2836
rect 23799 2805 23811 2808
rect 23753 2799 23811 2805
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 1104 2746 36524 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 36524 2746
rect 1104 2672 36524 2694
rect 14642 2592 14648 2644
rect 14700 2592 14706 2644
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 17552 2604 18705 2632
rect 17552 2592 17558 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19245 2635 19303 2641
rect 19245 2632 19257 2635
rect 19024 2604 19257 2632
rect 19024 2592 19030 2604
rect 19245 2601 19257 2604
rect 19291 2601 19303 2635
rect 19245 2595 19303 2601
rect 18414 2524 18420 2576
rect 18472 2524 18478 2576
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11388 2468 12388 2496
rect 11388 2456 11394 2468
rect 11882 2388 11888 2440
rect 11940 2428 11946 2440
rect 12360 2437 12388 2468
rect 15194 2456 15200 2508
rect 15252 2456 15258 2508
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 16669 2499 16727 2505
rect 16669 2496 16681 2499
rect 15528 2468 16681 2496
rect 15528 2456 15534 2468
rect 16669 2465 16681 2468
rect 16715 2465 16727 2499
rect 16669 2459 16727 2465
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17034 2496 17040 2508
rect 16991 2468 17040 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 19702 2456 19708 2508
rect 19760 2496 19766 2508
rect 19797 2499 19855 2505
rect 19797 2496 19809 2499
rect 19760 2468 19809 2496
rect 19760 2456 19766 2468
rect 19797 2465 19809 2468
rect 19843 2465 19855 2499
rect 19797 2459 19855 2465
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11940 2400 11989 2428
rect 11940 2388 11946 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12986 2388 12992 2440
rect 13044 2388 13050 2440
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13872 2400 14289 2428
rect 13872 2388 13878 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 15212 2428 15240 2456
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 15212 2400 15577 2428
rect 14277 2391 14335 2397
rect 15565 2397 15577 2400
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 16206 2388 16212 2440
rect 16264 2388 16270 2440
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24673 2431 24731 2437
rect 24673 2428 24685 2431
rect 24544 2400 24685 2428
rect 24544 2388 24550 2400
rect 24673 2397 24685 2400
rect 24719 2397 24731 2431
rect 24673 2391 24731 2397
rect 24857 2431 24915 2437
rect 24857 2397 24869 2431
rect 24903 2428 24915 2431
rect 24946 2428 24952 2440
rect 24903 2400 24952 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 24946 2388 24952 2400
rect 25004 2388 25010 2440
rect 25225 2431 25283 2437
rect 25225 2397 25237 2431
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 18230 2360 18236 2372
rect 18170 2332 18236 2360
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 25240 2360 25268 2391
rect 24811 2332 25268 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12529 2295 12587 2301
rect 12529 2292 12541 2295
rect 12308 2264 12541 2292
rect 12308 2252 12314 2264
rect 12529 2261 12541 2264
rect 12575 2261 12587 2295
rect 12529 2255 12587 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 13596 2264 13829 2292
rect 13596 2252 13602 2264
rect 13817 2261 13829 2264
rect 13863 2261 13875 2295
rect 13817 2255 13875 2261
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14461 2295 14519 2301
rect 14461 2292 14473 2295
rect 14240 2264 14473 2292
rect 14240 2252 14246 2264
rect 14461 2261 14473 2264
rect 14507 2261 14519 2295
rect 14461 2255 14519 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15528 2264 15761 2292
rect 15528 2252 15534 2264
rect 15749 2261 15761 2264
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16393 2295 16451 2301
rect 16393 2292 16405 2295
rect 16172 2264 16405 2292
rect 16172 2252 16178 2264
rect 16393 2261 16405 2264
rect 16439 2261 16451 2295
rect 16393 2255 16451 2261
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25409 2295 25467 2301
rect 25409 2292 25421 2295
rect 25188 2264 25421 2292
rect 25188 2252 25194 2264
rect 25409 2261 25421 2264
rect 25455 2261 25467 2295
rect 25409 2255 25467 2261
rect 1104 2202 36524 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 36524 2202
rect 1104 2128 36524 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 7564 37272 7616 37324
rect 9588 37272 9640 37324
rect 22284 37340 22336 37392
rect 17224 37315 17276 37324
rect 17224 37281 17233 37315
rect 17233 37281 17267 37315
rect 17267 37281 17276 37315
rect 17224 37272 17276 37281
rect 18144 37272 18196 37324
rect 5816 37204 5868 37256
rect 8392 37204 8444 37256
rect 8300 37136 8352 37188
rect 4436 37068 4488 37120
rect 7472 37111 7524 37120
rect 7472 37077 7481 37111
rect 7481 37077 7515 37111
rect 7515 37077 7524 37111
rect 7472 37068 7524 37077
rect 10968 37204 11020 37256
rect 11612 37204 11664 37256
rect 12256 37204 12308 37256
rect 17040 37204 17092 37256
rect 10784 37136 10836 37188
rect 9036 37068 9088 37120
rect 10048 37068 10100 37120
rect 10600 37111 10652 37120
rect 10600 37077 10609 37111
rect 10609 37077 10643 37111
rect 10643 37077 10652 37111
rect 10600 37068 10652 37077
rect 10876 37068 10928 37120
rect 11888 37068 11940 37120
rect 12348 37068 12400 37120
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 4436 36839 4488 36848
rect 4436 36805 4445 36839
rect 4445 36805 4479 36839
rect 4479 36805 4488 36839
rect 4436 36796 4488 36805
rect 7380 36796 7432 36848
rect 9680 36864 9732 36916
rect 5816 36728 5868 36780
rect 8024 36728 8076 36780
rect 10968 36796 11020 36848
rect 11888 36839 11940 36848
rect 11888 36805 11897 36839
rect 11897 36805 11931 36839
rect 11931 36805 11940 36839
rect 11888 36796 11940 36805
rect 12164 36796 12216 36848
rect 13820 36864 13872 36916
rect 14740 36796 14792 36848
rect 16948 36796 17000 36848
rect 17408 36771 17460 36780
rect 17408 36737 17417 36771
rect 17417 36737 17451 36771
rect 17451 36737 17460 36771
rect 17408 36728 17460 36737
rect 18144 36771 18196 36780
rect 18144 36737 18153 36771
rect 18153 36737 18187 36771
rect 18187 36737 18196 36771
rect 18144 36728 18196 36737
rect 19892 36796 19944 36848
rect 20168 36796 20220 36848
rect 20352 36796 20404 36848
rect 26608 36864 26660 36916
rect 19524 36728 19576 36780
rect 5540 36524 5592 36576
rect 6460 36524 6512 36576
rect 6920 36703 6972 36712
rect 6920 36669 6929 36703
rect 6929 36669 6963 36703
rect 6963 36669 6972 36703
rect 6920 36660 6972 36669
rect 8760 36703 8812 36712
rect 8760 36669 8769 36703
rect 8769 36669 8803 36703
rect 8803 36669 8812 36703
rect 8760 36660 8812 36669
rect 9036 36703 9088 36712
rect 9036 36669 9045 36703
rect 9045 36669 9079 36703
rect 9079 36669 9088 36703
rect 9036 36660 9088 36669
rect 10692 36660 10744 36712
rect 8300 36524 8352 36576
rect 9220 36524 9272 36576
rect 12256 36660 12308 36712
rect 14280 36703 14332 36712
rect 14280 36669 14289 36703
rect 14289 36669 14323 36703
rect 14323 36669 14332 36703
rect 14280 36660 14332 36669
rect 15016 36660 15068 36712
rect 17040 36660 17092 36712
rect 17500 36703 17552 36712
rect 17500 36669 17509 36703
rect 17509 36669 17543 36703
rect 17543 36669 17552 36703
rect 17500 36660 17552 36669
rect 18236 36703 18288 36712
rect 18236 36669 18245 36703
rect 18245 36669 18279 36703
rect 18279 36669 18288 36703
rect 18236 36660 18288 36669
rect 19340 36660 19392 36712
rect 14004 36524 14056 36576
rect 14648 36524 14700 36576
rect 16580 36524 16632 36576
rect 19984 36660 20036 36712
rect 20260 36660 20312 36712
rect 23204 36660 23256 36712
rect 24584 36660 24636 36712
rect 24952 36703 25004 36712
rect 24952 36669 24961 36703
rect 24961 36669 24995 36703
rect 24995 36669 25004 36703
rect 24952 36660 25004 36669
rect 25228 36703 25280 36712
rect 25228 36669 25237 36703
rect 25237 36669 25271 36703
rect 25271 36669 25280 36703
rect 25228 36660 25280 36669
rect 23112 36524 23164 36576
rect 25964 36524 26016 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 6920 36320 6972 36372
rect 8760 36252 8812 36304
rect 6460 36227 6512 36236
rect 6460 36193 6469 36227
rect 6469 36193 6503 36227
rect 6503 36193 6512 36227
rect 6460 36184 6512 36193
rect 7472 36184 7524 36236
rect 8392 36184 8444 36236
rect 9588 36227 9640 36236
rect 9588 36193 9597 36227
rect 9597 36193 9631 36227
rect 9631 36193 9640 36227
rect 9588 36184 9640 36193
rect 9680 36116 9732 36168
rect 11704 36252 11756 36304
rect 10600 36227 10652 36236
rect 10600 36193 10609 36227
rect 10609 36193 10643 36227
rect 10643 36193 10652 36227
rect 10600 36184 10652 36193
rect 13452 36320 13504 36372
rect 14740 36320 14792 36372
rect 13268 36252 13320 36304
rect 14004 36252 14056 36304
rect 8024 36048 8076 36100
rect 9772 36048 9824 36100
rect 12164 36116 12216 36168
rect 12624 36116 12676 36168
rect 14648 36159 14700 36168
rect 14648 36125 14657 36159
rect 14657 36125 14691 36159
rect 14691 36125 14700 36159
rect 14648 36116 14700 36125
rect 14740 36159 14792 36168
rect 14740 36125 14749 36159
rect 14749 36125 14783 36159
rect 14783 36125 14792 36159
rect 14740 36116 14792 36125
rect 14924 36227 14976 36236
rect 14924 36193 14933 36227
rect 14933 36193 14967 36227
rect 14967 36193 14976 36227
rect 14924 36184 14976 36193
rect 15016 36159 15068 36168
rect 15016 36125 15025 36159
rect 15025 36125 15059 36159
rect 15059 36125 15068 36159
rect 15016 36116 15068 36125
rect 17500 36320 17552 36372
rect 19984 36363 20036 36372
rect 19984 36329 19993 36363
rect 19993 36329 20027 36363
rect 20027 36329 20036 36363
rect 19984 36320 20036 36329
rect 18236 36252 18288 36304
rect 19616 36227 19668 36236
rect 19616 36193 19625 36227
rect 19625 36193 19659 36227
rect 19659 36193 19668 36227
rect 19616 36184 19668 36193
rect 16488 36116 16540 36168
rect 17040 36116 17092 36168
rect 17316 36159 17368 36168
rect 17316 36125 17325 36159
rect 17325 36125 17359 36159
rect 17359 36125 17368 36159
rect 17316 36116 17368 36125
rect 18144 36116 18196 36168
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 19340 36159 19392 36168
rect 19340 36125 19349 36159
rect 19349 36125 19383 36159
rect 19383 36125 19392 36159
rect 19340 36116 19392 36125
rect 19708 36116 19760 36168
rect 19892 36159 19944 36168
rect 19892 36125 19901 36159
rect 19901 36125 19935 36159
rect 19935 36125 19944 36159
rect 19892 36116 19944 36125
rect 10600 36048 10652 36100
rect 7380 35980 7432 36032
rect 15292 36048 15344 36100
rect 15384 36091 15436 36100
rect 15384 36057 15393 36091
rect 15393 36057 15427 36091
rect 15427 36057 15436 36091
rect 15384 36048 15436 36057
rect 16764 36048 16816 36100
rect 20996 36184 21048 36236
rect 23112 36184 23164 36236
rect 24952 36184 25004 36236
rect 25228 36320 25280 36372
rect 25688 36227 25740 36236
rect 25688 36193 25697 36227
rect 25697 36193 25731 36227
rect 25731 36193 25740 36227
rect 25688 36184 25740 36193
rect 25964 36184 26016 36236
rect 20352 36116 20404 36168
rect 23112 36091 23164 36100
rect 23112 36057 23121 36091
rect 23121 36057 23155 36091
rect 23155 36057 23164 36091
rect 23112 36048 23164 36057
rect 24216 36159 24268 36168
rect 24216 36125 24225 36159
rect 24225 36125 24259 36159
rect 24259 36125 24268 36159
rect 24584 36159 24636 36168
rect 24216 36116 24268 36125
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 25504 36116 25556 36168
rect 24124 36048 24176 36100
rect 26240 36159 26292 36168
rect 26240 36125 26249 36159
rect 26249 36125 26283 36159
rect 26283 36125 26292 36159
rect 26240 36116 26292 36125
rect 26332 36159 26384 36168
rect 26332 36125 26341 36159
rect 26341 36125 26375 36159
rect 26375 36125 26384 36159
rect 26332 36116 26384 36125
rect 14372 35980 14424 36032
rect 16856 36023 16908 36032
rect 16856 35989 16865 36023
rect 16865 35989 16899 36023
rect 16899 35989 16908 36023
rect 16856 35980 16908 35989
rect 19892 35980 19944 36032
rect 20444 36023 20496 36032
rect 20444 35989 20453 36023
rect 20453 35989 20487 36023
rect 20487 35989 20496 36023
rect 20444 35980 20496 35989
rect 22100 35980 22152 36032
rect 24676 35980 24728 36032
rect 24860 35980 24912 36032
rect 25320 35980 25372 36032
rect 26148 36023 26200 36032
rect 26148 35989 26157 36023
rect 26157 35989 26191 36023
rect 26191 35989 26200 36023
rect 26148 35980 26200 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 7380 35776 7432 35828
rect 12900 35776 12952 35828
rect 7932 35708 7984 35760
rect 13176 35776 13228 35828
rect 13636 35751 13688 35760
rect 13636 35717 13645 35751
rect 13645 35717 13679 35751
rect 13679 35717 13688 35751
rect 13636 35708 13688 35717
rect 9220 35683 9272 35692
rect 9220 35649 9229 35683
rect 9229 35649 9263 35683
rect 9263 35649 9272 35683
rect 9220 35640 9272 35649
rect 9496 35640 9548 35692
rect 9772 35640 9824 35692
rect 12164 35640 12216 35692
rect 12532 35640 12584 35692
rect 5540 35572 5592 35624
rect 7012 35572 7064 35624
rect 7104 35572 7156 35624
rect 9312 35615 9364 35624
rect 9312 35581 9321 35615
rect 9321 35581 9355 35615
rect 9355 35581 9364 35615
rect 9312 35572 9364 35581
rect 9956 35615 10008 35624
rect 9956 35581 9965 35615
rect 9965 35581 9999 35615
rect 9999 35581 10008 35615
rect 9956 35572 10008 35581
rect 12256 35572 12308 35624
rect 12992 35640 13044 35692
rect 15384 35776 15436 35828
rect 18052 35776 18104 35828
rect 19248 35776 19300 35828
rect 20444 35776 20496 35828
rect 23112 35776 23164 35828
rect 23204 35819 23256 35828
rect 23204 35785 23213 35819
rect 23213 35785 23247 35819
rect 23247 35785 23256 35819
rect 23204 35776 23256 35785
rect 14556 35708 14608 35760
rect 14924 35708 14976 35760
rect 16764 35708 16816 35760
rect 18236 35708 18288 35760
rect 20720 35708 20772 35760
rect 21640 35708 21692 35760
rect 10232 35547 10284 35556
rect 10232 35513 10241 35547
rect 10241 35513 10275 35547
rect 10275 35513 10284 35547
rect 10232 35504 10284 35513
rect 13728 35572 13780 35624
rect 14740 35640 14792 35692
rect 15200 35683 15252 35692
rect 15200 35649 15209 35683
rect 15209 35649 15243 35683
rect 15243 35649 15252 35683
rect 15200 35640 15252 35649
rect 15292 35640 15344 35692
rect 15936 35640 15988 35692
rect 14188 35615 14240 35624
rect 14188 35581 14197 35615
rect 14197 35581 14231 35615
rect 14231 35581 14240 35615
rect 14188 35572 14240 35581
rect 13452 35504 13504 35556
rect 15660 35572 15712 35624
rect 16856 35640 16908 35692
rect 17040 35683 17092 35692
rect 17040 35649 17049 35683
rect 17049 35649 17083 35683
rect 17083 35649 17092 35683
rect 17040 35640 17092 35649
rect 17224 35640 17276 35692
rect 17776 35640 17828 35692
rect 17868 35683 17920 35692
rect 17868 35649 17877 35683
rect 17877 35649 17911 35683
rect 17911 35649 17920 35683
rect 17868 35640 17920 35649
rect 19340 35640 19392 35692
rect 19616 35640 19668 35692
rect 20076 35640 20128 35692
rect 19708 35572 19760 35624
rect 20628 35615 20680 35624
rect 20628 35581 20637 35615
rect 20637 35581 20671 35615
rect 20671 35581 20680 35615
rect 20628 35572 20680 35581
rect 16580 35504 16632 35556
rect 21456 35640 21508 35692
rect 12808 35436 12860 35488
rect 14188 35436 14240 35488
rect 16856 35479 16908 35488
rect 16856 35445 16865 35479
rect 16865 35445 16899 35479
rect 16899 35445 16908 35479
rect 16856 35436 16908 35445
rect 17224 35436 17276 35488
rect 18328 35436 18380 35488
rect 19892 35436 19944 35488
rect 21364 35572 21416 35624
rect 22192 35683 22244 35692
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 22468 35640 22520 35692
rect 22560 35683 22612 35692
rect 22560 35649 22569 35683
rect 22569 35649 22603 35683
rect 22603 35649 22612 35683
rect 22560 35640 22612 35649
rect 23664 35776 23716 35828
rect 24216 35776 24268 35828
rect 24768 35776 24820 35828
rect 26240 35776 26292 35828
rect 22928 35683 22980 35692
rect 22928 35649 22937 35683
rect 22937 35649 22971 35683
rect 22971 35649 22980 35683
rect 22928 35640 22980 35649
rect 23020 35683 23072 35692
rect 23020 35649 23034 35683
rect 23034 35649 23068 35683
rect 23068 35649 23072 35683
rect 23020 35640 23072 35649
rect 22652 35504 22704 35556
rect 23940 35683 23992 35692
rect 23940 35649 23949 35683
rect 23949 35649 23983 35683
rect 23983 35649 23992 35683
rect 23940 35640 23992 35649
rect 24124 35640 24176 35692
rect 24860 35708 24912 35760
rect 24676 35640 24728 35692
rect 25044 35683 25096 35692
rect 25044 35649 25053 35683
rect 25053 35649 25087 35683
rect 25087 35649 25096 35683
rect 25044 35640 25096 35649
rect 25136 35572 25188 35624
rect 25412 35640 25464 35692
rect 26332 35683 26384 35692
rect 26332 35649 26341 35683
rect 26341 35649 26375 35683
rect 26375 35649 26384 35683
rect 26332 35640 26384 35649
rect 22100 35436 22152 35488
rect 22192 35436 22244 35488
rect 24124 35504 24176 35556
rect 23112 35436 23164 35488
rect 26516 35504 26568 35556
rect 25596 35479 25648 35488
rect 25596 35445 25605 35479
rect 25605 35445 25639 35479
rect 25639 35445 25648 35479
rect 25596 35436 25648 35445
rect 26148 35436 26200 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 7012 35275 7064 35284
rect 7012 35241 7021 35275
rect 7021 35241 7055 35275
rect 7055 35241 7064 35275
rect 7012 35232 7064 35241
rect 9312 35275 9364 35284
rect 9312 35241 9321 35275
rect 9321 35241 9355 35275
rect 9355 35241 9364 35275
rect 9312 35232 9364 35241
rect 9956 35232 10008 35284
rect 12532 35232 12584 35284
rect 12716 35232 12768 35284
rect 12992 35232 13044 35284
rect 10048 35164 10100 35216
rect 5540 35096 5592 35148
rect 6552 35096 6604 35148
rect 7104 35096 7156 35148
rect 7564 35139 7616 35148
rect 7564 35105 7573 35139
rect 7573 35105 7607 35139
rect 7607 35105 7616 35139
rect 7564 35096 7616 35105
rect 11520 35096 11572 35148
rect 11612 35096 11664 35148
rect 12256 35096 12308 35148
rect 9220 35071 9272 35080
rect 9220 35037 9229 35071
rect 9229 35037 9263 35071
rect 9263 35037 9272 35071
rect 9220 35028 9272 35037
rect 9404 35071 9456 35080
rect 9404 35037 9413 35071
rect 9413 35037 9447 35071
rect 9447 35037 9456 35071
rect 9404 35028 9456 35037
rect 5448 34960 5500 35012
rect 7932 34960 7984 35012
rect 9956 35028 10008 35080
rect 10232 35028 10284 35080
rect 10048 34960 10100 35012
rect 12348 35028 12400 35080
rect 12624 35071 12676 35080
rect 12624 35037 12633 35071
rect 12633 35037 12667 35071
rect 12667 35037 12676 35071
rect 12624 35028 12676 35037
rect 12440 34960 12492 35012
rect 14188 35275 14240 35284
rect 14188 35241 14197 35275
rect 14197 35241 14231 35275
rect 14231 35241 14240 35275
rect 14188 35232 14240 35241
rect 14280 35232 14332 35284
rect 20076 35275 20128 35284
rect 20076 35241 20085 35275
rect 20085 35241 20119 35275
rect 20119 35241 20128 35275
rect 20076 35232 20128 35241
rect 22560 35232 22612 35284
rect 22652 35275 22704 35284
rect 22652 35241 22661 35275
rect 22661 35241 22695 35275
rect 22695 35241 22704 35275
rect 22652 35232 22704 35241
rect 23940 35232 23992 35284
rect 25044 35232 25096 35284
rect 25504 35275 25556 35284
rect 25504 35241 25513 35275
rect 25513 35241 25547 35275
rect 25547 35241 25556 35275
rect 25504 35232 25556 35241
rect 26516 35275 26568 35284
rect 26516 35241 26525 35275
rect 26525 35241 26559 35275
rect 26559 35241 26568 35275
rect 26516 35232 26568 35241
rect 14740 35164 14792 35216
rect 12992 35071 13044 35080
rect 12992 35037 13001 35071
rect 13001 35037 13035 35071
rect 13035 35037 13044 35071
rect 12992 35028 13044 35037
rect 13728 35096 13780 35148
rect 14004 35028 14056 35080
rect 14372 35071 14424 35080
rect 14372 35037 14381 35071
rect 14381 35037 14415 35071
rect 14415 35037 14424 35071
rect 14372 35028 14424 35037
rect 15936 35028 15988 35080
rect 17408 35096 17460 35148
rect 17316 35028 17368 35080
rect 17868 35071 17920 35080
rect 17868 35037 17877 35071
rect 17877 35037 17911 35071
rect 17911 35037 17920 35071
rect 17868 35028 17920 35037
rect 18144 35071 18196 35080
rect 18144 35037 18153 35071
rect 18153 35037 18187 35071
rect 18187 35037 18196 35071
rect 18144 35028 18196 35037
rect 19892 35139 19944 35148
rect 19892 35105 19901 35139
rect 19901 35105 19935 35139
rect 19935 35105 19944 35139
rect 19892 35096 19944 35105
rect 21456 35164 21508 35216
rect 18328 35071 18380 35080
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 18512 35071 18564 35080
rect 18512 35037 18521 35071
rect 18521 35037 18555 35071
rect 18555 35037 18564 35071
rect 18512 35028 18564 35037
rect 18604 35071 18656 35080
rect 18604 35037 18613 35071
rect 18613 35037 18647 35071
rect 18647 35037 18656 35071
rect 18604 35028 18656 35037
rect 19340 35028 19392 35080
rect 21916 35071 21968 35080
rect 21916 35037 21925 35071
rect 21925 35037 21959 35071
rect 21959 35037 21968 35071
rect 21916 35028 21968 35037
rect 22008 35028 22060 35080
rect 21364 34960 21416 35012
rect 21548 34960 21600 35012
rect 22192 34960 22244 35012
rect 23112 35071 23164 35080
rect 23112 35037 23121 35071
rect 23121 35037 23155 35071
rect 23155 35037 23164 35071
rect 23112 35028 23164 35037
rect 24768 35071 24820 35080
rect 24768 35037 24777 35071
rect 24777 35037 24811 35071
rect 24811 35037 24820 35071
rect 24768 35028 24820 35037
rect 24860 35071 24912 35080
rect 24860 35037 24869 35071
rect 24869 35037 24903 35071
rect 24903 35037 24912 35071
rect 24860 35028 24912 35037
rect 26148 35164 26200 35216
rect 11704 34935 11756 34944
rect 11704 34901 11713 34935
rect 11713 34901 11747 34935
rect 11747 34901 11756 34935
rect 11704 34892 11756 34901
rect 11796 34892 11848 34944
rect 12716 34892 12768 34944
rect 12900 34892 12952 34944
rect 20628 34892 20680 34944
rect 20720 34892 20772 34944
rect 23848 34892 23900 34944
rect 25596 35139 25648 35148
rect 25596 35105 25605 35139
rect 25605 35105 25639 35139
rect 25639 35105 25648 35139
rect 25596 35096 25648 35105
rect 26240 35028 26292 35080
rect 26792 35139 26844 35148
rect 26792 35105 26801 35139
rect 26801 35105 26835 35139
rect 26835 35105 26844 35139
rect 26792 35096 26844 35105
rect 25872 35003 25924 35012
rect 25872 34969 25881 35003
rect 25881 34969 25915 35003
rect 25915 34969 25924 35003
rect 25872 34960 25924 34969
rect 26240 34935 26292 34944
rect 26240 34901 26249 34935
rect 26249 34901 26283 34935
rect 26283 34901 26292 34935
rect 26240 34892 26292 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 5448 34688 5500 34740
rect 6552 34688 6604 34740
rect 9220 34688 9272 34740
rect 11520 34731 11572 34740
rect 11520 34697 11529 34731
rect 11529 34697 11563 34731
rect 11563 34697 11572 34731
rect 11520 34688 11572 34697
rect 8300 34595 8352 34604
rect 8300 34561 8309 34595
rect 8309 34561 8343 34595
rect 8343 34561 8352 34595
rect 8300 34552 8352 34561
rect 9404 34620 9456 34672
rect 11704 34620 11756 34672
rect 12900 34688 12952 34740
rect 12992 34731 13044 34740
rect 12992 34697 13001 34731
rect 13001 34697 13035 34731
rect 13035 34697 13044 34731
rect 12992 34688 13044 34697
rect 14464 34688 14516 34740
rect 16856 34688 16908 34740
rect 12716 34620 12768 34672
rect 9772 34552 9824 34604
rect 10232 34595 10284 34604
rect 10232 34561 10241 34595
rect 10241 34561 10275 34595
rect 10275 34561 10284 34595
rect 10232 34552 10284 34561
rect 7564 34484 7616 34536
rect 8668 34459 8720 34468
rect 8668 34425 8677 34459
rect 8677 34425 8711 34459
rect 8711 34425 8720 34459
rect 8668 34416 8720 34425
rect 9496 34484 9548 34536
rect 10508 34484 10560 34536
rect 10048 34416 10100 34468
rect 9956 34391 10008 34400
rect 9956 34357 9965 34391
rect 9965 34357 9999 34391
rect 9999 34357 10008 34391
rect 11796 34552 11848 34604
rect 11888 34595 11940 34604
rect 11888 34561 11897 34595
rect 11897 34561 11931 34595
rect 11931 34561 11940 34595
rect 11888 34552 11940 34561
rect 12348 34595 12400 34604
rect 12348 34561 12357 34595
rect 12357 34561 12391 34595
rect 12391 34561 12400 34595
rect 12348 34552 12400 34561
rect 12808 34595 12860 34604
rect 12808 34561 12817 34595
rect 12817 34561 12851 34595
rect 12851 34561 12860 34595
rect 12808 34552 12860 34561
rect 15016 34595 15068 34604
rect 15016 34561 15025 34595
rect 15025 34561 15059 34595
rect 15059 34561 15068 34595
rect 15016 34552 15068 34561
rect 11060 34484 11112 34536
rect 16764 34595 16816 34604
rect 16764 34561 16773 34595
rect 16773 34561 16807 34595
rect 16807 34561 16816 34595
rect 16764 34552 16816 34561
rect 17960 34620 18012 34672
rect 18604 34688 18656 34740
rect 18972 34688 19024 34740
rect 19248 34731 19300 34740
rect 19248 34697 19257 34731
rect 19257 34697 19291 34731
rect 19291 34697 19300 34731
rect 19248 34688 19300 34697
rect 19616 34688 19668 34740
rect 19984 34688 20036 34740
rect 22192 34688 22244 34740
rect 17224 34552 17276 34604
rect 21732 34620 21784 34672
rect 21916 34620 21968 34672
rect 25872 34688 25924 34740
rect 10876 34416 10928 34468
rect 12532 34416 12584 34468
rect 14832 34416 14884 34468
rect 17316 34484 17368 34536
rect 18144 34484 18196 34536
rect 18788 34552 18840 34604
rect 18972 34595 19024 34604
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 19064 34552 19116 34604
rect 21548 34552 21600 34604
rect 22192 34595 22244 34604
rect 22192 34561 22201 34595
rect 22201 34561 22235 34595
rect 22235 34561 22244 34595
rect 22192 34552 22244 34561
rect 22008 34484 22060 34536
rect 22468 34595 22520 34604
rect 22468 34561 22477 34595
rect 22477 34561 22511 34595
rect 22511 34561 22520 34595
rect 22468 34552 22520 34561
rect 22836 34552 22888 34604
rect 23204 34595 23256 34604
rect 23204 34561 23213 34595
rect 23213 34561 23247 34595
rect 23247 34561 23256 34595
rect 23204 34552 23256 34561
rect 23480 34595 23532 34604
rect 23480 34561 23489 34595
rect 23489 34561 23523 34595
rect 23523 34561 23532 34595
rect 23480 34552 23532 34561
rect 26332 34620 26384 34672
rect 25136 34484 25188 34536
rect 26240 34552 26292 34604
rect 9956 34348 10008 34357
rect 11888 34348 11940 34400
rect 12624 34348 12676 34400
rect 13360 34348 13412 34400
rect 15384 34391 15436 34400
rect 15384 34357 15393 34391
rect 15393 34357 15427 34391
rect 15427 34357 15436 34391
rect 15384 34348 15436 34357
rect 15476 34391 15528 34400
rect 15476 34357 15485 34391
rect 15485 34357 15519 34391
rect 15519 34357 15528 34391
rect 15476 34348 15528 34357
rect 18604 34459 18656 34468
rect 18604 34425 18613 34459
rect 18613 34425 18647 34459
rect 18647 34425 18656 34459
rect 18604 34416 18656 34425
rect 19156 34416 19208 34468
rect 25688 34459 25740 34468
rect 25688 34425 25697 34459
rect 25697 34425 25731 34459
rect 25731 34425 25740 34459
rect 25688 34416 25740 34425
rect 26792 34527 26844 34536
rect 26792 34493 26801 34527
rect 26801 34493 26835 34527
rect 26835 34493 26844 34527
rect 26792 34484 26844 34493
rect 27528 34416 27580 34468
rect 18420 34348 18472 34400
rect 23664 34391 23716 34400
rect 23664 34357 23673 34391
rect 23673 34357 23707 34391
rect 23707 34357 23716 34391
rect 23664 34348 23716 34357
rect 26056 34348 26108 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 10232 34144 10284 34196
rect 12440 34144 12492 34196
rect 5540 34008 5592 34060
rect 6368 34008 6420 34060
rect 8668 34008 8720 34060
rect 8944 34076 8996 34128
rect 10876 34076 10928 34128
rect 9496 34008 9548 34060
rect 8852 33940 8904 33992
rect 7012 33915 7064 33924
rect 7012 33881 7021 33915
rect 7021 33881 7055 33915
rect 7055 33881 7064 33915
rect 7012 33872 7064 33881
rect 10048 33940 10100 33992
rect 10140 33983 10192 33992
rect 10140 33949 10149 33983
rect 10149 33949 10183 33983
rect 10183 33949 10192 33983
rect 10140 33940 10192 33949
rect 10784 33940 10836 33992
rect 7932 33804 7984 33856
rect 9680 33847 9732 33856
rect 9680 33813 9689 33847
rect 9689 33813 9723 33847
rect 9723 33813 9732 33847
rect 9680 33804 9732 33813
rect 9772 33847 9824 33856
rect 9772 33813 9781 33847
rect 9781 33813 9815 33847
rect 9815 33813 9824 33847
rect 9772 33804 9824 33813
rect 10232 33804 10284 33856
rect 11612 33940 11664 33992
rect 11888 33983 11940 33992
rect 11888 33949 11897 33983
rect 11897 33949 11931 33983
rect 11931 33949 11940 33983
rect 11888 33940 11940 33949
rect 12072 33983 12124 33992
rect 12072 33949 12081 33983
rect 12081 33949 12115 33983
rect 12115 33949 12124 33983
rect 12072 33940 12124 33949
rect 14740 33940 14792 33992
rect 14924 33983 14976 33992
rect 14924 33949 14933 33983
rect 14933 33949 14967 33983
rect 14967 33949 14976 33983
rect 14924 33940 14976 33949
rect 15108 33940 15160 33992
rect 15200 33983 15252 33992
rect 15200 33949 15209 33983
rect 15209 33949 15243 33983
rect 15243 33949 15252 33983
rect 15200 33940 15252 33949
rect 17224 34144 17276 34196
rect 17960 34187 18012 34196
rect 17960 34153 17969 34187
rect 17969 34153 18003 34187
rect 18003 34153 18012 34187
rect 17960 34144 18012 34153
rect 18328 34144 18380 34196
rect 19064 34144 19116 34196
rect 19708 34144 19760 34196
rect 20812 34144 20864 34196
rect 23204 34144 23256 34196
rect 27528 34187 27580 34196
rect 27528 34153 27537 34187
rect 27537 34153 27571 34187
rect 27571 34153 27580 34187
rect 27528 34144 27580 34153
rect 18328 34008 18380 34060
rect 11336 33915 11388 33924
rect 11336 33881 11370 33915
rect 11370 33881 11388 33915
rect 11336 33872 11388 33881
rect 11980 33872 12032 33924
rect 12348 33872 12400 33924
rect 13360 33872 13412 33924
rect 11244 33847 11296 33856
rect 11244 33813 11253 33847
rect 11253 33813 11287 33847
rect 11287 33813 11296 33847
rect 11244 33804 11296 33813
rect 14556 33915 14608 33924
rect 14556 33881 14565 33915
rect 14565 33881 14599 33915
rect 14599 33881 14608 33915
rect 14556 33872 14608 33881
rect 15844 33872 15896 33924
rect 17592 33983 17644 33992
rect 17592 33949 17601 33983
rect 17601 33949 17635 33983
rect 17635 33949 17644 33983
rect 17592 33940 17644 33949
rect 17776 33983 17828 33992
rect 17776 33949 17785 33983
rect 17785 33949 17819 33983
rect 17819 33949 17828 33983
rect 17776 33940 17828 33949
rect 18420 33983 18472 33992
rect 18420 33949 18429 33983
rect 18429 33949 18463 33983
rect 18463 33949 18472 33983
rect 18420 33940 18472 33949
rect 18512 33983 18564 33992
rect 18512 33949 18522 33983
rect 18522 33949 18556 33983
rect 18556 33949 18564 33983
rect 19064 34008 19116 34060
rect 21180 34076 21232 34128
rect 21640 34119 21692 34128
rect 21640 34085 21649 34119
rect 21649 34085 21683 34119
rect 21683 34085 21692 34119
rect 21640 34076 21692 34085
rect 23020 34076 23072 34128
rect 22468 34008 22520 34060
rect 18512 33940 18564 33949
rect 16488 33872 16540 33924
rect 20812 33940 20864 33992
rect 21732 33940 21784 33992
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 22560 33940 22612 33992
rect 24952 34076 25004 34128
rect 26056 34051 26108 34060
rect 26056 34017 26065 34051
rect 26065 34017 26099 34051
rect 26099 34017 26108 34051
rect 26056 34008 26108 34017
rect 17500 33804 17552 33856
rect 19432 33872 19484 33924
rect 19800 33872 19852 33924
rect 20260 33872 20312 33924
rect 21548 33872 21600 33924
rect 24124 33915 24176 33924
rect 24124 33881 24133 33915
rect 24133 33881 24167 33915
rect 24167 33881 24176 33915
rect 24124 33872 24176 33881
rect 26608 33872 26660 33924
rect 19340 33804 19392 33856
rect 22192 33804 22244 33856
rect 23572 33804 23624 33856
rect 23848 33804 23900 33856
rect 24032 33847 24084 33856
rect 24032 33813 24041 33847
rect 24041 33813 24075 33847
rect 24075 33813 24084 33847
rect 24032 33804 24084 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 7012 33600 7064 33652
rect 9772 33600 9824 33652
rect 11060 33600 11112 33652
rect 12072 33600 12124 33652
rect 7932 33532 7984 33584
rect 9496 33532 9548 33584
rect 10876 33532 10928 33584
rect 6368 33507 6420 33516
rect 6368 33473 6377 33507
rect 6377 33473 6411 33507
rect 6411 33473 6420 33507
rect 6368 33464 6420 33473
rect 8484 33507 8536 33516
rect 8484 33473 8493 33507
rect 8493 33473 8527 33507
rect 8527 33473 8536 33507
rect 8484 33464 8536 33473
rect 8668 33507 8720 33516
rect 8668 33473 8677 33507
rect 8677 33473 8711 33507
rect 8711 33473 8720 33507
rect 8668 33464 8720 33473
rect 7012 33396 7064 33448
rect 7840 33396 7892 33448
rect 10232 33396 10284 33448
rect 11060 33507 11112 33516
rect 11060 33473 11069 33507
rect 11069 33473 11103 33507
rect 11103 33473 11112 33507
rect 11060 33464 11112 33473
rect 11152 33328 11204 33380
rect 10968 33260 11020 33312
rect 11336 33507 11388 33516
rect 11336 33473 11345 33507
rect 11345 33473 11379 33507
rect 11379 33473 11388 33507
rect 11336 33464 11388 33473
rect 11520 33575 11572 33584
rect 11520 33541 11529 33575
rect 11529 33541 11563 33575
rect 11563 33541 11572 33575
rect 11520 33532 11572 33541
rect 12624 33532 12676 33584
rect 13728 33532 13780 33584
rect 12348 33464 12400 33516
rect 14556 33464 14608 33516
rect 14832 33643 14884 33652
rect 14832 33609 14841 33643
rect 14841 33609 14875 33643
rect 14875 33609 14884 33643
rect 14832 33600 14884 33609
rect 15108 33643 15160 33652
rect 15108 33609 15117 33643
rect 15117 33609 15151 33643
rect 15151 33609 15160 33643
rect 15108 33600 15160 33609
rect 16764 33600 16816 33652
rect 17040 33600 17092 33652
rect 17776 33600 17828 33652
rect 18512 33600 18564 33652
rect 15384 33532 15436 33584
rect 18604 33532 18656 33584
rect 20904 33532 20956 33584
rect 16028 33464 16080 33516
rect 16948 33464 17000 33516
rect 14004 33439 14056 33448
rect 14004 33405 14013 33439
rect 14013 33405 14047 33439
rect 14047 33405 14056 33439
rect 14004 33396 14056 33405
rect 15200 33396 15252 33448
rect 15844 33396 15896 33448
rect 17592 33464 17644 33516
rect 21548 33532 21600 33584
rect 22008 33600 22060 33652
rect 23480 33600 23532 33652
rect 21916 33532 21968 33584
rect 11888 33328 11940 33380
rect 14648 33328 14700 33380
rect 15476 33328 15528 33380
rect 15568 33328 15620 33380
rect 16120 33328 16172 33380
rect 21732 33396 21784 33448
rect 22376 33464 22428 33516
rect 22652 33507 22704 33516
rect 22652 33473 22661 33507
rect 22661 33473 22695 33507
rect 22695 33473 22704 33507
rect 22652 33464 22704 33473
rect 22836 33507 22888 33516
rect 22836 33473 22845 33507
rect 22845 33473 22879 33507
rect 22879 33473 22888 33507
rect 22836 33464 22888 33473
rect 22744 33396 22796 33448
rect 23664 33532 23716 33584
rect 24676 33532 24728 33584
rect 25136 33532 25188 33584
rect 25688 33532 25740 33584
rect 23020 33464 23072 33516
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 25044 33464 25096 33473
rect 24400 33396 24452 33448
rect 25688 33396 25740 33448
rect 11796 33260 11848 33312
rect 14924 33260 14976 33312
rect 15660 33260 15712 33312
rect 18144 33260 18196 33312
rect 20904 33260 20956 33312
rect 21824 33328 21876 33380
rect 22192 33260 22244 33312
rect 22744 33260 22796 33312
rect 25044 33260 25096 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 7012 33099 7064 33108
rect 7012 33065 7021 33099
rect 7021 33065 7055 33099
rect 7055 33065 7064 33099
rect 7012 33056 7064 33065
rect 9680 33056 9732 33108
rect 10692 33056 10744 33108
rect 10876 33099 10928 33108
rect 10876 33065 10885 33099
rect 10885 33065 10919 33099
rect 10919 33065 10928 33099
rect 10876 33056 10928 33065
rect 11060 33056 11112 33108
rect 11244 33099 11296 33108
rect 11244 33065 11253 33099
rect 11253 33065 11287 33099
rect 11287 33065 11296 33099
rect 11244 33056 11296 33065
rect 14004 33056 14056 33108
rect 8300 32988 8352 33040
rect 8484 32988 8536 33040
rect 18328 33056 18380 33108
rect 7840 32852 7892 32904
rect 10876 32895 10928 32904
rect 10876 32861 10885 32895
rect 10885 32861 10919 32895
rect 10919 32861 10928 32895
rect 10876 32852 10928 32861
rect 12624 32920 12676 32972
rect 15016 32988 15068 33040
rect 11060 32784 11112 32836
rect 9128 32716 9180 32768
rect 14556 32895 14608 32904
rect 14556 32861 14565 32895
rect 14565 32861 14599 32895
rect 14599 32861 14608 32895
rect 14556 32852 14608 32861
rect 14832 32895 14884 32904
rect 14832 32861 14841 32895
rect 14841 32861 14875 32895
rect 14875 32861 14884 32895
rect 14832 32852 14884 32861
rect 15016 32852 15068 32904
rect 15568 32920 15620 32972
rect 15200 32784 15252 32836
rect 15384 32895 15436 32904
rect 15384 32861 15393 32895
rect 15393 32861 15427 32895
rect 15427 32861 15436 32895
rect 15384 32852 15436 32861
rect 15476 32895 15528 32904
rect 15476 32861 15485 32895
rect 15485 32861 15519 32895
rect 15519 32861 15528 32895
rect 15476 32852 15528 32861
rect 16580 32784 16632 32836
rect 14648 32716 14700 32768
rect 15108 32716 15160 32768
rect 15660 32716 15712 32768
rect 18512 32988 18564 33040
rect 17960 32920 18012 32972
rect 18788 33056 18840 33108
rect 21180 33056 21232 33108
rect 21732 33056 21784 33108
rect 22468 33099 22520 33108
rect 22468 33065 22477 33099
rect 22477 33065 22511 33099
rect 22511 33065 22520 33099
rect 22468 33056 22520 33065
rect 19432 32988 19484 33040
rect 18788 32920 18840 32972
rect 19156 32920 19208 32972
rect 17868 32895 17920 32904
rect 17868 32861 17877 32895
rect 17877 32861 17911 32895
rect 17911 32861 17920 32895
rect 17868 32852 17920 32861
rect 18052 32895 18104 32904
rect 18052 32861 18061 32895
rect 18061 32861 18095 32895
rect 18095 32861 18104 32895
rect 18052 32852 18104 32861
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 18144 32716 18196 32768
rect 18420 32895 18472 32904
rect 18420 32861 18429 32895
rect 18429 32861 18463 32895
rect 18463 32861 18472 32895
rect 18420 32852 18472 32861
rect 18972 32895 19024 32904
rect 18972 32861 18981 32895
rect 18981 32861 19015 32895
rect 19015 32861 19024 32895
rect 18972 32852 19024 32861
rect 22744 32920 22796 32972
rect 23572 32852 23624 32904
rect 18696 32827 18748 32836
rect 18696 32793 18705 32827
rect 18705 32793 18739 32827
rect 18739 32793 18748 32827
rect 18696 32784 18748 32793
rect 20536 32784 20588 32836
rect 24676 32920 24728 32972
rect 25136 32920 25188 32972
rect 30196 32920 30248 32972
rect 23848 32852 23900 32904
rect 28816 32852 28868 32904
rect 29920 32895 29972 32904
rect 29920 32861 29929 32895
rect 29929 32861 29963 32895
rect 29963 32861 29972 32895
rect 29920 32852 29972 32861
rect 18604 32759 18656 32768
rect 18604 32725 18613 32759
rect 18613 32725 18647 32759
rect 18647 32725 18656 32759
rect 18604 32716 18656 32725
rect 18880 32716 18932 32768
rect 20720 32716 20772 32768
rect 20812 32716 20864 32768
rect 24216 32827 24268 32836
rect 24216 32793 24225 32827
rect 24225 32793 24259 32827
rect 24259 32793 24268 32827
rect 24216 32784 24268 32793
rect 24308 32784 24360 32836
rect 25964 32784 26016 32836
rect 26608 32784 26660 32836
rect 27344 32827 27396 32836
rect 27344 32793 27353 32827
rect 27353 32793 27387 32827
rect 27387 32793 27396 32827
rect 27344 32784 27396 32793
rect 30840 32784 30892 32836
rect 21824 32716 21876 32768
rect 22560 32716 22612 32768
rect 24860 32716 24912 32768
rect 25504 32716 25556 32768
rect 28172 32716 28224 32768
rect 30012 32716 30064 32768
rect 30656 32716 30708 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 6552 32512 6604 32564
rect 8484 32512 8536 32564
rect 8852 32512 8904 32564
rect 2688 32444 2740 32496
rect 7288 32444 7340 32496
rect 7932 32444 7984 32496
rect 10324 32444 10376 32496
rect 11060 32555 11112 32564
rect 11060 32521 11069 32555
rect 11069 32521 11103 32555
rect 11103 32521 11112 32555
rect 11060 32512 11112 32521
rect 11796 32512 11848 32564
rect 14740 32512 14792 32564
rect 13820 32444 13872 32496
rect 14648 32444 14700 32496
rect 17316 32512 17368 32564
rect 18420 32512 18472 32564
rect 18696 32512 18748 32564
rect 20536 32555 20588 32564
rect 20536 32521 20545 32555
rect 20545 32521 20579 32555
rect 20579 32521 20588 32555
rect 20536 32512 20588 32521
rect 15384 32444 15436 32496
rect 4896 32419 4948 32428
rect 4896 32385 4905 32419
rect 4905 32385 4939 32419
rect 4939 32385 4948 32419
rect 4896 32376 4948 32385
rect 5356 32376 5408 32428
rect 8208 32376 8260 32428
rect 9404 32419 9456 32428
rect 9404 32385 9413 32419
rect 9413 32385 9447 32419
rect 9447 32385 9456 32419
rect 9404 32376 9456 32385
rect 9588 32419 9640 32428
rect 9588 32385 9597 32419
rect 9597 32385 9631 32419
rect 9631 32385 9640 32419
rect 9588 32376 9640 32385
rect 10140 32376 10192 32428
rect 11060 32376 11112 32428
rect 11244 32376 11296 32428
rect 11520 32419 11572 32428
rect 11520 32385 11529 32419
rect 11529 32385 11563 32419
rect 11563 32385 11572 32419
rect 11520 32376 11572 32385
rect 11704 32419 11756 32428
rect 11704 32385 11713 32419
rect 11713 32385 11747 32419
rect 11747 32385 11756 32419
rect 11704 32376 11756 32385
rect 13176 32376 13228 32428
rect 14740 32419 14792 32428
rect 14740 32385 14749 32419
rect 14749 32385 14783 32419
rect 14783 32385 14792 32419
rect 14740 32376 14792 32385
rect 15108 32419 15160 32428
rect 15108 32385 15117 32419
rect 15117 32385 15151 32419
rect 15151 32385 15160 32419
rect 15108 32376 15160 32385
rect 15200 32376 15252 32428
rect 15752 32444 15804 32496
rect 5540 32172 5592 32224
rect 7104 32308 7156 32360
rect 10324 32308 10376 32360
rect 9312 32283 9364 32292
rect 9312 32249 9321 32283
rect 9321 32249 9355 32283
rect 9355 32249 9364 32283
rect 9312 32240 9364 32249
rect 9680 32240 9732 32292
rect 11980 32308 12032 32360
rect 7196 32172 7248 32224
rect 10416 32172 10468 32224
rect 11336 32240 11388 32292
rect 12900 32351 12952 32360
rect 12900 32317 12909 32351
rect 12909 32317 12943 32351
rect 12943 32317 12952 32351
rect 12900 32308 12952 32317
rect 15844 32419 15896 32428
rect 15844 32385 15853 32419
rect 15853 32385 15887 32419
rect 15887 32385 15896 32419
rect 15844 32376 15896 32385
rect 16120 32419 16172 32428
rect 16120 32385 16129 32419
rect 16129 32385 16163 32419
rect 16163 32385 16172 32419
rect 16120 32376 16172 32385
rect 16672 32419 16724 32428
rect 16672 32385 16681 32419
rect 16681 32385 16715 32419
rect 16715 32385 16724 32419
rect 16672 32376 16724 32385
rect 16856 32376 16908 32428
rect 16304 32308 16356 32360
rect 16948 32351 17000 32360
rect 16948 32317 16957 32351
rect 16957 32317 16991 32351
rect 16991 32317 17000 32351
rect 16948 32308 17000 32317
rect 17776 32419 17828 32428
rect 17776 32385 17785 32419
rect 17785 32385 17819 32419
rect 17819 32385 17828 32419
rect 17776 32376 17828 32385
rect 11152 32172 11204 32224
rect 12532 32172 12584 32224
rect 13176 32172 13228 32224
rect 15384 32215 15436 32224
rect 15384 32181 15393 32215
rect 15393 32181 15427 32215
rect 15427 32181 15436 32215
rect 15384 32172 15436 32181
rect 15660 32172 15712 32224
rect 15752 32172 15804 32224
rect 16120 32215 16172 32224
rect 16120 32181 16129 32215
rect 16129 32181 16163 32215
rect 16163 32181 16172 32215
rect 16120 32172 16172 32181
rect 16764 32215 16816 32224
rect 16764 32181 16773 32215
rect 16773 32181 16807 32215
rect 16807 32181 16816 32215
rect 16764 32172 16816 32181
rect 17592 32172 17644 32224
rect 17776 32240 17828 32292
rect 18788 32444 18840 32496
rect 20444 32444 20496 32496
rect 21640 32512 21692 32564
rect 21732 32512 21784 32564
rect 22652 32512 22704 32564
rect 24952 32512 25004 32564
rect 27344 32512 27396 32564
rect 20812 32376 20864 32428
rect 20904 32419 20956 32428
rect 20904 32385 20913 32419
rect 20913 32385 20947 32419
rect 20947 32385 20956 32419
rect 20904 32376 20956 32385
rect 21640 32376 21692 32428
rect 20076 32240 20128 32292
rect 21732 32308 21784 32360
rect 22008 32419 22060 32428
rect 22008 32385 22017 32419
rect 22017 32385 22051 32419
rect 22051 32385 22060 32419
rect 22008 32376 22060 32385
rect 22100 32419 22152 32428
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 22100 32376 22152 32385
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 23020 32419 23072 32428
rect 23020 32385 23029 32419
rect 23029 32385 23063 32419
rect 23063 32385 23072 32419
rect 23020 32376 23072 32385
rect 24216 32419 24268 32428
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 24400 32419 24452 32428
rect 24400 32385 24409 32419
rect 24409 32385 24443 32419
rect 24443 32385 24452 32419
rect 24400 32376 24452 32385
rect 22652 32308 22704 32360
rect 24032 32308 24084 32360
rect 24584 32376 24636 32428
rect 25044 32376 25096 32428
rect 25412 32419 25464 32428
rect 25412 32385 25421 32419
rect 25421 32385 25455 32419
rect 25455 32385 25464 32419
rect 25412 32376 25464 32385
rect 28908 32444 28960 32496
rect 30932 32512 30984 32564
rect 30196 32444 30248 32496
rect 33324 32512 33376 32564
rect 25688 32419 25740 32428
rect 25688 32385 25697 32419
rect 25697 32385 25731 32419
rect 25731 32385 25740 32419
rect 25688 32376 25740 32385
rect 25964 32419 26016 32428
rect 25964 32385 25973 32419
rect 25973 32385 26007 32419
rect 26007 32385 26016 32419
rect 25964 32376 26016 32385
rect 30656 32419 30708 32428
rect 30656 32385 30665 32419
rect 30665 32385 30699 32419
rect 30699 32385 30708 32419
rect 30656 32376 30708 32385
rect 31116 32419 31168 32428
rect 31116 32385 31125 32419
rect 31125 32385 31159 32419
rect 31159 32385 31168 32419
rect 31116 32376 31168 32385
rect 31300 32419 31352 32428
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 31484 32419 31536 32428
rect 31484 32385 31493 32419
rect 31493 32385 31527 32419
rect 31527 32385 31536 32419
rect 31484 32376 31536 32385
rect 24860 32351 24912 32360
rect 24860 32317 24869 32351
rect 24869 32317 24903 32351
rect 24903 32317 24912 32351
rect 24860 32308 24912 32317
rect 25780 32308 25832 32360
rect 27252 32351 27304 32360
rect 27252 32317 27261 32351
rect 27261 32317 27295 32351
rect 27295 32317 27304 32351
rect 27252 32308 27304 32317
rect 29092 32308 29144 32360
rect 32312 32308 32364 32360
rect 32496 32351 32548 32360
rect 32496 32317 32505 32351
rect 32505 32317 32539 32351
rect 32539 32317 32548 32351
rect 32496 32308 32548 32317
rect 34428 32308 34480 32360
rect 18144 32172 18196 32224
rect 18604 32172 18656 32224
rect 19524 32172 19576 32224
rect 20628 32172 20680 32224
rect 21456 32172 21508 32224
rect 24124 32240 24176 32292
rect 24400 32240 24452 32292
rect 28816 32283 28868 32292
rect 23204 32172 23256 32224
rect 25504 32172 25556 32224
rect 26240 32172 26292 32224
rect 28816 32249 28825 32283
rect 28825 32249 28859 32283
rect 28859 32249 28868 32283
rect 28816 32240 28868 32249
rect 30564 32240 30616 32292
rect 28724 32215 28776 32224
rect 28724 32181 28733 32215
rect 28733 32181 28767 32215
rect 28767 32181 28776 32215
rect 28724 32172 28776 32181
rect 29000 32172 29052 32224
rect 31300 32172 31352 32224
rect 34060 32215 34112 32224
rect 34060 32181 34069 32215
rect 34069 32181 34103 32215
rect 34103 32181 34112 32215
rect 34060 32172 34112 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4896 31968 4948 32020
rect 6920 31900 6972 31952
rect 7104 32011 7156 32020
rect 7104 31977 7113 32011
rect 7113 31977 7147 32011
rect 7147 31977 7156 32011
rect 7104 31968 7156 31977
rect 5540 31875 5592 31884
rect 5540 31841 5549 31875
rect 5549 31841 5583 31875
rect 5583 31841 5592 31875
rect 5540 31832 5592 31841
rect 7196 31832 7248 31884
rect 7932 31900 7984 31952
rect 9496 32011 9548 32020
rect 9496 31977 9505 32011
rect 9505 31977 9539 32011
rect 9539 31977 9548 32011
rect 9496 31968 9548 31977
rect 9588 32011 9640 32020
rect 9588 31977 9597 32011
rect 9597 31977 9631 32011
rect 9631 31977 9640 32011
rect 9588 31968 9640 31977
rect 10048 31968 10100 32020
rect 10784 31968 10836 32020
rect 11336 31968 11388 32020
rect 11980 32011 12032 32020
rect 11980 31977 11989 32011
rect 11989 31977 12023 32011
rect 12023 31977 12032 32011
rect 11980 31968 12032 31977
rect 12532 31968 12584 32020
rect 14648 31968 14700 32020
rect 15384 32011 15436 32020
rect 15384 31977 15393 32011
rect 15393 31977 15427 32011
rect 15427 31977 15436 32011
rect 15384 31968 15436 31977
rect 9680 31900 9732 31952
rect 2688 31764 2740 31816
rect 4068 31696 4120 31748
rect 5264 31696 5316 31748
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 8300 31832 8352 31884
rect 8484 31832 8536 31884
rect 5356 31628 5408 31680
rect 8208 31764 8260 31816
rect 10324 31807 10376 31816
rect 10324 31773 10333 31807
rect 10333 31773 10367 31807
rect 10367 31773 10376 31807
rect 10324 31764 10376 31773
rect 10416 31807 10468 31816
rect 10416 31773 10425 31807
rect 10425 31773 10459 31807
rect 10459 31773 10468 31807
rect 10416 31764 10468 31773
rect 16304 31943 16356 31952
rect 16304 31909 16313 31943
rect 16313 31909 16347 31943
rect 16347 31909 16356 31943
rect 16304 31900 16356 31909
rect 16764 31968 16816 32020
rect 18972 31968 19024 32020
rect 19064 31968 19116 32020
rect 16856 31943 16908 31952
rect 11152 31832 11204 31884
rect 11520 31875 11572 31884
rect 11520 31841 11529 31875
rect 11529 31841 11563 31875
rect 11563 31841 11572 31875
rect 11520 31832 11572 31841
rect 14556 31832 14608 31884
rect 11612 31807 11664 31816
rect 8024 31671 8076 31680
rect 8024 31637 8033 31671
rect 8033 31637 8067 31671
rect 8067 31637 8076 31671
rect 8024 31628 8076 31637
rect 10048 31696 10100 31748
rect 10140 31739 10192 31748
rect 10140 31705 10149 31739
rect 10149 31705 10183 31739
rect 10183 31705 10192 31739
rect 10140 31696 10192 31705
rect 11612 31773 11621 31807
rect 11621 31773 11655 31807
rect 11655 31773 11664 31807
rect 11612 31764 11664 31773
rect 12072 31807 12124 31816
rect 12072 31773 12081 31807
rect 12081 31773 12115 31807
rect 12115 31773 12124 31807
rect 12072 31764 12124 31773
rect 13820 31764 13872 31816
rect 14004 31764 14056 31816
rect 15016 31807 15068 31816
rect 15016 31773 15025 31807
rect 15025 31773 15059 31807
rect 15059 31773 15068 31807
rect 15016 31764 15068 31773
rect 15292 31764 15344 31816
rect 15752 31764 15804 31816
rect 11060 31696 11112 31748
rect 15108 31696 15160 31748
rect 16120 31807 16172 31816
rect 16120 31773 16129 31807
rect 16129 31773 16163 31807
rect 16163 31773 16172 31807
rect 16120 31764 16172 31773
rect 16672 31875 16724 31884
rect 16672 31841 16681 31875
rect 16681 31841 16715 31875
rect 16715 31841 16724 31875
rect 16672 31832 16724 31841
rect 16856 31909 16865 31943
rect 16865 31909 16899 31943
rect 16899 31909 16908 31943
rect 16856 31900 16908 31909
rect 17684 31900 17736 31952
rect 17868 31900 17920 31952
rect 16856 31764 16908 31816
rect 17132 31807 17184 31816
rect 17132 31773 17141 31807
rect 17141 31773 17175 31807
rect 17175 31773 17184 31807
rect 17132 31764 17184 31773
rect 17316 31764 17368 31816
rect 17592 31764 17644 31816
rect 17960 31764 18012 31816
rect 18880 31875 18932 31884
rect 18880 31841 18889 31875
rect 18889 31841 18923 31875
rect 18923 31841 18932 31875
rect 18880 31832 18932 31841
rect 19248 31900 19300 31952
rect 8760 31628 8812 31680
rect 9128 31671 9180 31680
rect 9128 31637 9137 31671
rect 9137 31637 9171 31671
rect 9171 31637 9180 31671
rect 9128 31628 9180 31637
rect 9220 31671 9272 31680
rect 9220 31637 9229 31671
rect 9229 31637 9263 31671
rect 9263 31637 9272 31671
rect 9220 31628 9272 31637
rect 9404 31628 9456 31680
rect 11888 31628 11940 31680
rect 14740 31628 14792 31680
rect 15660 31671 15712 31680
rect 15660 31637 15669 31671
rect 15669 31637 15703 31671
rect 15703 31637 15712 31671
rect 15660 31628 15712 31637
rect 17776 31696 17828 31748
rect 19524 31764 19576 31816
rect 18880 31696 18932 31748
rect 17500 31628 17552 31680
rect 19340 31628 19392 31680
rect 19984 31807 20036 31816
rect 19984 31773 19993 31807
rect 19993 31773 20027 31807
rect 20027 31773 20036 31807
rect 19984 31764 20036 31773
rect 20076 31807 20128 31816
rect 20076 31773 20085 31807
rect 20085 31773 20119 31807
rect 20119 31773 20128 31807
rect 20076 31764 20128 31773
rect 20812 32011 20864 32020
rect 20812 31977 20821 32011
rect 20821 31977 20855 32011
rect 20855 31977 20864 32011
rect 20812 31968 20864 31977
rect 22652 31968 22704 32020
rect 22836 31968 22888 32020
rect 23848 31968 23900 32020
rect 23940 31968 23992 32020
rect 24768 31968 24820 32020
rect 27252 31968 27304 32020
rect 27528 31968 27580 32020
rect 29000 32011 29052 32020
rect 29000 31977 29009 32011
rect 29009 31977 29043 32011
rect 29043 31977 29052 32011
rect 29000 31968 29052 31977
rect 20628 31900 20680 31952
rect 22192 31900 22244 31952
rect 22376 31900 22428 31952
rect 19892 31696 19944 31748
rect 20996 31807 21048 31816
rect 20996 31773 21005 31807
rect 21005 31773 21039 31807
rect 21039 31773 21048 31807
rect 20996 31764 21048 31773
rect 21364 31807 21416 31816
rect 21364 31773 21373 31807
rect 21373 31773 21407 31807
rect 21407 31773 21416 31807
rect 21364 31764 21416 31773
rect 21456 31807 21508 31816
rect 21456 31773 21465 31807
rect 21465 31773 21499 31807
rect 21499 31773 21508 31807
rect 21456 31764 21508 31773
rect 21640 31807 21692 31816
rect 21640 31773 21649 31807
rect 21649 31773 21683 31807
rect 21683 31773 21692 31807
rect 21640 31764 21692 31773
rect 22836 31832 22888 31884
rect 25412 31900 25464 31952
rect 23940 31875 23992 31884
rect 23940 31841 23949 31875
rect 23949 31841 23983 31875
rect 23983 31841 23992 31875
rect 23940 31832 23992 31841
rect 22468 31807 22520 31816
rect 22468 31773 22477 31807
rect 22477 31773 22511 31807
rect 22511 31773 22520 31807
rect 22468 31764 22520 31773
rect 22744 31764 22796 31816
rect 23112 31764 23164 31816
rect 23204 31807 23256 31816
rect 23204 31773 23213 31807
rect 23213 31773 23247 31807
rect 23247 31773 23256 31807
rect 23204 31764 23256 31773
rect 23572 31807 23624 31816
rect 23572 31773 23581 31807
rect 23581 31773 23615 31807
rect 23615 31773 23624 31807
rect 25780 31832 25832 31884
rect 28264 31900 28316 31952
rect 23572 31764 23624 31773
rect 24308 31764 24360 31816
rect 21088 31739 21140 31748
rect 21088 31705 21097 31739
rect 21097 31705 21131 31739
rect 21131 31705 21140 31739
rect 21088 31696 21140 31705
rect 21548 31696 21600 31748
rect 19984 31628 20036 31680
rect 22928 31739 22980 31748
rect 22928 31705 22937 31739
rect 22937 31705 22971 31739
rect 22971 31705 22980 31739
rect 22928 31696 22980 31705
rect 24860 31807 24912 31816
rect 24860 31773 24869 31807
rect 24869 31773 24903 31807
rect 24903 31773 24912 31807
rect 24860 31764 24912 31773
rect 27620 31807 27672 31816
rect 27620 31773 27629 31807
rect 27629 31773 27663 31807
rect 27663 31773 27672 31807
rect 27620 31764 27672 31773
rect 25504 31696 25556 31748
rect 24400 31628 24452 31680
rect 24768 31671 24820 31680
rect 24768 31637 24777 31671
rect 24777 31637 24811 31671
rect 24811 31637 24820 31671
rect 24768 31628 24820 31637
rect 24860 31628 24912 31680
rect 27804 31739 27856 31748
rect 27804 31705 27813 31739
rect 27813 31705 27847 31739
rect 27847 31705 27856 31739
rect 27804 31696 27856 31705
rect 28448 31832 28500 31884
rect 28540 31730 28592 31782
rect 28080 31628 28132 31680
rect 28448 31628 28500 31680
rect 30748 31968 30800 32020
rect 31484 31968 31536 32020
rect 30656 31900 30708 31952
rect 29736 31832 29788 31884
rect 30196 31832 30248 31884
rect 31392 31832 31444 31884
rect 32312 31875 32364 31884
rect 32312 31841 32321 31875
rect 32321 31841 32355 31875
rect 32355 31841 32364 31875
rect 32312 31832 32364 31841
rect 33416 31832 33468 31884
rect 34520 31875 34572 31884
rect 34520 31841 34529 31875
rect 34529 31841 34563 31875
rect 34563 31841 34572 31875
rect 34520 31832 34572 31841
rect 29552 31807 29604 31816
rect 29552 31773 29561 31807
rect 29561 31773 29595 31807
rect 29595 31773 29604 31807
rect 29552 31764 29604 31773
rect 30012 31628 30064 31680
rect 30104 31628 30156 31680
rect 30564 31628 30616 31680
rect 30932 31764 30984 31816
rect 32588 31764 32640 31816
rect 34336 31696 34388 31748
rect 31116 31628 31168 31680
rect 32404 31628 32456 31680
rect 33968 31628 34020 31680
rect 34704 31671 34756 31680
rect 34704 31637 34713 31671
rect 34713 31637 34747 31671
rect 34747 31637 34756 31671
rect 34704 31628 34756 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 6736 31424 6788 31476
rect 9496 31424 9548 31476
rect 11888 31467 11940 31476
rect 11888 31433 11897 31467
rect 11897 31433 11931 31467
rect 11931 31433 11940 31467
rect 11888 31424 11940 31433
rect 5356 31356 5408 31408
rect 6368 31356 6420 31408
rect 7196 31356 7248 31408
rect 7656 31288 7708 31340
rect 3700 31152 3752 31204
rect 8208 31288 8260 31340
rect 9220 31331 9272 31340
rect 9220 31297 9229 31331
rect 9229 31297 9263 31331
rect 9263 31297 9272 31331
rect 9220 31288 9272 31297
rect 9312 31288 9364 31340
rect 8944 31220 8996 31272
rect 10140 31356 10192 31408
rect 10784 31399 10836 31408
rect 10784 31365 10793 31399
rect 10793 31365 10827 31399
rect 10827 31365 10836 31399
rect 10784 31356 10836 31365
rect 9956 31331 10008 31340
rect 9956 31297 9965 31331
rect 9965 31297 9999 31331
rect 9999 31297 10008 31331
rect 9956 31288 10008 31297
rect 10508 31288 10560 31340
rect 11336 31356 11388 31408
rect 11520 31399 11572 31408
rect 11520 31365 11529 31399
rect 11529 31365 11563 31399
rect 11563 31365 11572 31399
rect 11520 31356 11572 31365
rect 11612 31356 11664 31408
rect 11060 31288 11112 31340
rect 11244 31288 11296 31340
rect 11888 31331 11940 31340
rect 11888 31297 11897 31331
rect 11897 31297 11931 31331
rect 11931 31297 11940 31331
rect 11888 31288 11940 31297
rect 12072 31331 12124 31340
rect 12072 31297 12081 31331
rect 12081 31297 12115 31331
rect 12115 31297 12124 31331
rect 12072 31288 12124 31297
rect 13176 31288 13228 31340
rect 14740 31424 14792 31476
rect 15844 31424 15896 31476
rect 16028 31424 16080 31476
rect 17316 31424 17368 31476
rect 18880 31467 18932 31476
rect 18880 31433 18889 31467
rect 18889 31433 18923 31467
rect 18923 31433 18932 31467
rect 18880 31424 18932 31433
rect 19432 31467 19484 31476
rect 19432 31433 19441 31467
rect 19441 31433 19475 31467
rect 19475 31433 19484 31467
rect 19432 31424 19484 31433
rect 19892 31424 19944 31476
rect 20720 31424 20772 31476
rect 24216 31424 24268 31476
rect 14004 31356 14056 31408
rect 15292 31356 15344 31408
rect 13728 31331 13780 31340
rect 13728 31297 13737 31331
rect 13737 31297 13771 31331
rect 13771 31297 13780 31331
rect 13728 31288 13780 31297
rect 15108 31288 15160 31340
rect 17684 31356 17736 31408
rect 18144 31399 18196 31408
rect 18144 31365 18153 31399
rect 18153 31365 18187 31399
rect 18187 31365 18196 31399
rect 18144 31356 18196 31365
rect 8484 31152 8536 31204
rect 9312 31195 9364 31204
rect 9312 31161 9321 31195
rect 9321 31161 9355 31195
rect 9355 31161 9364 31195
rect 9312 31152 9364 31161
rect 14556 31220 14608 31272
rect 15016 31220 15068 31272
rect 16856 31288 16908 31340
rect 18604 31356 18656 31408
rect 19156 31356 19208 31408
rect 19340 31331 19392 31340
rect 19340 31297 19349 31331
rect 19349 31297 19383 31331
rect 19383 31297 19392 31331
rect 19340 31288 19392 31297
rect 19432 31331 19484 31340
rect 19432 31297 19441 31331
rect 19441 31297 19475 31331
rect 19475 31297 19484 31331
rect 19432 31288 19484 31297
rect 19984 31356 20036 31408
rect 12900 31152 12952 31204
rect 15108 31152 15160 31204
rect 17684 31220 17736 31272
rect 18052 31220 18104 31272
rect 19248 31220 19300 31272
rect 18696 31152 18748 31204
rect 19892 31288 19944 31340
rect 20812 31331 20864 31340
rect 20812 31297 20821 31331
rect 20821 31297 20855 31331
rect 20855 31297 20864 31331
rect 20812 31288 20864 31297
rect 21364 31288 21416 31340
rect 21456 31331 21508 31340
rect 21456 31297 21465 31331
rect 21465 31297 21499 31331
rect 21499 31297 21508 31331
rect 21456 31288 21508 31297
rect 21548 31220 21600 31272
rect 22100 31356 22152 31408
rect 23848 31399 23900 31408
rect 23848 31365 23857 31399
rect 23857 31365 23891 31399
rect 23891 31365 23900 31399
rect 23848 31356 23900 31365
rect 24124 31356 24176 31408
rect 24768 31424 24820 31476
rect 24584 31399 24636 31408
rect 24584 31365 24593 31399
rect 24593 31365 24627 31399
rect 24627 31365 24636 31399
rect 24584 31356 24636 31365
rect 22468 31331 22520 31340
rect 20076 31152 20128 31204
rect 22468 31297 22477 31331
rect 22477 31297 22511 31331
rect 22511 31297 22520 31331
rect 22468 31288 22520 31297
rect 22836 31288 22888 31340
rect 24216 31331 24268 31340
rect 24216 31297 24225 31331
rect 24225 31297 24259 31331
rect 24259 31297 24268 31331
rect 24216 31288 24268 31297
rect 24400 31331 24452 31340
rect 24400 31297 24409 31331
rect 24409 31297 24443 31331
rect 24443 31297 24452 31331
rect 24400 31288 24452 31297
rect 24860 31331 24912 31340
rect 24860 31297 24869 31331
rect 24869 31297 24903 31331
rect 24903 31297 24912 31331
rect 24860 31288 24912 31297
rect 26148 31288 26200 31340
rect 27988 31399 28040 31408
rect 27988 31365 27997 31399
rect 27997 31365 28031 31399
rect 28031 31365 28040 31399
rect 27988 31356 28040 31365
rect 28080 31399 28132 31408
rect 28080 31365 28089 31399
rect 28089 31365 28123 31399
rect 28123 31365 28132 31399
rect 28080 31356 28132 31365
rect 29092 31424 29144 31476
rect 22560 31220 22612 31272
rect 25596 31220 25648 31272
rect 25688 31263 25740 31272
rect 25688 31229 25697 31263
rect 25697 31229 25731 31263
rect 25731 31229 25740 31263
rect 25688 31220 25740 31229
rect 5540 31084 5592 31136
rect 9036 31127 9088 31136
rect 9036 31093 9045 31127
rect 9045 31093 9079 31127
rect 9079 31093 9088 31127
rect 9036 31084 9088 31093
rect 9220 31084 9272 31136
rect 9956 31084 10008 31136
rect 14188 31084 14240 31136
rect 16672 31127 16724 31136
rect 16672 31093 16681 31127
rect 16681 31093 16715 31127
rect 16715 31093 16724 31127
rect 16672 31084 16724 31093
rect 16764 31084 16816 31136
rect 21272 31084 21324 31136
rect 21456 31084 21508 31136
rect 25964 31084 26016 31136
rect 26608 31084 26660 31136
rect 26976 31084 27028 31136
rect 27620 31220 27672 31272
rect 28356 31288 28408 31340
rect 28264 31220 28316 31272
rect 28724 31288 28776 31340
rect 29184 31331 29236 31340
rect 29184 31297 29193 31331
rect 29193 31297 29227 31331
rect 29227 31297 29236 31331
rect 29184 31288 29236 31297
rect 28816 31220 28868 31272
rect 29460 31220 29512 31272
rect 29736 31356 29788 31408
rect 30840 31424 30892 31476
rect 32496 31424 32548 31476
rect 33416 31424 33468 31476
rect 34704 31424 34756 31476
rect 34060 31356 34112 31408
rect 34428 31399 34480 31408
rect 34428 31365 34437 31399
rect 34437 31365 34471 31399
rect 34471 31365 34480 31399
rect 34428 31356 34480 31365
rect 29828 31263 29880 31272
rect 29828 31229 29837 31263
rect 29837 31229 29871 31263
rect 29871 31229 29880 31263
rect 29828 31220 29880 31229
rect 30840 31220 30892 31272
rect 32404 31288 32456 31340
rect 32680 31331 32732 31340
rect 32680 31297 32689 31331
rect 32689 31297 32723 31331
rect 32723 31297 32732 31331
rect 32680 31288 32732 31297
rect 33048 31288 33100 31340
rect 33876 31288 33928 31340
rect 33968 31331 34020 31340
rect 33968 31297 33977 31331
rect 33977 31297 34011 31331
rect 34011 31297 34020 31331
rect 33968 31288 34020 31297
rect 34520 31288 34572 31340
rect 34152 31220 34204 31272
rect 29092 31152 29144 31204
rect 31116 31152 31168 31204
rect 27620 31084 27672 31136
rect 27712 31084 27764 31136
rect 30196 31084 30248 31136
rect 31300 31127 31352 31136
rect 31300 31093 31309 31127
rect 31309 31093 31343 31127
rect 31343 31093 31352 31127
rect 31300 31084 31352 31093
rect 31668 31084 31720 31136
rect 33324 31084 33376 31136
rect 34428 31084 34480 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 8944 30880 8996 30932
rect 8392 30812 8444 30864
rect 8576 30812 8628 30864
rect 9128 30812 9180 30864
rect 9312 30880 9364 30932
rect 6920 30787 6972 30796
rect 6920 30753 6929 30787
rect 6929 30753 6963 30787
rect 6963 30753 6972 30787
rect 6920 30744 6972 30753
rect 10968 30880 11020 30932
rect 11704 30880 11756 30932
rect 11888 30880 11940 30932
rect 14464 30880 14516 30932
rect 14556 30923 14608 30932
rect 14556 30889 14565 30923
rect 14565 30889 14599 30923
rect 14599 30889 14608 30923
rect 14556 30880 14608 30889
rect 10784 30812 10836 30864
rect 12072 30812 12124 30864
rect 17040 30880 17092 30932
rect 17684 30880 17736 30932
rect 17868 30880 17920 30932
rect 5172 30719 5224 30728
rect 5172 30685 5181 30719
rect 5181 30685 5215 30719
rect 5215 30685 5224 30719
rect 5172 30676 5224 30685
rect 7196 30719 7248 30728
rect 7196 30685 7205 30719
rect 7205 30685 7239 30719
rect 7239 30685 7248 30719
rect 10048 30744 10100 30796
rect 14556 30744 14608 30796
rect 18236 30812 18288 30864
rect 20812 30812 20864 30864
rect 20996 30923 21048 30932
rect 20996 30889 21005 30923
rect 21005 30889 21039 30923
rect 21039 30889 21048 30923
rect 20996 30880 21048 30889
rect 21088 30880 21140 30932
rect 22284 30880 22336 30932
rect 24860 30880 24912 30932
rect 28816 30880 28868 30932
rect 21456 30812 21508 30864
rect 23572 30812 23624 30864
rect 27804 30812 27856 30864
rect 29276 30812 29328 30864
rect 29920 30880 29972 30932
rect 30932 30880 30984 30932
rect 34336 30880 34388 30932
rect 7196 30676 7248 30685
rect 4068 30608 4120 30660
rect 5632 30608 5684 30660
rect 7104 30540 7156 30592
rect 7288 30540 7340 30592
rect 7840 30651 7892 30660
rect 7840 30617 7849 30651
rect 7849 30617 7883 30651
rect 7883 30617 7892 30651
rect 7840 30608 7892 30617
rect 8208 30608 8260 30660
rect 9128 30676 9180 30728
rect 9588 30719 9640 30728
rect 9588 30685 9597 30719
rect 9597 30685 9631 30719
rect 9631 30685 9640 30719
rect 9588 30676 9640 30685
rect 9772 30719 9824 30728
rect 9772 30685 9781 30719
rect 9781 30685 9815 30719
rect 9815 30685 9824 30719
rect 9772 30676 9824 30685
rect 9680 30608 9732 30660
rect 11152 30719 11204 30728
rect 11152 30685 11161 30719
rect 11161 30685 11195 30719
rect 11195 30685 11204 30719
rect 11152 30676 11204 30685
rect 14188 30719 14240 30728
rect 14188 30685 14197 30719
rect 14197 30685 14231 30719
rect 14231 30685 14240 30719
rect 14188 30676 14240 30685
rect 15660 30676 15712 30728
rect 16672 30676 16724 30728
rect 17132 30676 17184 30728
rect 17316 30676 17368 30728
rect 21364 30744 21416 30796
rect 22928 30744 22980 30796
rect 25780 30744 25832 30796
rect 25964 30787 26016 30796
rect 25964 30753 25973 30787
rect 25973 30753 26007 30787
rect 26007 30753 26016 30787
rect 25964 30744 26016 30753
rect 26148 30744 26200 30796
rect 9956 30608 10008 30660
rect 10324 30608 10376 30660
rect 16764 30608 16816 30660
rect 8852 30540 8904 30592
rect 11244 30583 11296 30592
rect 11244 30549 11253 30583
rect 11253 30549 11287 30583
rect 11287 30549 11296 30583
rect 11244 30540 11296 30549
rect 13912 30540 13964 30592
rect 17500 30540 17552 30592
rect 19892 30608 19944 30660
rect 21272 30719 21324 30728
rect 21272 30685 21281 30719
rect 21281 30685 21315 30719
rect 21315 30685 21324 30719
rect 21272 30676 21324 30685
rect 23112 30719 23164 30728
rect 23112 30685 23121 30719
rect 23121 30685 23155 30719
rect 23155 30685 23164 30719
rect 23112 30676 23164 30685
rect 23204 30676 23256 30728
rect 22928 30608 22980 30660
rect 24676 30719 24728 30728
rect 24676 30685 24685 30719
rect 24685 30685 24719 30719
rect 24719 30685 24728 30719
rect 24676 30676 24728 30685
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 25228 30719 25280 30728
rect 25228 30685 25237 30719
rect 25237 30685 25271 30719
rect 25271 30685 25280 30719
rect 25228 30676 25280 30685
rect 23756 30608 23808 30660
rect 25688 30676 25740 30728
rect 27712 30719 27764 30728
rect 27712 30685 27721 30719
rect 27721 30685 27755 30719
rect 27755 30685 27764 30719
rect 27712 30676 27764 30685
rect 23020 30540 23072 30592
rect 23664 30540 23716 30592
rect 26976 30608 27028 30660
rect 27344 30540 27396 30592
rect 28172 30744 28224 30796
rect 31024 30812 31076 30864
rect 32496 30812 32548 30864
rect 28080 30676 28132 30728
rect 30840 30744 30892 30796
rect 32312 30744 32364 30796
rect 30012 30676 30064 30728
rect 30656 30676 30708 30728
rect 29460 30608 29512 30660
rect 29644 30608 29696 30660
rect 32864 30651 32916 30660
rect 32864 30617 32873 30651
rect 32873 30617 32907 30651
rect 32907 30617 32916 30651
rect 32864 30608 32916 30617
rect 34428 30608 34480 30660
rect 31024 30540 31076 30592
rect 31116 30583 31168 30592
rect 31116 30549 31125 30583
rect 31125 30549 31159 30583
rect 31159 30549 31168 30583
rect 31116 30540 31168 30549
rect 33232 30540 33284 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 5632 30336 5684 30388
rect 8024 30336 8076 30388
rect 3700 30311 3752 30320
rect 3700 30277 3709 30311
rect 3709 30277 3743 30311
rect 3743 30277 3752 30311
rect 3700 30268 3752 30277
rect 4068 30268 4120 30320
rect 5540 30268 5592 30320
rect 7104 30268 7156 30320
rect 8760 30336 8812 30388
rect 9220 30336 9272 30388
rect 11152 30336 11204 30388
rect 14464 30336 14516 30388
rect 5816 30200 5868 30252
rect 6276 30200 6328 30252
rect 9404 30268 9456 30320
rect 19892 30336 19944 30388
rect 20352 30336 20404 30388
rect 23296 30336 23348 30388
rect 23664 30336 23716 30388
rect 24768 30336 24820 30388
rect 6644 30175 6696 30184
rect 6644 30141 6653 30175
rect 6653 30141 6687 30175
rect 6687 30141 6696 30175
rect 6644 30132 6696 30141
rect 6736 30132 6788 30184
rect 8300 30132 8352 30184
rect 8484 30200 8536 30252
rect 8852 30200 8904 30252
rect 9496 30200 9548 30252
rect 10048 30200 10100 30252
rect 10876 30200 10928 30252
rect 18788 30268 18840 30320
rect 20260 30268 20312 30320
rect 26240 30268 26292 30320
rect 26608 30268 26660 30320
rect 28632 30336 28684 30388
rect 29184 30336 29236 30388
rect 29276 30336 29328 30388
rect 29920 30336 29972 30388
rect 29736 30268 29788 30320
rect 18144 30200 18196 30252
rect 18512 30200 18564 30252
rect 18604 30243 18656 30252
rect 18604 30209 18613 30243
rect 18613 30209 18647 30243
rect 18647 30209 18656 30243
rect 18604 30200 18656 30209
rect 22928 30243 22980 30252
rect 22928 30209 22937 30243
rect 22937 30209 22971 30243
rect 22971 30209 22980 30243
rect 22928 30200 22980 30209
rect 8116 30039 8168 30048
rect 8116 30005 8125 30039
rect 8125 30005 8159 30039
rect 8159 30005 8168 30039
rect 8116 29996 8168 30005
rect 9128 29996 9180 30048
rect 9496 29996 9548 30048
rect 10140 30064 10192 30116
rect 16948 30064 17000 30116
rect 17684 30132 17736 30184
rect 18420 30175 18472 30184
rect 18420 30141 18429 30175
rect 18429 30141 18463 30175
rect 18463 30141 18472 30175
rect 18420 30132 18472 30141
rect 17960 30064 18012 30116
rect 19892 30132 19944 30184
rect 11796 29996 11848 30048
rect 12716 29996 12768 30048
rect 13176 29996 13228 30048
rect 13452 29996 13504 30048
rect 18236 29996 18288 30048
rect 21180 30132 21232 30184
rect 23204 30200 23256 30252
rect 23664 30243 23716 30252
rect 23664 30209 23673 30243
rect 23673 30209 23707 30243
rect 23707 30209 23716 30243
rect 23664 30200 23716 30209
rect 23480 30132 23532 30184
rect 23112 30064 23164 30116
rect 27344 30243 27396 30252
rect 27344 30209 27353 30243
rect 27353 30209 27387 30243
rect 27387 30209 27396 30243
rect 27344 30200 27396 30209
rect 27528 30243 27580 30252
rect 27528 30209 27537 30243
rect 27537 30209 27571 30243
rect 27571 30209 27580 30243
rect 27528 30200 27580 30209
rect 24952 30132 25004 30184
rect 28264 30175 28316 30184
rect 28264 30141 28273 30175
rect 28273 30141 28307 30175
rect 28307 30141 28316 30175
rect 28264 30132 28316 30141
rect 28540 30200 28592 30252
rect 28908 30200 28960 30252
rect 30288 30243 30340 30252
rect 30288 30209 30297 30243
rect 30297 30209 30331 30243
rect 30331 30209 30340 30243
rect 30288 30200 30340 30209
rect 30748 30311 30800 30320
rect 30748 30277 30757 30311
rect 30757 30277 30791 30311
rect 30791 30277 30800 30311
rect 30748 30268 30800 30277
rect 29000 30132 29052 30184
rect 29368 30132 29420 30184
rect 30656 30243 30708 30252
rect 30656 30209 30665 30243
rect 30665 30209 30699 30243
rect 30699 30209 30708 30243
rect 30656 30200 30708 30209
rect 30932 30200 30984 30252
rect 32404 30336 32456 30388
rect 31392 30268 31444 30320
rect 32220 30268 32272 30320
rect 32680 30379 32732 30388
rect 32680 30345 32689 30379
rect 32689 30345 32723 30379
rect 32723 30345 32732 30379
rect 32680 30336 32732 30345
rect 31484 30243 31536 30252
rect 31484 30209 31493 30243
rect 31493 30209 31527 30243
rect 31527 30209 31536 30243
rect 31484 30200 31536 30209
rect 30564 30132 30616 30184
rect 31760 30243 31812 30252
rect 31760 30209 31769 30243
rect 31769 30209 31803 30243
rect 31803 30209 31812 30243
rect 31760 30200 31812 30209
rect 32128 30243 32180 30252
rect 32128 30209 32137 30243
rect 32137 30209 32171 30243
rect 32171 30209 32180 30243
rect 32128 30200 32180 30209
rect 32312 30243 32364 30252
rect 32312 30209 32321 30243
rect 32321 30209 32355 30243
rect 32355 30209 32364 30243
rect 32312 30200 32364 30209
rect 32404 30243 32456 30252
rect 32404 30209 32413 30243
rect 32413 30209 32447 30243
rect 32447 30209 32456 30243
rect 32404 30200 32456 30209
rect 32864 30268 32916 30320
rect 32772 30243 32824 30252
rect 32772 30209 32781 30243
rect 32781 30209 32815 30243
rect 32815 30209 32824 30243
rect 32772 30200 32824 30209
rect 32956 30243 33008 30252
rect 32956 30209 32965 30243
rect 32965 30209 32999 30243
rect 32999 30209 33008 30243
rect 32956 30200 33008 30209
rect 33600 30268 33652 30320
rect 33416 30243 33468 30252
rect 33416 30209 33425 30243
rect 33425 30209 33459 30243
rect 33459 30209 33468 30243
rect 33416 30200 33468 30209
rect 33692 30243 33744 30252
rect 33692 30209 33701 30243
rect 33701 30209 33735 30243
rect 33735 30209 33744 30243
rect 33692 30200 33744 30209
rect 23572 29996 23624 30048
rect 24216 30039 24268 30048
rect 24216 30005 24225 30039
rect 24225 30005 24259 30039
rect 24259 30005 24268 30039
rect 24216 29996 24268 30005
rect 25320 29996 25372 30048
rect 26332 30039 26384 30048
rect 26332 30005 26341 30039
rect 26341 30005 26375 30039
rect 26375 30005 26384 30039
rect 26332 29996 26384 30005
rect 27620 30107 27672 30116
rect 27620 30073 27629 30107
rect 27629 30073 27663 30107
rect 27663 30073 27672 30107
rect 27620 30064 27672 30073
rect 27896 30064 27948 30116
rect 27988 30064 28040 30116
rect 28632 30064 28684 30116
rect 28908 30064 28960 30116
rect 28172 29996 28224 30048
rect 28724 29996 28776 30048
rect 31944 30064 31996 30116
rect 32588 29996 32640 30048
rect 32864 29996 32916 30048
rect 34152 30175 34204 30184
rect 34152 30141 34161 30175
rect 34161 30141 34195 30175
rect 34195 30141 34204 30175
rect 34152 30132 34204 30141
rect 34428 29996 34480 30048
rect 36084 30200 36136 30252
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6644 29792 6696 29844
rect 3056 29699 3108 29708
rect 3056 29665 3065 29699
rect 3065 29665 3099 29699
rect 3099 29665 3108 29699
rect 3056 29656 3108 29665
rect 6276 29656 6328 29708
rect 9680 29792 9732 29844
rect 10692 29792 10744 29844
rect 8024 29724 8076 29776
rect 8208 29699 8260 29708
rect 8208 29665 8217 29699
rect 8217 29665 8251 29699
rect 8251 29665 8260 29699
rect 8208 29656 8260 29665
rect 4344 29588 4396 29640
rect 5264 29588 5316 29640
rect 6920 29588 6972 29640
rect 7656 29631 7708 29640
rect 7656 29597 7665 29631
rect 7665 29597 7699 29631
rect 7699 29597 7708 29631
rect 7656 29588 7708 29597
rect 7932 29588 7984 29640
rect 8300 29588 8352 29640
rect 8392 29631 8444 29640
rect 8392 29597 8401 29631
rect 8401 29597 8435 29631
rect 8435 29597 8444 29631
rect 8392 29588 8444 29597
rect 8668 29588 8720 29640
rect 10048 29724 10100 29776
rect 17500 29835 17552 29844
rect 17500 29801 17509 29835
rect 17509 29801 17543 29835
rect 17543 29801 17552 29835
rect 17500 29792 17552 29801
rect 9312 29631 9364 29640
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 11060 29699 11112 29708
rect 11060 29665 11069 29699
rect 11069 29665 11103 29699
rect 11103 29665 11112 29699
rect 11060 29656 11112 29665
rect 12440 29656 12492 29708
rect 13360 29656 13412 29708
rect 13452 29656 13504 29708
rect 10324 29631 10376 29640
rect 10324 29597 10333 29631
rect 10333 29597 10367 29631
rect 10367 29597 10376 29631
rect 10324 29588 10376 29597
rect 5448 29520 5500 29572
rect 7564 29520 7616 29572
rect 8116 29520 8168 29572
rect 10508 29588 10560 29640
rect 10876 29588 10928 29640
rect 12716 29631 12768 29640
rect 12716 29597 12720 29631
rect 12720 29597 12754 29631
rect 12754 29597 12768 29631
rect 12716 29588 12768 29597
rect 13084 29631 13136 29640
rect 13084 29597 13092 29631
rect 13092 29597 13126 29631
rect 13126 29597 13136 29631
rect 13084 29588 13136 29597
rect 13636 29588 13688 29640
rect 15200 29656 15252 29708
rect 15936 29656 15988 29708
rect 17224 29724 17276 29776
rect 17408 29656 17460 29708
rect 1768 29452 1820 29504
rect 2872 29452 2924 29504
rect 4160 29452 4212 29504
rect 4620 29495 4672 29504
rect 4620 29461 4629 29495
rect 4629 29461 4663 29495
rect 4663 29461 4672 29495
rect 4620 29452 4672 29461
rect 5724 29495 5776 29504
rect 5724 29461 5733 29495
rect 5733 29461 5767 29495
rect 5767 29461 5776 29495
rect 5724 29452 5776 29461
rect 7104 29495 7156 29504
rect 7104 29461 7113 29495
rect 7113 29461 7147 29495
rect 7147 29461 7156 29495
rect 7104 29452 7156 29461
rect 7288 29452 7340 29504
rect 10140 29452 10192 29504
rect 10600 29520 10652 29572
rect 10968 29520 11020 29572
rect 11244 29520 11296 29572
rect 12624 29520 12676 29572
rect 13728 29520 13780 29572
rect 11336 29452 11388 29504
rect 12532 29495 12584 29504
rect 12532 29461 12541 29495
rect 12541 29461 12575 29495
rect 12575 29461 12584 29495
rect 12532 29452 12584 29461
rect 13820 29452 13872 29504
rect 14464 29452 14516 29504
rect 15292 29563 15344 29572
rect 15292 29529 15301 29563
rect 15301 29529 15335 29563
rect 15335 29529 15344 29563
rect 15292 29520 15344 29529
rect 15568 29631 15620 29640
rect 15568 29597 15577 29631
rect 15577 29597 15611 29631
rect 15611 29597 15620 29631
rect 15568 29588 15620 29597
rect 15752 29588 15804 29640
rect 17500 29588 17552 29640
rect 17684 29631 17736 29640
rect 17684 29597 17693 29631
rect 17693 29597 17727 29631
rect 17727 29597 17736 29631
rect 17684 29588 17736 29597
rect 18604 29792 18656 29844
rect 17960 29724 18012 29776
rect 18788 29835 18840 29844
rect 18788 29801 18797 29835
rect 18797 29801 18831 29835
rect 18831 29801 18840 29835
rect 18788 29792 18840 29801
rect 19892 29792 19944 29844
rect 17960 29631 18012 29640
rect 17960 29597 17969 29631
rect 17969 29597 18003 29631
rect 18003 29597 18012 29631
rect 17960 29588 18012 29597
rect 18420 29656 18472 29708
rect 21824 29724 21876 29776
rect 21916 29724 21968 29776
rect 22560 29724 22612 29776
rect 24952 29835 25004 29844
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 24952 29792 25004 29801
rect 27620 29792 27672 29844
rect 28264 29792 28316 29844
rect 29276 29792 29328 29844
rect 29368 29835 29420 29844
rect 29368 29801 29377 29835
rect 29377 29801 29411 29835
rect 29411 29801 29420 29835
rect 29368 29792 29420 29801
rect 29828 29792 29880 29844
rect 31484 29792 31536 29844
rect 33692 29792 33744 29844
rect 26332 29724 26384 29776
rect 18696 29656 18748 29708
rect 22100 29656 22152 29708
rect 18144 29631 18196 29640
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 18236 29631 18288 29640
rect 18236 29597 18246 29631
rect 18246 29597 18280 29631
rect 18280 29597 18288 29631
rect 18236 29588 18288 29597
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 21640 29631 21692 29640
rect 21640 29597 21649 29631
rect 21649 29597 21683 29631
rect 21683 29597 21692 29631
rect 21640 29588 21692 29597
rect 15660 29520 15712 29572
rect 16212 29520 16264 29572
rect 16856 29563 16908 29572
rect 16856 29529 16865 29563
rect 16865 29529 16899 29563
rect 16899 29529 16908 29563
rect 16856 29520 16908 29529
rect 15384 29452 15436 29504
rect 18052 29452 18104 29504
rect 18328 29452 18380 29504
rect 18512 29563 18564 29572
rect 18512 29529 18521 29563
rect 18521 29529 18555 29563
rect 18555 29529 18564 29563
rect 18512 29520 18564 29529
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 22284 29631 22336 29640
rect 22284 29597 22293 29631
rect 22293 29597 22327 29631
rect 22327 29597 22336 29631
rect 22284 29588 22336 29597
rect 22468 29699 22520 29708
rect 22468 29665 22477 29699
rect 22477 29665 22511 29699
rect 22511 29665 22520 29699
rect 22468 29656 22520 29665
rect 22744 29699 22796 29708
rect 22744 29665 22753 29699
rect 22753 29665 22787 29699
rect 22787 29665 22796 29699
rect 22744 29656 22796 29665
rect 24216 29656 24268 29708
rect 22468 29520 22520 29572
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 22836 29588 22888 29597
rect 24308 29588 24360 29640
rect 24860 29656 24912 29708
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 26884 29656 26936 29708
rect 27988 29656 28040 29708
rect 24768 29588 24820 29597
rect 26608 29588 26660 29640
rect 23664 29520 23716 29572
rect 26056 29563 26108 29572
rect 26056 29529 26065 29563
rect 26065 29529 26099 29563
rect 26099 29529 26108 29563
rect 26056 29520 26108 29529
rect 20628 29452 20680 29504
rect 21824 29452 21876 29504
rect 22100 29452 22152 29504
rect 22192 29452 22244 29504
rect 23940 29452 23992 29504
rect 26884 29563 26936 29572
rect 26884 29529 26893 29563
rect 26893 29529 26927 29563
rect 26927 29529 26936 29563
rect 26884 29520 26936 29529
rect 27252 29563 27304 29572
rect 27252 29529 27261 29563
rect 27261 29529 27295 29563
rect 27295 29529 27304 29563
rect 27252 29520 27304 29529
rect 28540 29520 28592 29572
rect 27160 29452 27212 29504
rect 29000 29656 29052 29708
rect 30012 29656 30064 29708
rect 30472 29699 30524 29708
rect 30472 29665 30481 29699
rect 30481 29665 30515 29699
rect 30515 29665 30524 29699
rect 30472 29656 30524 29665
rect 31576 29724 31628 29776
rect 32312 29724 32364 29776
rect 34704 29724 34756 29776
rect 31668 29699 31720 29708
rect 31668 29665 31677 29699
rect 31677 29665 31711 29699
rect 31711 29665 31720 29699
rect 31668 29656 31720 29665
rect 28724 29588 28776 29640
rect 28908 29588 28960 29640
rect 30196 29588 30248 29640
rect 30748 29588 30800 29640
rect 30840 29588 30892 29640
rect 29000 29563 29052 29572
rect 29000 29529 29009 29563
rect 29009 29529 29043 29563
rect 29043 29529 29052 29563
rect 29000 29520 29052 29529
rect 29276 29520 29328 29572
rect 31208 29631 31260 29640
rect 31208 29597 31217 29631
rect 31217 29597 31251 29631
rect 31251 29597 31260 29631
rect 31208 29588 31260 29597
rect 31392 29631 31444 29640
rect 31392 29597 31401 29631
rect 31401 29597 31435 29631
rect 31435 29597 31444 29631
rect 31392 29588 31444 29597
rect 32128 29631 32180 29640
rect 32128 29597 32137 29631
rect 32137 29597 32171 29631
rect 32171 29597 32180 29631
rect 32128 29588 32180 29597
rect 32404 29588 32456 29640
rect 32680 29588 32732 29640
rect 34520 29631 34572 29640
rect 34520 29597 34529 29631
rect 34529 29597 34563 29631
rect 34563 29597 34572 29631
rect 34520 29588 34572 29597
rect 34612 29588 34664 29640
rect 35624 29631 35676 29640
rect 35624 29597 35633 29631
rect 35633 29597 35667 29631
rect 35667 29597 35676 29631
rect 35624 29588 35676 29597
rect 32588 29520 32640 29572
rect 33784 29520 33836 29572
rect 28816 29452 28868 29504
rect 30288 29452 30340 29504
rect 30748 29452 30800 29504
rect 31668 29452 31720 29504
rect 32128 29452 32180 29504
rect 32220 29495 32272 29504
rect 32220 29461 32229 29495
rect 32229 29461 32263 29495
rect 32263 29461 32272 29495
rect 32220 29452 32272 29461
rect 32404 29452 32456 29504
rect 33048 29452 33100 29504
rect 34060 29452 34112 29504
rect 34336 29452 34388 29504
rect 36084 29495 36136 29504
rect 36084 29461 36093 29495
rect 36093 29461 36127 29495
rect 36127 29461 36136 29495
rect 36084 29452 36136 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 1768 29223 1820 29232
rect 1768 29189 1777 29223
rect 1777 29189 1811 29223
rect 1811 29189 1820 29223
rect 1768 29180 1820 29189
rect 4068 29248 4120 29300
rect 4160 29180 4212 29232
rect 4804 29248 4856 29300
rect 5724 29248 5776 29300
rect 7104 29248 7156 29300
rect 6644 29180 6696 29232
rect 6920 29180 6972 29232
rect 7656 29180 7708 29232
rect 8024 29248 8076 29300
rect 5264 29112 5316 29164
rect 1400 29044 1452 29096
rect 4344 29044 4396 29096
rect 6276 29044 6328 29096
rect 7288 29112 7340 29164
rect 7380 29155 7432 29164
rect 7380 29121 7389 29155
rect 7389 29121 7423 29155
rect 7423 29121 7432 29155
rect 7380 29112 7432 29121
rect 7748 29112 7800 29164
rect 5264 28976 5316 29028
rect 7380 28976 7432 29028
rect 8024 28976 8076 29028
rect 8300 29155 8352 29164
rect 9036 29248 9088 29300
rect 9312 29291 9364 29300
rect 9312 29257 9321 29291
rect 9321 29257 9355 29291
rect 9355 29257 9364 29291
rect 9312 29248 9364 29257
rect 10232 29248 10284 29300
rect 10324 29248 10376 29300
rect 11612 29248 11664 29300
rect 9404 29180 9456 29232
rect 8300 29121 8345 29155
rect 8345 29121 8352 29155
rect 8300 29112 8352 29121
rect 8944 29155 8996 29164
rect 8944 29121 8953 29155
rect 8953 29121 8987 29155
rect 8987 29121 8996 29155
rect 8944 29112 8996 29121
rect 9128 29112 9180 29164
rect 9588 29155 9640 29164
rect 9588 29121 9597 29155
rect 9597 29121 9631 29155
rect 9631 29121 9640 29155
rect 9588 29112 9640 29121
rect 11244 29180 11296 29232
rect 11336 29180 11388 29232
rect 13084 29248 13136 29300
rect 10048 29112 10100 29164
rect 10140 29044 10192 29096
rect 9220 28976 9272 29028
rect 10232 28976 10284 29028
rect 5356 28951 5408 28960
rect 5356 28917 5365 28951
rect 5365 28917 5399 28951
rect 5399 28917 5408 28951
rect 5356 28908 5408 28917
rect 6092 28908 6144 28960
rect 8668 28908 8720 28960
rect 10324 28908 10376 28960
rect 10600 29112 10652 29164
rect 10876 29155 10928 29164
rect 10876 29121 10885 29155
rect 10885 29121 10919 29155
rect 10919 29121 10928 29155
rect 10876 29112 10928 29121
rect 11520 29112 11572 29164
rect 12992 29180 13044 29232
rect 13820 29248 13872 29300
rect 13728 29180 13780 29232
rect 10784 29087 10836 29096
rect 10784 29053 10793 29087
rect 10793 29053 10827 29087
rect 10827 29053 10836 29087
rect 10784 29044 10836 29053
rect 10968 29044 11020 29096
rect 10692 28976 10744 29028
rect 12072 29112 12124 29164
rect 11888 29044 11940 29096
rect 12348 29155 12400 29164
rect 12348 29121 12358 29155
rect 12358 29121 12392 29155
rect 12392 29121 12400 29155
rect 12348 29112 12400 29121
rect 12900 29112 12952 29164
rect 13176 29155 13228 29164
rect 13176 29121 13180 29155
rect 13180 29121 13214 29155
rect 13214 29121 13228 29155
rect 13176 29112 13228 29121
rect 13452 29112 13504 29164
rect 13636 29155 13688 29164
rect 13636 29121 13645 29155
rect 13645 29121 13679 29155
rect 13679 29121 13688 29155
rect 15568 29248 15620 29300
rect 15200 29180 15252 29232
rect 13636 29112 13688 29121
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14096 29112 14148 29121
rect 13820 29044 13872 29096
rect 14188 29044 14240 29096
rect 13452 28976 13504 29028
rect 13544 28976 13596 29028
rect 14464 29155 14516 29164
rect 14464 29121 14473 29155
rect 14473 29121 14507 29155
rect 14507 29121 14516 29155
rect 14464 29112 14516 29121
rect 14740 29155 14792 29164
rect 14740 29121 14749 29155
rect 14749 29121 14783 29155
rect 14783 29121 14792 29155
rect 14740 29112 14792 29121
rect 14832 29112 14884 29164
rect 15384 29180 15436 29232
rect 16856 29180 16908 29232
rect 15476 29155 15528 29164
rect 15476 29121 15485 29155
rect 15485 29121 15519 29155
rect 15519 29121 15528 29155
rect 15476 29112 15528 29121
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 16304 29155 16356 29164
rect 16304 29121 16313 29155
rect 16313 29121 16347 29155
rect 16347 29121 16356 29155
rect 16304 29112 16356 29121
rect 15384 29044 15436 29096
rect 15660 29044 15712 29096
rect 16580 29112 16632 29164
rect 17592 29248 17644 29300
rect 17960 29248 18012 29300
rect 17500 29180 17552 29232
rect 18512 29180 18564 29232
rect 22100 29248 22152 29300
rect 20444 29180 20496 29232
rect 12164 28951 12216 28960
rect 12164 28917 12173 28951
rect 12173 28917 12207 28951
rect 12207 28917 12216 28951
rect 12164 28908 12216 28917
rect 12808 28908 12860 28960
rect 15936 28951 15988 28960
rect 15936 28917 15945 28951
rect 15945 28917 15979 28951
rect 15979 28917 15988 28951
rect 15936 28908 15988 28917
rect 17132 29044 17184 29096
rect 19432 29112 19484 29164
rect 19892 29155 19944 29164
rect 19892 29121 19901 29155
rect 19901 29121 19935 29155
rect 19935 29121 19944 29155
rect 19892 29112 19944 29121
rect 19984 29155 20036 29164
rect 19984 29121 19993 29155
rect 19993 29121 20027 29155
rect 20027 29121 20036 29155
rect 19984 29112 20036 29121
rect 20352 29112 20404 29164
rect 18236 29044 18288 29096
rect 20628 29155 20680 29164
rect 20628 29121 20637 29155
rect 20637 29121 20671 29155
rect 20671 29121 20680 29155
rect 20628 29112 20680 29121
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 21180 29155 21232 29164
rect 21180 29121 21189 29155
rect 21189 29121 21223 29155
rect 21223 29121 21232 29155
rect 21180 29112 21232 29121
rect 21824 29180 21876 29232
rect 22560 29248 22612 29300
rect 23112 29248 23164 29300
rect 17316 28976 17368 29028
rect 17408 29019 17460 29028
rect 17408 28985 17417 29019
rect 17417 28985 17451 29019
rect 17451 28985 17460 29019
rect 17408 28976 17460 28985
rect 17868 28976 17920 29028
rect 18144 29019 18196 29028
rect 18144 28985 18153 29019
rect 18153 28985 18187 29019
rect 18187 28985 18196 29019
rect 18144 28976 18196 28985
rect 18420 29019 18472 29028
rect 18420 28985 18429 29019
rect 18429 28985 18463 29019
rect 18463 28985 18472 29019
rect 18420 28976 18472 28985
rect 20260 29019 20312 29028
rect 20260 28985 20269 29019
rect 20269 28985 20303 29019
rect 20303 28985 20312 29019
rect 20260 28976 20312 28985
rect 21272 28976 21324 29028
rect 19156 28908 19208 28960
rect 20628 28908 20680 28960
rect 22008 29112 22060 29164
rect 22652 29180 22704 29232
rect 24308 29248 24360 29300
rect 25136 29248 25188 29300
rect 26516 29248 26568 29300
rect 27252 29248 27304 29300
rect 28172 29248 28224 29300
rect 28356 29248 28408 29300
rect 28448 29248 28500 29300
rect 28908 29248 28960 29300
rect 22192 29044 22244 29096
rect 23296 29112 23348 29164
rect 23112 29044 23164 29096
rect 23940 29155 23992 29164
rect 23940 29121 23949 29155
rect 23949 29121 23983 29155
rect 23983 29121 23992 29155
rect 23940 29112 23992 29121
rect 24124 29180 24176 29232
rect 26056 29180 26108 29232
rect 24492 29155 24544 29164
rect 24492 29121 24501 29155
rect 24501 29121 24535 29155
rect 24535 29121 24544 29155
rect 24492 29112 24544 29121
rect 24584 29155 24636 29164
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 24768 29155 24820 29164
rect 24768 29121 24777 29155
rect 24777 29121 24811 29155
rect 24811 29121 24820 29155
rect 24768 29112 24820 29121
rect 25228 29112 25280 29164
rect 25320 29155 25372 29164
rect 25320 29121 25329 29155
rect 25329 29121 25363 29155
rect 25363 29121 25372 29155
rect 25320 29112 25372 29121
rect 26240 29112 26292 29164
rect 26332 29155 26384 29164
rect 26332 29121 26341 29155
rect 26341 29121 26375 29155
rect 26375 29121 26384 29155
rect 26332 29112 26384 29121
rect 27160 29155 27212 29164
rect 27160 29121 27164 29155
rect 27164 29121 27198 29155
rect 27198 29121 27212 29155
rect 22284 28976 22336 29028
rect 22560 28976 22612 29028
rect 23020 28976 23072 29028
rect 25044 29044 25096 29096
rect 22376 28908 22428 28960
rect 24032 28976 24084 29028
rect 27160 29112 27212 29121
rect 26976 29044 27028 29096
rect 27344 29155 27396 29164
rect 27344 29121 27353 29155
rect 27353 29121 27387 29155
rect 27387 29121 27396 29155
rect 27344 29112 27396 29121
rect 27528 29155 27580 29164
rect 27528 29121 27536 29155
rect 27536 29121 27570 29155
rect 27570 29121 27580 29155
rect 27528 29112 27580 29121
rect 27804 29223 27856 29232
rect 27804 29189 27813 29223
rect 27813 29189 27847 29223
rect 27847 29189 27856 29223
rect 27804 29180 27856 29189
rect 30196 29248 30248 29300
rect 30656 29248 30708 29300
rect 27712 29155 27764 29164
rect 27712 29121 27721 29155
rect 27721 29121 27755 29155
rect 27755 29121 27764 29155
rect 27712 29112 27764 29121
rect 26792 28976 26844 29028
rect 26884 28976 26936 29028
rect 28356 29155 28408 29164
rect 28356 29121 28365 29155
rect 28365 29121 28399 29155
rect 28399 29121 28408 29155
rect 28356 29112 28408 29121
rect 28448 29155 28500 29164
rect 28448 29121 28483 29155
rect 28483 29121 28500 29155
rect 28448 29112 28500 29121
rect 28816 29112 28868 29164
rect 28908 29155 28960 29164
rect 28908 29121 28917 29155
rect 28917 29121 28951 29155
rect 28951 29121 28960 29155
rect 28908 29112 28960 29121
rect 29552 29112 29604 29164
rect 29736 29112 29788 29164
rect 29184 29044 29236 29096
rect 29368 29087 29420 29096
rect 29368 29053 29377 29087
rect 29377 29053 29411 29087
rect 29411 29053 29420 29087
rect 30196 29112 30248 29164
rect 30380 29155 30432 29164
rect 30380 29121 30389 29155
rect 30389 29121 30423 29155
rect 30423 29121 30432 29155
rect 30380 29112 30432 29121
rect 30932 29248 30984 29300
rect 31208 29180 31260 29232
rect 31024 29112 31076 29164
rect 31668 29248 31720 29300
rect 31576 29180 31628 29232
rect 32036 29248 32088 29300
rect 32312 29248 32364 29300
rect 32772 29291 32824 29300
rect 32772 29257 32781 29291
rect 32781 29257 32815 29291
rect 32815 29257 32824 29291
rect 32772 29248 32824 29257
rect 32128 29180 32180 29232
rect 29368 29044 29420 29053
rect 31392 29044 31444 29096
rect 31576 29087 31628 29096
rect 31576 29053 31585 29087
rect 31585 29053 31619 29087
rect 31619 29053 31628 29087
rect 31576 29044 31628 29053
rect 23480 28951 23532 28960
rect 23480 28917 23489 28951
rect 23489 28917 23523 28951
rect 23523 28917 23532 28951
rect 23480 28908 23532 28917
rect 24584 28908 24636 28960
rect 24952 28908 25004 28960
rect 26240 28908 26292 28960
rect 27804 28908 27856 28960
rect 28540 28976 28592 29028
rect 29460 28976 29512 29028
rect 31944 29112 31996 29164
rect 32404 29155 32456 29164
rect 32404 29121 32413 29155
rect 32413 29121 32447 29155
rect 32447 29121 32456 29155
rect 32404 29112 32456 29121
rect 32588 29155 32640 29164
rect 32588 29121 32597 29155
rect 32597 29121 32631 29155
rect 32631 29121 32640 29155
rect 32588 29112 32640 29121
rect 33048 29248 33100 29300
rect 34520 29248 34572 29300
rect 33416 29223 33468 29232
rect 33416 29189 33425 29223
rect 33425 29189 33459 29223
rect 33459 29189 33468 29223
rect 33416 29180 33468 29189
rect 35348 29248 35400 29300
rect 36084 29180 36136 29232
rect 31944 28976 31996 29028
rect 32772 29044 32824 29096
rect 32864 29044 32916 29096
rect 33784 29155 33836 29164
rect 33784 29121 33793 29155
rect 33793 29121 33827 29155
rect 33827 29121 33836 29155
rect 33784 29112 33836 29121
rect 33324 29044 33376 29096
rect 33232 28976 33284 29028
rect 28816 28908 28868 28960
rect 29276 28908 29328 28960
rect 29552 28908 29604 28960
rect 30472 28908 30524 28960
rect 32312 28908 32364 28960
rect 33048 28908 33100 28960
rect 34152 29087 34204 29096
rect 34152 29053 34161 29087
rect 34161 29053 34195 29087
rect 34195 29053 34204 29087
rect 34152 29044 34204 29053
rect 34428 29087 34480 29096
rect 34428 29053 34437 29087
rect 34437 29053 34471 29087
rect 34471 29053 34480 29087
rect 34428 29044 34480 29053
rect 36176 29087 36228 29096
rect 36176 29053 36185 29087
rect 36185 29053 36219 29087
rect 36219 29053 36228 29087
rect 36176 29044 36228 29053
rect 34796 28908 34848 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4252 28704 4304 28756
rect 5172 28704 5224 28756
rect 5448 28704 5500 28756
rect 7656 28704 7708 28756
rect 7748 28704 7800 28756
rect 8116 28704 8168 28756
rect 8392 28704 8444 28756
rect 4528 28568 4580 28620
rect 4712 28568 4764 28620
rect 5264 28611 5316 28620
rect 5264 28577 5273 28611
rect 5273 28577 5307 28611
rect 5307 28577 5316 28611
rect 5264 28568 5316 28577
rect 5816 28611 5868 28620
rect 5816 28577 5825 28611
rect 5825 28577 5859 28611
rect 5859 28577 5868 28611
rect 5816 28568 5868 28577
rect 6092 28611 6144 28620
rect 6092 28577 6101 28611
rect 6101 28577 6135 28611
rect 6135 28577 6144 28611
rect 6092 28568 6144 28577
rect 6644 28568 6696 28620
rect 15936 28704 15988 28756
rect 16580 28704 16632 28756
rect 17224 28747 17276 28756
rect 17224 28713 17233 28747
rect 17233 28713 17267 28747
rect 17267 28713 17276 28747
rect 17224 28704 17276 28713
rect 18420 28704 18472 28756
rect 20444 28747 20496 28756
rect 20444 28713 20453 28747
rect 20453 28713 20487 28747
rect 20487 28713 20496 28747
rect 20444 28704 20496 28713
rect 10232 28679 10284 28688
rect 10232 28645 10241 28679
rect 10241 28645 10275 28679
rect 10275 28645 10284 28679
rect 10232 28636 10284 28645
rect 11244 28636 11296 28688
rect 12256 28636 12308 28688
rect 12532 28679 12584 28688
rect 12532 28645 12541 28679
rect 12541 28645 12575 28679
rect 12575 28645 12584 28679
rect 12532 28636 12584 28645
rect 14556 28636 14608 28688
rect 21732 28704 21784 28756
rect 25044 28704 25096 28756
rect 1400 28543 1452 28552
rect 1400 28509 1409 28543
rect 1409 28509 1443 28543
rect 1443 28509 1452 28543
rect 1400 28500 1452 28509
rect 1676 28475 1728 28484
rect 1676 28441 1685 28475
rect 1685 28441 1719 28475
rect 1719 28441 1728 28475
rect 1676 28432 1728 28441
rect 3148 28407 3200 28416
rect 3148 28373 3157 28407
rect 3157 28373 3191 28407
rect 3191 28373 3200 28407
rect 3148 28364 3200 28373
rect 4804 28432 4856 28484
rect 10784 28568 10836 28620
rect 11152 28611 11204 28620
rect 11152 28577 11161 28611
rect 11161 28577 11195 28611
rect 11195 28577 11204 28611
rect 11152 28568 11204 28577
rect 11520 28568 11572 28620
rect 12164 28611 12216 28620
rect 12164 28577 12173 28611
rect 12173 28577 12207 28611
rect 12207 28577 12216 28611
rect 12164 28568 12216 28577
rect 5448 28364 5500 28416
rect 8116 28543 8168 28552
rect 8116 28509 8130 28543
rect 8130 28509 8164 28543
rect 8164 28509 8168 28543
rect 8116 28500 8168 28509
rect 8300 28500 8352 28552
rect 9588 28500 9640 28552
rect 11888 28500 11940 28552
rect 12256 28543 12308 28552
rect 12256 28509 12265 28543
rect 12265 28509 12299 28543
rect 12299 28509 12308 28543
rect 12256 28500 12308 28509
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 12716 28543 12768 28552
rect 12716 28509 12720 28543
rect 12720 28509 12754 28543
rect 12754 28509 12768 28543
rect 12716 28500 12768 28509
rect 13268 28568 13320 28620
rect 14188 28568 14240 28620
rect 16856 28568 16908 28620
rect 16948 28568 17000 28620
rect 13636 28500 13688 28552
rect 9036 28432 9088 28484
rect 9680 28475 9732 28484
rect 9680 28441 9689 28475
rect 9689 28441 9723 28475
rect 9723 28441 9732 28475
rect 9680 28432 9732 28441
rect 10232 28432 10284 28484
rect 11520 28475 11572 28484
rect 11520 28441 11529 28475
rect 11529 28441 11563 28475
rect 11563 28441 11572 28475
rect 11520 28432 11572 28441
rect 11612 28432 11664 28484
rect 9772 28364 9824 28416
rect 10324 28364 10376 28416
rect 11428 28364 11480 28416
rect 12164 28364 12216 28416
rect 13728 28432 13780 28484
rect 16212 28432 16264 28484
rect 15292 28364 15344 28416
rect 16948 28475 17000 28484
rect 16948 28441 16957 28475
rect 16957 28441 16991 28475
rect 16991 28441 17000 28475
rect 16948 28432 17000 28441
rect 26240 28704 26292 28756
rect 26332 28704 26384 28756
rect 27528 28704 27580 28756
rect 28816 28747 28868 28756
rect 28816 28713 28825 28747
rect 28825 28713 28859 28747
rect 28859 28713 28868 28747
rect 28816 28704 28868 28713
rect 28908 28704 28960 28756
rect 33232 28704 33284 28756
rect 33968 28704 34020 28756
rect 17224 28500 17276 28552
rect 17776 28500 17828 28552
rect 18052 28543 18104 28552
rect 18052 28509 18061 28543
rect 18061 28509 18095 28543
rect 18095 28509 18104 28543
rect 18052 28500 18104 28509
rect 19708 28543 19760 28552
rect 19708 28509 19717 28543
rect 19717 28509 19751 28543
rect 19751 28509 19760 28543
rect 19708 28500 19760 28509
rect 17592 28432 17644 28484
rect 18880 28432 18932 28484
rect 20904 28500 20956 28552
rect 21180 28568 21232 28620
rect 21272 28568 21324 28620
rect 21456 28543 21508 28552
rect 21456 28509 21464 28543
rect 21464 28509 21498 28543
rect 21498 28509 21508 28543
rect 21456 28500 21508 28509
rect 21732 28568 21784 28620
rect 22008 28568 22060 28620
rect 20352 28432 20404 28484
rect 21180 28475 21232 28484
rect 21180 28441 21189 28475
rect 21189 28441 21223 28475
rect 21223 28441 21232 28475
rect 21180 28432 21232 28441
rect 22192 28543 22244 28552
rect 22192 28509 22196 28543
rect 22196 28509 22230 28543
rect 22230 28509 22244 28543
rect 22192 28500 22244 28509
rect 24492 28568 24544 28620
rect 25136 28568 25188 28620
rect 26884 28679 26936 28688
rect 26884 28645 26893 28679
rect 26893 28645 26927 28679
rect 26927 28645 26936 28679
rect 26884 28636 26936 28645
rect 27712 28636 27764 28688
rect 31944 28636 31996 28688
rect 26608 28568 26660 28620
rect 22560 28543 22612 28552
rect 22560 28509 22568 28543
rect 22568 28509 22602 28543
rect 22602 28509 22612 28543
rect 22560 28500 22612 28509
rect 17408 28407 17460 28416
rect 17408 28373 17417 28407
rect 17417 28373 17451 28407
rect 17451 28373 17460 28407
rect 17408 28364 17460 28373
rect 17776 28364 17828 28416
rect 21364 28364 21416 28416
rect 22192 28364 22244 28416
rect 23388 28500 23440 28552
rect 25872 28500 25924 28552
rect 26056 28500 26108 28552
rect 26240 28543 26292 28552
rect 26240 28509 26249 28543
rect 26249 28509 26283 28543
rect 26283 28509 26292 28543
rect 26240 28500 26292 28509
rect 26424 28432 26476 28484
rect 26700 28543 26752 28552
rect 26700 28509 26709 28543
rect 26709 28509 26743 28543
rect 26743 28509 26752 28543
rect 26700 28500 26752 28509
rect 26792 28543 26844 28552
rect 26792 28509 26801 28543
rect 26801 28509 26835 28543
rect 26835 28509 26844 28543
rect 26792 28500 26844 28509
rect 26976 28543 27028 28552
rect 26976 28509 26985 28543
rect 26985 28509 27019 28543
rect 27019 28509 27028 28543
rect 26976 28500 27028 28509
rect 27620 28500 27672 28552
rect 31024 28568 31076 28620
rect 29184 28500 29236 28552
rect 30472 28500 30524 28552
rect 31116 28500 31168 28552
rect 32036 28500 32088 28552
rect 32128 28543 32180 28552
rect 32128 28509 32137 28543
rect 32137 28509 32171 28543
rect 32171 28509 32180 28543
rect 32128 28500 32180 28509
rect 32680 28636 32732 28688
rect 33140 28636 33192 28688
rect 33600 28679 33652 28688
rect 33600 28645 33609 28679
rect 33609 28645 33643 28679
rect 33643 28645 33652 28679
rect 33600 28636 33652 28645
rect 22560 28364 22612 28416
rect 23112 28407 23164 28416
rect 23112 28373 23121 28407
rect 23121 28373 23155 28407
rect 23155 28373 23164 28407
rect 23112 28364 23164 28373
rect 23388 28364 23440 28416
rect 23848 28364 23900 28416
rect 25596 28407 25648 28416
rect 25596 28373 25605 28407
rect 25605 28373 25639 28407
rect 25639 28373 25648 28407
rect 25596 28364 25648 28373
rect 25780 28407 25832 28416
rect 25780 28373 25789 28407
rect 25789 28373 25823 28407
rect 25823 28373 25832 28407
rect 25780 28364 25832 28373
rect 26516 28407 26568 28416
rect 26516 28373 26525 28407
rect 26525 28373 26559 28407
rect 26559 28373 26568 28407
rect 26516 28364 26568 28373
rect 26792 28364 26844 28416
rect 28264 28432 28316 28484
rect 28356 28432 28408 28484
rect 31392 28432 31444 28484
rect 32680 28543 32732 28552
rect 32680 28509 32689 28543
rect 32689 28509 32723 28543
rect 32723 28509 32732 28543
rect 32680 28500 32732 28509
rect 34060 28611 34112 28620
rect 34060 28577 34069 28611
rect 34069 28577 34103 28611
rect 34103 28577 34112 28611
rect 34060 28568 34112 28577
rect 34612 28568 34664 28620
rect 33232 28543 33284 28552
rect 33232 28509 33241 28543
rect 33241 28509 33275 28543
rect 33275 28509 33284 28543
rect 33232 28500 33284 28509
rect 33416 28543 33468 28552
rect 33416 28509 33425 28543
rect 33425 28509 33459 28543
rect 33459 28509 33468 28543
rect 33416 28500 33468 28509
rect 33784 28543 33836 28552
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 34704 28500 34756 28552
rect 34796 28500 34848 28552
rect 34980 28543 35032 28552
rect 34980 28509 34989 28543
rect 34989 28509 35023 28543
rect 35023 28509 35032 28543
rect 34980 28500 35032 28509
rect 35072 28543 35124 28552
rect 35072 28509 35081 28543
rect 35081 28509 35115 28543
rect 35115 28509 35124 28543
rect 35072 28500 35124 28509
rect 35256 28543 35308 28552
rect 35256 28509 35265 28543
rect 35265 28509 35299 28543
rect 35299 28509 35308 28543
rect 35256 28500 35308 28509
rect 35440 28432 35492 28484
rect 27804 28407 27856 28416
rect 27804 28373 27813 28407
rect 27813 28373 27847 28407
rect 27847 28373 27856 28407
rect 27804 28364 27856 28373
rect 28816 28407 28868 28416
rect 28816 28373 28834 28407
rect 28834 28373 28868 28407
rect 28816 28364 28868 28373
rect 29184 28364 29236 28416
rect 29736 28364 29788 28416
rect 30840 28364 30892 28416
rect 31576 28364 31628 28416
rect 32036 28407 32088 28416
rect 32036 28373 32045 28407
rect 32045 28373 32079 28407
rect 32079 28373 32088 28407
rect 32036 28364 32088 28373
rect 32864 28364 32916 28416
rect 33416 28364 33468 28416
rect 34336 28364 34388 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 1676 28160 1728 28212
rect 4252 28092 4304 28144
rect 4804 28160 4856 28212
rect 2780 28067 2832 28076
rect 2780 28033 2789 28067
rect 2789 28033 2823 28067
rect 2823 28033 2832 28067
rect 2780 28024 2832 28033
rect 3148 28024 3200 28076
rect 3056 27999 3108 28008
rect 3056 27965 3065 27999
rect 3065 27965 3099 27999
rect 3099 27965 3108 27999
rect 3056 27956 3108 27965
rect 4160 28067 4212 28076
rect 4160 28033 4169 28067
rect 4169 28033 4203 28067
rect 4203 28033 4212 28067
rect 4160 28024 4212 28033
rect 4436 28067 4488 28076
rect 4436 28033 4445 28067
rect 4445 28033 4479 28067
rect 4479 28033 4488 28067
rect 4436 28024 4488 28033
rect 4620 28067 4672 28076
rect 4620 28033 4629 28067
rect 4629 28033 4663 28067
rect 4663 28033 4672 28067
rect 4620 28024 4672 28033
rect 4988 28024 5040 28076
rect 5448 28024 5500 28076
rect 5724 28024 5776 28076
rect 7656 28092 7708 28144
rect 8484 28203 8536 28212
rect 8484 28169 8493 28203
rect 8493 28169 8527 28203
rect 8527 28169 8536 28203
rect 8484 28160 8536 28169
rect 9680 28160 9732 28212
rect 5816 27888 5868 27940
rect 7564 28067 7616 28076
rect 7564 28033 7573 28067
rect 7573 28033 7607 28067
rect 7607 28033 7616 28067
rect 7564 28024 7616 28033
rect 8392 28067 8444 28076
rect 8392 28033 8401 28067
rect 8401 28033 8435 28067
rect 8435 28033 8444 28067
rect 8392 28024 8444 28033
rect 8944 28024 8996 28076
rect 10508 28067 10560 28076
rect 10508 28033 10517 28067
rect 10517 28033 10551 28067
rect 10551 28033 10560 28067
rect 10508 28024 10560 28033
rect 10692 28092 10744 28144
rect 11520 28160 11572 28212
rect 12256 28160 12308 28212
rect 17684 28160 17736 28212
rect 18052 28160 18104 28212
rect 19156 28160 19208 28212
rect 28816 28160 28868 28212
rect 29092 28203 29144 28212
rect 29092 28169 29101 28203
rect 29101 28169 29135 28203
rect 29135 28169 29144 28203
rect 29092 28160 29144 28169
rect 11060 28092 11112 28144
rect 11244 28024 11296 28076
rect 12348 28024 12400 28076
rect 14832 28092 14884 28144
rect 16672 28024 16724 28076
rect 10140 27956 10192 28008
rect 11152 27956 11204 28008
rect 11704 27956 11756 28008
rect 12808 27956 12860 28008
rect 12900 27999 12952 28008
rect 12900 27965 12909 27999
rect 12909 27965 12943 27999
rect 12943 27965 12952 27999
rect 12900 27956 12952 27965
rect 7380 27931 7432 27940
rect 7380 27897 7389 27931
rect 7389 27897 7423 27931
rect 7423 27897 7432 27931
rect 7380 27888 7432 27897
rect 11612 27888 11664 27940
rect 17224 28067 17276 28076
rect 2504 27820 2556 27872
rect 4712 27820 4764 27872
rect 11244 27820 11296 27872
rect 16396 27820 16448 27872
rect 16856 27820 16908 27872
rect 17224 28033 17232 28067
rect 17232 28033 17266 28067
rect 17266 28033 17276 28067
rect 17224 28024 17276 28033
rect 17408 28024 17460 28076
rect 18052 28024 18104 28076
rect 18328 28067 18380 28076
rect 18328 28033 18337 28067
rect 18337 28033 18371 28067
rect 18371 28033 18380 28067
rect 18328 28024 18380 28033
rect 18420 28067 18472 28076
rect 18420 28033 18429 28067
rect 18429 28033 18463 28067
rect 18463 28033 18472 28067
rect 18420 28024 18472 28033
rect 18696 27999 18748 28008
rect 18696 27965 18705 27999
rect 18705 27965 18739 27999
rect 18739 27965 18748 27999
rect 18696 27956 18748 27965
rect 18144 27888 18196 27940
rect 17960 27820 18012 27872
rect 18972 27956 19024 28008
rect 19524 27863 19576 27872
rect 19524 27829 19533 27863
rect 19533 27829 19567 27863
rect 19567 27829 19576 27863
rect 19524 27820 19576 27829
rect 19616 27820 19668 27872
rect 19892 28024 19944 28076
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 20628 27956 20680 28008
rect 21548 28024 21600 28076
rect 22744 28024 22796 28076
rect 28356 28092 28408 28144
rect 29000 28092 29052 28144
rect 29920 28135 29972 28144
rect 29920 28101 29929 28135
rect 29929 28101 29963 28135
rect 29963 28101 29972 28135
rect 29920 28092 29972 28101
rect 30012 28092 30064 28144
rect 23940 28024 23992 28076
rect 24308 28024 24360 28076
rect 23388 27956 23440 28008
rect 25596 28024 25648 28076
rect 25964 28024 26016 28076
rect 27804 28024 27856 28076
rect 28908 28067 28960 28076
rect 28908 28033 28917 28067
rect 28917 28033 28951 28067
rect 28951 28033 28960 28067
rect 28908 28024 28960 28033
rect 29184 28024 29236 28076
rect 29276 28024 29328 28076
rect 30472 28160 30524 28212
rect 31576 28160 31628 28212
rect 32128 28160 32180 28212
rect 31300 28092 31352 28144
rect 32496 28203 32548 28212
rect 32496 28169 32505 28203
rect 32505 28169 32539 28203
rect 32539 28169 32548 28203
rect 32496 28160 32548 28169
rect 33876 28160 33928 28212
rect 24584 27956 24636 28008
rect 25320 27956 25372 28008
rect 25872 27956 25924 28008
rect 23664 27888 23716 27940
rect 21548 27820 21600 27872
rect 22284 27820 22336 27872
rect 25412 27888 25464 27940
rect 26884 27956 26936 28008
rect 28356 27999 28408 28008
rect 28356 27965 28365 27999
rect 28365 27965 28399 27999
rect 28399 27965 28408 27999
rect 28356 27956 28408 27965
rect 30104 27956 30156 28008
rect 30472 27956 30524 28008
rect 29460 27888 29512 27940
rect 31484 28067 31536 28076
rect 31484 28033 31493 28067
rect 31493 28033 31527 28067
rect 31527 28033 31536 28067
rect 31484 28024 31536 28033
rect 31576 28024 31628 28076
rect 30932 27999 30984 28008
rect 30932 27965 30941 27999
rect 30941 27965 30975 27999
rect 30975 27965 30984 27999
rect 30932 27956 30984 27965
rect 24308 27820 24360 27872
rect 24860 27820 24912 27872
rect 25872 27863 25924 27872
rect 25872 27829 25881 27863
rect 25881 27829 25915 27863
rect 25915 27829 25924 27863
rect 25872 27820 25924 27829
rect 26424 27820 26476 27872
rect 28172 27863 28224 27872
rect 28172 27829 28181 27863
rect 28181 27829 28215 27863
rect 28215 27829 28224 27863
rect 28172 27820 28224 27829
rect 29092 27820 29144 27872
rect 31668 27888 31720 27940
rect 31760 27888 31812 27940
rect 30288 27820 30340 27872
rect 30564 27820 30616 27872
rect 30840 27820 30892 27872
rect 31300 27820 31352 27872
rect 32128 27956 32180 28008
rect 32496 28024 32548 28076
rect 33416 28135 33468 28144
rect 33416 28101 33422 28135
rect 33422 28101 33456 28135
rect 33456 28101 33468 28135
rect 33416 28092 33468 28101
rect 33232 27956 33284 28008
rect 33692 28067 33744 28076
rect 33692 28033 33701 28067
rect 33701 28033 33735 28067
rect 33735 28033 33744 28067
rect 34612 28067 34664 28076
rect 33692 28024 33744 28033
rect 34612 28033 34621 28067
rect 34621 28033 34655 28067
rect 34655 28033 34664 28067
rect 34612 28024 34664 28033
rect 34980 28067 35032 28076
rect 34980 28033 34989 28067
rect 34989 28033 35023 28067
rect 35023 28033 35032 28067
rect 34980 28024 35032 28033
rect 35072 28067 35124 28076
rect 35072 28033 35081 28067
rect 35081 28033 35115 28067
rect 35115 28033 35124 28067
rect 35072 28024 35124 28033
rect 35256 28067 35308 28076
rect 35256 28033 35265 28067
rect 35265 28033 35299 28067
rect 35299 28033 35308 28067
rect 35256 28024 35308 28033
rect 35532 28024 35584 28076
rect 36176 28067 36228 28076
rect 36176 28033 36185 28067
rect 36185 28033 36219 28067
rect 36219 28033 36228 28067
rect 36176 28024 36228 28033
rect 33508 27888 33560 27940
rect 32588 27820 32640 27872
rect 32680 27820 32732 27872
rect 32956 27863 33008 27872
rect 32956 27829 32965 27863
rect 32965 27829 32999 27863
rect 32999 27829 33008 27863
rect 32956 27820 33008 27829
rect 33140 27863 33192 27872
rect 33140 27829 33149 27863
rect 33149 27829 33183 27863
rect 33183 27829 33192 27863
rect 33140 27820 33192 27829
rect 33968 27820 34020 27872
rect 34336 27820 34388 27872
rect 34980 27888 35032 27940
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2780 27616 2832 27668
rect 6920 27616 6972 27668
rect 8024 27616 8076 27668
rect 8852 27616 8904 27668
rect 8944 27659 8996 27668
rect 8944 27625 8953 27659
rect 8953 27625 8987 27659
rect 8987 27625 8996 27659
rect 8944 27616 8996 27625
rect 2688 27480 2740 27532
rect 10416 27548 10468 27600
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 7196 27480 7248 27532
rect 7472 27480 7524 27532
rect 7932 27480 7984 27532
rect 4988 27455 5040 27464
rect 4988 27421 4997 27455
rect 4997 27421 5031 27455
rect 5031 27421 5040 27455
rect 4988 27412 5040 27421
rect 5448 27412 5500 27464
rect 1676 27387 1728 27396
rect 1676 27353 1685 27387
rect 1685 27353 1719 27387
rect 1719 27353 1728 27387
rect 1676 27344 1728 27353
rect 3792 27387 3844 27396
rect 3792 27353 3801 27387
rect 3801 27353 3835 27387
rect 3835 27353 3844 27387
rect 3792 27344 3844 27353
rect 4804 27387 4856 27396
rect 4804 27353 4813 27387
rect 4813 27353 4847 27387
rect 4847 27353 4856 27387
rect 4804 27344 4856 27353
rect 4068 27276 4120 27328
rect 5172 27319 5224 27328
rect 5172 27285 5181 27319
rect 5181 27285 5215 27319
rect 5215 27285 5224 27319
rect 5172 27276 5224 27285
rect 6184 27344 6236 27396
rect 6460 27344 6512 27396
rect 8116 27412 8168 27464
rect 8208 27455 8260 27464
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 8760 27480 8812 27532
rect 8576 27412 8628 27464
rect 10048 27480 10100 27532
rect 9956 27412 10008 27464
rect 10968 27480 11020 27532
rect 12900 27616 12952 27668
rect 15936 27616 15988 27668
rect 16580 27616 16632 27668
rect 17408 27616 17460 27668
rect 18420 27616 18472 27668
rect 24860 27659 24912 27668
rect 24860 27625 24869 27659
rect 24869 27625 24903 27659
rect 24903 27625 24912 27659
rect 24860 27616 24912 27625
rect 15384 27591 15436 27600
rect 15384 27557 15393 27591
rect 15393 27557 15427 27591
rect 15427 27557 15436 27591
rect 15384 27548 15436 27557
rect 10324 27412 10376 27464
rect 10416 27455 10468 27464
rect 10416 27421 10425 27455
rect 10425 27421 10459 27455
rect 10459 27421 10468 27455
rect 10416 27412 10468 27421
rect 10600 27412 10652 27464
rect 10784 27455 10836 27464
rect 10784 27421 10793 27455
rect 10793 27421 10827 27455
rect 10827 27421 10836 27455
rect 10784 27412 10836 27421
rect 11336 27412 11388 27464
rect 12532 27455 12584 27464
rect 12532 27421 12541 27455
rect 12541 27421 12575 27455
rect 12575 27421 12584 27455
rect 12532 27412 12584 27421
rect 7104 27319 7156 27328
rect 7104 27285 7113 27319
rect 7113 27285 7147 27319
rect 7147 27285 7156 27319
rect 7104 27276 7156 27285
rect 7564 27276 7616 27328
rect 8484 27276 8536 27328
rect 8852 27276 8904 27328
rect 11152 27344 11204 27396
rect 12900 27455 12952 27464
rect 12900 27421 12909 27455
rect 12909 27421 12943 27455
rect 12943 27421 12952 27455
rect 12900 27412 12952 27421
rect 13176 27412 13228 27464
rect 13268 27412 13320 27464
rect 15568 27480 15620 27532
rect 16396 27480 16448 27532
rect 17500 27548 17552 27600
rect 16580 27480 16632 27532
rect 18328 27548 18380 27600
rect 18696 27548 18748 27600
rect 14740 27412 14792 27464
rect 14924 27412 14976 27464
rect 16672 27455 16724 27464
rect 16672 27421 16676 27455
rect 16676 27421 16710 27455
rect 16710 27421 16724 27455
rect 16672 27412 16724 27421
rect 16764 27455 16816 27464
rect 16764 27421 16773 27455
rect 16773 27421 16807 27455
rect 16807 27421 16816 27455
rect 16764 27412 16816 27421
rect 16856 27455 16908 27464
rect 16856 27421 16865 27455
rect 16865 27421 16899 27455
rect 16899 27421 16908 27455
rect 16856 27412 16908 27421
rect 16948 27455 17000 27464
rect 16948 27421 16993 27455
rect 16993 27421 17000 27455
rect 16948 27412 17000 27421
rect 17316 27412 17368 27464
rect 17408 27455 17460 27464
rect 17408 27421 17417 27455
rect 17417 27421 17451 27455
rect 17451 27421 17460 27455
rect 17408 27412 17460 27421
rect 9404 27276 9456 27328
rect 10324 27319 10376 27328
rect 10324 27285 10333 27319
rect 10333 27285 10367 27319
rect 10367 27285 10376 27319
rect 10324 27276 10376 27285
rect 12716 27276 12768 27328
rect 13544 27387 13596 27396
rect 13544 27353 13553 27387
rect 13553 27353 13587 27387
rect 13587 27353 13596 27387
rect 13544 27344 13596 27353
rect 15016 27387 15068 27396
rect 15016 27353 15025 27387
rect 15025 27353 15059 27387
rect 15059 27353 15068 27387
rect 15016 27344 15068 27353
rect 15660 27344 15712 27396
rect 15844 27344 15896 27396
rect 18052 27412 18104 27464
rect 18236 27387 18288 27396
rect 18236 27353 18245 27387
rect 18245 27353 18279 27387
rect 18279 27353 18288 27387
rect 18236 27344 18288 27353
rect 19708 27480 19760 27532
rect 13636 27276 13688 27328
rect 16212 27319 16264 27328
rect 16212 27285 16237 27319
rect 16237 27285 16264 27319
rect 16212 27276 16264 27285
rect 16396 27319 16448 27328
rect 16396 27285 16405 27319
rect 16405 27285 16439 27319
rect 16439 27285 16448 27319
rect 16396 27276 16448 27285
rect 17132 27276 17184 27328
rect 17224 27319 17276 27328
rect 17224 27285 17233 27319
rect 17233 27285 17267 27319
rect 17267 27285 17276 27319
rect 17224 27276 17276 27285
rect 17868 27276 17920 27328
rect 18420 27276 18472 27328
rect 19248 27344 19300 27396
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 18880 27319 18932 27328
rect 18880 27285 18889 27319
rect 18889 27285 18923 27319
rect 18923 27285 18932 27319
rect 18880 27276 18932 27285
rect 20904 27548 20956 27600
rect 21180 27548 21232 27600
rect 21732 27548 21784 27600
rect 23112 27548 23164 27600
rect 24308 27548 24360 27600
rect 21272 27412 21324 27464
rect 21364 27455 21416 27464
rect 21364 27421 21373 27455
rect 21373 27421 21407 27455
rect 21407 27421 21416 27455
rect 21364 27412 21416 27421
rect 21456 27412 21508 27464
rect 23480 27480 23532 27532
rect 23020 27455 23072 27464
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 19708 27387 19760 27396
rect 19708 27353 19717 27387
rect 19717 27353 19751 27387
rect 19751 27353 19760 27387
rect 19708 27344 19760 27353
rect 19984 27276 20036 27328
rect 20536 27276 20588 27328
rect 21456 27319 21508 27328
rect 21456 27285 21465 27319
rect 21465 27285 21499 27319
rect 21499 27285 21508 27319
rect 21456 27276 21508 27285
rect 21732 27344 21784 27396
rect 22468 27344 22520 27396
rect 23388 27412 23440 27464
rect 24216 27480 24268 27532
rect 24032 27412 24084 27464
rect 24676 27455 24728 27464
rect 24676 27421 24685 27455
rect 24685 27421 24719 27455
rect 24719 27421 24728 27455
rect 24676 27412 24728 27421
rect 24860 27412 24912 27464
rect 25136 27412 25188 27464
rect 23756 27344 23808 27396
rect 24124 27387 24176 27396
rect 24124 27353 24133 27387
rect 24133 27353 24167 27387
rect 24167 27353 24176 27387
rect 24124 27344 24176 27353
rect 25780 27616 25832 27668
rect 26884 27659 26936 27668
rect 26884 27625 26893 27659
rect 26893 27625 26927 27659
rect 26927 27625 26936 27659
rect 26884 27616 26936 27625
rect 28172 27616 28224 27668
rect 29552 27616 29604 27668
rect 29828 27616 29880 27668
rect 30104 27616 30156 27668
rect 28264 27480 28316 27532
rect 28632 27523 28684 27532
rect 28632 27489 28641 27523
rect 28641 27489 28675 27523
rect 28675 27489 28684 27523
rect 28632 27480 28684 27489
rect 30380 27548 30432 27600
rect 30748 27616 30800 27668
rect 31852 27616 31904 27668
rect 32128 27616 32180 27668
rect 33968 27616 34020 27668
rect 25504 27455 25556 27464
rect 25504 27421 25513 27455
rect 25513 27421 25547 27455
rect 25547 27421 25556 27455
rect 25504 27412 25556 27421
rect 22284 27276 22336 27328
rect 22744 27276 22796 27328
rect 23388 27319 23440 27328
rect 23388 27285 23397 27319
rect 23397 27285 23431 27319
rect 23431 27285 23440 27319
rect 23388 27276 23440 27285
rect 23480 27276 23532 27328
rect 24768 27276 24820 27328
rect 26792 27412 26844 27464
rect 25780 27344 25832 27396
rect 26056 27387 26108 27396
rect 26056 27353 26065 27387
rect 26065 27353 26099 27387
rect 26099 27353 26108 27387
rect 26056 27344 26108 27353
rect 27068 27344 27120 27396
rect 29000 27387 29052 27396
rect 29000 27353 29009 27387
rect 29009 27353 29043 27387
rect 29043 27353 29052 27387
rect 29000 27344 29052 27353
rect 25688 27319 25740 27328
rect 25688 27285 25697 27319
rect 25697 27285 25731 27319
rect 25731 27285 25740 27319
rect 25688 27276 25740 27285
rect 26240 27319 26292 27328
rect 26240 27285 26249 27319
rect 26249 27285 26283 27319
rect 26283 27285 26292 27319
rect 26240 27276 26292 27285
rect 27436 27276 27488 27328
rect 29276 27276 29328 27328
rect 29460 27276 29512 27328
rect 30380 27455 30432 27464
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 32312 27548 32364 27600
rect 29736 27387 29788 27396
rect 29736 27353 29745 27387
rect 29745 27353 29779 27387
rect 29779 27353 29788 27387
rect 29736 27344 29788 27353
rect 29920 27387 29972 27396
rect 29920 27353 29929 27387
rect 29929 27353 29963 27387
rect 29963 27353 29972 27387
rect 29920 27344 29972 27353
rect 30288 27344 30340 27396
rect 30932 27412 30984 27464
rect 31484 27480 31536 27532
rect 31760 27412 31812 27464
rect 31852 27455 31904 27464
rect 31852 27421 31861 27455
rect 31861 27421 31895 27455
rect 31895 27421 31904 27455
rect 31852 27412 31904 27421
rect 33140 27480 33192 27532
rect 34336 27616 34388 27668
rect 34428 27616 34480 27668
rect 35348 27616 35400 27668
rect 34336 27523 34388 27532
rect 34336 27489 34345 27523
rect 34345 27489 34379 27523
rect 34379 27489 34388 27523
rect 34336 27480 34388 27489
rect 34060 27455 34112 27464
rect 34060 27421 34069 27455
rect 34069 27421 34103 27455
rect 34103 27421 34112 27455
rect 34060 27412 34112 27421
rect 31668 27387 31720 27396
rect 31668 27353 31677 27387
rect 31677 27353 31711 27387
rect 31711 27353 31720 27387
rect 31668 27344 31720 27353
rect 30564 27276 30616 27328
rect 31484 27276 31536 27328
rect 32772 27344 32824 27396
rect 35256 27455 35308 27464
rect 35256 27421 35265 27455
rect 35265 27421 35299 27455
rect 35299 27421 35308 27455
rect 35256 27412 35308 27421
rect 35348 27412 35400 27464
rect 35992 27412 36044 27464
rect 36268 27412 36320 27464
rect 36084 27344 36136 27396
rect 32036 27319 32088 27328
rect 32036 27285 32045 27319
rect 32045 27285 32079 27319
rect 32079 27285 32088 27319
rect 32036 27276 32088 27285
rect 33600 27276 33652 27328
rect 34336 27276 34388 27328
rect 35256 27276 35308 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 1676 27072 1728 27124
rect 2688 27115 2740 27124
rect 2688 27081 2697 27115
rect 2697 27081 2731 27115
rect 2731 27081 2740 27115
rect 2688 27072 2740 27081
rect 3700 27072 3752 27124
rect 4804 27072 4856 27124
rect 5816 27072 5868 27124
rect 6460 27072 6512 27124
rect 7104 27072 7156 27124
rect 7564 27115 7616 27124
rect 7564 27081 7573 27115
rect 7573 27081 7607 27115
rect 7607 27081 7616 27115
rect 7564 27072 7616 27081
rect 8024 27072 8076 27124
rect 3792 27004 3844 27056
rect 4068 27004 4120 27056
rect 3056 26868 3108 26920
rect 1400 26800 1452 26852
rect 4804 26868 4856 26920
rect 5908 26936 5960 26988
rect 6184 26936 6236 26988
rect 7104 26936 7156 26988
rect 7472 26979 7524 26988
rect 7472 26945 7481 26979
rect 7481 26945 7515 26979
rect 7515 26945 7524 26979
rect 7472 26936 7524 26945
rect 7748 26936 7800 26988
rect 6828 26911 6880 26920
rect 6828 26877 6837 26911
rect 6837 26877 6871 26911
rect 6871 26877 6880 26911
rect 6828 26868 6880 26877
rect 3700 26732 3752 26784
rect 6276 26800 6328 26852
rect 7656 26868 7708 26920
rect 8576 26936 8628 26988
rect 8760 26979 8812 26988
rect 8760 26945 8769 26979
rect 8769 26945 8803 26979
rect 8803 26945 8812 26979
rect 8760 26936 8812 26945
rect 9956 26936 10008 26988
rect 5172 26775 5224 26784
rect 5172 26741 5181 26775
rect 5181 26741 5215 26775
rect 5215 26741 5224 26775
rect 5172 26732 5224 26741
rect 8024 26732 8076 26784
rect 8852 26732 8904 26784
rect 10692 27072 10744 27124
rect 10876 27072 10928 27124
rect 10324 27004 10376 27056
rect 12716 27072 12768 27124
rect 10232 26936 10284 26988
rect 11336 27047 11388 27056
rect 11336 27013 11345 27047
rect 11345 27013 11379 27047
rect 11379 27013 11388 27047
rect 11336 27004 11388 27013
rect 10692 26936 10744 26988
rect 11152 26936 11204 26988
rect 12164 26936 12216 26988
rect 12532 26979 12584 26988
rect 12532 26945 12541 26979
rect 12541 26945 12575 26979
rect 12575 26945 12584 26979
rect 12532 26936 12584 26945
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 13912 27072 13964 27124
rect 14096 27072 14148 27124
rect 18052 27072 18104 27124
rect 21456 27072 21508 27124
rect 18512 27004 18564 27056
rect 19248 27004 19300 27056
rect 11336 26800 11388 26852
rect 12900 26800 12952 26852
rect 13268 26936 13320 26988
rect 13544 26979 13596 26988
rect 13544 26945 13554 26979
rect 13554 26945 13588 26979
rect 13588 26945 13596 26979
rect 13544 26936 13596 26945
rect 13636 26936 13688 26988
rect 13912 26979 13964 26988
rect 13912 26945 13926 26979
rect 13926 26945 13960 26979
rect 13960 26945 13964 26979
rect 13912 26936 13964 26945
rect 15752 26936 15804 26988
rect 16212 26936 16264 26988
rect 16672 26936 16724 26988
rect 17408 26936 17460 26988
rect 18328 26936 18380 26988
rect 19524 26936 19576 26988
rect 19708 26979 19760 26988
rect 19708 26945 19717 26979
rect 19717 26945 19751 26979
rect 19751 26945 19760 26979
rect 19708 26936 19760 26945
rect 19892 26936 19944 26988
rect 20444 26979 20496 26988
rect 20444 26945 20453 26979
rect 20453 26945 20487 26979
rect 20487 26945 20496 26979
rect 20444 26936 20496 26945
rect 20904 26979 20956 26988
rect 20904 26945 20913 26979
rect 20913 26945 20947 26979
rect 20947 26945 20956 26979
rect 20904 26936 20956 26945
rect 21088 26936 21140 26988
rect 14464 26868 14516 26920
rect 15016 26868 15068 26920
rect 16488 26868 16540 26920
rect 17776 26868 17828 26920
rect 11060 26732 11112 26784
rect 11244 26732 11296 26784
rect 12808 26732 12860 26784
rect 13912 26732 13964 26784
rect 14096 26775 14148 26784
rect 14096 26741 14105 26775
rect 14105 26741 14139 26775
rect 14139 26741 14148 26775
rect 14096 26732 14148 26741
rect 14372 26800 14424 26852
rect 18144 26843 18196 26852
rect 18144 26809 18153 26843
rect 18153 26809 18187 26843
rect 18187 26809 18196 26843
rect 18144 26800 18196 26809
rect 18236 26800 18288 26852
rect 20076 26843 20128 26852
rect 20076 26809 20085 26843
rect 20085 26809 20119 26843
rect 20119 26809 20128 26843
rect 20076 26800 20128 26809
rect 21548 27004 21600 27056
rect 22468 27072 22520 27124
rect 23480 27072 23532 27124
rect 24032 27115 24084 27124
rect 24032 27081 24041 27115
rect 24041 27081 24075 27115
rect 24075 27081 24084 27115
rect 24032 27072 24084 27081
rect 24216 27115 24268 27124
rect 24216 27081 24225 27115
rect 24225 27081 24259 27115
rect 24259 27081 24268 27115
rect 24216 27072 24268 27081
rect 24492 27072 24544 27124
rect 25964 27115 26016 27124
rect 25964 27081 25973 27115
rect 25973 27081 26007 27115
rect 26007 27081 26016 27115
rect 25964 27072 26016 27081
rect 28356 27072 28408 27124
rect 28908 27072 28960 27124
rect 29000 27072 29052 27124
rect 29368 27072 29420 27124
rect 22744 27004 22796 27056
rect 24584 27047 24636 27056
rect 22284 26979 22336 26988
rect 22284 26945 22293 26979
rect 22293 26945 22327 26979
rect 22327 26945 22336 26979
rect 22284 26936 22336 26945
rect 24584 27013 24593 27047
rect 24593 27013 24627 27047
rect 24627 27013 24636 27047
rect 24584 27004 24636 27013
rect 24216 26936 24268 26988
rect 24308 26936 24360 26988
rect 24676 26979 24728 26988
rect 24676 26945 24685 26979
rect 24685 26945 24719 26979
rect 24719 26945 24728 26979
rect 24676 26936 24728 26945
rect 25136 27004 25188 27056
rect 26332 27004 26384 27056
rect 26976 27004 27028 27056
rect 26792 26979 26844 26988
rect 26792 26945 26801 26979
rect 26801 26945 26835 26979
rect 26835 26945 26844 26979
rect 26792 26936 26844 26945
rect 28264 26936 28316 26988
rect 30104 27004 30156 27056
rect 30656 27004 30708 27056
rect 29000 26936 29052 26988
rect 29460 26936 29512 26988
rect 30756 26979 30808 26988
rect 30756 26945 30803 26979
rect 30803 26945 30808 26979
rect 30756 26936 30808 26945
rect 31024 26979 31076 26988
rect 31024 26945 31033 26979
rect 31033 26945 31067 26979
rect 31067 26945 31076 26979
rect 31024 26936 31076 26945
rect 22560 26911 22612 26920
rect 22560 26877 22569 26911
rect 22569 26877 22603 26911
rect 22603 26877 22612 26911
rect 22560 26868 22612 26877
rect 24032 26868 24084 26920
rect 25596 26868 25648 26920
rect 17224 26732 17276 26784
rect 17500 26732 17552 26784
rect 17776 26732 17828 26784
rect 18052 26775 18104 26784
rect 18052 26741 18061 26775
rect 18061 26741 18095 26775
rect 18095 26741 18104 26775
rect 18052 26732 18104 26741
rect 20444 26732 20496 26784
rect 21548 26732 21600 26784
rect 21732 26732 21784 26784
rect 23848 26800 23900 26852
rect 24216 26800 24268 26852
rect 25504 26800 25556 26852
rect 27436 26868 27488 26920
rect 29552 26868 29604 26920
rect 29000 26800 29052 26852
rect 30380 26800 30432 26852
rect 30656 26800 30708 26852
rect 31484 27115 31536 27124
rect 31484 27081 31493 27115
rect 31493 27081 31527 27115
rect 31527 27081 31536 27115
rect 31484 27072 31536 27081
rect 32220 27072 32272 27124
rect 32772 27072 32824 27124
rect 31576 27004 31628 27056
rect 31852 27004 31904 27056
rect 32404 27004 32456 27056
rect 32588 27004 32640 27056
rect 33140 27047 33192 27056
rect 33140 27013 33149 27047
rect 33149 27013 33183 27047
rect 33183 27013 33192 27047
rect 33140 27004 33192 27013
rect 34244 27004 34296 27056
rect 33232 26979 33284 26988
rect 33232 26945 33241 26979
rect 33241 26945 33275 26979
rect 33275 26945 33284 26979
rect 33232 26936 33284 26945
rect 33600 26936 33652 26988
rect 34336 26979 34388 26988
rect 34336 26945 34345 26979
rect 34345 26945 34379 26979
rect 34379 26945 34388 26979
rect 34336 26936 34388 26945
rect 34428 26979 34480 26988
rect 34428 26945 34437 26979
rect 34437 26945 34471 26979
rect 34471 26945 34480 26979
rect 34428 26936 34480 26945
rect 34796 26979 34848 26988
rect 34796 26945 34805 26979
rect 34805 26945 34839 26979
rect 34839 26945 34848 26979
rect 34796 26936 34848 26945
rect 35072 27004 35124 27056
rect 35348 27004 35400 27056
rect 35532 26979 35584 26988
rect 35532 26945 35541 26979
rect 35541 26945 35575 26979
rect 35575 26945 35584 26979
rect 35532 26936 35584 26945
rect 35716 26979 35768 26988
rect 35716 26945 35725 26979
rect 35725 26945 35759 26979
rect 35759 26945 35768 26979
rect 35716 26936 35768 26945
rect 36084 26936 36136 26988
rect 22652 26732 22704 26784
rect 26240 26732 26292 26784
rect 30104 26775 30156 26784
rect 30104 26741 30113 26775
rect 30113 26741 30147 26775
rect 30147 26741 30156 26775
rect 30104 26732 30156 26741
rect 30288 26732 30340 26784
rect 32404 26732 32456 26784
rect 32864 26732 32916 26784
rect 33968 26800 34020 26852
rect 34060 26800 34112 26852
rect 34796 26800 34848 26852
rect 33048 26732 33100 26784
rect 35992 26732 36044 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4804 26571 4856 26580
rect 4804 26537 4813 26571
rect 4813 26537 4847 26571
rect 4847 26537 4856 26571
rect 4804 26528 4856 26537
rect 3792 26392 3844 26444
rect 6276 26528 6328 26580
rect 7748 26528 7800 26580
rect 8392 26528 8444 26580
rect 9864 26528 9916 26580
rect 9956 26528 10008 26580
rect 14372 26528 14424 26580
rect 5448 26460 5500 26512
rect 6000 26392 6052 26444
rect 5172 26299 5224 26308
rect 5172 26265 5181 26299
rect 5181 26265 5215 26299
rect 5215 26265 5224 26299
rect 5172 26256 5224 26265
rect 5724 26256 5776 26308
rect 5908 26367 5960 26376
rect 5908 26333 5917 26367
rect 5917 26333 5951 26367
rect 5951 26333 5960 26367
rect 5908 26324 5960 26333
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 9220 26460 9272 26512
rect 9404 26460 9456 26512
rect 13268 26460 13320 26512
rect 7656 26392 7708 26444
rect 8024 26392 8076 26444
rect 7932 26367 7984 26376
rect 7932 26333 7941 26367
rect 7941 26333 7975 26367
rect 7975 26333 7984 26367
rect 7932 26324 7984 26333
rect 8300 26392 8352 26444
rect 14280 26460 14332 26512
rect 14924 26528 14976 26580
rect 17776 26571 17828 26580
rect 17776 26537 17785 26571
rect 17785 26537 17819 26571
rect 17819 26537 17828 26571
rect 17776 26528 17828 26537
rect 20996 26528 21048 26580
rect 21916 26571 21968 26580
rect 21916 26537 21925 26571
rect 21925 26537 21959 26571
rect 21959 26537 21968 26571
rect 21916 26528 21968 26537
rect 26148 26528 26200 26580
rect 26608 26528 26660 26580
rect 26976 26571 27028 26580
rect 26976 26537 26985 26571
rect 26985 26537 27019 26571
rect 27019 26537 27028 26571
rect 26976 26528 27028 26537
rect 27896 26528 27948 26580
rect 29460 26528 29512 26580
rect 29736 26528 29788 26580
rect 30472 26528 30524 26580
rect 32772 26528 32824 26580
rect 33600 26528 33652 26580
rect 33876 26528 33928 26580
rect 8576 26367 8628 26376
rect 4160 26188 4212 26240
rect 5816 26188 5868 26240
rect 6736 26299 6788 26308
rect 6736 26265 6745 26299
rect 6745 26265 6779 26299
rect 6779 26265 6788 26299
rect 6736 26256 6788 26265
rect 8576 26333 8584 26367
rect 8584 26333 8618 26367
rect 8618 26333 8628 26367
rect 8576 26324 8628 26333
rect 8944 26256 8996 26308
rect 9772 26324 9824 26376
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 10416 26324 10468 26376
rect 10784 26324 10836 26376
rect 12532 26367 12584 26376
rect 12532 26333 12541 26367
rect 12541 26333 12575 26367
rect 12575 26333 12584 26367
rect 12532 26324 12584 26333
rect 12716 26367 12768 26376
rect 12716 26333 12725 26367
rect 12725 26333 12759 26367
rect 12759 26333 12768 26367
rect 12716 26324 12768 26333
rect 7012 26188 7064 26240
rect 8852 26188 8904 26240
rect 9312 26299 9364 26308
rect 9312 26265 9321 26299
rect 9321 26265 9355 26299
rect 9355 26265 9364 26299
rect 9312 26256 9364 26265
rect 9956 26256 10008 26308
rect 11060 26256 11112 26308
rect 12624 26256 12676 26308
rect 12900 26367 12952 26376
rect 12900 26333 12909 26367
rect 12909 26333 12943 26367
rect 12943 26333 12952 26367
rect 12900 26324 12952 26333
rect 13084 26367 13136 26376
rect 13084 26333 13093 26367
rect 13093 26333 13127 26367
rect 13127 26333 13136 26367
rect 13084 26324 13136 26333
rect 13268 26324 13320 26376
rect 13912 26367 13964 26376
rect 13912 26333 13921 26367
rect 13921 26333 13955 26367
rect 13955 26333 13964 26367
rect 13912 26324 13964 26333
rect 14096 26324 14148 26376
rect 14372 26367 14424 26376
rect 14372 26333 14379 26367
rect 14379 26333 14424 26367
rect 14372 26324 14424 26333
rect 14924 26435 14976 26444
rect 14924 26401 14933 26435
rect 14933 26401 14967 26435
rect 14967 26401 14976 26435
rect 14924 26392 14976 26401
rect 15844 26392 15896 26444
rect 14648 26367 14700 26376
rect 14648 26333 14662 26367
rect 14662 26333 14696 26367
rect 14696 26333 14700 26367
rect 14648 26324 14700 26333
rect 9772 26188 9824 26240
rect 10600 26188 10652 26240
rect 11152 26188 11204 26240
rect 13268 26188 13320 26240
rect 14004 26256 14056 26308
rect 14924 26256 14976 26308
rect 15568 26324 15620 26376
rect 16672 26324 16724 26376
rect 17132 26324 17184 26376
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 17408 26367 17460 26376
rect 17408 26333 17412 26367
rect 17412 26333 17446 26367
rect 17446 26333 17460 26367
rect 17408 26324 17460 26333
rect 17592 26392 17644 26444
rect 21180 26460 21232 26512
rect 20076 26392 20128 26444
rect 21732 26435 21784 26444
rect 21732 26401 21741 26435
rect 21741 26401 21775 26435
rect 21775 26401 21784 26435
rect 21732 26392 21784 26401
rect 21824 26392 21876 26444
rect 20168 26324 20220 26376
rect 22100 26324 22152 26376
rect 22468 26367 22520 26376
rect 22468 26333 22477 26367
rect 22477 26333 22511 26367
rect 22511 26333 22520 26367
rect 22468 26324 22520 26333
rect 17684 26256 17736 26308
rect 18144 26256 18196 26308
rect 20444 26256 20496 26308
rect 21088 26299 21140 26308
rect 21088 26265 21113 26299
rect 21113 26265 21140 26299
rect 21088 26256 21140 26265
rect 21456 26256 21508 26308
rect 24308 26460 24360 26512
rect 26332 26435 26384 26444
rect 26332 26401 26341 26435
rect 26341 26401 26375 26435
rect 26375 26401 26384 26435
rect 26332 26392 26384 26401
rect 22928 26324 22980 26376
rect 25872 26367 25924 26376
rect 25872 26333 25881 26367
rect 25881 26333 25915 26367
rect 25915 26333 25924 26367
rect 25872 26324 25924 26333
rect 26424 26324 26476 26376
rect 26884 26392 26936 26444
rect 29828 26460 29880 26512
rect 32128 26460 32180 26512
rect 27436 26367 27488 26376
rect 27436 26333 27445 26367
rect 27445 26333 27479 26367
rect 27479 26333 27488 26367
rect 27436 26324 27488 26333
rect 24768 26256 24820 26308
rect 26608 26256 26660 26308
rect 26700 26256 26752 26308
rect 27896 26367 27948 26376
rect 27896 26333 27905 26367
rect 27905 26333 27939 26367
rect 27939 26333 27948 26367
rect 27896 26324 27948 26333
rect 28356 26367 28408 26376
rect 28356 26333 28365 26367
rect 28365 26333 28399 26367
rect 28399 26333 28408 26367
rect 28356 26324 28408 26333
rect 16304 26188 16356 26240
rect 16764 26188 16816 26240
rect 17316 26188 17368 26240
rect 18880 26188 18932 26240
rect 24676 26188 24728 26240
rect 28080 26256 28132 26308
rect 28264 26299 28316 26308
rect 28264 26265 28273 26299
rect 28273 26265 28307 26299
rect 28307 26265 28316 26299
rect 28264 26256 28316 26265
rect 29920 26392 29972 26444
rect 30196 26392 30248 26444
rect 30380 26392 30432 26444
rect 34060 26460 34112 26512
rect 31760 26324 31812 26376
rect 33048 26392 33100 26444
rect 33140 26392 33192 26444
rect 34336 26528 34388 26580
rect 34520 26460 34572 26512
rect 32864 26367 32916 26376
rect 32864 26333 32873 26367
rect 32873 26333 32907 26367
rect 32907 26333 32916 26367
rect 32864 26324 32916 26333
rect 34796 26392 34848 26444
rect 35164 26392 35216 26444
rect 31024 26256 31076 26308
rect 32128 26256 32180 26308
rect 33324 26367 33376 26376
rect 33324 26333 33333 26367
rect 33333 26333 33367 26367
rect 33367 26333 33376 26367
rect 33324 26324 33376 26333
rect 33600 26367 33652 26376
rect 33600 26333 33609 26367
rect 33609 26333 33643 26367
rect 33643 26333 33652 26367
rect 33600 26324 33652 26333
rect 33876 26367 33928 26376
rect 33876 26333 33885 26367
rect 33885 26333 33919 26367
rect 33919 26333 33928 26367
rect 33876 26324 33928 26333
rect 34060 26367 34112 26376
rect 34060 26333 34069 26367
rect 34069 26333 34103 26367
rect 34103 26333 34112 26367
rect 34060 26324 34112 26333
rect 34244 26324 34296 26376
rect 35256 26367 35308 26376
rect 35256 26333 35265 26367
rect 35265 26333 35299 26367
rect 35299 26333 35308 26367
rect 35256 26324 35308 26333
rect 34612 26256 34664 26308
rect 35624 26256 35676 26308
rect 36176 26367 36228 26376
rect 36176 26333 36185 26367
rect 36185 26333 36219 26367
rect 36219 26333 36228 26367
rect 36176 26324 36228 26333
rect 36360 26256 36412 26308
rect 27988 26231 28040 26240
rect 27988 26197 27997 26231
rect 27997 26197 28031 26231
rect 28031 26197 28040 26231
rect 27988 26188 28040 26197
rect 28908 26188 28960 26240
rect 30748 26231 30800 26240
rect 30748 26197 30757 26231
rect 30757 26197 30791 26231
rect 30791 26197 30800 26231
rect 30748 26188 30800 26197
rect 31944 26188 31996 26240
rect 32404 26188 32456 26240
rect 32496 26188 32548 26240
rect 35072 26188 35124 26240
rect 35348 26188 35400 26240
rect 35532 26188 35584 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 3148 26027 3200 26036
rect 3148 25993 3157 26027
rect 3157 25993 3191 26027
rect 3191 25993 3200 26027
rect 3148 25984 3200 25993
rect 6184 25984 6236 26036
rect 2964 25916 3016 25968
rect 3976 25916 4028 25968
rect 6000 25959 6052 25968
rect 6000 25925 6009 25959
rect 6009 25925 6043 25959
rect 6043 25925 6052 25959
rect 6000 25916 6052 25925
rect 6736 25916 6788 25968
rect 8208 26027 8260 26036
rect 8208 25993 8217 26027
rect 8217 25993 8251 26027
rect 8251 25993 8260 26027
rect 8208 25984 8260 25993
rect 9772 26027 9824 26036
rect 9772 25993 9781 26027
rect 9781 25993 9815 26027
rect 9815 25993 9824 26027
rect 9772 25984 9824 25993
rect 10324 25984 10376 26036
rect 1400 25823 1452 25832
rect 1400 25789 1409 25823
rect 1409 25789 1443 25823
rect 1443 25789 1452 25823
rect 1400 25780 1452 25789
rect 2228 25780 2280 25832
rect 2412 25780 2464 25832
rect 3884 25780 3936 25832
rect 4068 25780 4120 25832
rect 8300 25848 8352 25900
rect 4712 25780 4764 25832
rect 6644 25823 6696 25832
rect 6644 25789 6653 25823
rect 6653 25789 6687 25823
rect 6687 25789 6696 25823
rect 6644 25780 6696 25789
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 9312 25780 9364 25832
rect 8668 25712 8720 25764
rect 1400 25644 1452 25696
rect 2412 25644 2464 25696
rect 7196 25644 7248 25696
rect 7932 25644 7984 25696
rect 9312 25687 9364 25696
rect 9312 25653 9321 25687
rect 9321 25653 9355 25687
rect 9355 25653 9364 25687
rect 9312 25644 9364 25653
rect 10232 25916 10284 25968
rect 11244 25984 11296 26036
rect 11888 25984 11940 26036
rect 9956 25848 10008 25900
rect 10416 25780 10468 25832
rect 10784 25959 10836 25968
rect 10784 25925 10793 25959
rect 10793 25925 10827 25959
rect 10827 25925 10836 25959
rect 10784 25916 10836 25925
rect 10876 25848 10928 25900
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 11152 25823 11204 25832
rect 11152 25789 11161 25823
rect 11161 25789 11195 25823
rect 11195 25789 11204 25823
rect 11152 25780 11204 25789
rect 10140 25712 10192 25764
rect 10692 25712 10744 25764
rect 12072 25891 12124 25900
rect 12072 25857 12081 25891
rect 12081 25857 12115 25891
rect 12115 25857 12124 25891
rect 12072 25848 12124 25857
rect 12164 25848 12216 25900
rect 12624 25916 12676 25968
rect 11888 25823 11940 25832
rect 11888 25789 11897 25823
rect 11897 25789 11931 25823
rect 11931 25789 11940 25823
rect 11888 25780 11940 25789
rect 12532 25891 12584 25900
rect 12532 25857 12542 25891
rect 12542 25857 12576 25891
rect 12576 25857 12584 25891
rect 12532 25848 12584 25857
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 12992 25848 13044 25900
rect 13636 25848 13688 25900
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 15936 25891 15988 25900
rect 15936 25857 15945 25891
rect 15945 25857 15979 25891
rect 15979 25857 15988 25891
rect 15936 25848 15988 25857
rect 16120 25848 16172 25900
rect 16580 25984 16632 26036
rect 16304 25891 16356 25900
rect 16304 25857 16313 25891
rect 16313 25857 16347 25891
rect 16347 25857 16356 25891
rect 16304 25848 16356 25857
rect 17776 25916 17828 25968
rect 18236 25959 18288 25968
rect 17408 25848 17460 25900
rect 17592 25848 17644 25900
rect 17868 25848 17920 25900
rect 18236 25925 18270 25959
rect 18270 25925 18288 25959
rect 18236 25916 18288 25925
rect 18788 25848 18840 25900
rect 12624 25780 12676 25832
rect 12164 25712 12216 25764
rect 12716 25712 12768 25764
rect 13544 25712 13596 25764
rect 12532 25644 12584 25696
rect 13360 25644 13412 25696
rect 14648 25644 14700 25696
rect 15108 25644 15160 25696
rect 17040 25823 17092 25832
rect 17040 25789 17049 25823
rect 17049 25789 17083 25823
rect 17083 25789 17092 25823
rect 17040 25780 17092 25789
rect 17776 25780 17828 25832
rect 18144 25780 18196 25832
rect 16396 25712 16448 25764
rect 19524 25984 19576 26036
rect 20352 25984 20404 26036
rect 22100 25984 22152 26036
rect 23296 25984 23348 26036
rect 23572 26027 23624 26036
rect 23572 25993 23581 26027
rect 23581 25993 23615 26027
rect 23615 25993 23624 26027
rect 23572 25984 23624 25993
rect 23848 25984 23900 26036
rect 19064 25848 19116 25900
rect 19708 25848 19760 25900
rect 23204 25925 23213 25934
rect 23213 25925 23247 25934
rect 23247 25925 23256 25934
rect 23204 25882 23256 25925
rect 25136 25984 25188 26036
rect 25780 25984 25832 26036
rect 32036 25984 32088 26036
rect 32128 25984 32180 26036
rect 32496 25984 32548 26036
rect 23848 25891 23900 25900
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 19432 25823 19484 25832
rect 19432 25789 19441 25823
rect 19441 25789 19475 25823
rect 19475 25789 19484 25823
rect 19432 25780 19484 25789
rect 19984 25823 20036 25832
rect 19984 25789 19993 25823
rect 19993 25789 20027 25823
rect 20027 25789 20036 25823
rect 19984 25780 20036 25789
rect 24308 25891 24360 25900
rect 24308 25857 24322 25891
rect 24322 25857 24356 25891
rect 24356 25857 24360 25891
rect 24308 25848 24360 25857
rect 24492 25848 24544 25900
rect 17868 25644 17920 25696
rect 19156 25712 19208 25764
rect 21548 25712 21600 25764
rect 23756 25712 23808 25764
rect 24584 25780 24636 25832
rect 24492 25755 24544 25764
rect 24492 25721 24501 25755
rect 24501 25721 24535 25755
rect 24535 25721 24544 25755
rect 24492 25712 24544 25721
rect 24768 25712 24820 25764
rect 25320 25848 25372 25900
rect 25688 25848 25740 25900
rect 25964 25848 26016 25900
rect 26424 25916 26476 25968
rect 26884 25916 26936 25968
rect 26240 25891 26292 25900
rect 26240 25857 26249 25891
rect 26249 25857 26283 25891
rect 26283 25857 26292 25891
rect 26240 25848 26292 25857
rect 25412 25780 25464 25832
rect 26976 25848 27028 25900
rect 25136 25712 25188 25764
rect 27620 25916 27672 25968
rect 27988 25916 28040 25968
rect 29276 25916 29328 25968
rect 29460 25916 29512 25968
rect 27528 25891 27580 25900
rect 27528 25857 27537 25891
rect 27537 25857 27571 25891
rect 27571 25857 27580 25891
rect 27528 25848 27580 25857
rect 28724 25848 28776 25900
rect 30196 25916 30248 25968
rect 29000 25780 29052 25832
rect 28172 25712 28224 25764
rect 29920 25848 29972 25900
rect 30012 25848 30064 25900
rect 32312 25916 32364 25968
rect 31760 25891 31812 25900
rect 31760 25857 31769 25891
rect 31769 25857 31803 25891
rect 31803 25857 31812 25891
rect 31760 25848 31812 25857
rect 31944 25891 31996 25900
rect 31944 25857 31953 25891
rect 31953 25857 31987 25891
rect 31987 25857 31996 25891
rect 31944 25848 31996 25857
rect 32128 25848 32180 25900
rect 33232 25984 33284 26036
rect 33600 25984 33652 26036
rect 34520 25984 34572 26036
rect 33968 25959 34020 25968
rect 33968 25925 33977 25959
rect 33977 25925 34011 25959
rect 34011 25925 34020 25959
rect 33968 25916 34020 25925
rect 33140 25891 33192 25900
rect 33140 25857 33149 25891
rect 33149 25857 33183 25891
rect 33183 25857 33192 25891
rect 33140 25848 33192 25857
rect 33324 25891 33376 25900
rect 33324 25857 33333 25891
rect 33333 25857 33367 25891
rect 33367 25857 33376 25891
rect 33324 25848 33376 25857
rect 34060 25848 34112 25900
rect 34244 25848 34296 25900
rect 34520 25891 34572 25900
rect 34520 25857 34529 25891
rect 34529 25857 34563 25891
rect 34563 25857 34572 25891
rect 34520 25848 34572 25857
rect 35072 25916 35124 25968
rect 35624 25916 35676 25968
rect 35256 25848 35308 25900
rect 35716 25848 35768 25900
rect 31024 25780 31076 25832
rect 33048 25823 33100 25832
rect 33048 25789 33057 25823
rect 33057 25789 33091 25823
rect 33091 25789 33100 25823
rect 33048 25780 33100 25789
rect 33600 25780 33652 25832
rect 18696 25687 18748 25696
rect 18696 25653 18705 25687
rect 18705 25653 18739 25687
rect 18739 25653 18748 25687
rect 18696 25644 18748 25653
rect 19800 25644 19852 25696
rect 23296 25644 23348 25696
rect 23388 25687 23440 25696
rect 23388 25653 23397 25687
rect 23397 25653 23431 25687
rect 23431 25653 23440 25687
rect 23388 25644 23440 25653
rect 23664 25644 23716 25696
rect 27344 25644 27396 25696
rect 29276 25687 29328 25696
rect 29276 25653 29285 25687
rect 29285 25653 29319 25687
rect 29319 25653 29328 25687
rect 29276 25644 29328 25653
rect 29460 25755 29512 25764
rect 29460 25721 29469 25755
rect 29469 25721 29503 25755
rect 29503 25721 29512 25755
rect 29460 25712 29512 25721
rect 29552 25712 29604 25764
rect 32496 25712 32548 25764
rect 32680 25712 32732 25764
rect 32864 25712 32916 25764
rect 33416 25712 33468 25764
rect 33968 25780 34020 25832
rect 35348 25780 35400 25832
rect 29736 25644 29788 25696
rect 29920 25687 29972 25696
rect 29920 25653 29929 25687
rect 29929 25653 29963 25687
rect 29963 25653 29972 25687
rect 29920 25644 29972 25653
rect 30748 25644 30800 25696
rect 31852 25644 31904 25696
rect 32220 25644 32272 25696
rect 34428 25712 34480 25764
rect 35164 25712 35216 25764
rect 35532 25712 35584 25764
rect 34060 25687 34112 25696
rect 34060 25653 34069 25687
rect 34069 25653 34103 25687
rect 34103 25653 34112 25687
rect 34060 25644 34112 25653
rect 34244 25687 34296 25696
rect 34244 25653 34253 25687
rect 34253 25653 34287 25687
rect 34287 25653 34296 25687
rect 34244 25644 34296 25653
rect 34796 25644 34848 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2228 25483 2280 25492
rect 2228 25449 2237 25483
rect 2237 25449 2271 25483
rect 2271 25449 2280 25483
rect 2228 25440 2280 25449
rect 3884 25483 3936 25492
rect 3884 25449 3893 25483
rect 3893 25449 3927 25483
rect 3927 25449 3936 25483
rect 3884 25440 3936 25449
rect 6644 25440 6696 25492
rect 2412 25100 2464 25152
rect 3056 25304 3108 25356
rect 3792 25304 3844 25356
rect 6184 25304 6236 25356
rect 6276 25347 6328 25356
rect 6276 25313 6285 25347
rect 6285 25313 6319 25347
rect 6319 25313 6328 25347
rect 6276 25304 6328 25313
rect 9312 25440 9364 25492
rect 9864 25440 9916 25492
rect 10600 25440 10652 25492
rect 13636 25440 13688 25492
rect 15200 25440 15252 25492
rect 15476 25440 15528 25492
rect 17500 25440 17552 25492
rect 17868 25440 17920 25492
rect 3148 25236 3200 25288
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 6000 25279 6052 25288
rect 6000 25245 6009 25279
rect 6009 25245 6043 25279
rect 6043 25245 6052 25279
rect 6000 25236 6052 25245
rect 7012 25236 7064 25288
rect 7656 25304 7708 25356
rect 8208 25304 8260 25356
rect 8484 25415 8536 25424
rect 8484 25381 8493 25415
rect 8493 25381 8527 25415
rect 8527 25381 8536 25415
rect 8484 25372 8536 25381
rect 8944 25415 8996 25424
rect 8944 25381 8953 25415
rect 8953 25381 8987 25415
rect 8987 25381 8996 25415
rect 8944 25372 8996 25381
rect 11612 25372 11664 25424
rect 5816 25211 5868 25220
rect 5816 25177 5825 25211
rect 5825 25177 5859 25211
rect 5859 25177 5868 25211
rect 5816 25168 5868 25177
rect 5908 25168 5960 25220
rect 8024 25211 8076 25220
rect 8024 25177 8041 25211
rect 8041 25177 8076 25211
rect 3976 25100 4028 25152
rect 5632 25100 5684 25152
rect 6460 25100 6512 25152
rect 8024 25168 8076 25177
rect 8116 25211 8168 25220
rect 8116 25177 8125 25211
rect 8125 25177 8159 25211
rect 8159 25177 8168 25211
rect 8116 25168 8168 25177
rect 9128 25279 9180 25288
rect 9128 25245 9137 25279
rect 9137 25245 9171 25279
rect 9171 25245 9180 25279
rect 9128 25236 9180 25245
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 12532 25304 12584 25356
rect 9956 25279 10008 25288
rect 9956 25245 9965 25279
rect 9965 25245 9999 25279
rect 9999 25245 10008 25279
rect 9956 25236 10008 25245
rect 10232 25236 10284 25288
rect 10140 25168 10192 25220
rect 11612 25236 11664 25288
rect 11888 25279 11940 25288
rect 11888 25245 11897 25279
rect 11897 25245 11931 25279
rect 11931 25245 11940 25279
rect 11888 25236 11940 25245
rect 12072 25279 12124 25288
rect 12072 25245 12081 25279
rect 12081 25245 12115 25279
rect 12115 25245 12124 25279
rect 12072 25236 12124 25245
rect 12992 25236 13044 25288
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 7748 25143 7800 25152
rect 7748 25109 7757 25143
rect 7757 25109 7791 25143
rect 7791 25109 7800 25143
rect 7748 25100 7800 25109
rect 7840 25100 7892 25152
rect 10600 25100 10652 25152
rect 10784 25100 10836 25152
rect 11152 25168 11204 25220
rect 12716 25168 12768 25220
rect 13360 25279 13412 25288
rect 13360 25245 13369 25279
rect 13369 25245 13403 25279
rect 13403 25245 13412 25279
rect 13360 25236 13412 25245
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 14648 25279 14700 25288
rect 14648 25245 14657 25279
rect 14657 25245 14691 25279
rect 14691 25245 14700 25279
rect 14648 25236 14700 25245
rect 15384 25372 15436 25424
rect 16580 25372 16632 25424
rect 17040 25304 17092 25356
rect 13728 25168 13780 25220
rect 11796 25100 11848 25152
rect 12440 25100 12492 25152
rect 12808 25100 12860 25152
rect 13360 25100 13412 25152
rect 15476 25279 15528 25288
rect 15476 25245 15485 25279
rect 15485 25245 15519 25279
rect 15519 25245 15528 25279
rect 15476 25236 15528 25245
rect 16764 25236 16816 25288
rect 18236 25372 18288 25424
rect 18972 25372 19024 25424
rect 19432 25440 19484 25492
rect 23848 25440 23900 25492
rect 24400 25440 24452 25492
rect 24676 25440 24728 25492
rect 21364 25372 21416 25424
rect 22192 25372 22244 25424
rect 22744 25372 22796 25424
rect 18512 25279 18564 25288
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 19524 25236 19576 25288
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 19984 25236 20036 25288
rect 20444 25236 20496 25288
rect 16856 25211 16908 25220
rect 16856 25177 16865 25211
rect 16865 25177 16899 25211
rect 16899 25177 16908 25211
rect 16856 25168 16908 25177
rect 18144 25168 18196 25220
rect 21364 25236 21416 25288
rect 23020 25304 23072 25356
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 24768 25372 24820 25424
rect 23664 25347 23716 25356
rect 23664 25313 23673 25347
rect 23673 25313 23707 25347
rect 23707 25313 23716 25347
rect 23664 25304 23716 25313
rect 28172 25440 28224 25492
rect 29736 25483 29788 25492
rect 29736 25449 29745 25483
rect 29745 25449 29779 25483
rect 29779 25449 29788 25483
rect 29736 25440 29788 25449
rect 33048 25440 33100 25492
rect 33232 25440 33284 25492
rect 34244 25440 34296 25492
rect 34336 25440 34388 25492
rect 25780 25415 25832 25424
rect 25780 25381 25789 25415
rect 25789 25381 25823 25415
rect 25823 25381 25832 25415
rect 25780 25372 25832 25381
rect 28908 25372 28960 25424
rect 29920 25372 29972 25424
rect 23480 25236 23532 25288
rect 24492 25236 24544 25288
rect 24860 25236 24912 25288
rect 25320 25236 25372 25288
rect 25964 25236 26016 25288
rect 22928 25211 22980 25220
rect 22928 25177 22937 25211
rect 22937 25177 22971 25211
rect 22971 25177 22980 25211
rect 22928 25168 22980 25177
rect 25412 25168 25464 25220
rect 26424 25236 26476 25288
rect 27344 25347 27396 25356
rect 27344 25313 27353 25347
rect 27353 25313 27387 25347
rect 27387 25313 27396 25347
rect 27344 25304 27396 25313
rect 28632 25304 28684 25356
rect 29000 25304 29052 25356
rect 27804 25236 27856 25288
rect 15660 25143 15712 25152
rect 15660 25109 15669 25143
rect 15669 25109 15703 25143
rect 15703 25109 15712 25143
rect 15660 25100 15712 25109
rect 17408 25100 17460 25152
rect 17500 25100 17552 25152
rect 23204 25143 23256 25152
rect 23204 25109 23213 25143
rect 23213 25109 23247 25143
rect 23247 25109 23256 25143
rect 23204 25100 23256 25109
rect 23388 25100 23440 25152
rect 29000 25168 29052 25220
rect 31024 25236 31076 25288
rect 31208 25279 31260 25288
rect 31208 25245 31217 25279
rect 31217 25245 31251 25279
rect 31251 25245 31260 25279
rect 31208 25236 31260 25245
rect 31300 25279 31352 25288
rect 31300 25245 31309 25279
rect 31309 25245 31343 25279
rect 31343 25245 31352 25279
rect 31300 25236 31352 25245
rect 32036 25347 32088 25356
rect 32036 25313 32045 25347
rect 32045 25313 32079 25347
rect 32079 25313 32088 25347
rect 32036 25304 32088 25313
rect 32220 25372 32272 25424
rect 33416 25372 33468 25424
rect 33692 25372 33744 25424
rect 34520 25372 34572 25424
rect 35348 25440 35400 25492
rect 35532 25483 35584 25492
rect 35532 25449 35541 25483
rect 35541 25449 35575 25483
rect 35575 25449 35584 25483
rect 35532 25440 35584 25449
rect 36544 25440 36596 25492
rect 35716 25372 35768 25424
rect 35808 25372 35860 25424
rect 32404 25304 32456 25356
rect 31760 25236 31812 25288
rect 31852 25279 31904 25288
rect 31852 25245 31861 25279
rect 31861 25245 31895 25279
rect 31895 25245 31904 25279
rect 31852 25236 31904 25245
rect 32496 25279 32548 25288
rect 32496 25245 32505 25279
rect 32505 25245 32539 25279
rect 32539 25245 32548 25279
rect 32496 25236 32548 25245
rect 26056 25100 26108 25152
rect 26792 25100 26844 25152
rect 27068 25100 27120 25152
rect 28356 25100 28408 25152
rect 28632 25100 28684 25152
rect 30748 25143 30800 25152
rect 30748 25109 30757 25143
rect 30757 25109 30791 25143
rect 30791 25109 30800 25143
rect 30748 25100 30800 25109
rect 32404 25168 32456 25220
rect 34060 25304 34112 25356
rect 33692 25279 33744 25288
rect 33692 25245 33701 25279
rect 33701 25245 33735 25279
rect 33735 25245 33744 25279
rect 33692 25236 33744 25245
rect 33784 25279 33836 25288
rect 33784 25245 33793 25279
rect 33793 25245 33827 25279
rect 33827 25245 33836 25279
rect 33784 25236 33836 25245
rect 34796 25236 34848 25288
rect 33876 25168 33928 25220
rect 35256 25279 35308 25288
rect 35256 25245 35265 25279
rect 35265 25245 35299 25279
rect 35299 25245 35308 25279
rect 35256 25236 35308 25245
rect 35624 25236 35676 25288
rect 35716 25279 35768 25288
rect 35716 25245 35725 25279
rect 35725 25245 35759 25279
rect 35759 25245 35768 25279
rect 35716 25236 35768 25245
rect 35992 25236 36044 25288
rect 35348 25168 35400 25220
rect 32956 25100 33008 25152
rect 33232 25143 33284 25152
rect 33232 25109 33241 25143
rect 33241 25109 33275 25143
rect 33275 25109 33284 25143
rect 33232 25100 33284 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 2964 24828 3016 24880
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 3608 24871 3660 24880
rect 3608 24837 3617 24871
rect 3617 24837 3651 24871
rect 3651 24837 3660 24871
rect 3608 24828 3660 24837
rect 2780 24624 2832 24676
rect 3792 24735 3844 24744
rect 3792 24701 3801 24735
rect 3801 24701 3835 24735
rect 3835 24701 3844 24735
rect 3792 24692 3844 24701
rect 4068 24760 4120 24812
rect 4712 24828 4764 24880
rect 5908 24939 5960 24948
rect 5908 24905 5917 24939
rect 5917 24905 5951 24939
rect 5951 24905 5960 24939
rect 5908 24896 5960 24905
rect 6000 24896 6052 24948
rect 5724 24828 5776 24880
rect 6460 24828 6512 24880
rect 7012 24828 7064 24880
rect 9036 24896 9088 24948
rect 9588 24896 9640 24948
rect 10048 24896 10100 24948
rect 11888 24896 11940 24948
rect 13360 24896 13412 24948
rect 13544 24896 13596 24948
rect 15384 24896 15436 24948
rect 15844 24939 15896 24948
rect 15844 24905 15853 24939
rect 15853 24905 15887 24939
rect 15887 24905 15896 24939
rect 15844 24896 15896 24905
rect 17408 24939 17460 24948
rect 17408 24905 17417 24939
rect 17417 24905 17451 24939
rect 17451 24905 17460 24939
rect 17408 24896 17460 24905
rect 18880 24896 18932 24948
rect 13084 24828 13136 24880
rect 9680 24803 9732 24812
rect 9680 24769 9686 24803
rect 9686 24769 9720 24803
rect 9720 24769 9732 24803
rect 9680 24760 9732 24769
rect 9772 24760 9824 24812
rect 11152 24760 11204 24812
rect 4528 24692 4580 24744
rect 4804 24692 4856 24744
rect 7288 24692 7340 24744
rect 8208 24735 8260 24744
rect 8208 24701 8217 24735
rect 8217 24701 8251 24735
rect 8251 24701 8260 24735
rect 8208 24692 8260 24701
rect 9220 24692 9272 24744
rect 10232 24692 10284 24744
rect 9128 24624 9180 24676
rect 11428 24692 11480 24744
rect 11796 24735 11848 24744
rect 11796 24701 11805 24735
rect 11805 24701 11839 24735
rect 11839 24701 11848 24735
rect 11796 24692 11848 24701
rect 11888 24735 11940 24744
rect 11888 24701 11897 24735
rect 11897 24701 11931 24735
rect 11931 24701 11940 24735
rect 11888 24692 11940 24701
rect 11980 24692 12032 24744
rect 12164 24624 12216 24676
rect 12348 24803 12400 24812
rect 12348 24769 12357 24803
rect 12357 24769 12391 24803
rect 12391 24769 12400 24803
rect 12348 24760 12400 24769
rect 12440 24803 12492 24812
rect 12440 24769 12449 24803
rect 12449 24769 12483 24803
rect 12483 24769 12492 24803
rect 12440 24760 12492 24769
rect 12716 24803 12768 24812
rect 12716 24769 12725 24803
rect 12725 24769 12759 24803
rect 12759 24769 12768 24803
rect 12716 24760 12768 24769
rect 15108 24828 15160 24880
rect 13360 24803 13412 24812
rect 13360 24769 13369 24803
rect 13369 24769 13403 24803
rect 13403 24769 13412 24803
rect 13360 24760 13412 24769
rect 13452 24760 13504 24812
rect 14096 24760 14148 24812
rect 15660 24760 15712 24812
rect 17684 24760 17736 24812
rect 17868 24803 17920 24812
rect 17868 24769 17877 24803
rect 17877 24769 17911 24803
rect 17911 24769 17920 24803
rect 17868 24760 17920 24769
rect 18512 24803 18564 24812
rect 18512 24769 18521 24803
rect 18521 24769 18555 24803
rect 18555 24769 18564 24803
rect 18512 24760 18564 24769
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 19432 24828 19484 24880
rect 18972 24760 19024 24769
rect 19892 24803 19944 24812
rect 19892 24769 19901 24803
rect 19901 24769 19935 24803
rect 19935 24769 19944 24803
rect 19892 24760 19944 24769
rect 12900 24692 12952 24744
rect 18696 24692 18748 24744
rect 19524 24692 19576 24744
rect 19248 24624 19300 24676
rect 20812 24828 20864 24880
rect 20168 24760 20220 24812
rect 20628 24760 20680 24812
rect 20720 24760 20772 24812
rect 21732 24828 21784 24880
rect 21824 24828 21876 24880
rect 26976 24896 27028 24948
rect 28816 24939 28868 24948
rect 28816 24905 28825 24939
rect 28825 24905 28859 24939
rect 28859 24905 28868 24939
rect 28816 24896 28868 24905
rect 24768 24828 24820 24880
rect 26240 24828 26292 24880
rect 23296 24803 23348 24812
rect 23296 24769 23305 24803
rect 23305 24769 23339 24803
rect 23339 24769 23348 24803
rect 23296 24760 23348 24769
rect 23388 24803 23440 24812
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 23572 24760 23624 24812
rect 20352 24692 20404 24744
rect 21364 24692 21416 24744
rect 21732 24692 21784 24744
rect 22744 24692 22796 24744
rect 23020 24692 23072 24744
rect 24124 24692 24176 24744
rect 25228 24760 25280 24812
rect 28724 24828 28776 24880
rect 30196 24896 30248 24948
rect 30932 24896 30984 24948
rect 26608 24760 26660 24812
rect 26700 24760 26752 24812
rect 22376 24624 22428 24676
rect 25872 24692 25924 24744
rect 27160 24735 27212 24744
rect 27160 24701 27169 24735
rect 27169 24701 27203 24735
rect 27203 24701 27212 24735
rect 27160 24692 27212 24701
rect 26240 24624 26292 24676
rect 27528 24624 27580 24676
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 28264 24803 28316 24812
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 28540 24803 28592 24812
rect 28540 24769 28549 24803
rect 28549 24769 28583 24803
rect 28583 24769 28592 24803
rect 28540 24760 28592 24769
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 29184 24803 29236 24812
rect 29184 24769 29193 24803
rect 29193 24769 29227 24803
rect 29227 24769 29236 24803
rect 29184 24760 29236 24769
rect 29736 24828 29788 24880
rect 31852 24896 31904 24948
rect 32496 24896 32548 24948
rect 33140 24896 33192 24948
rect 35256 24896 35308 24948
rect 35808 24896 35860 24948
rect 31300 24871 31352 24880
rect 31300 24837 31309 24871
rect 31309 24837 31343 24871
rect 31343 24837 31352 24871
rect 31300 24828 31352 24837
rect 28172 24735 28224 24744
rect 28172 24701 28181 24735
rect 28181 24701 28215 24735
rect 28215 24701 28224 24735
rect 30380 24760 30432 24812
rect 28172 24692 28224 24701
rect 30932 24803 30984 24812
rect 30932 24769 30941 24803
rect 30941 24769 30975 24803
rect 30975 24769 30984 24803
rect 30932 24760 30984 24769
rect 31944 24828 31996 24880
rect 32128 24760 32180 24812
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32312 24760 32364 24769
rect 32404 24803 32456 24812
rect 32404 24769 32413 24803
rect 32413 24769 32447 24803
rect 32447 24769 32456 24803
rect 32404 24760 32456 24769
rect 31484 24692 31536 24744
rect 32588 24760 32640 24812
rect 32864 24803 32916 24812
rect 32864 24769 32873 24803
rect 32873 24769 32907 24803
rect 32907 24769 32916 24803
rect 32864 24760 32916 24769
rect 35164 24828 35216 24880
rect 33324 24760 33376 24812
rect 33692 24803 33744 24812
rect 33692 24769 33701 24803
rect 33701 24769 33735 24803
rect 33735 24769 33744 24803
rect 33692 24760 33744 24769
rect 33968 24760 34020 24812
rect 34152 24803 34204 24812
rect 34152 24769 34161 24803
rect 34161 24769 34195 24803
rect 34195 24769 34204 24803
rect 34152 24760 34204 24769
rect 6000 24556 6052 24608
rect 6184 24556 6236 24608
rect 7840 24556 7892 24608
rect 8024 24556 8076 24608
rect 8484 24556 8536 24608
rect 10416 24556 10468 24608
rect 11704 24556 11756 24608
rect 11980 24556 12032 24608
rect 12256 24556 12308 24608
rect 12992 24556 13044 24608
rect 15476 24599 15528 24608
rect 15476 24565 15485 24599
rect 15485 24565 15519 24599
rect 15519 24565 15528 24599
rect 15476 24556 15528 24565
rect 15660 24599 15712 24608
rect 15660 24565 15669 24599
rect 15669 24565 15703 24599
rect 15703 24565 15712 24599
rect 15660 24556 15712 24565
rect 17960 24599 18012 24608
rect 17960 24565 17969 24599
rect 17969 24565 18003 24599
rect 18003 24565 18012 24599
rect 17960 24556 18012 24565
rect 18144 24599 18196 24608
rect 18144 24565 18153 24599
rect 18153 24565 18187 24599
rect 18187 24565 18196 24599
rect 18144 24556 18196 24565
rect 18696 24556 18748 24608
rect 19616 24556 19668 24608
rect 19708 24599 19760 24608
rect 19708 24565 19717 24599
rect 19717 24565 19751 24599
rect 19751 24565 19760 24599
rect 19708 24556 19760 24565
rect 19800 24556 19852 24608
rect 21364 24556 21416 24608
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 21548 24556 21600 24608
rect 24124 24556 24176 24608
rect 25044 24556 25096 24608
rect 25872 24556 25924 24608
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 27160 24556 27212 24608
rect 28356 24556 28408 24608
rect 29276 24556 29328 24608
rect 30932 24556 30984 24608
rect 31024 24556 31076 24608
rect 31300 24556 31352 24608
rect 31760 24556 31812 24608
rect 31944 24556 31996 24608
rect 32128 24556 32180 24608
rect 32404 24556 32456 24608
rect 32588 24556 32640 24608
rect 33232 24556 33284 24608
rect 34060 24599 34112 24608
rect 34060 24565 34069 24599
rect 34069 24565 34103 24599
rect 34103 24565 34112 24599
rect 34060 24556 34112 24565
rect 34428 24735 34480 24744
rect 34428 24701 34437 24735
rect 34437 24701 34471 24735
rect 34471 24701 34480 24735
rect 34428 24692 34480 24701
rect 36176 24735 36228 24744
rect 36176 24701 36185 24735
rect 36185 24701 36219 24735
rect 36219 24701 36228 24735
rect 36176 24692 36228 24701
rect 34612 24556 34664 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4620 24352 4672 24404
rect 4068 24284 4120 24336
rect 7104 24352 7156 24404
rect 7288 24395 7340 24404
rect 7288 24361 7297 24395
rect 7297 24361 7331 24395
rect 7331 24361 7340 24395
rect 7288 24352 7340 24361
rect 11428 24395 11480 24404
rect 11428 24361 11437 24395
rect 11437 24361 11471 24395
rect 11471 24361 11480 24395
rect 11428 24352 11480 24361
rect 11612 24352 11664 24404
rect 12532 24352 12584 24404
rect 14096 24395 14148 24404
rect 14096 24361 14105 24395
rect 14105 24361 14139 24395
rect 14139 24361 14148 24395
rect 14096 24352 14148 24361
rect 14464 24352 14516 24404
rect 3608 24216 3660 24268
rect 6276 24284 6328 24336
rect 8392 24327 8444 24336
rect 8392 24293 8401 24327
rect 8401 24293 8435 24327
rect 8435 24293 8444 24327
rect 8392 24284 8444 24293
rect 10140 24284 10192 24336
rect 10324 24284 10376 24336
rect 3424 24191 3476 24200
rect 3424 24157 3433 24191
rect 3433 24157 3467 24191
rect 3467 24157 3476 24191
rect 3424 24148 3476 24157
rect 4528 24191 4580 24200
rect 4528 24157 4537 24191
rect 4537 24157 4571 24191
rect 4571 24157 4580 24191
rect 4528 24148 4580 24157
rect 5908 24216 5960 24268
rect 6184 24148 6236 24200
rect 6460 24191 6512 24200
rect 6460 24157 6469 24191
rect 6469 24157 6503 24191
rect 6503 24157 6512 24191
rect 6460 24148 6512 24157
rect 7196 24216 7248 24268
rect 7840 24259 7892 24268
rect 7840 24225 7849 24259
rect 7849 24225 7883 24259
rect 7883 24225 7892 24259
rect 7840 24216 7892 24225
rect 6828 24191 6880 24200
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 8024 24148 8076 24200
rect 6644 24123 6696 24132
rect 6644 24089 6653 24123
rect 6653 24089 6687 24123
rect 6687 24089 6696 24123
rect 6644 24080 6696 24089
rect 8484 24080 8536 24132
rect 2320 24012 2372 24064
rect 4620 24012 4672 24064
rect 6276 24055 6328 24064
rect 6276 24021 6285 24055
rect 6285 24021 6319 24055
rect 6319 24021 6328 24055
rect 6276 24012 6328 24021
rect 8392 24012 8444 24064
rect 9772 24148 9824 24200
rect 10140 24148 10192 24200
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 10324 24148 10376 24157
rect 12716 24284 12768 24336
rect 10876 24216 10928 24268
rect 11980 24259 12032 24268
rect 11980 24225 11989 24259
rect 11989 24225 12023 24259
rect 12023 24225 12032 24259
rect 11980 24216 12032 24225
rect 9864 24080 9916 24132
rect 10048 24012 10100 24064
rect 10600 24012 10652 24064
rect 10784 24012 10836 24064
rect 11704 24191 11756 24200
rect 11704 24157 11713 24191
rect 11713 24157 11747 24191
rect 11747 24157 11756 24191
rect 11704 24148 11756 24157
rect 12348 24148 12400 24200
rect 11888 24012 11940 24064
rect 11980 24012 12032 24064
rect 12164 24080 12216 24132
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 13544 24216 13596 24268
rect 16396 24352 16448 24404
rect 17040 24352 17092 24404
rect 19708 24352 19760 24404
rect 15476 24284 15528 24336
rect 19432 24284 19484 24336
rect 19892 24284 19944 24336
rect 22376 24395 22428 24404
rect 22376 24361 22385 24395
rect 22385 24361 22419 24395
rect 22419 24361 22428 24395
rect 22376 24352 22428 24361
rect 22928 24352 22980 24404
rect 23388 24395 23440 24404
rect 23388 24361 23397 24395
rect 23397 24361 23431 24395
rect 23431 24361 23440 24395
rect 23388 24352 23440 24361
rect 25964 24352 26016 24404
rect 26516 24352 26568 24404
rect 28356 24352 28408 24404
rect 29000 24395 29052 24404
rect 29000 24361 29009 24395
rect 29009 24361 29043 24395
rect 29043 24361 29052 24395
rect 29000 24352 29052 24361
rect 29184 24395 29236 24404
rect 29184 24361 29193 24395
rect 29193 24361 29227 24395
rect 29227 24361 29236 24395
rect 29184 24352 29236 24361
rect 30380 24352 30432 24404
rect 31668 24352 31720 24404
rect 33048 24284 33100 24336
rect 33324 24395 33376 24404
rect 33324 24361 33333 24395
rect 33333 24361 33367 24395
rect 33367 24361 33376 24395
rect 33324 24352 33376 24361
rect 33784 24395 33836 24404
rect 33784 24361 33793 24395
rect 33793 24361 33827 24395
rect 33827 24361 33836 24395
rect 33784 24352 33836 24361
rect 34428 24352 34480 24404
rect 35164 24352 35216 24404
rect 35808 24395 35860 24404
rect 35808 24361 35817 24395
rect 35817 24361 35851 24395
rect 35851 24361 35860 24395
rect 35808 24352 35860 24361
rect 13636 24148 13688 24200
rect 14280 24191 14332 24200
rect 14280 24157 14289 24191
rect 14289 24157 14323 24191
rect 14323 24157 14332 24191
rect 14280 24148 14332 24157
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 14648 24191 14700 24200
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 18144 24216 18196 24268
rect 19064 24216 19116 24268
rect 23296 24216 23348 24268
rect 27344 24216 27396 24268
rect 13820 24080 13872 24132
rect 15016 24080 15068 24132
rect 16120 24123 16172 24132
rect 16120 24089 16129 24123
rect 16129 24089 16163 24123
rect 16163 24089 16172 24123
rect 16120 24080 16172 24089
rect 12716 24012 12768 24064
rect 12900 24012 12952 24064
rect 13176 24012 13228 24064
rect 16028 24012 16080 24064
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 17224 24148 17276 24200
rect 17684 24148 17736 24200
rect 19616 24148 19668 24200
rect 20352 24191 20404 24200
rect 17592 24080 17644 24132
rect 19432 24080 19484 24132
rect 20352 24157 20361 24191
rect 20361 24157 20395 24191
rect 20395 24157 20404 24191
rect 20352 24148 20404 24157
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 22744 24191 22796 24200
rect 22744 24157 22753 24191
rect 22753 24157 22787 24191
rect 22787 24157 22796 24191
rect 22744 24148 22796 24157
rect 20628 24080 20680 24132
rect 23020 24191 23072 24200
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 23020 24148 23072 24157
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 24860 24148 24912 24200
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25044 24191 25096 24200
rect 25044 24157 25053 24191
rect 25053 24157 25087 24191
rect 25087 24157 25096 24191
rect 25044 24148 25096 24157
rect 25136 24191 25188 24200
rect 25136 24157 25145 24191
rect 25145 24157 25179 24191
rect 25179 24157 25188 24191
rect 25136 24148 25188 24157
rect 25780 24148 25832 24200
rect 25872 24191 25924 24200
rect 25872 24157 25881 24191
rect 25881 24157 25915 24191
rect 25915 24157 25924 24191
rect 25872 24148 25924 24157
rect 26332 24191 26384 24200
rect 26332 24157 26341 24191
rect 26341 24157 26375 24191
rect 26375 24157 26384 24191
rect 26332 24148 26384 24157
rect 27160 24148 27212 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 28724 24148 28776 24200
rect 22928 24080 22980 24132
rect 23756 24080 23808 24132
rect 25504 24123 25556 24132
rect 25504 24089 25513 24123
rect 25513 24089 25547 24123
rect 25547 24089 25556 24123
rect 25504 24080 25556 24089
rect 27712 24080 27764 24132
rect 29276 24148 29328 24200
rect 31116 24148 31168 24200
rect 32496 24191 32548 24200
rect 32496 24157 32505 24191
rect 32505 24157 32539 24191
rect 32539 24157 32548 24191
rect 32496 24148 32548 24157
rect 32864 24216 32916 24268
rect 36360 24284 36412 24336
rect 33876 24259 33928 24268
rect 33876 24225 33885 24259
rect 33885 24225 33919 24259
rect 33919 24225 33928 24259
rect 33876 24216 33928 24225
rect 36176 24216 36228 24268
rect 32772 24148 32824 24200
rect 17316 24012 17368 24064
rect 19524 24055 19576 24064
rect 19524 24021 19533 24055
rect 19533 24021 19567 24055
rect 19567 24021 19576 24055
rect 19524 24012 19576 24021
rect 19800 24012 19852 24064
rect 20168 24012 20220 24064
rect 21824 24012 21876 24064
rect 22468 24012 22520 24064
rect 23664 24012 23716 24064
rect 25136 24012 25188 24064
rect 25596 24012 25648 24064
rect 28080 24012 28132 24064
rect 28172 24012 28224 24064
rect 29736 24080 29788 24132
rect 28724 24012 28776 24064
rect 29920 24012 29972 24064
rect 31760 24080 31812 24132
rect 31944 24080 31996 24132
rect 32588 24080 32640 24132
rect 31668 24012 31720 24064
rect 32772 24012 32824 24064
rect 33416 24080 33468 24132
rect 33784 24080 33836 24132
rect 33876 24080 33928 24132
rect 33600 24012 33652 24064
rect 34244 24012 34296 24064
rect 34796 24148 34848 24200
rect 34980 24191 35032 24200
rect 34980 24157 34989 24191
rect 34989 24157 35023 24191
rect 35023 24157 35032 24191
rect 34980 24148 35032 24157
rect 35256 24191 35308 24200
rect 35256 24157 35265 24191
rect 35265 24157 35299 24191
rect 35299 24157 35308 24191
rect 35256 24148 35308 24157
rect 36084 24191 36136 24200
rect 36084 24157 36093 24191
rect 36093 24157 36127 24191
rect 36127 24157 36136 24191
rect 36084 24148 36136 24157
rect 34612 24080 34664 24132
rect 35532 24123 35584 24132
rect 35532 24089 35541 24123
rect 35541 24089 35575 24123
rect 35575 24089 35584 24123
rect 35532 24080 35584 24089
rect 35348 24012 35400 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 2320 23851 2372 23860
rect 2320 23817 2329 23851
rect 2329 23817 2363 23851
rect 2363 23817 2372 23851
rect 2320 23808 2372 23817
rect 3148 23740 3200 23792
rect 4068 23808 4120 23860
rect 4528 23851 4580 23860
rect 4528 23817 4537 23851
rect 4537 23817 4571 23851
rect 4571 23817 4580 23851
rect 4528 23808 4580 23817
rect 5172 23808 5224 23860
rect 5448 23808 5500 23860
rect 6000 23808 6052 23860
rect 8668 23808 8720 23860
rect 9680 23808 9732 23860
rect 10140 23808 10192 23860
rect 10324 23808 10376 23860
rect 2688 23672 2740 23724
rect 2780 23715 2832 23724
rect 2780 23681 2789 23715
rect 2789 23681 2823 23715
rect 2823 23681 2832 23715
rect 2780 23672 2832 23681
rect 5172 23715 5224 23724
rect 5172 23681 5181 23715
rect 5181 23681 5215 23715
rect 5215 23681 5224 23715
rect 5172 23672 5224 23681
rect 5356 23672 5408 23724
rect 6644 23740 6696 23792
rect 7104 23740 7156 23792
rect 9220 23783 9272 23792
rect 9220 23749 9229 23783
rect 9229 23749 9263 23783
rect 9263 23749 9272 23783
rect 9220 23740 9272 23749
rect 2320 23604 2372 23656
rect 2596 23647 2648 23656
rect 2596 23613 2605 23647
rect 2605 23613 2639 23647
rect 2639 23613 2648 23647
rect 2596 23604 2648 23613
rect 3056 23647 3108 23656
rect 3056 23613 3065 23647
rect 3065 23613 3099 23647
rect 3099 23613 3108 23647
rect 3056 23604 3108 23613
rect 4712 23604 4764 23656
rect 7012 23604 7064 23656
rect 9128 23715 9180 23724
rect 9128 23681 9137 23715
rect 9137 23681 9171 23715
rect 9171 23681 9180 23715
rect 9128 23672 9180 23681
rect 9220 23604 9272 23656
rect 10600 23672 10652 23724
rect 11428 23672 11480 23724
rect 11888 23715 11940 23724
rect 11888 23681 11897 23715
rect 11897 23681 11931 23715
rect 11931 23681 11940 23715
rect 11888 23672 11940 23681
rect 12440 23672 12492 23724
rect 12900 23672 12952 23724
rect 10416 23604 10468 23656
rect 12072 23604 12124 23656
rect 12164 23647 12216 23656
rect 12164 23613 12173 23647
rect 12173 23613 12207 23647
rect 12207 23613 12216 23647
rect 12164 23604 12216 23613
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 13360 23715 13412 23724
rect 13360 23681 13369 23715
rect 13369 23681 13403 23715
rect 13403 23681 13412 23715
rect 13360 23672 13412 23681
rect 14280 23808 14332 23860
rect 15660 23808 15712 23860
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 13820 23783 13872 23792
rect 13820 23749 13829 23783
rect 13829 23749 13863 23783
rect 13863 23749 13872 23783
rect 13820 23740 13872 23749
rect 14464 23740 14516 23792
rect 16120 23740 16172 23792
rect 16948 23808 17000 23860
rect 17960 23808 18012 23860
rect 14096 23715 14148 23724
rect 14096 23681 14105 23715
rect 14105 23681 14139 23715
rect 14139 23681 14148 23715
rect 14096 23672 14148 23681
rect 15200 23672 15252 23724
rect 15660 23672 15712 23724
rect 16304 23715 16356 23724
rect 16304 23681 16313 23715
rect 16313 23681 16347 23715
rect 16347 23681 16356 23715
rect 16304 23672 16356 23681
rect 16396 23672 16448 23724
rect 16948 23672 17000 23724
rect 17316 23715 17368 23724
rect 17316 23681 17325 23715
rect 17325 23681 17359 23715
rect 17359 23681 17368 23715
rect 17316 23672 17368 23681
rect 18052 23672 18104 23724
rect 18328 23672 18380 23724
rect 19156 23740 19208 23792
rect 21548 23808 21600 23860
rect 21640 23808 21692 23860
rect 22008 23740 22060 23792
rect 18696 23715 18748 23724
rect 18696 23681 18705 23715
rect 18705 23681 18739 23715
rect 18739 23681 18748 23715
rect 18696 23672 18748 23681
rect 18788 23672 18840 23724
rect 21548 23672 21600 23724
rect 21640 23672 21692 23724
rect 22376 23672 22428 23724
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 25688 23808 25740 23860
rect 26516 23808 26568 23860
rect 28172 23808 28224 23860
rect 28540 23808 28592 23860
rect 30196 23808 30248 23860
rect 23296 23740 23348 23792
rect 23756 23740 23808 23792
rect 24492 23783 24544 23792
rect 24492 23749 24501 23783
rect 24501 23749 24535 23783
rect 24535 23749 24544 23783
rect 24492 23740 24544 23749
rect 22560 23672 22612 23681
rect 23388 23715 23440 23724
rect 23388 23681 23397 23715
rect 23397 23681 23431 23715
rect 23431 23681 23440 23715
rect 23388 23672 23440 23681
rect 24676 23715 24728 23724
rect 24676 23681 24685 23715
rect 24685 23681 24719 23715
rect 24719 23681 24728 23715
rect 24676 23672 24728 23681
rect 24860 23672 24912 23724
rect 24952 23715 25004 23724
rect 24952 23681 24961 23715
rect 24961 23681 24995 23715
rect 24995 23681 25004 23715
rect 24952 23672 25004 23681
rect 25228 23672 25280 23724
rect 25320 23715 25372 23724
rect 25320 23681 25329 23715
rect 25329 23681 25363 23715
rect 25363 23681 25372 23715
rect 25320 23672 25372 23681
rect 25504 23740 25556 23792
rect 27252 23740 27304 23792
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 7748 23536 7800 23588
rect 9864 23536 9916 23588
rect 10140 23536 10192 23588
rect 11060 23536 11112 23588
rect 15292 23604 15344 23656
rect 15476 23647 15528 23656
rect 15476 23613 15485 23647
rect 15485 23613 15519 23647
rect 15519 23613 15528 23647
rect 15476 23604 15528 23613
rect 15568 23604 15620 23656
rect 15844 23604 15896 23656
rect 17684 23647 17736 23656
rect 17684 23613 17693 23647
rect 17693 23613 17727 23647
rect 17727 23613 17736 23647
rect 17684 23604 17736 23613
rect 15936 23536 15988 23588
rect 16304 23536 16356 23588
rect 1676 23468 1728 23520
rect 3240 23468 3292 23520
rect 4988 23468 5040 23520
rect 6000 23468 6052 23520
rect 7196 23468 7248 23520
rect 8024 23468 8076 23520
rect 8208 23511 8260 23520
rect 8208 23477 8217 23511
rect 8217 23477 8251 23511
rect 8251 23477 8260 23511
rect 8208 23468 8260 23477
rect 8392 23468 8444 23520
rect 11796 23468 11848 23520
rect 12348 23468 12400 23520
rect 16028 23468 16080 23520
rect 18972 23647 19024 23656
rect 18972 23613 18981 23647
rect 18981 23613 19015 23647
rect 19015 23613 19024 23647
rect 18972 23604 19024 23613
rect 19248 23604 19300 23656
rect 18604 23536 18656 23588
rect 19800 23604 19852 23656
rect 21824 23604 21876 23656
rect 22192 23647 22244 23656
rect 22192 23613 22201 23647
rect 22201 23613 22235 23647
rect 22235 23613 22244 23647
rect 22192 23604 22244 23613
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 28080 23715 28132 23724
rect 28080 23681 28089 23715
rect 28089 23681 28123 23715
rect 28123 23681 28132 23715
rect 28080 23672 28132 23681
rect 28172 23672 28224 23724
rect 28540 23672 28592 23724
rect 29092 23740 29144 23792
rect 33324 23808 33376 23860
rect 34520 23808 34572 23860
rect 35256 23808 35308 23860
rect 27804 23604 27856 23656
rect 19892 23536 19944 23588
rect 20260 23536 20312 23588
rect 31300 23715 31352 23724
rect 31300 23681 31309 23715
rect 31309 23681 31343 23715
rect 31343 23681 31352 23715
rect 31300 23672 31352 23681
rect 31576 23783 31628 23792
rect 31576 23749 31585 23783
rect 31585 23749 31619 23783
rect 31619 23749 31628 23783
rect 31576 23740 31628 23749
rect 32312 23672 32364 23724
rect 28816 23536 28868 23588
rect 29736 23536 29788 23588
rect 18420 23468 18472 23520
rect 18696 23468 18748 23520
rect 19156 23468 19208 23520
rect 19340 23468 19392 23520
rect 19616 23468 19668 23520
rect 20352 23468 20404 23520
rect 22008 23468 22060 23520
rect 22284 23468 22336 23520
rect 27988 23468 28040 23520
rect 28448 23511 28500 23520
rect 28448 23477 28457 23511
rect 28457 23477 28491 23511
rect 28491 23477 28500 23511
rect 28448 23468 28500 23477
rect 28540 23468 28592 23520
rect 30288 23511 30340 23520
rect 30288 23477 30297 23511
rect 30297 23477 30331 23511
rect 30331 23477 30340 23511
rect 30288 23468 30340 23477
rect 31392 23536 31444 23588
rect 31668 23536 31720 23588
rect 33600 23647 33652 23656
rect 33600 23613 33609 23647
rect 33609 23613 33643 23647
rect 33643 23613 33652 23647
rect 33600 23604 33652 23613
rect 33784 23715 33836 23724
rect 33784 23681 33793 23715
rect 33793 23681 33827 23715
rect 33827 23681 33836 23715
rect 33784 23672 33836 23681
rect 35348 23672 35400 23724
rect 36176 23715 36228 23724
rect 36176 23681 36185 23715
rect 36185 23681 36219 23715
rect 36219 23681 36228 23715
rect 36176 23672 36228 23681
rect 33876 23604 33928 23656
rect 33232 23536 33284 23588
rect 33416 23579 33468 23588
rect 33416 23545 33425 23579
rect 33425 23545 33459 23579
rect 33459 23545 33468 23579
rect 33416 23536 33468 23545
rect 33968 23536 34020 23588
rect 30564 23468 30616 23520
rect 31116 23468 31168 23520
rect 32036 23468 32088 23520
rect 32588 23468 32640 23520
rect 33876 23468 33928 23520
rect 35164 23511 35216 23520
rect 35164 23477 35173 23511
rect 35173 23477 35207 23511
rect 35207 23477 35216 23511
rect 35164 23468 35216 23477
rect 35348 23468 35400 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3056 23264 3108 23316
rect 3976 23264 4028 23316
rect 9680 23307 9732 23316
rect 9680 23273 9689 23307
rect 9689 23273 9723 23307
rect 9723 23273 9732 23307
rect 9680 23264 9732 23273
rect 9772 23264 9824 23316
rect 12072 23264 12124 23316
rect 3424 23196 3476 23248
rect 4712 23196 4764 23248
rect 4896 23196 4948 23248
rect 5356 23196 5408 23248
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 1676 23171 1728 23180
rect 1676 23137 1685 23171
rect 1685 23137 1719 23171
rect 1719 23137 1728 23171
rect 1676 23128 1728 23137
rect 4068 23128 4120 23180
rect 4528 23060 4580 23112
rect 6276 23128 6328 23180
rect 7012 23128 7064 23180
rect 4712 23103 4764 23112
rect 4712 23069 4722 23103
rect 4722 23069 4756 23103
rect 4756 23069 4764 23103
rect 4712 23060 4764 23069
rect 4896 23103 4948 23112
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 5816 23060 5868 23112
rect 3148 22992 3200 23044
rect 3424 22992 3476 23044
rect 3976 22992 4028 23044
rect 4988 23035 5040 23044
rect 4988 23001 4997 23035
rect 4997 23001 5031 23035
rect 5031 23001 5040 23035
rect 4988 22992 5040 23001
rect 4620 22924 4672 22976
rect 6460 23060 6512 23112
rect 7564 23128 7616 23180
rect 8024 23239 8076 23248
rect 8024 23205 8033 23239
rect 8033 23205 8067 23239
rect 8067 23205 8076 23239
rect 8024 23196 8076 23205
rect 8852 23128 8904 23180
rect 8208 23060 8260 23112
rect 9404 23103 9456 23112
rect 9404 23069 9413 23103
rect 9413 23069 9447 23103
rect 9447 23069 9456 23103
rect 9404 23060 9456 23069
rect 8024 22924 8076 22976
rect 9312 22992 9364 23044
rect 10140 23196 10192 23248
rect 11980 23196 12032 23248
rect 13544 23264 13596 23316
rect 15476 23264 15528 23316
rect 15660 23264 15712 23316
rect 10048 23171 10100 23180
rect 10048 23137 10057 23171
rect 10057 23137 10091 23171
rect 10091 23137 10100 23171
rect 10048 23128 10100 23137
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 10048 22992 10100 23044
rect 11612 23128 11664 23180
rect 11796 23128 11848 23180
rect 10784 23060 10836 23112
rect 11244 23060 11296 23112
rect 11428 23060 11480 23112
rect 12532 23196 12584 23248
rect 12808 23128 12860 23180
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 12992 23103 13044 23112
rect 12992 23069 13001 23103
rect 13001 23069 13035 23103
rect 13035 23069 13044 23103
rect 12992 23060 13044 23069
rect 13360 23128 13412 23180
rect 13912 23103 13964 23112
rect 13912 23069 13921 23103
rect 13921 23069 13955 23103
rect 13955 23069 13964 23103
rect 13912 23060 13964 23069
rect 15108 23196 15160 23248
rect 15936 23196 15988 23248
rect 16396 23196 16448 23248
rect 15200 23128 15252 23180
rect 14372 23060 14424 23112
rect 15660 23060 15712 23112
rect 15752 23103 15804 23112
rect 15752 23069 15761 23103
rect 15761 23069 15795 23103
rect 15795 23069 15804 23103
rect 15752 23060 15804 23069
rect 8392 22924 8444 22976
rect 8668 22924 8720 22976
rect 10232 22924 10284 22976
rect 11612 22924 11664 22976
rect 11888 22924 11940 22976
rect 12440 22924 12492 22976
rect 12992 22967 13044 22976
rect 12992 22933 13001 22967
rect 13001 22933 13035 22967
rect 13035 22933 13044 22967
rect 12992 22924 13044 22933
rect 14280 22924 14332 22976
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 15384 22992 15436 23044
rect 15844 22992 15896 23044
rect 16120 23060 16172 23112
rect 17868 23264 17920 23316
rect 18972 23264 19024 23316
rect 18604 23196 18656 23248
rect 16304 22992 16356 23044
rect 14924 22967 14976 22976
rect 14924 22933 14933 22967
rect 14933 22933 14967 22967
rect 14967 22933 14976 22967
rect 14924 22924 14976 22933
rect 15016 22924 15068 22976
rect 16856 23103 16908 23112
rect 16856 23069 16866 23103
rect 16866 23069 16900 23103
rect 16900 23069 16908 23103
rect 18144 23128 18196 23180
rect 19248 23171 19300 23180
rect 19248 23137 19257 23171
rect 19257 23137 19291 23171
rect 19291 23137 19300 23171
rect 19248 23128 19300 23137
rect 16856 23060 16908 23069
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 18972 23060 19024 23112
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 19524 23103 19576 23112
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 19892 23128 19944 23180
rect 20536 23171 20588 23180
rect 20536 23137 20545 23171
rect 20545 23137 20579 23171
rect 20579 23137 20588 23171
rect 20536 23128 20588 23137
rect 20076 23060 20128 23112
rect 20352 23060 20404 23112
rect 16764 22924 16816 22976
rect 17776 22992 17828 23044
rect 19156 22992 19208 23044
rect 21180 23196 21232 23248
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 21272 23060 21324 23112
rect 21916 23196 21968 23248
rect 22008 23196 22060 23248
rect 21640 23171 21692 23180
rect 21640 23137 21649 23171
rect 21649 23137 21683 23171
rect 21683 23137 21692 23171
rect 21640 23128 21692 23137
rect 22468 23196 22520 23248
rect 22836 23307 22888 23316
rect 22836 23273 22845 23307
rect 22845 23273 22879 23307
rect 22879 23273 22888 23307
rect 22836 23264 22888 23273
rect 23388 23264 23440 23316
rect 26148 23264 26200 23316
rect 26332 23264 26384 23316
rect 27344 23307 27396 23316
rect 27344 23273 27353 23307
rect 27353 23273 27387 23307
rect 27387 23273 27396 23307
rect 27344 23264 27396 23273
rect 22376 23128 22428 23180
rect 23480 23196 23532 23248
rect 25136 23196 25188 23248
rect 25596 23196 25648 23248
rect 22284 23060 22336 23112
rect 23756 23103 23808 23112
rect 23756 23069 23765 23103
rect 23765 23069 23799 23103
rect 23799 23069 23808 23103
rect 23756 23060 23808 23069
rect 25044 23103 25096 23112
rect 25044 23069 25053 23103
rect 25053 23069 25087 23103
rect 25087 23069 25096 23103
rect 25044 23060 25096 23069
rect 25320 23103 25372 23112
rect 25320 23069 25329 23103
rect 25329 23069 25363 23103
rect 25363 23069 25372 23103
rect 25320 23060 25372 23069
rect 25688 23060 25740 23112
rect 28540 23264 28592 23316
rect 29092 23264 29144 23316
rect 28356 23239 28408 23248
rect 28356 23205 28365 23239
rect 28365 23205 28399 23239
rect 28399 23205 28408 23239
rect 28356 23196 28408 23205
rect 30012 23264 30064 23316
rect 31576 23264 31628 23316
rect 33232 23264 33284 23316
rect 34796 23264 34848 23316
rect 30380 23196 30432 23248
rect 31116 23196 31168 23248
rect 28816 23128 28868 23180
rect 18052 22924 18104 22976
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 19708 22967 19760 22976
rect 19708 22933 19717 22967
rect 19717 22933 19751 22967
rect 19751 22933 19760 22967
rect 19708 22924 19760 22933
rect 19800 22924 19852 22976
rect 20996 22924 21048 22976
rect 21364 22924 21416 22976
rect 22376 22992 22428 23044
rect 22836 22992 22888 23044
rect 23572 22992 23624 23044
rect 25136 22992 25188 23044
rect 25504 22992 25556 23044
rect 26148 23103 26200 23112
rect 26148 23069 26157 23103
rect 26157 23069 26191 23103
rect 26191 23069 26200 23103
rect 26148 23060 26200 23069
rect 26424 23060 26476 23112
rect 26700 23060 26752 23112
rect 22744 22924 22796 22976
rect 23388 22967 23440 22976
rect 23388 22933 23397 22967
rect 23397 22933 23431 22967
rect 23431 22933 23440 22967
rect 23388 22924 23440 22933
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 25320 22924 25372 22976
rect 26976 23060 27028 23112
rect 28448 23103 28500 23112
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 26884 22924 26936 22976
rect 27160 22992 27212 23044
rect 27528 23035 27580 23044
rect 27528 23001 27537 23035
rect 27537 23001 27571 23035
rect 27571 23001 27580 23035
rect 27528 22992 27580 23001
rect 28540 22992 28592 23044
rect 29184 22992 29236 23044
rect 30196 23060 30248 23112
rect 30288 23103 30340 23112
rect 30288 23069 30297 23103
rect 30297 23069 30331 23103
rect 30331 23069 30340 23103
rect 30288 23060 30340 23069
rect 30380 23103 30432 23112
rect 30380 23069 30389 23103
rect 30389 23069 30423 23103
rect 30423 23069 30432 23103
rect 30380 23060 30432 23069
rect 30564 23103 30616 23112
rect 30564 23069 30573 23103
rect 30573 23069 30607 23103
rect 30607 23069 30616 23103
rect 30564 23060 30616 23069
rect 30840 23060 30892 23112
rect 27896 22924 27948 22976
rect 29092 22924 29144 22976
rect 29552 22924 29604 22976
rect 29828 22924 29880 22976
rect 30012 22924 30064 22976
rect 31208 23103 31260 23112
rect 31208 23069 31217 23103
rect 31217 23069 31251 23103
rect 31251 23069 31260 23103
rect 31208 23060 31260 23069
rect 32036 23196 32088 23248
rect 31668 23171 31720 23180
rect 31668 23137 31677 23171
rect 31677 23137 31711 23171
rect 31711 23137 31720 23171
rect 31668 23128 31720 23137
rect 31484 23103 31536 23112
rect 31484 23069 31519 23103
rect 31519 23069 31536 23103
rect 31484 23060 31536 23069
rect 31760 23103 31812 23112
rect 31760 23069 31769 23103
rect 31769 23069 31803 23103
rect 31803 23069 31812 23103
rect 31760 23060 31812 23069
rect 32312 23103 32364 23112
rect 32312 23069 32321 23103
rect 32321 23069 32355 23103
rect 32355 23069 32364 23103
rect 32312 23060 32364 23069
rect 35256 23103 35308 23112
rect 35256 23069 35265 23103
rect 35265 23069 35299 23103
rect 35299 23069 35308 23103
rect 35256 23060 35308 23069
rect 30196 22967 30248 22976
rect 30196 22933 30205 22967
rect 30205 22933 30239 22967
rect 30239 22933 30248 22967
rect 30196 22924 30248 22933
rect 30656 22924 30708 22976
rect 30932 22924 30984 22976
rect 31208 22924 31260 22976
rect 32496 22992 32548 23044
rect 33048 22992 33100 23044
rect 35072 23035 35124 23044
rect 35072 23001 35081 23035
rect 35081 23001 35115 23035
rect 35115 23001 35124 23035
rect 35072 22992 35124 23001
rect 32956 22924 33008 22976
rect 34428 22924 34480 22976
rect 34796 22924 34848 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 3240 22720 3292 22772
rect 3608 22720 3660 22772
rect 7288 22720 7340 22772
rect 7564 22720 7616 22772
rect 8116 22720 8168 22772
rect 8300 22720 8352 22772
rect 8944 22720 8996 22772
rect 9404 22720 9456 22772
rect 10600 22720 10652 22772
rect 3884 22584 3936 22636
rect 4436 22627 4488 22636
rect 4436 22593 4445 22627
rect 4445 22593 4479 22627
rect 4479 22593 4488 22627
rect 4436 22584 4488 22593
rect 2596 22516 2648 22568
rect 3976 22559 4028 22568
rect 3976 22525 3985 22559
rect 3985 22525 4019 22559
rect 4019 22525 4028 22559
rect 3976 22516 4028 22525
rect 4712 22627 4764 22636
rect 4712 22593 4721 22627
rect 4721 22593 4755 22627
rect 4755 22593 4764 22627
rect 4712 22584 4764 22593
rect 5540 22652 5592 22704
rect 5172 22627 5224 22636
rect 5172 22593 5181 22627
rect 5181 22593 5215 22627
rect 5215 22593 5224 22627
rect 5172 22584 5224 22593
rect 5356 22584 5408 22636
rect 5448 22627 5500 22636
rect 5448 22593 5457 22627
rect 5457 22593 5491 22627
rect 5491 22593 5500 22627
rect 5448 22584 5500 22593
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 5816 22627 5868 22636
rect 5816 22593 5825 22627
rect 5825 22593 5859 22627
rect 5859 22593 5868 22627
rect 5816 22584 5868 22593
rect 6828 22652 6880 22704
rect 7656 22695 7708 22704
rect 7656 22661 7665 22695
rect 7665 22661 7699 22695
rect 7699 22661 7708 22695
rect 7656 22652 7708 22661
rect 7932 22695 7984 22704
rect 7932 22661 7941 22695
rect 7941 22661 7975 22695
rect 7975 22661 7984 22695
rect 7932 22652 7984 22661
rect 8484 22652 8536 22704
rect 12256 22720 12308 22772
rect 12532 22720 12584 22772
rect 12716 22720 12768 22772
rect 15200 22720 15252 22772
rect 17684 22720 17736 22772
rect 18788 22720 18840 22772
rect 19156 22720 19208 22772
rect 20904 22720 20956 22772
rect 11888 22652 11940 22704
rect 5724 22516 5776 22568
rect 6644 22584 6696 22636
rect 8024 22627 8076 22636
rect 8024 22593 8038 22627
rect 8038 22593 8072 22627
rect 8072 22593 8076 22627
rect 8024 22584 8076 22593
rect 6736 22516 6788 22568
rect 10232 22584 10284 22636
rect 12164 22584 12216 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 13360 22584 13412 22636
rect 13912 22584 13964 22636
rect 14188 22584 14240 22636
rect 9864 22516 9916 22568
rect 11060 22516 11112 22568
rect 4068 22448 4120 22500
rect 4436 22448 4488 22500
rect 5356 22448 5408 22500
rect 5632 22448 5684 22500
rect 7472 22448 7524 22500
rect 1676 22380 1728 22432
rect 10692 22448 10744 22500
rect 10968 22448 11020 22500
rect 12072 22516 12124 22568
rect 12256 22448 12308 22500
rect 7656 22423 7708 22432
rect 7656 22389 7665 22423
rect 7665 22389 7699 22423
rect 7699 22389 7708 22423
rect 7656 22380 7708 22389
rect 7932 22380 7984 22432
rect 10324 22380 10376 22432
rect 10784 22380 10836 22432
rect 11060 22380 11112 22432
rect 11704 22380 11756 22432
rect 19248 22652 19300 22704
rect 15568 22627 15620 22636
rect 15568 22593 15577 22627
rect 15577 22593 15611 22627
rect 15611 22593 15620 22627
rect 15568 22584 15620 22593
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 15936 22584 15988 22636
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 17224 22584 17276 22636
rect 17592 22627 17644 22636
rect 17592 22593 17600 22627
rect 17600 22593 17634 22627
rect 17634 22593 17644 22627
rect 17592 22584 17644 22593
rect 15844 22516 15896 22568
rect 16672 22516 16724 22568
rect 17776 22627 17828 22636
rect 17776 22593 17785 22627
rect 17785 22593 17819 22627
rect 17819 22593 17828 22627
rect 17776 22584 17828 22593
rect 18328 22584 18380 22636
rect 18972 22584 19024 22636
rect 19800 22584 19852 22636
rect 19892 22627 19944 22636
rect 19892 22593 19901 22627
rect 19901 22593 19935 22627
rect 19935 22593 19944 22627
rect 19892 22584 19944 22593
rect 20076 22627 20128 22636
rect 20076 22593 20085 22627
rect 20085 22593 20119 22627
rect 20119 22593 20128 22627
rect 20076 22584 20128 22593
rect 20168 22627 20220 22636
rect 20168 22593 20177 22627
rect 20177 22593 20211 22627
rect 20211 22593 20220 22627
rect 20168 22584 20220 22593
rect 20536 22652 20588 22704
rect 21272 22652 21324 22704
rect 22008 22695 22060 22704
rect 22008 22661 22017 22695
rect 22017 22661 22051 22695
rect 22051 22661 22060 22695
rect 22008 22652 22060 22661
rect 22652 22720 22704 22772
rect 23388 22720 23440 22772
rect 25504 22720 25556 22772
rect 26148 22720 26200 22772
rect 26884 22720 26936 22772
rect 26976 22763 27028 22772
rect 26976 22729 26985 22763
rect 26985 22729 27019 22763
rect 27019 22729 27028 22763
rect 26976 22720 27028 22729
rect 30564 22720 30616 22772
rect 30840 22720 30892 22772
rect 31484 22720 31536 22772
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 21180 22627 21232 22636
rect 21180 22593 21189 22627
rect 21189 22593 21223 22627
rect 21223 22593 21232 22627
rect 21180 22584 21232 22593
rect 21456 22584 21508 22636
rect 21732 22584 21784 22636
rect 21916 22584 21968 22636
rect 18144 22516 18196 22568
rect 19248 22559 19300 22568
rect 19248 22525 19257 22559
rect 19257 22525 19291 22559
rect 19291 22525 19300 22559
rect 19248 22516 19300 22525
rect 12808 22448 12860 22500
rect 13084 22448 13136 22500
rect 12716 22380 12768 22432
rect 14280 22448 14332 22500
rect 14556 22448 14608 22500
rect 16304 22448 16356 22500
rect 18512 22448 18564 22500
rect 18788 22448 18840 22500
rect 19064 22448 19116 22500
rect 19156 22448 19208 22500
rect 22100 22448 22152 22500
rect 14188 22423 14240 22432
rect 14188 22389 14197 22423
rect 14197 22389 14231 22423
rect 14231 22389 14240 22423
rect 14188 22380 14240 22389
rect 18144 22380 18196 22432
rect 19616 22380 19668 22432
rect 20260 22423 20312 22432
rect 20260 22389 20269 22423
rect 20269 22389 20303 22423
rect 20303 22389 20312 22423
rect 20260 22380 20312 22389
rect 20628 22380 20680 22432
rect 22652 22627 22704 22636
rect 22652 22593 22661 22627
rect 22661 22593 22695 22627
rect 22695 22593 22704 22627
rect 22652 22584 22704 22593
rect 23204 22584 23256 22636
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24216 22584 24268 22636
rect 24400 22627 24452 22636
rect 24400 22593 24409 22627
rect 24409 22593 24443 22627
rect 24443 22593 24452 22627
rect 24400 22584 24452 22593
rect 24676 22584 24728 22636
rect 22744 22559 22796 22568
rect 22744 22525 22753 22559
rect 22753 22525 22787 22559
rect 22787 22525 22796 22559
rect 22744 22516 22796 22525
rect 22376 22448 22428 22500
rect 24124 22380 24176 22432
rect 24492 22380 24544 22432
rect 24768 22423 24820 22432
rect 24768 22389 24777 22423
rect 24777 22389 24811 22423
rect 24811 22389 24820 22423
rect 24768 22380 24820 22389
rect 27068 22652 27120 22704
rect 28356 22695 28408 22704
rect 28356 22661 28365 22695
rect 28365 22661 28399 22695
rect 28399 22661 28408 22695
rect 28356 22652 28408 22661
rect 26976 22584 27028 22636
rect 27344 22627 27396 22636
rect 27344 22593 27353 22627
rect 27353 22593 27387 22627
rect 27387 22593 27396 22627
rect 27344 22584 27396 22593
rect 26608 22516 26660 22568
rect 27160 22516 27212 22568
rect 27528 22584 27580 22636
rect 27528 22448 27580 22500
rect 29368 22627 29420 22636
rect 29368 22593 29377 22627
rect 29377 22593 29411 22627
rect 29411 22593 29420 22627
rect 29368 22584 29420 22593
rect 29552 22652 29604 22704
rect 29920 22627 29972 22636
rect 29920 22593 29929 22627
rect 29929 22593 29963 22627
rect 29963 22593 29972 22627
rect 29920 22584 29972 22593
rect 30012 22627 30064 22636
rect 30012 22593 30021 22627
rect 30021 22593 30055 22627
rect 30055 22593 30064 22627
rect 30012 22584 30064 22593
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 30288 22584 30340 22636
rect 28540 22448 28592 22500
rect 29276 22559 29328 22568
rect 29276 22525 29285 22559
rect 29285 22525 29319 22559
rect 29319 22525 29328 22559
rect 29276 22516 29328 22525
rect 30196 22448 30248 22500
rect 26884 22380 26936 22432
rect 28080 22380 28132 22432
rect 28908 22380 28960 22432
rect 29552 22380 29604 22432
rect 30840 22584 30892 22636
rect 31116 22652 31168 22704
rect 31852 22652 31904 22704
rect 31576 22584 31628 22636
rect 31116 22559 31168 22568
rect 31116 22525 31125 22559
rect 31125 22525 31159 22559
rect 31159 22525 31168 22559
rect 31116 22516 31168 22525
rect 31392 22559 31444 22568
rect 31392 22525 31401 22559
rect 31401 22525 31435 22559
rect 31435 22525 31444 22559
rect 31392 22516 31444 22525
rect 32220 22559 32272 22568
rect 32220 22525 32229 22559
rect 32229 22525 32263 22559
rect 32263 22525 32272 22559
rect 32220 22516 32272 22525
rect 32956 22652 33008 22704
rect 34428 22720 34480 22772
rect 34336 22695 34388 22704
rect 34336 22661 34345 22695
rect 34345 22661 34379 22695
rect 34379 22661 34388 22695
rect 34336 22652 34388 22661
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 33048 22627 33100 22636
rect 33048 22593 33057 22627
rect 33057 22593 33091 22627
rect 33091 22593 33100 22627
rect 33048 22584 33100 22593
rect 33232 22627 33284 22636
rect 33232 22593 33241 22627
rect 33241 22593 33275 22627
rect 33275 22593 33284 22627
rect 33232 22584 33284 22593
rect 34888 22627 34940 22636
rect 34888 22593 34897 22627
rect 34897 22593 34931 22627
rect 34931 22593 34940 22627
rect 34888 22584 34940 22593
rect 35348 22584 35400 22636
rect 36176 22559 36228 22568
rect 36176 22525 36185 22559
rect 36185 22525 36219 22559
rect 36219 22525 36228 22559
rect 36176 22516 36228 22525
rect 34612 22448 34664 22500
rect 31576 22423 31628 22432
rect 31576 22389 31585 22423
rect 31585 22389 31619 22423
rect 31619 22389 31628 22423
rect 31576 22380 31628 22389
rect 31668 22380 31720 22432
rect 32404 22380 32456 22432
rect 33508 22380 33560 22432
rect 33968 22423 34020 22432
rect 33968 22389 33977 22423
rect 33977 22389 34011 22423
rect 34011 22389 34020 22423
rect 33968 22380 34020 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1676 22219 1728 22228
rect 1676 22185 1706 22219
rect 1706 22185 1728 22219
rect 1676 22176 1728 22185
rect 3700 22176 3752 22228
rect 3976 22176 4028 22228
rect 2780 22108 2832 22160
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 2688 22040 2740 22092
rect 3976 22040 4028 22092
rect 4344 22083 4396 22092
rect 4344 22049 4353 22083
rect 4353 22049 4387 22083
rect 4387 22049 4396 22083
rect 4344 22040 4396 22049
rect 4712 22176 4764 22228
rect 8024 22176 8076 22228
rect 8300 22219 8352 22228
rect 8300 22185 8309 22219
rect 8309 22185 8343 22219
rect 8343 22185 8352 22219
rect 8300 22176 8352 22185
rect 9588 22176 9640 22228
rect 14188 22176 14240 22228
rect 14280 22219 14332 22228
rect 14280 22185 14289 22219
rect 14289 22185 14323 22219
rect 14323 22185 14332 22219
rect 14280 22176 14332 22185
rect 15476 22219 15528 22228
rect 15476 22185 15485 22219
rect 15485 22185 15519 22219
rect 15519 22185 15528 22219
rect 15476 22176 15528 22185
rect 5172 22108 5224 22160
rect 5080 21972 5132 22024
rect 5172 22015 5224 22024
rect 5172 21981 5180 22015
rect 5180 21981 5214 22015
rect 5214 21981 5224 22015
rect 5172 21972 5224 21981
rect 5264 22015 5316 22024
rect 5264 21981 5273 22015
rect 5273 21981 5307 22015
rect 5307 21981 5316 22015
rect 5264 21972 5316 21981
rect 5632 22040 5684 22092
rect 6644 22108 6696 22160
rect 7472 22108 7524 22160
rect 8484 22108 8536 22160
rect 9312 22108 9364 22160
rect 9864 22108 9916 22160
rect 2964 21904 3016 21956
rect 2412 21836 2464 21888
rect 4620 21904 4672 21956
rect 5724 22015 5776 22024
rect 5724 21981 5733 22015
rect 5733 21981 5767 22015
rect 5767 21981 5776 22015
rect 5724 21972 5776 21981
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 6092 22015 6144 22024
rect 6092 21981 6101 22015
rect 6101 21981 6135 22015
rect 6135 21981 6144 22015
rect 6092 21972 6144 21981
rect 6184 21972 6236 22024
rect 6736 22083 6788 22092
rect 6736 22049 6745 22083
rect 6745 22049 6779 22083
rect 6779 22049 6788 22083
rect 6736 22040 6788 22049
rect 7656 22083 7708 22092
rect 7656 22049 7665 22083
rect 7665 22049 7699 22083
rect 7699 22049 7708 22083
rect 7656 22040 7708 22049
rect 7748 22083 7800 22092
rect 7748 22049 7757 22083
rect 7757 22049 7791 22083
rect 7791 22049 7800 22083
rect 7748 22040 7800 22049
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 7564 22015 7616 22024
rect 7564 21981 7573 22015
rect 7573 21981 7607 22015
rect 7607 21981 7616 22015
rect 7564 21972 7616 21981
rect 8760 21972 8812 22024
rect 3792 21879 3844 21888
rect 3792 21845 3801 21879
rect 3801 21845 3835 21879
rect 3835 21845 3844 21879
rect 3792 21836 3844 21845
rect 4436 21836 4488 21888
rect 4712 21836 4764 21888
rect 6460 21904 6512 21956
rect 9220 21904 9272 21956
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 9588 22015 9640 22024
rect 9588 21981 9597 22015
rect 9597 21981 9631 22015
rect 9631 21981 9640 22015
rect 9588 21972 9640 21981
rect 9864 22015 9916 22024
rect 9864 21981 9873 22015
rect 9873 21981 9907 22015
rect 9907 21981 9916 22015
rect 9864 21972 9916 21981
rect 10048 21972 10100 22024
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 11152 22015 11204 22024
rect 11152 21981 11161 22015
rect 11161 21981 11195 22015
rect 11195 21981 11204 22015
rect 11152 21972 11204 21981
rect 12164 22108 12216 22160
rect 12808 22040 12860 22092
rect 14372 22108 14424 22160
rect 14556 22108 14608 22160
rect 20260 22176 20312 22228
rect 24860 22176 24912 22228
rect 27160 22176 27212 22228
rect 29368 22176 29420 22228
rect 30012 22176 30064 22228
rect 30380 22176 30432 22228
rect 15752 22108 15804 22160
rect 10600 21904 10652 21956
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 13084 22015 13136 22024
rect 13084 21981 13093 22015
rect 13093 21981 13127 22015
rect 13127 21981 13136 22015
rect 13084 21972 13136 21981
rect 12440 21904 12492 21956
rect 5448 21836 5500 21888
rect 6276 21836 6328 21888
rect 7932 21879 7984 21888
rect 7932 21845 7941 21879
rect 7941 21845 7975 21879
rect 7975 21845 7984 21879
rect 7932 21836 7984 21845
rect 8760 21836 8812 21888
rect 9404 21836 9456 21888
rect 10140 21836 10192 21888
rect 11060 21836 11112 21888
rect 11152 21836 11204 21888
rect 11612 21836 11664 21888
rect 13544 22015 13596 22024
rect 13544 21981 13553 22015
rect 13553 21981 13587 22015
rect 13587 21981 13596 22015
rect 13544 21972 13596 21981
rect 13912 21972 13964 22024
rect 14556 21972 14608 22024
rect 16028 22083 16080 22092
rect 16028 22049 16037 22083
rect 16037 22049 16071 22083
rect 16071 22049 16080 22083
rect 16028 22040 16080 22049
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 16120 22015 16172 22024
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 16764 22108 16816 22160
rect 18144 22108 18196 22160
rect 16856 22040 16908 22092
rect 17408 22040 17460 22092
rect 18972 22108 19024 22160
rect 16948 21972 17000 22024
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 18144 21972 18196 22024
rect 13820 21836 13872 21888
rect 16304 21904 16356 21956
rect 20628 22040 20680 22092
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 18788 21972 18840 21981
rect 18604 21836 18656 21888
rect 19432 21972 19484 22024
rect 22008 21904 22060 21956
rect 22928 21972 22980 22024
rect 24584 22040 24636 22092
rect 26240 22108 26292 22160
rect 24032 21972 24084 22024
rect 24124 21972 24176 22024
rect 23848 21904 23900 21956
rect 24860 22015 24912 22024
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 24860 21972 24912 21981
rect 25044 22015 25096 22024
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 24952 21904 25004 21956
rect 19340 21836 19392 21888
rect 20076 21836 20128 21888
rect 20260 21836 20312 21888
rect 23572 21836 23624 21888
rect 24032 21879 24084 21888
rect 24032 21845 24041 21879
rect 24041 21845 24075 21879
rect 24075 21845 24084 21879
rect 24032 21836 24084 21845
rect 24308 21836 24360 21888
rect 24400 21836 24452 21888
rect 25688 22015 25740 22024
rect 25688 21981 25697 22015
rect 25697 21981 25731 22015
rect 25731 21981 25740 22015
rect 25688 21972 25740 21981
rect 26148 22083 26200 22092
rect 26148 22049 26157 22083
rect 26157 22049 26191 22083
rect 26191 22049 26200 22083
rect 26148 22040 26200 22049
rect 27344 22108 27396 22160
rect 30196 22108 30248 22160
rect 31116 22176 31168 22228
rect 32220 22176 32272 22228
rect 32772 22176 32824 22228
rect 33140 22176 33192 22228
rect 36176 22176 36228 22228
rect 26884 22083 26936 22092
rect 26884 22049 26893 22083
rect 26893 22049 26927 22083
rect 26927 22049 26936 22083
rect 26884 22040 26936 22049
rect 26516 22015 26568 22024
rect 26516 21981 26525 22015
rect 26525 21981 26559 22015
rect 26559 21981 26568 22015
rect 26516 21972 26568 21981
rect 26608 22015 26660 22024
rect 26608 21981 26617 22015
rect 26617 21981 26651 22015
rect 26651 21981 26660 22015
rect 26608 21972 26660 21981
rect 26884 21904 26936 21956
rect 27160 22015 27212 22024
rect 27160 21981 27169 22015
rect 27169 21981 27203 22015
rect 27203 21981 27212 22015
rect 27160 21972 27212 21981
rect 27620 22015 27672 22024
rect 27620 21981 27629 22015
rect 27629 21981 27663 22015
rect 27663 21981 27672 22015
rect 27620 21972 27672 21981
rect 28724 21972 28776 22024
rect 30196 21972 30248 22024
rect 29368 21904 29420 21956
rect 30564 21904 30616 21956
rect 30840 22040 30892 22092
rect 34612 22040 34664 22092
rect 30932 21972 30984 22024
rect 31208 21972 31260 22024
rect 32036 21972 32088 22024
rect 35992 21972 36044 22024
rect 26056 21836 26108 21888
rect 26608 21836 26660 21888
rect 26792 21836 26844 21888
rect 28172 21836 28224 21888
rect 28356 21836 28408 21888
rect 29000 21836 29052 21888
rect 29920 21879 29972 21888
rect 29920 21845 29945 21879
rect 29945 21845 29972 21879
rect 29920 21836 29972 21845
rect 30288 21836 30340 21888
rect 31116 21836 31168 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 3792 21632 3844 21684
rect 4436 21675 4488 21684
rect 4436 21641 4445 21675
rect 4445 21641 4479 21675
rect 4479 21641 4488 21675
rect 4436 21632 4488 21641
rect 4620 21632 4672 21684
rect 6368 21632 6420 21684
rect 7932 21632 7984 21684
rect 9772 21632 9824 21684
rect 10692 21632 10744 21684
rect 12072 21632 12124 21684
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 14372 21632 14424 21684
rect 15844 21632 15896 21684
rect 16488 21632 16540 21684
rect 19432 21632 19484 21684
rect 19616 21632 19668 21684
rect 20720 21632 20772 21684
rect 21824 21675 21876 21684
rect 21824 21641 21833 21675
rect 21833 21641 21867 21675
rect 21867 21641 21876 21675
rect 21824 21632 21876 21641
rect 22284 21632 22336 21684
rect 22744 21675 22796 21684
rect 22744 21641 22753 21675
rect 22753 21641 22787 21675
rect 22787 21641 22796 21675
rect 22744 21632 22796 21641
rect 24492 21632 24544 21684
rect 1400 21496 1452 21548
rect 5264 21564 5316 21616
rect 2964 21428 3016 21480
rect 4528 21539 4580 21548
rect 4528 21505 4537 21539
rect 4537 21505 4571 21539
rect 4571 21505 4580 21539
rect 4528 21496 4580 21505
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 3332 21428 3384 21480
rect 3884 21360 3936 21412
rect 5540 21496 5592 21548
rect 5632 21496 5684 21548
rect 7104 21496 7156 21548
rect 9128 21564 9180 21616
rect 8300 21496 8352 21548
rect 8760 21539 8812 21548
rect 8760 21505 8769 21539
rect 8769 21505 8803 21539
rect 8803 21505 8812 21539
rect 8760 21496 8812 21505
rect 9220 21539 9272 21548
rect 9220 21505 9229 21539
rect 9229 21505 9263 21539
rect 9263 21505 9272 21539
rect 9220 21496 9272 21505
rect 9312 21496 9364 21548
rect 9956 21564 10008 21616
rect 6644 21360 6696 21412
rect 9588 21360 9640 21412
rect 10600 21496 10652 21548
rect 10876 21564 10928 21616
rect 11060 21539 11112 21548
rect 11060 21505 11069 21539
rect 11069 21505 11103 21539
rect 11103 21505 11112 21539
rect 11060 21496 11112 21505
rect 16948 21607 17000 21616
rect 11336 21539 11388 21546
rect 11336 21505 11339 21539
rect 11339 21505 11373 21539
rect 11373 21505 11388 21539
rect 11336 21494 11388 21505
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 14096 21496 14148 21548
rect 10600 21360 10652 21412
rect 12072 21471 12124 21480
rect 12072 21437 12081 21471
rect 12081 21437 12115 21471
rect 12115 21437 12124 21471
rect 12072 21428 12124 21437
rect 11612 21403 11664 21412
rect 11612 21369 11621 21403
rect 11621 21369 11655 21403
rect 11655 21369 11664 21403
rect 11612 21360 11664 21369
rect 16948 21573 16957 21607
rect 16957 21573 16991 21607
rect 16991 21573 17000 21607
rect 16948 21564 17000 21573
rect 17040 21607 17092 21616
rect 17040 21573 17049 21607
rect 17049 21573 17083 21607
rect 17083 21573 17092 21607
rect 17040 21564 17092 21573
rect 17408 21564 17460 21616
rect 14556 21496 14608 21548
rect 15108 21496 15160 21548
rect 16212 21496 16264 21548
rect 16672 21496 16724 21548
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17316 21496 17368 21548
rect 19248 21564 19300 21616
rect 17868 21496 17920 21548
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18236 21496 18288 21505
rect 18788 21496 18840 21548
rect 13084 21428 13136 21480
rect 14372 21428 14424 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 16304 21360 16356 21412
rect 17040 21360 17092 21412
rect 17316 21360 17368 21412
rect 18420 21428 18472 21480
rect 21272 21564 21324 21616
rect 22192 21607 22244 21616
rect 22192 21573 22201 21607
rect 22201 21573 22235 21607
rect 22235 21573 22244 21607
rect 22192 21564 22244 21573
rect 23572 21564 23624 21616
rect 23848 21564 23900 21616
rect 25596 21632 25648 21684
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 20352 21496 20404 21505
rect 20536 21496 20588 21548
rect 20996 21496 21048 21548
rect 22560 21496 22612 21548
rect 24216 21496 24268 21548
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 24676 21496 24728 21548
rect 19524 21428 19576 21480
rect 10232 21292 10284 21344
rect 14924 21292 14976 21344
rect 15660 21292 15712 21344
rect 16948 21292 17000 21344
rect 18328 21292 18380 21344
rect 18788 21335 18840 21344
rect 18788 21301 18797 21335
rect 18797 21301 18831 21335
rect 18831 21301 18840 21335
rect 18788 21292 18840 21301
rect 19156 21292 19208 21344
rect 19432 21292 19484 21344
rect 20444 21428 20496 21480
rect 23112 21360 23164 21412
rect 23848 21471 23900 21480
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 20352 21292 20404 21344
rect 20444 21292 20496 21344
rect 20628 21292 20680 21344
rect 24032 21292 24084 21344
rect 24492 21335 24544 21344
rect 24492 21301 24501 21335
rect 24501 21301 24535 21335
rect 24535 21301 24544 21335
rect 24492 21292 24544 21301
rect 24952 21292 25004 21344
rect 25228 21360 25280 21412
rect 27344 21564 27396 21616
rect 28080 21564 28132 21616
rect 28632 21632 28684 21684
rect 30288 21632 30340 21684
rect 31760 21632 31812 21684
rect 30564 21564 30616 21616
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 27252 21428 27304 21480
rect 27436 21428 27488 21480
rect 29000 21496 29052 21548
rect 29184 21496 29236 21548
rect 29920 21496 29972 21548
rect 35532 21496 35584 21548
rect 30656 21428 30708 21480
rect 31392 21428 31444 21480
rect 29552 21360 29604 21412
rect 30840 21360 30892 21412
rect 31024 21360 31076 21412
rect 31300 21360 31352 21412
rect 33416 21360 33468 21412
rect 26976 21335 27028 21344
rect 26976 21301 26985 21335
rect 26985 21301 27019 21335
rect 27019 21301 27028 21335
rect 26976 21292 27028 21301
rect 31116 21292 31168 21344
rect 32036 21292 32088 21344
rect 32864 21292 32916 21344
rect 35348 21292 35400 21344
rect 35716 21292 35768 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5724 21131 5776 21140
rect 5724 21097 5733 21131
rect 5733 21097 5767 21131
rect 5767 21097 5776 21131
rect 5724 21088 5776 21097
rect 7012 21088 7064 21140
rect 7472 21088 7524 21140
rect 4068 20952 4120 21004
rect 2872 20884 2924 20936
rect 1676 20748 1728 20800
rect 2872 20791 2924 20800
rect 2872 20757 2881 20791
rect 2881 20757 2915 20791
rect 2915 20757 2924 20791
rect 2872 20748 2924 20757
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 4620 20884 4672 20936
rect 4712 20927 4764 20936
rect 4712 20893 4721 20927
rect 4721 20893 4755 20927
rect 4755 20893 4764 20927
rect 4712 20884 4764 20893
rect 4896 21020 4948 21072
rect 6552 21020 6604 21072
rect 5356 20927 5408 20936
rect 5356 20893 5365 20927
rect 5365 20893 5399 20927
rect 5399 20893 5408 20927
rect 5356 20884 5408 20893
rect 7380 20952 7432 21004
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 5632 20927 5684 20936
rect 5632 20893 5641 20927
rect 5641 20893 5675 20927
rect 5675 20893 5684 20927
rect 5632 20884 5684 20893
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 7012 20927 7064 20936
rect 7012 20893 7021 20927
rect 7021 20893 7055 20927
rect 7055 20893 7064 20927
rect 7012 20884 7064 20893
rect 7196 20927 7248 20936
rect 7196 20893 7205 20927
rect 7205 20893 7239 20927
rect 7239 20893 7248 20927
rect 7196 20884 7248 20893
rect 7748 20995 7800 21004
rect 7748 20961 7757 20995
rect 7757 20961 7791 20995
rect 7791 20961 7800 20995
rect 7748 20952 7800 20961
rect 8024 21088 8076 21140
rect 10508 21088 10560 21140
rect 11060 21088 11112 21140
rect 11612 21088 11664 21140
rect 13360 21088 13412 21140
rect 15568 21088 15620 21140
rect 8300 20952 8352 21004
rect 8760 20952 8812 21004
rect 9036 20952 9088 21004
rect 10232 20995 10284 21004
rect 10232 20961 10241 20995
rect 10241 20961 10275 20995
rect 10275 20961 10284 20995
rect 10232 20952 10284 20961
rect 10508 20952 10560 21004
rect 11152 20995 11204 21004
rect 11152 20961 11161 20995
rect 11161 20961 11195 20995
rect 11195 20961 11204 20995
rect 11152 20952 11204 20961
rect 11520 21020 11572 21072
rect 12256 21020 12308 21072
rect 13452 21020 13504 21072
rect 17776 21088 17828 21140
rect 18144 21088 18196 21140
rect 18328 21088 18380 21140
rect 18880 21088 18932 21140
rect 19524 21088 19576 21140
rect 19800 21088 19852 21140
rect 20536 21131 20588 21140
rect 20536 21097 20545 21131
rect 20545 21097 20579 21131
rect 20579 21097 20588 21131
rect 20536 21088 20588 21097
rect 5908 20816 5960 20868
rect 3516 20748 3568 20800
rect 3792 20791 3844 20800
rect 3792 20757 3801 20791
rect 3801 20757 3835 20791
rect 3835 20757 3844 20791
rect 3792 20748 3844 20757
rect 5264 20748 5316 20800
rect 7380 20748 7432 20800
rect 8760 20816 8812 20868
rect 9220 20884 9272 20936
rect 9864 20884 9916 20936
rect 10048 20927 10100 20936
rect 10048 20893 10057 20927
rect 10057 20893 10091 20927
rect 10091 20893 10100 20927
rect 10048 20884 10100 20893
rect 10876 20884 10928 20936
rect 11612 20884 11664 20936
rect 14004 20952 14056 21004
rect 10416 20816 10468 20868
rect 12992 20884 13044 20936
rect 13268 20884 13320 20936
rect 13360 20884 13412 20936
rect 15476 20927 15528 20936
rect 15476 20893 15485 20927
rect 15485 20893 15519 20927
rect 15519 20893 15528 20927
rect 15476 20884 15528 20893
rect 16212 20995 16264 21004
rect 16212 20961 16221 20995
rect 16221 20961 16255 20995
rect 16255 20961 16264 20995
rect 16212 20952 16264 20961
rect 13084 20816 13136 20868
rect 14924 20816 14976 20868
rect 15568 20859 15620 20868
rect 15568 20825 15577 20859
rect 15577 20825 15611 20859
rect 15611 20825 15620 20859
rect 15568 20816 15620 20825
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 18052 20952 18104 21004
rect 17224 20927 17276 20936
rect 17224 20893 17233 20927
rect 17233 20893 17267 20927
rect 17267 20893 17276 20927
rect 17224 20884 17276 20893
rect 18420 21020 18472 21072
rect 22652 21088 22704 21140
rect 22836 21088 22888 21140
rect 23480 21088 23532 21140
rect 24124 21088 24176 21140
rect 26976 21088 27028 21140
rect 28724 21088 28776 21140
rect 20812 21020 20864 21072
rect 17500 20859 17552 20868
rect 17500 20825 17509 20859
rect 17509 20825 17543 20859
rect 17543 20825 17552 20859
rect 17500 20816 17552 20825
rect 17592 20859 17644 20868
rect 17592 20825 17601 20859
rect 17601 20825 17635 20859
rect 17635 20825 17644 20859
rect 17592 20816 17644 20825
rect 18144 20927 18196 20936
rect 18144 20893 18153 20927
rect 18153 20893 18187 20927
rect 18187 20893 18196 20927
rect 18144 20884 18196 20893
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 18328 20927 18380 20936
rect 18328 20893 18337 20927
rect 18337 20893 18371 20927
rect 18371 20893 18380 20927
rect 18328 20884 18380 20893
rect 19248 20995 19300 21004
rect 19248 20961 19257 20995
rect 19257 20961 19291 20995
rect 19291 20961 19300 20995
rect 19248 20952 19300 20961
rect 18972 20884 19024 20936
rect 19340 20884 19392 20936
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 19616 20927 19668 20936
rect 19616 20893 19625 20927
rect 19625 20893 19659 20927
rect 19659 20893 19668 20927
rect 19616 20884 19668 20893
rect 19708 20927 19760 20936
rect 19708 20893 19717 20927
rect 19717 20893 19751 20927
rect 19751 20893 19760 20927
rect 19708 20884 19760 20893
rect 20628 20952 20680 21004
rect 20076 20927 20128 20936
rect 20076 20893 20083 20927
rect 20083 20893 20128 20927
rect 20076 20884 20128 20893
rect 21640 20952 21692 21004
rect 22008 20995 22060 21004
rect 22008 20961 22017 20995
rect 22017 20961 22051 20995
rect 22051 20961 22060 20995
rect 22008 20952 22060 20961
rect 20904 20884 20956 20936
rect 21916 20884 21968 20936
rect 22376 20884 22428 20936
rect 22560 20927 22612 20936
rect 26516 21020 26568 21072
rect 22560 20893 22594 20927
rect 22594 20893 22612 20927
rect 22560 20884 22612 20893
rect 18788 20816 18840 20868
rect 8024 20791 8076 20800
rect 8024 20757 8033 20791
rect 8033 20757 8067 20791
rect 8067 20757 8076 20791
rect 8024 20748 8076 20757
rect 8208 20748 8260 20800
rect 9312 20748 9364 20800
rect 9496 20791 9548 20800
rect 9496 20757 9505 20791
rect 9505 20757 9539 20791
rect 9539 20757 9548 20791
rect 9496 20748 9548 20757
rect 9588 20791 9640 20800
rect 9588 20757 9597 20791
rect 9597 20757 9631 20791
rect 9631 20757 9640 20791
rect 9588 20748 9640 20757
rect 11152 20748 11204 20800
rect 11796 20748 11848 20800
rect 13636 20748 13688 20800
rect 14188 20748 14240 20800
rect 14372 20791 14424 20800
rect 14372 20757 14381 20791
rect 14381 20757 14415 20791
rect 14415 20757 14424 20791
rect 14372 20748 14424 20757
rect 14832 20748 14884 20800
rect 15200 20748 15252 20800
rect 15752 20748 15804 20800
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 16396 20791 16448 20800
rect 16396 20757 16405 20791
rect 16405 20757 16439 20791
rect 16439 20757 16448 20791
rect 16396 20748 16448 20757
rect 17868 20748 17920 20800
rect 20168 20859 20220 20868
rect 20168 20825 20177 20859
rect 20177 20825 20211 20859
rect 20211 20825 20220 20859
rect 20168 20816 20220 20825
rect 21180 20816 21232 20868
rect 20352 20748 20404 20800
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 27896 20884 27948 20936
rect 29184 21020 29236 21072
rect 28448 20952 28500 21004
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 28724 20884 28776 20936
rect 29000 20884 29052 20936
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 29736 20927 29788 20936
rect 29736 20893 29753 20927
rect 29753 20893 29788 20927
rect 29736 20884 29788 20893
rect 31024 21088 31076 21140
rect 31392 21088 31444 21140
rect 33416 21088 33468 21140
rect 29920 21020 29972 21072
rect 30380 20952 30432 21004
rect 31484 20952 31536 21004
rect 28448 20859 28500 20868
rect 28448 20825 28483 20859
rect 28483 20825 28500 20859
rect 28448 20816 28500 20825
rect 23020 20791 23072 20800
rect 23020 20757 23029 20791
rect 23029 20757 23063 20791
rect 23063 20757 23072 20791
rect 23020 20748 23072 20757
rect 23112 20791 23164 20800
rect 23112 20757 23121 20791
rect 23121 20757 23155 20791
rect 23155 20757 23164 20791
rect 23112 20748 23164 20757
rect 27988 20791 28040 20800
rect 27988 20757 27997 20791
rect 27997 20757 28031 20791
rect 28031 20757 28040 20791
rect 27988 20748 28040 20757
rect 29368 20748 29420 20800
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 30196 20816 30248 20868
rect 30564 20859 30616 20868
rect 30564 20825 30573 20859
rect 30573 20825 30607 20859
rect 30607 20825 30616 20859
rect 30564 20816 30616 20825
rect 30840 20816 30892 20868
rect 31576 20884 31628 20936
rect 31760 20884 31812 20936
rect 31024 20748 31076 20800
rect 32128 20816 32180 20868
rect 33692 21020 33744 21072
rect 32680 20952 32732 21004
rect 33416 20952 33468 21004
rect 33784 20952 33836 21004
rect 34244 20952 34296 21004
rect 34520 20952 34572 21004
rect 34796 20952 34848 21004
rect 33232 20884 33284 20936
rect 35348 20952 35400 21004
rect 34980 20927 35032 20936
rect 34980 20893 34989 20927
rect 34989 20893 35023 20927
rect 35023 20893 35032 20927
rect 34980 20884 35032 20893
rect 33140 20816 33192 20868
rect 31576 20748 31628 20800
rect 31668 20791 31720 20800
rect 31668 20757 31677 20791
rect 31677 20757 31711 20791
rect 31711 20757 31720 20791
rect 31668 20748 31720 20757
rect 32864 20791 32916 20800
rect 32864 20757 32873 20791
rect 32873 20757 32907 20791
rect 32907 20757 32916 20791
rect 32864 20748 32916 20757
rect 34520 20816 34572 20868
rect 35716 20927 35768 20936
rect 35716 20893 35725 20927
rect 35725 20893 35759 20927
rect 35759 20893 35768 20927
rect 35716 20884 35768 20893
rect 33600 20748 33652 20800
rect 34704 20791 34756 20800
rect 34704 20757 34713 20791
rect 34713 20757 34747 20791
rect 34747 20757 34756 20791
rect 34704 20748 34756 20757
rect 35440 20748 35492 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 2504 20544 2556 20596
rect 3792 20587 3844 20596
rect 3792 20553 3801 20587
rect 3801 20553 3835 20587
rect 3835 20553 3844 20587
rect 3792 20544 3844 20553
rect 4344 20544 4396 20596
rect 5080 20544 5132 20596
rect 5632 20544 5684 20596
rect 5816 20544 5868 20596
rect 7564 20544 7616 20596
rect 8024 20544 8076 20596
rect 1400 20408 1452 20460
rect 2964 20408 3016 20460
rect 3884 20383 3936 20392
rect 3884 20349 3893 20383
rect 3893 20349 3927 20383
rect 3927 20349 3936 20383
rect 3884 20340 3936 20349
rect 4068 20383 4120 20392
rect 4068 20349 4077 20383
rect 4077 20349 4111 20383
rect 4111 20349 4120 20383
rect 4068 20340 4120 20349
rect 4712 20451 4764 20460
rect 4712 20417 4721 20451
rect 4721 20417 4755 20451
rect 4755 20417 4764 20451
rect 4712 20408 4764 20417
rect 4804 20408 4856 20460
rect 5264 20408 5316 20460
rect 5724 20519 5776 20528
rect 5724 20485 5733 20519
rect 5733 20485 5767 20519
rect 5767 20485 5776 20519
rect 5724 20476 5776 20485
rect 6552 20476 6604 20528
rect 6736 20476 6788 20528
rect 7104 20519 7156 20528
rect 7104 20485 7113 20519
rect 7113 20485 7147 20519
rect 7147 20485 7156 20519
rect 7104 20476 7156 20485
rect 7472 20476 7524 20528
rect 8300 20476 8352 20528
rect 5080 20340 5132 20392
rect 4896 20272 4948 20324
rect 5908 20408 5960 20460
rect 6644 20451 6696 20460
rect 6644 20417 6653 20451
rect 6653 20417 6687 20451
rect 6687 20417 6696 20451
rect 6644 20408 6696 20417
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 6920 20451 6972 20460
rect 6920 20417 6929 20451
rect 6929 20417 6963 20451
rect 6963 20417 6972 20451
rect 6920 20408 6972 20417
rect 8576 20408 8628 20460
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 9496 20476 9548 20528
rect 13268 20519 13320 20528
rect 13268 20485 13277 20519
rect 13277 20485 13311 20519
rect 13311 20485 13320 20519
rect 13268 20476 13320 20485
rect 13728 20476 13780 20528
rect 15200 20544 15252 20596
rect 15568 20544 15620 20596
rect 17040 20587 17092 20596
rect 17040 20553 17049 20587
rect 17049 20553 17083 20587
rect 17083 20553 17092 20587
rect 17040 20544 17092 20553
rect 17592 20544 17644 20596
rect 16304 20476 16356 20528
rect 17776 20544 17828 20596
rect 18236 20544 18288 20596
rect 20812 20587 20864 20596
rect 20812 20553 20821 20587
rect 20821 20553 20855 20587
rect 20855 20553 20864 20587
rect 20812 20544 20864 20553
rect 22192 20544 22244 20596
rect 9772 20408 9824 20460
rect 10968 20408 11020 20460
rect 11612 20408 11664 20460
rect 13636 20451 13688 20460
rect 13636 20417 13645 20451
rect 13645 20417 13679 20451
rect 13679 20417 13688 20451
rect 13636 20408 13688 20417
rect 15568 20408 15620 20460
rect 16028 20451 16080 20460
rect 16028 20417 16037 20451
rect 16037 20417 16071 20451
rect 16071 20417 16080 20451
rect 16028 20408 16080 20417
rect 16120 20408 16172 20460
rect 8208 20340 8260 20392
rect 6736 20272 6788 20324
rect 7196 20272 7248 20324
rect 8116 20272 8168 20324
rect 12532 20383 12584 20392
rect 12532 20349 12541 20383
rect 12541 20349 12575 20383
rect 12575 20349 12584 20383
rect 12532 20340 12584 20349
rect 13820 20340 13872 20392
rect 14004 20383 14056 20392
rect 14004 20349 14013 20383
rect 14013 20349 14047 20383
rect 14047 20349 14056 20383
rect 14004 20340 14056 20349
rect 14648 20340 14700 20392
rect 15752 20340 15804 20392
rect 18052 20408 18104 20460
rect 18512 20519 18564 20528
rect 18512 20485 18537 20519
rect 18537 20485 18564 20519
rect 18512 20476 18564 20485
rect 18788 20519 18840 20528
rect 18788 20485 18797 20519
rect 18797 20485 18831 20519
rect 18831 20485 18840 20519
rect 18788 20476 18840 20485
rect 20168 20476 20220 20528
rect 19064 20408 19116 20460
rect 20076 20408 20128 20460
rect 20352 20408 20404 20460
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 17224 20272 17276 20324
rect 19708 20340 19760 20392
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 4344 20204 4396 20256
rect 4528 20204 4580 20256
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 7104 20204 7156 20256
rect 9588 20204 9640 20256
rect 11428 20204 11480 20256
rect 13636 20204 13688 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 18788 20272 18840 20324
rect 20720 20272 20772 20324
rect 21180 20408 21232 20460
rect 21548 20451 21600 20460
rect 21548 20417 21557 20451
rect 21557 20417 21591 20451
rect 21591 20417 21600 20451
rect 21548 20408 21600 20417
rect 22008 20408 22060 20460
rect 21640 20340 21692 20392
rect 23112 20544 23164 20596
rect 22836 20476 22888 20528
rect 23296 20476 23348 20528
rect 22652 20408 22704 20460
rect 23480 20408 23532 20460
rect 23020 20340 23072 20392
rect 23296 20340 23348 20392
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 24768 20451 24820 20460
rect 24768 20417 24777 20451
rect 24777 20417 24811 20451
rect 24811 20417 24820 20451
rect 24768 20408 24820 20417
rect 25044 20451 25096 20460
rect 25044 20417 25053 20451
rect 25053 20417 25087 20451
rect 25087 20417 25096 20451
rect 25044 20408 25096 20417
rect 26608 20544 26660 20596
rect 27896 20544 27948 20596
rect 28724 20544 28776 20596
rect 26884 20476 26936 20528
rect 26608 20408 26660 20460
rect 27344 20408 27396 20460
rect 27896 20408 27948 20460
rect 28264 20476 28316 20528
rect 28724 20408 28776 20460
rect 24216 20340 24268 20392
rect 21088 20272 21140 20324
rect 21272 20315 21324 20324
rect 21272 20281 21281 20315
rect 21281 20281 21315 20315
rect 21315 20281 21324 20315
rect 21272 20272 21324 20281
rect 21456 20272 21508 20324
rect 19432 20204 19484 20256
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 23296 20204 23348 20256
rect 23480 20204 23532 20256
rect 23664 20204 23716 20256
rect 24032 20272 24084 20324
rect 25320 20340 25372 20392
rect 27436 20383 27488 20392
rect 27436 20349 27445 20383
rect 27445 20349 27479 20383
rect 27479 20349 27488 20383
rect 27436 20340 27488 20349
rect 28632 20340 28684 20392
rect 29644 20476 29696 20528
rect 29092 20408 29144 20460
rect 29828 20451 29880 20460
rect 29828 20417 29837 20451
rect 29837 20417 29871 20451
rect 29871 20417 29880 20451
rect 29828 20408 29880 20417
rect 30288 20476 30340 20528
rect 30196 20408 30248 20460
rect 30840 20451 30892 20460
rect 30840 20417 30849 20451
rect 30849 20417 30883 20451
rect 30883 20417 30892 20451
rect 30840 20408 30892 20417
rect 30288 20340 30340 20392
rect 30748 20340 30800 20392
rect 31116 20383 31168 20392
rect 31116 20349 31125 20383
rect 31125 20349 31159 20383
rect 31159 20349 31168 20383
rect 31116 20340 31168 20349
rect 31392 20340 31444 20392
rect 25136 20315 25188 20324
rect 25136 20281 25145 20315
rect 25145 20281 25179 20315
rect 25179 20281 25188 20315
rect 25136 20272 25188 20281
rect 25780 20272 25832 20324
rect 28816 20272 28868 20324
rect 29092 20272 29144 20324
rect 29828 20272 29880 20324
rect 24860 20204 24912 20256
rect 26240 20204 26292 20256
rect 27620 20247 27672 20256
rect 27620 20213 27629 20247
rect 27629 20213 27663 20247
rect 27663 20213 27672 20247
rect 27620 20204 27672 20213
rect 27804 20204 27856 20256
rect 28448 20204 28500 20256
rect 29184 20204 29236 20256
rect 30840 20272 30892 20324
rect 30104 20247 30156 20256
rect 30104 20213 30113 20247
rect 30113 20213 30147 20247
rect 30147 20213 30156 20247
rect 30104 20204 30156 20213
rect 30656 20247 30708 20256
rect 30656 20213 30665 20247
rect 30665 20213 30699 20247
rect 30699 20213 30708 20247
rect 30656 20204 30708 20213
rect 31484 20204 31536 20256
rect 32312 20408 32364 20460
rect 33232 20476 33284 20528
rect 32864 20451 32916 20460
rect 32864 20417 32873 20451
rect 32873 20417 32907 20451
rect 32907 20417 32916 20451
rect 32864 20408 32916 20417
rect 31668 20340 31720 20392
rect 33692 20408 33744 20460
rect 33876 20451 33928 20460
rect 33876 20417 33885 20451
rect 33885 20417 33919 20451
rect 33919 20417 33928 20451
rect 33876 20408 33928 20417
rect 34428 20408 34480 20460
rect 34796 20451 34848 20460
rect 34796 20417 34805 20451
rect 34805 20417 34839 20451
rect 34839 20417 34848 20451
rect 34796 20408 34848 20417
rect 35256 20340 35308 20392
rect 35532 20340 35584 20392
rect 33140 20272 33192 20324
rect 33692 20272 33744 20324
rect 31668 20204 31720 20256
rect 31852 20204 31904 20256
rect 32404 20247 32456 20256
rect 32404 20213 32413 20247
rect 32413 20213 32447 20247
rect 32447 20213 32456 20247
rect 32404 20204 32456 20213
rect 32588 20247 32640 20256
rect 32588 20213 32597 20247
rect 32597 20213 32631 20247
rect 32631 20213 32640 20247
rect 32588 20204 32640 20213
rect 34704 20247 34756 20256
rect 34704 20213 34713 20247
rect 34713 20213 34747 20247
rect 34747 20213 34756 20247
rect 34704 20204 34756 20213
rect 35348 20204 35400 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2872 20000 2924 20052
rect 4620 20000 4672 20052
rect 5356 20000 5408 20052
rect 5908 20000 5960 20052
rect 7012 20000 7064 20052
rect 7748 20000 7800 20052
rect 12532 20000 12584 20052
rect 13268 20000 13320 20052
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 1676 19907 1728 19916
rect 1676 19873 1685 19907
rect 1685 19873 1719 19907
rect 1719 19873 1728 19907
rect 1676 19864 1728 19873
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 4804 19932 4856 19984
rect 6092 19932 6144 19984
rect 6276 19932 6328 19984
rect 9680 19932 9732 19984
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 15292 20000 15344 20052
rect 17132 20000 17184 20052
rect 18052 20000 18104 20052
rect 18512 20000 18564 20052
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 20168 20000 20220 20052
rect 23940 20000 23992 20052
rect 24860 20000 24912 20052
rect 2964 19728 3016 19780
rect 4252 19728 4304 19780
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 7104 19864 7156 19916
rect 8024 19864 8076 19916
rect 8116 19907 8168 19916
rect 8116 19873 8125 19907
rect 8125 19873 8159 19907
rect 8159 19873 8168 19907
rect 8116 19864 8168 19873
rect 11244 19907 11296 19916
rect 11244 19873 11253 19907
rect 11253 19873 11287 19907
rect 11287 19873 11296 19907
rect 11244 19864 11296 19873
rect 13636 19907 13688 19916
rect 13636 19873 13645 19907
rect 13645 19873 13679 19907
rect 13679 19873 13688 19907
rect 13636 19864 13688 19873
rect 6828 19796 6880 19848
rect 10416 19796 10468 19848
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 12348 19796 12400 19848
rect 14004 19796 14056 19848
rect 6644 19728 6696 19780
rect 8300 19728 8352 19780
rect 9036 19728 9088 19780
rect 13728 19728 13780 19780
rect 14188 19796 14240 19848
rect 14924 19932 14976 19984
rect 16672 19932 16724 19984
rect 17960 19932 18012 19984
rect 18144 19932 18196 19984
rect 20536 19932 20588 19984
rect 20628 19932 20680 19984
rect 21180 19932 21232 19984
rect 23664 19932 23716 19984
rect 14648 19796 14700 19848
rect 14832 19796 14884 19848
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15568 19796 15620 19848
rect 16304 19839 16356 19848
rect 16304 19805 16335 19839
rect 16335 19805 16356 19839
rect 16304 19796 16356 19805
rect 3884 19660 3936 19712
rect 6276 19660 6328 19712
rect 7104 19660 7156 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 11980 19660 12032 19712
rect 13820 19660 13872 19712
rect 15752 19728 15804 19780
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 17500 19796 17552 19848
rect 17868 19796 17920 19848
rect 18512 19796 18564 19848
rect 23664 19796 23716 19848
rect 25872 19932 25924 19984
rect 29828 20000 29880 20052
rect 29920 20000 29972 20052
rect 31668 20000 31720 20052
rect 35348 20000 35400 20052
rect 35532 20000 35584 20052
rect 25412 19907 25464 19916
rect 25412 19873 25421 19907
rect 25421 19873 25455 19907
rect 25455 19873 25464 19907
rect 25412 19864 25464 19873
rect 27712 19864 27764 19916
rect 28264 19932 28316 19984
rect 18052 19728 18104 19780
rect 19800 19771 19852 19780
rect 19800 19737 19809 19771
rect 19809 19737 19843 19771
rect 19843 19737 19852 19771
rect 19800 19728 19852 19737
rect 14832 19660 14884 19712
rect 19708 19660 19760 19712
rect 20812 19728 20864 19780
rect 21180 19728 21232 19780
rect 21640 19728 21692 19780
rect 24216 19796 24268 19848
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 24584 19839 24636 19848
rect 24584 19805 24593 19839
rect 24593 19805 24627 19839
rect 24627 19805 24636 19839
rect 24584 19796 24636 19805
rect 24952 19796 25004 19848
rect 26240 19796 26292 19848
rect 26884 19839 26936 19848
rect 26884 19805 26893 19839
rect 26893 19805 26927 19839
rect 26927 19805 26936 19839
rect 26884 19796 26936 19805
rect 27528 19796 27580 19848
rect 29736 19796 29788 19848
rect 30472 19796 30524 19848
rect 31300 19839 31352 19848
rect 31300 19805 31309 19839
rect 31309 19805 31343 19839
rect 31343 19805 31352 19839
rect 31300 19796 31352 19805
rect 34704 19796 34756 19848
rect 21088 19660 21140 19712
rect 21272 19660 21324 19712
rect 21824 19660 21876 19712
rect 25228 19728 25280 19780
rect 25780 19660 25832 19712
rect 26516 19703 26568 19712
rect 26516 19669 26525 19703
rect 26525 19669 26559 19703
rect 26559 19669 26568 19703
rect 26516 19660 26568 19669
rect 32680 19728 32732 19780
rect 28724 19660 28776 19712
rect 31300 19660 31352 19712
rect 34428 19660 34480 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 2688 19456 2740 19508
rect 8484 19456 8536 19508
rect 9404 19456 9456 19508
rect 10416 19456 10468 19508
rect 17224 19456 17276 19508
rect 3240 19431 3292 19440
rect 3240 19397 3249 19431
rect 3249 19397 3283 19431
rect 3283 19397 3292 19431
rect 3240 19388 3292 19397
rect 3424 19388 3476 19440
rect 5172 19388 5224 19440
rect 10048 19388 10100 19440
rect 11428 19388 11480 19440
rect 12348 19431 12400 19440
rect 12348 19397 12357 19431
rect 12357 19397 12391 19431
rect 12391 19397 12400 19431
rect 12348 19388 12400 19397
rect 13544 19388 13596 19440
rect 16580 19388 16632 19440
rect 4252 19363 4304 19372
rect 4252 19329 4261 19363
rect 4261 19329 4295 19363
rect 4295 19329 4304 19363
rect 4252 19320 4304 19329
rect 4712 19320 4764 19372
rect 5264 19320 5316 19372
rect 7012 19320 7064 19372
rect 10692 19320 10744 19372
rect 2964 19252 3016 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 10324 19252 10376 19304
rect 3700 19184 3752 19236
rect 8392 19184 8444 19236
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 16488 19320 16540 19372
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 17592 19388 17644 19440
rect 18328 19456 18380 19508
rect 19432 19456 19484 19508
rect 20812 19456 20864 19508
rect 21548 19456 21600 19508
rect 23756 19499 23808 19508
rect 23756 19465 23765 19499
rect 23765 19465 23799 19499
rect 23799 19465 23808 19499
rect 23756 19456 23808 19465
rect 24400 19456 24452 19508
rect 24768 19456 24820 19508
rect 27436 19456 27488 19508
rect 27712 19456 27764 19508
rect 12624 19252 12676 19304
rect 14648 19252 14700 19304
rect 17408 19252 17460 19304
rect 2780 19159 2832 19168
rect 2780 19125 2789 19159
rect 2789 19125 2823 19159
rect 2823 19125 2832 19159
rect 2780 19116 2832 19125
rect 4620 19116 4672 19168
rect 12164 19116 12216 19168
rect 16948 19116 17000 19168
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 17960 19252 18012 19304
rect 18144 19363 18196 19372
rect 18144 19329 18153 19363
rect 18153 19329 18187 19363
rect 18187 19329 18196 19363
rect 18144 19320 18196 19329
rect 18328 19363 18380 19372
rect 18328 19329 18335 19363
rect 18335 19329 18380 19363
rect 18328 19320 18380 19329
rect 18144 19184 18196 19236
rect 18236 19184 18288 19236
rect 18512 19363 18564 19372
rect 18512 19329 18521 19363
rect 18521 19329 18555 19363
rect 18555 19329 18564 19363
rect 18512 19320 18564 19329
rect 18788 19320 18840 19372
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19064 19363 19116 19372
rect 19064 19329 19073 19363
rect 19073 19329 19107 19363
rect 19107 19329 19116 19363
rect 19064 19320 19116 19329
rect 19248 19388 19300 19440
rect 19248 19252 19300 19304
rect 19524 19320 19576 19372
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 20904 19388 20956 19440
rect 21732 19388 21784 19440
rect 22836 19388 22888 19440
rect 20628 19252 20680 19304
rect 21456 19320 21508 19372
rect 21824 19320 21876 19372
rect 23940 19320 23992 19372
rect 24400 19363 24452 19372
rect 24400 19329 24409 19363
rect 24409 19329 24443 19363
rect 24443 19329 24452 19363
rect 24400 19320 24452 19329
rect 24492 19320 24544 19372
rect 25320 19388 25372 19440
rect 25596 19388 25648 19440
rect 24860 19363 24912 19372
rect 24860 19329 24869 19363
rect 24869 19329 24903 19363
rect 24903 19329 24912 19363
rect 24860 19320 24912 19329
rect 25044 19320 25096 19372
rect 25228 19363 25280 19372
rect 25228 19329 25237 19363
rect 25237 19329 25271 19363
rect 25271 19329 25280 19363
rect 25228 19320 25280 19329
rect 25412 19363 25464 19372
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 25504 19363 25556 19372
rect 25504 19329 25513 19363
rect 25513 19329 25547 19363
rect 25547 19329 25556 19363
rect 25504 19320 25556 19329
rect 25780 19320 25832 19372
rect 26884 19320 26936 19372
rect 27988 19320 28040 19372
rect 28356 19363 28408 19372
rect 28356 19329 28366 19363
rect 28366 19329 28400 19363
rect 28400 19329 28408 19363
rect 28356 19320 28408 19329
rect 25136 19252 25188 19304
rect 27252 19295 27304 19304
rect 27252 19261 27261 19295
rect 27261 19261 27295 19295
rect 27295 19261 27304 19295
rect 27252 19252 27304 19261
rect 27896 19252 27948 19304
rect 28172 19252 28224 19304
rect 21456 19184 21508 19236
rect 23480 19184 23532 19236
rect 26240 19184 26292 19236
rect 26332 19184 26384 19236
rect 28540 19184 28592 19236
rect 28724 19363 28776 19372
rect 29736 19431 29788 19440
rect 29736 19397 29745 19431
rect 29745 19397 29779 19431
rect 29779 19397 29788 19431
rect 29736 19388 29788 19397
rect 30748 19456 30800 19508
rect 32128 19456 32180 19508
rect 30472 19431 30524 19440
rect 30472 19397 30481 19431
rect 30481 19397 30515 19431
rect 30515 19397 30524 19431
rect 30472 19388 30524 19397
rect 31300 19388 31352 19440
rect 28724 19329 28738 19363
rect 28738 19329 28772 19363
rect 28772 19329 28776 19363
rect 28724 19320 28776 19329
rect 29552 19363 29604 19372
rect 29552 19329 29562 19363
rect 29562 19329 29596 19363
rect 29596 19329 29604 19363
rect 29552 19320 29604 19329
rect 29184 19252 29236 19304
rect 29920 19363 29972 19372
rect 29920 19329 29934 19363
rect 29934 19329 29968 19363
rect 29968 19329 29972 19363
rect 29920 19320 29972 19329
rect 30196 19363 30248 19372
rect 30196 19329 30205 19363
rect 30205 19329 30239 19363
rect 30239 19329 30248 19363
rect 30196 19320 30248 19329
rect 30288 19363 30340 19372
rect 30288 19329 30298 19363
rect 30298 19329 30332 19363
rect 30332 19329 30340 19363
rect 30288 19320 30340 19329
rect 32496 19184 32548 19236
rect 33048 19184 33100 19236
rect 18328 19116 18380 19168
rect 20076 19116 20128 19168
rect 22100 19116 22152 19168
rect 24400 19116 24452 19168
rect 26056 19116 26108 19168
rect 26148 19159 26200 19168
rect 26148 19125 26157 19159
rect 26157 19125 26191 19159
rect 26191 19125 26200 19159
rect 26148 19116 26200 19125
rect 26424 19159 26476 19168
rect 26424 19125 26433 19159
rect 26433 19125 26467 19159
rect 26467 19125 26476 19159
rect 26424 19116 26476 19125
rect 27160 19116 27212 19168
rect 27528 19159 27580 19168
rect 27528 19125 27537 19159
rect 27537 19125 27571 19159
rect 27571 19125 27580 19159
rect 27528 19116 27580 19125
rect 27620 19116 27672 19168
rect 34520 19116 34572 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4068 18912 4120 18964
rect 5172 18912 5224 18964
rect 5540 18912 5592 18964
rect 6920 18912 6972 18964
rect 7840 18912 7892 18964
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 8576 18955 8628 18964
rect 8576 18921 8585 18955
rect 8585 18921 8619 18955
rect 8619 18921 8628 18955
rect 8576 18912 8628 18921
rect 8760 18912 8812 18964
rect 12072 18912 12124 18964
rect 16488 18912 16540 18964
rect 18328 18912 18380 18964
rect 1400 18776 1452 18828
rect 2688 18776 2740 18828
rect 4436 18776 4488 18828
rect 7288 18819 7340 18828
rect 7288 18785 7297 18819
rect 7297 18785 7331 18819
rect 7331 18785 7340 18819
rect 7288 18776 7340 18785
rect 7564 18776 7616 18828
rect 10416 18844 10468 18896
rect 16856 18844 16908 18896
rect 17224 18844 17276 18896
rect 17316 18844 17368 18896
rect 8392 18776 8444 18828
rect 4712 18708 4764 18760
rect 3424 18640 3476 18692
rect 3516 18640 3568 18692
rect 2780 18572 2832 18624
rect 3700 18572 3752 18624
rect 4620 18640 4672 18692
rect 4528 18572 4580 18624
rect 5356 18572 5408 18624
rect 7104 18708 7156 18760
rect 8116 18708 8168 18760
rect 8760 18708 8812 18760
rect 9404 18819 9456 18828
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 11060 18776 11112 18828
rect 11520 18776 11572 18828
rect 12256 18776 12308 18828
rect 12624 18819 12676 18828
rect 12624 18785 12633 18819
rect 12633 18785 12667 18819
rect 12667 18785 12676 18819
rect 12624 18776 12676 18785
rect 17132 18776 17184 18828
rect 18972 18776 19024 18828
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 19616 18912 19668 18964
rect 20812 18844 20864 18896
rect 21364 18844 21416 18896
rect 10048 18708 10100 18760
rect 10416 18708 10468 18760
rect 11244 18708 11296 18760
rect 12072 18708 12124 18760
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 7104 18615 7156 18624
rect 7104 18581 7113 18615
rect 7113 18581 7147 18615
rect 7147 18581 7156 18615
rect 9772 18640 9824 18692
rect 9956 18683 10008 18692
rect 9956 18649 9965 18683
rect 9965 18649 9999 18683
rect 9999 18649 10008 18683
rect 9956 18640 10008 18649
rect 11704 18640 11756 18692
rect 14372 18683 14424 18692
rect 14372 18649 14381 18683
rect 14381 18649 14415 18683
rect 14415 18649 14424 18683
rect 14372 18640 14424 18649
rect 15384 18640 15436 18692
rect 17224 18708 17276 18760
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 17776 18708 17828 18760
rect 19248 18708 19300 18760
rect 7104 18572 7156 18581
rect 8668 18572 8720 18624
rect 10232 18572 10284 18624
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 10876 18572 10928 18624
rect 11796 18572 11848 18624
rect 12348 18615 12400 18624
rect 12348 18581 12357 18615
rect 12357 18581 12391 18615
rect 12391 18581 12400 18615
rect 12348 18572 12400 18581
rect 14096 18572 14148 18624
rect 15016 18572 15068 18624
rect 15936 18615 15988 18624
rect 15936 18581 15945 18615
rect 15945 18581 15979 18615
rect 15979 18581 15988 18615
rect 15936 18572 15988 18581
rect 16028 18572 16080 18624
rect 18972 18640 19024 18692
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 19708 18776 19760 18828
rect 20352 18776 20404 18828
rect 20628 18776 20680 18828
rect 22192 18912 22244 18964
rect 25044 18955 25096 18964
rect 25044 18921 25053 18955
rect 25053 18921 25087 18955
rect 25087 18921 25096 18955
rect 25044 18912 25096 18921
rect 21732 18844 21784 18896
rect 19708 18683 19760 18692
rect 19708 18649 19717 18683
rect 19717 18649 19751 18683
rect 19751 18649 19760 18683
rect 19708 18640 19760 18649
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 22192 18776 22244 18828
rect 24952 18776 25004 18828
rect 25412 18912 25464 18964
rect 27620 18912 27672 18964
rect 31208 18912 31260 18964
rect 32864 18955 32916 18964
rect 32864 18921 32873 18955
rect 32873 18921 32907 18955
rect 32907 18921 32916 18955
rect 32864 18912 32916 18921
rect 32956 18912 33008 18964
rect 34704 18912 34756 18964
rect 28724 18844 28776 18896
rect 29368 18844 29420 18896
rect 31576 18844 31628 18896
rect 25872 18776 25924 18828
rect 32404 18776 32456 18828
rect 33508 18819 33560 18828
rect 33508 18785 33517 18819
rect 33517 18785 33551 18819
rect 33551 18785 33560 18819
rect 33508 18776 33560 18785
rect 34152 18776 34204 18828
rect 34428 18776 34480 18828
rect 21088 18751 21140 18760
rect 21088 18717 21097 18751
rect 21097 18717 21131 18751
rect 21131 18717 21140 18751
rect 21088 18708 21140 18717
rect 20720 18640 20772 18692
rect 19432 18572 19484 18624
rect 19524 18572 19576 18624
rect 20444 18572 20496 18624
rect 20904 18572 20956 18624
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 21732 18708 21784 18760
rect 22100 18708 22152 18760
rect 24400 18708 24452 18760
rect 24676 18708 24728 18760
rect 21548 18683 21600 18692
rect 21548 18649 21557 18683
rect 21557 18649 21591 18683
rect 21591 18649 21600 18683
rect 21548 18640 21600 18649
rect 22468 18683 22520 18692
rect 22468 18649 22477 18683
rect 22477 18649 22511 18683
rect 22511 18649 22520 18683
rect 22468 18640 22520 18649
rect 22652 18640 22704 18692
rect 22928 18640 22980 18692
rect 25228 18683 25280 18692
rect 25228 18649 25255 18683
rect 25255 18649 25280 18683
rect 25228 18640 25280 18649
rect 26240 18708 26292 18760
rect 26332 18751 26384 18760
rect 26332 18717 26341 18751
rect 26341 18717 26375 18751
rect 26375 18717 26384 18751
rect 26332 18708 26384 18717
rect 25688 18640 25740 18692
rect 23756 18572 23808 18624
rect 24492 18572 24544 18624
rect 25504 18572 25556 18624
rect 26424 18640 26476 18692
rect 26332 18572 26384 18624
rect 26976 18708 27028 18760
rect 29184 18708 29236 18760
rect 32220 18751 32272 18760
rect 32220 18717 32229 18751
rect 32229 18717 32263 18751
rect 32263 18717 32272 18751
rect 32220 18708 32272 18717
rect 32496 18751 32548 18760
rect 32496 18717 32505 18751
rect 32505 18717 32539 18751
rect 32539 18717 32548 18751
rect 32496 18708 32548 18717
rect 32680 18708 32732 18760
rect 34704 18708 34756 18760
rect 27252 18640 27304 18692
rect 29552 18640 29604 18692
rect 31024 18640 31076 18692
rect 31208 18640 31260 18692
rect 34888 18751 34940 18760
rect 34888 18717 34898 18751
rect 34898 18717 34932 18751
rect 34932 18717 34940 18751
rect 34888 18708 34940 18717
rect 30104 18572 30156 18624
rect 35072 18683 35124 18692
rect 35072 18649 35081 18683
rect 35081 18649 35115 18683
rect 35115 18649 35124 18683
rect 35072 18640 35124 18649
rect 33968 18572 34020 18624
rect 34520 18572 34572 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 3332 18368 3384 18420
rect 3424 18368 3476 18420
rect 3700 18343 3752 18352
rect 3700 18309 3709 18343
rect 3709 18309 3743 18343
rect 3743 18309 3752 18343
rect 3700 18300 3752 18309
rect 5264 18368 5316 18420
rect 7104 18368 7156 18420
rect 8208 18368 8260 18420
rect 10324 18368 10376 18420
rect 10876 18411 10928 18420
rect 10876 18377 10885 18411
rect 10885 18377 10919 18411
rect 10919 18377 10928 18411
rect 10876 18368 10928 18377
rect 10968 18411 11020 18420
rect 10968 18377 10977 18411
rect 10977 18377 11011 18411
rect 11011 18377 11020 18411
rect 10968 18368 11020 18377
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 12348 18368 12400 18420
rect 14372 18368 14424 18420
rect 15936 18368 15988 18420
rect 16580 18368 16632 18420
rect 17500 18368 17552 18420
rect 18880 18411 18932 18420
rect 18880 18377 18889 18411
rect 18889 18377 18923 18411
rect 18923 18377 18932 18411
rect 18880 18368 18932 18377
rect 19984 18368 20036 18420
rect 21456 18368 21508 18420
rect 21732 18368 21784 18420
rect 22008 18368 22060 18420
rect 5356 18300 5408 18352
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 6644 18232 6696 18284
rect 7012 18275 7064 18284
rect 7012 18241 7021 18275
rect 7021 18241 7055 18275
rect 7055 18241 7064 18275
rect 7012 18232 7064 18241
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 2688 18164 2740 18216
rect 4068 18164 4120 18216
rect 4436 18164 4488 18216
rect 6828 18164 6880 18216
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 7380 18164 7432 18216
rect 9036 18300 9088 18352
rect 9496 18300 9548 18352
rect 10232 18300 10284 18352
rect 10416 18232 10468 18284
rect 11428 18232 11480 18284
rect 11704 18343 11756 18352
rect 11704 18309 11713 18343
rect 11713 18309 11747 18343
rect 11747 18309 11756 18343
rect 11704 18300 11756 18309
rect 13820 18300 13872 18352
rect 15016 18300 15068 18352
rect 18144 18300 18196 18352
rect 9956 18207 10008 18216
rect 9956 18173 9965 18207
rect 9965 18173 9999 18207
rect 9999 18173 10008 18207
rect 9956 18164 10008 18173
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 12992 18207 13044 18216
rect 10048 18096 10100 18148
rect 11612 18096 11664 18148
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 13176 18164 13228 18216
rect 17960 18232 18012 18284
rect 18420 18275 18472 18284
rect 18420 18241 18427 18275
rect 18427 18241 18472 18275
rect 18420 18232 18472 18241
rect 14832 18164 14884 18216
rect 15660 18164 15712 18216
rect 12624 18096 12676 18148
rect 14280 18096 14332 18148
rect 18236 18096 18288 18148
rect 18512 18096 18564 18148
rect 18788 18232 18840 18284
rect 19156 18300 19208 18352
rect 19524 18300 19576 18352
rect 20168 18300 20220 18352
rect 22836 18368 22888 18420
rect 22928 18368 22980 18420
rect 23756 18368 23808 18420
rect 24492 18368 24544 18420
rect 19708 18232 19760 18284
rect 20444 18275 20496 18284
rect 20444 18241 20453 18275
rect 20453 18241 20487 18275
rect 20487 18241 20496 18275
rect 20444 18232 20496 18241
rect 22468 18300 22520 18352
rect 22744 18300 22796 18352
rect 21364 18232 21416 18284
rect 21456 18275 21508 18284
rect 21456 18241 21465 18275
rect 21465 18241 21499 18275
rect 21499 18241 21508 18275
rect 21456 18232 21508 18241
rect 18788 18096 18840 18148
rect 19156 18096 19208 18148
rect 5816 18028 5868 18080
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 10140 18028 10192 18080
rect 17592 18028 17644 18080
rect 21180 18164 21232 18216
rect 19432 18096 19484 18148
rect 22284 18232 22336 18284
rect 22560 18232 22612 18284
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 22928 18164 22980 18216
rect 23756 18232 23808 18284
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 23296 18164 23348 18216
rect 23848 18164 23900 18216
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 25136 18275 25188 18284
rect 25136 18241 25145 18275
rect 25145 18241 25179 18275
rect 25179 18241 25188 18275
rect 25136 18232 25188 18241
rect 24768 18164 24820 18216
rect 21824 18096 21876 18148
rect 25320 18343 25372 18352
rect 25320 18309 25329 18343
rect 25329 18309 25363 18343
rect 25363 18309 25372 18343
rect 25320 18300 25372 18309
rect 25688 18300 25740 18352
rect 26240 18411 26292 18420
rect 26240 18377 26249 18411
rect 26249 18377 26283 18411
rect 26283 18377 26292 18411
rect 26240 18368 26292 18377
rect 26424 18368 26476 18420
rect 26056 18232 26108 18284
rect 27804 18232 27856 18284
rect 27988 18232 28040 18284
rect 28264 18343 28316 18352
rect 28264 18309 28273 18343
rect 28273 18309 28307 18343
rect 28307 18309 28316 18343
rect 28264 18300 28316 18309
rect 29368 18368 29420 18420
rect 29920 18368 29972 18420
rect 31208 18411 31260 18420
rect 31208 18377 31217 18411
rect 31217 18377 31251 18411
rect 31251 18377 31260 18411
rect 31208 18368 31260 18377
rect 30748 18343 30800 18352
rect 30748 18309 30757 18343
rect 30757 18309 30791 18343
rect 30791 18309 30800 18343
rect 30748 18300 30800 18309
rect 30012 18232 30064 18284
rect 30288 18232 30340 18284
rect 25320 18096 25372 18148
rect 27804 18096 27856 18148
rect 29184 18164 29236 18216
rect 30840 18207 30892 18216
rect 30840 18173 30849 18207
rect 30849 18173 30883 18207
rect 30883 18173 30892 18207
rect 30840 18164 30892 18173
rect 29460 18096 29512 18148
rect 19524 18028 19576 18080
rect 20076 18028 20128 18080
rect 21640 18028 21692 18080
rect 22652 18028 22704 18080
rect 23204 18028 23256 18080
rect 23756 18071 23808 18080
rect 23756 18037 23765 18071
rect 23765 18037 23799 18071
rect 23799 18037 23808 18071
rect 23756 18028 23808 18037
rect 24216 18028 24268 18080
rect 25228 18028 25280 18080
rect 25688 18071 25740 18080
rect 25688 18037 25697 18071
rect 25697 18037 25731 18071
rect 25731 18037 25740 18071
rect 25688 18028 25740 18037
rect 26148 18028 26200 18080
rect 28264 18028 28316 18080
rect 30472 18028 30524 18080
rect 30932 18028 30984 18080
rect 34244 18028 34296 18080
rect 35072 18028 35124 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1676 17824 1728 17876
rect 4620 17824 4672 17876
rect 7104 17824 7156 17876
rect 7288 17824 7340 17876
rect 2320 17688 2372 17740
rect 2504 17688 2556 17740
rect 2964 17756 3016 17808
rect 6828 17756 6880 17808
rect 12900 17824 12952 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15936 17867 15988 17876
rect 15936 17833 15945 17867
rect 15945 17833 15979 17867
rect 15979 17833 15988 17867
rect 15936 17824 15988 17833
rect 3332 17688 3384 17740
rect 4712 17688 4764 17740
rect 5816 17731 5868 17740
rect 5816 17697 5825 17731
rect 5825 17697 5859 17731
rect 5859 17697 5868 17731
rect 5816 17688 5868 17697
rect 7288 17731 7340 17740
rect 7288 17697 7297 17731
rect 7297 17697 7331 17731
rect 7331 17697 7340 17731
rect 7288 17688 7340 17697
rect 8116 17688 8168 17740
rect 13728 17756 13780 17808
rect 14924 17756 14976 17808
rect 16672 17756 16724 17808
rect 8760 17688 8812 17740
rect 5448 17620 5500 17672
rect 12348 17688 12400 17740
rect 2688 17484 2740 17536
rect 4712 17552 4764 17604
rect 7196 17552 7248 17604
rect 7380 17552 7432 17604
rect 3240 17484 3292 17536
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 11152 17663 11204 17672
rect 11152 17629 11161 17663
rect 11161 17629 11195 17663
rect 11195 17629 11204 17663
rect 11152 17620 11204 17629
rect 12164 17620 12216 17672
rect 12624 17620 12676 17672
rect 13544 17688 13596 17740
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 13820 17688 13872 17740
rect 13912 17620 13964 17672
rect 16396 17688 16448 17740
rect 16488 17688 16540 17740
rect 14924 17620 14976 17672
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 15200 17663 15252 17672
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 14648 17595 14700 17604
rect 14648 17561 14657 17595
rect 14657 17561 14691 17595
rect 14691 17561 14700 17595
rect 14648 17552 14700 17561
rect 16212 17620 16264 17672
rect 21088 17824 21140 17876
rect 22376 17867 22428 17876
rect 22376 17833 22385 17867
rect 22385 17833 22419 17867
rect 22419 17833 22428 17867
rect 22376 17824 22428 17833
rect 22468 17824 22520 17876
rect 18236 17756 18288 17808
rect 18144 17688 18196 17740
rect 18512 17756 18564 17808
rect 20720 17756 20772 17808
rect 21456 17756 21508 17808
rect 22284 17756 22336 17808
rect 23664 17799 23716 17808
rect 23664 17765 23673 17799
rect 23673 17765 23707 17799
rect 23707 17765 23716 17799
rect 23664 17756 23716 17765
rect 24032 17824 24084 17876
rect 25228 17867 25280 17876
rect 25228 17833 25237 17867
rect 25237 17833 25271 17867
rect 25271 17833 25280 17867
rect 25228 17824 25280 17833
rect 17868 17620 17920 17672
rect 17960 17620 18012 17672
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 18880 17663 18932 17672
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 20260 17688 20312 17740
rect 20628 17620 20680 17672
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 16120 17595 16172 17604
rect 8668 17484 8720 17536
rect 9588 17484 9640 17536
rect 11060 17527 11112 17536
rect 11060 17493 11069 17527
rect 11069 17493 11103 17527
rect 11103 17493 11112 17527
rect 11060 17484 11112 17493
rect 12532 17484 12584 17536
rect 12808 17527 12860 17536
rect 12808 17493 12817 17527
rect 12817 17493 12851 17527
rect 12851 17493 12860 17527
rect 12808 17484 12860 17493
rect 13268 17484 13320 17536
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 14924 17527 14976 17536
rect 14924 17493 14933 17527
rect 14933 17493 14967 17527
rect 14967 17493 14976 17527
rect 14924 17484 14976 17493
rect 15016 17484 15068 17536
rect 16120 17561 16129 17595
rect 16129 17561 16163 17595
rect 16163 17561 16172 17595
rect 16120 17552 16172 17561
rect 17132 17552 17184 17604
rect 15568 17484 15620 17536
rect 17040 17527 17092 17536
rect 17040 17493 17049 17527
rect 17049 17493 17083 17527
rect 17083 17493 17092 17527
rect 17040 17484 17092 17493
rect 17500 17552 17552 17604
rect 18144 17552 18196 17604
rect 19340 17552 19392 17604
rect 20536 17552 20588 17604
rect 21180 17552 21232 17604
rect 22652 17620 22704 17672
rect 23572 17620 23624 17672
rect 21640 17552 21692 17604
rect 21732 17595 21784 17604
rect 21732 17561 21741 17595
rect 21741 17561 21775 17595
rect 21775 17561 21784 17595
rect 21732 17552 21784 17561
rect 22744 17595 22796 17604
rect 22744 17561 22753 17595
rect 22753 17561 22787 17595
rect 22787 17561 22796 17595
rect 22744 17552 22796 17561
rect 23296 17552 23348 17604
rect 17592 17484 17644 17536
rect 18420 17484 18472 17536
rect 18512 17527 18564 17536
rect 18512 17493 18521 17527
rect 18521 17493 18555 17527
rect 18555 17493 18564 17527
rect 18512 17484 18564 17493
rect 19800 17527 19852 17536
rect 19800 17493 19809 17527
rect 19809 17493 19843 17527
rect 19843 17493 19852 17527
rect 19800 17484 19852 17493
rect 20720 17484 20772 17536
rect 22284 17484 22336 17536
rect 22560 17527 22612 17536
rect 22560 17493 22587 17527
rect 22587 17493 22612 17527
rect 22560 17484 22612 17493
rect 26240 17731 26292 17740
rect 26240 17697 26249 17731
rect 26249 17697 26283 17731
rect 26283 17697 26292 17731
rect 26240 17688 26292 17697
rect 24216 17620 24268 17672
rect 24952 17620 25004 17672
rect 25044 17595 25096 17604
rect 25044 17561 25053 17595
rect 25053 17561 25087 17595
rect 25087 17561 25096 17595
rect 25044 17552 25096 17561
rect 25688 17663 25740 17672
rect 25688 17629 25697 17663
rect 25697 17629 25731 17663
rect 25731 17629 25740 17663
rect 25688 17620 25740 17629
rect 25872 17620 25924 17672
rect 27068 17688 27120 17740
rect 29644 17552 29696 17604
rect 31024 17552 31076 17604
rect 32312 17552 32364 17604
rect 33416 17552 33468 17604
rect 29184 17484 29236 17536
rect 34060 17484 34112 17536
rect 36452 17484 36504 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 6644 17323 6696 17332
rect 6644 17289 6653 17323
rect 6653 17289 6687 17323
rect 6687 17289 6696 17323
rect 6644 17280 6696 17289
rect 8852 17280 8904 17332
rect 8944 17280 8996 17332
rect 2596 17212 2648 17264
rect 2964 17212 3016 17264
rect 3976 17212 4028 17264
rect 5356 17212 5408 17264
rect 3608 17119 3660 17128
rect 3608 17085 3617 17119
rect 3617 17085 3651 17119
rect 3651 17085 3660 17119
rect 3608 17076 3660 17085
rect 4620 17076 4672 17128
rect 6184 17144 6236 17196
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 1676 16940 1728 16992
rect 2504 16940 2556 16992
rect 8668 17008 8720 17060
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 9956 17144 10008 17196
rect 10968 17280 11020 17332
rect 10232 17212 10284 17264
rect 10876 17255 10928 17264
rect 10876 17221 10885 17255
rect 10885 17221 10919 17255
rect 10919 17221 10928 17255
rect 10876 17212 10928 17221
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 12900 17280 12952 17332
rect 13636 17280 13688 17332
rect 12348 17212 12400 17264
rect 12624 17212 12676 17264
rect 14188 17280 14240 17332
rect 14464 17280 14516 17332
rect 15936 17280 15988 17332
rect 21180 17280 21232 17332
rect 21364 17280 21416 17332
rect 22560 17323 22612 17332
rect 22560 17289 22569 17323
rect 22569 17289 22603 17323
rect 22603 17289 22612 17323
rect 22560 17280 22612 17289
rect 22744 17323 22796 17332
rect 22744 17289 22753 17323
rect 22753 17289 22787 17323
rect 22787 17289 22796 17323
rect 22744 17280 22796 17289
rect 23296 17323 23348 17332
rect 23296 17289 23305 17323
rect 23305 17289 23339 17323
rect 23339 17289 23348 17323
rect 23296 17280 23348 17289
rect 23572 17280 23624 17332
rect 24768 17280 24820 17332
rect 25228 17280 25280 17332
rect 25872 17323 25924 17332
rect 25872 17289 25881 17323
rect 25881 17289 25915 17323
rect 25915 17289 25924 17323
rect 25872 17280 25924 17289
rect 27068 17323 27120 17332
rect 27068 17289 27077 17323
rect 27077 17289 27111 17323
rect 27111 17289 27120 17323
rect 27068 17280 27120 17289
rect 29368 17280 29420 17332
rect 10784 17144 10836 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 11152 17076 11204 17128
rect 12440 17008 12492 17060
rect 12716 17076 12768 17128
rect 16120 17212 16172 17264
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 14740 17144 14792 17196
rect 15108 17144 15160 17196
rect 15384 17144 15436 17196
rect 12992 17008 13044 17060
rect 15660 17144 15712 17196
rect 16672 17144 16724 17196
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 17316 17144 17368 17196
rect 18236 17144 18288 17196
rect 15844 17076 15896 17128
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 16396 17076 16448 17128
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 8576 16940 8628 16992
rect 9036 16940 9088 16992
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 13176 16983 13228 16992
rect 13176 16949 13185 16983
rect 13185 16949 13219 16983
rect 13219 16949 13228 16983
rect 13176 16940 13228 16949
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 14924 17008 14976 17060
rect 15108 17008 15160 17060
rect 15384 17051 15436 17060
rect 15384 17017 15393 17051
rect 15393 17017 15427 17051
rect 15427 17017 15436 17051
rect 15384 17008 15436 17017
rect 15476 17008 15528 17060
rect 17868 17076 17920 17128
rect 17040 17008 17092 17060
rect 14740 16983 14792 16992
rect 14740 16949 14749 16983
rect 14749 16949 14783 16983
rect 14783 16949 14792 16983
rect 14740 16940 14792 16949
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 17316 16940 17368 16992
rect 17960 17051 18012 17060
rect 17960 17017 17969 17051
rect 17969 17017 18003 17051
rect 18003 17017 18012 17051
rect 17960 17008 18012 17017
rect 20720 17212 20772 17264
rect 19340 17144 19392 17196
rect 19616 17144 19668 17196
rect 19800 17144 19852 17196
rect 19156 17076 19208 17128
rect 20076 17076 20128 17128
rect 20168 17119 20220 17128
rect 20168 17085 20177 17119
rect 20177 17085 20211 17119
rect 20211 17085 20220 17119
rect 20168 17076 20220 17085
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 21088 17187 21140 17196
rect 21088 17153 21095 17187
rect 21095 17153 21140 17187
rect 21088 17144 21140 17153
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 21272 17187 21324 17196
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 21548 17144 21600 17196
rect 22284 17187 22336 17196
rect 22284 17153 22293 17187
rect 22293 17153 22327 17187
rect 22327 17153 22336 17187
rect 22284 17144 22336 17153
rect 21732 17076 21784 17128
rect 19708 17008 19760 17060
rect 20444 17008 20496 17060
rect 21088 17008 21140 17060
rect 22192 17008 22244 17060
rect 22744 17144 22796 17196
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 23664 17187 23716 17196
rect 23664 17153 23673 17187
rect 23673 17153 23707 17187
rect 23707 17153 23716 17187
rect 23664 17144 23716 17153
rect 24400 17187 24452 17196
rect 24400 17153 24409 17187
rect 24409 17153 24443 17187
rect 24443 17153 24452 17187
rect 24400 17144 24452 17153
rect 25320 17212 25372 17264
rect 27712 17212 27764 17264
rect 25688 17144 25740 17196
rect 26148 17144 26200 17196
rect 26976 17187 27028 17196
rect 26976 17153 26985 17187
rect 26985 17153 27019 17187
rect 27019 17153 27028 17187
rect 26976 17144 27028 17153
rect 27528 17144 27580 17196
rect 30288 17280 30340 17332
rect 31208 17144 31260 17196
rect 32036 17144 32088 17196
rect 32312 17144 32364 17196
rect 33232 17280 33284 17332
rect 33508 17280 33560 17332
rect 34060 17212 34112 17264
rect 34796 17212 34848 17264
rect 26792 17076 26844 17128
rect 29276 17076 29328 17128
rect 29368 17076 29420 17128
rect 23296 17008 23348 17060
rect 19156 16983 19208 16992
rect 19156 16949 19165 16983
rect 19165 16949 19199 16983
rect 19199 16949 19208 16983
rect 19156 16940 19208 16949
rect 19340 16940 19392 16992
rect 20352 16940 20404 16992
rect 22652 16940 22704 16992
rect 23480 16940 23532 16992
rect 24032 17051 24084 17060
rect 24032 17017 24041 17051
rect 24041 17017 24075 17051
rect 24075 17017 24084 17051
rect 24032 17008 24084 17017
rect 24124 17051 24176 17060
rect 24124 17017 24133 17051
rect 24133 17017 24167 17051
rect 24167 17017 24176 17051
rect 24124 17008 24176 17017
rect 24676 17008 24728 17060
rect 25596 17008 25648 17060
rect 32036 17008 32088 17060
rect 34152 17187 34204 17196
rect 34152 17153 34161 17187
rect 34161 17153 34195 17187
rect 34195 17153 34204 17187
rect 34152 17144 34204 17153
rect 36452 17144 36504 17196
rect 33416 17076 33468 17128
rect 25044 16940 25096 16992
rect 27712 16940 27764 16992
rect 29000 16940 29052 16992
rect 29184 16940 29236 16992
rect 32588 16983 32640 16992
rect 32588 16949 32597 16983
rect 32597 16949 32631 16983
rect 32631 16949 32640 16983
rect 32588 16940 32640 16949
rect 32680 16983 32732 16992
rect 32680 16949 32689 16983
rect 32689 16949 32723 16983
rect 32723 16949 32732 16983
rect 32680 16940 32732 16949
rect 32772 16940 32824 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2688 16736 2740 16788
rect 4620 16736 4672 16788
rect 7104 16736 7156 16788
rect 9404 16736 9456 16788
rect 9680 16736 9732 16788
rect 10508 16736 10560 16788
rect 4068 16668 4120 16720
rect 2596 16600 2648 16652
rect 2688 16600 2740 16652
rect 3424 16600 3476 16652
rect 8024 16668 8076 16720
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 6276 16600 6328 16652
rect 5448 16532 5500 16584
rect 3056 16396 3108 16448
rect 5356 16464 5408 16516
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 8944 16532 8996 16541
rect 10048 16668 10100 16720
rect 10600 16668 10652 16720
rect 14004 16736 14056 16788
rect 14188 16736 14240 16788
rect 15200 16736 15252 16788
rect 15476 16736 15528 16788
rect 16212 16736 16264 16788
rect 17132 16779 17184 16788
rect 17132 16745 17141 16779
rect 17141 16745 17175 16779
rect 17175 16745 17184 16779
rect 17132 16736 17184 16745
rect 17316 16736 17368 16788
rect 19248 16779 19300 16788
rect 19248 16745 19257 16779
rect 19257 16745 19291 16779
rect 19291 16745 19300 16779
rect 19248 16736 19300 16745
rect 19984 16736 20036 16788
rect 9956 16600 10008 16652
rect 9404 16575 9456 16584
rect 9404 16541 9413 16575
rect 9413 16541 9447 16575
rect 9447 16541 9456 16575
rect 9404 16532 9456 16541
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 9772 16532 9824 16584
rect 10508 16600 10560 16652
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 13912 16668 13964 16720
rect 14648 16668 14700 16720
rect 12164 16600 12216 16652
rect 4712 16396 4764 16448
rect 4896 16396 4948 16448
rect 7472 16396 7524 16448
rect 7748 16439 7800 16448
rect 7748 16405 7757 16439
rect 7757 16405 7791 16439
rect 7791 16405 7800 16439
rect 7748 16396 7800 16405
rect 8024 16396 8076 16448
rect 9588 16464 9640 16516
rect 10784 16575 10836 16584
rect 10784 16541 10793 16575
rect 10793 16541 10827 16575
rect 10827 16541 10836 16575
rect 10784 16532 10836 16541
rect 11060 16532 11112 16584
rect 11520 16532 11572 16584
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 12532 16532 12584 16584
rect 12900 16532 12952 16584
rect 13176 16532 13228 16584
rect 12716 16464 12768 16516
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 13820 16532 13872 16584
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 9128 16439 9180 16448
rect 9128 16405 9137 16439
rect 9137 16405 9171 16439
rect 9171 16405 9180 16439
rect 9128 16396 9180 16405
rect 9220 16439 9272 16448
rect 9220 16405 9229 16439
rect 9229 16405 9263 16439
rect 9263 16405 9272 16439
rect 9220 16396 9272 16405
rect 9956 16396 10008 16448
rect 10968 16396 11020 16448
rect 11980 16396 12032 16448
rect 15200 16439 15252 16448
rect 15200 16405 15209 16439
rect 15209 16405 15243 16439
rect 15243 16405 15252 16439
rect 15200 16396 15252 16405
rect 15752 16668 15804 16720
rect 20352 16668 20404 16720
rect 21180 16736 21232 16788
rect 24032 16736 24084 16788
rect 21732 16668 21784 16720
rect 25964 16668 26016 16720
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 15936 16532 15988 16584
rect 17040 16575 17092 16584
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 17040 16532 17092 16541
rect 16120 16507 16172 16516
rect 16120 16473 16129 16507
rect 16129 16473 16163 16507
rect 16163 16473 16172 16507
rect 16120 16464 16172 16473
rect 16948 16464 17000 16516
rect 17316 16575 17368 16584
rect 17316 16541 17325 16575
rect 17325 16541 17359 16575
rect 17359 16541 17368 16575
rect 17316 16532 17368 16541
rect 17500 16532 17552 16584
rect 17868 16532 17920 16584
rect 18696 16532 18748 16584
rect 18972 16532 19024 16584
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 20260 16600 20312 16652
rect 19800 16575 19852 16584
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 16212 16396 16264 16448
rect 16856 16439 16908 16448
rect 16856 16405 16865 16439
rect 16865 16405 16899 16439
rect 16899 16405 16908 16439
rect 16856 16396 16908 16405
rect 17776 16464 17828 16516
rect 17960 16507 18012 16516
rect 17960 16473 17969 16507
rect 17969 16473 18003 16507
rect 18003 16473 18012 16507
rect 17960 16464 18012 16473
rect 17224 16396 17276 16448
rect 17684 16396 17736 16448
rect 18512 16464 18564 16516
rect 19156 16464 19208 16516
rect 19708 16464 19760 16516
rect 20076 16575 20128 16584
rect 20076 16541 20085 16575
rect 20085 16541 20119 16575
rect 20119 16541 20128 16575
rect 20076 16532 20128 16541
rect 20168 16575 20220 16584
rect 20168 16541 20177 16575
rect 20177 16541 20211 16575
rect 20211 16541 20220 16575
rect 20168 16532 20220 16541
rect 20628 16532 20680 16584
rect 23296 16575 23348 16584
rect 23296 16541 23305 16575
rect 23305 16541 23339 16575
rect 23339 16541 23348 16575
rect 23296 16532 23348 16541
rect 20536 16439 20588 16448
rect 20536 16405 20545 16439
rect 20545 16405 20579 16439
rect 20579 16405 20588 16439
rect 20536 16396 20588 16405
rect 20628 16396 20680 16448
rect 22744 16464 22796 16516
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 23572 16532 23624 16541
rect 23664 16575 23716 16584
rect 23664 16541 23673 16575
rect 23673 16541 23707 16575
rect 23707 16541 23716 16575
rect 23664 16532 23716 16541
rect 24860 16532 24912 16584
rect 21272 16396 21324 16448
rect 21456 16396 21508 16448
rect 21732 16396 21784 16448
rect 24032 16464 24084 16516
rect 24400 16507 24452 16516
rect 24400 16473 24409 16507
rect 24409 16473 24443 16507
rect 24443 16473 24452 16507
rect 24400 16464 24452 16473
rect 25412 16575 25464 16584
rect 25412 16541 25421 16575
rect 25421 16541 25455 16575
rect 25455 16541 25464 16575
rect 25412 16532 25464 16541
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 25964 16575 26016 16584
rect 25964 16541 25973 16575
rect 25973 16541 26007 16575
rect 26007 16541 26016 16575
rect 25964 16532 26016 16541
rect 32588 16736 32640 16788
rect 33416 16779 33468 16788
rect 33416 16745 33425 16779
rect 33425 16745 33459 16779
rect 33459 16745 33468 16779
rect 33416 16736 33468 16745
rect 28356 16600 28408 16652
rect 28908 16600 28960 16652
rect 27620 16575 27672 16584
rect 27620 16541 27629 16575
rect 27629 16541 27663 16575
rect 27663 16541 27672 16575
rect 27620 16532 27672 16541
rect 27804 16575 27856 16584
rect 27804 16541 27811 16575
rect 27811 16541 27856 16575
rect 27804 16532 27856 16541
rect 27896 16575 27948 16584
rect 27896 16541 27905 16575
rect 27905 16541 27939 16575
rect 27939 16541 27948 16575
rect 27896 16532 27948 16541
rect 28080 16532 28132 16584
rect 29368 16532 29420 16584
rect 29828 16643 29880 16652
rect 29828 16609 29837 16643
rect 29837 16609 29871 16643
rect 29871 16609 29880 16643
rect 29828 16600 29880 16609
rect 30104 16532 30156 16584
rect 27436 16464 27488 16516
rect 30288 16464 30340 16516
rect 31852 16464 31904 16516
rect 32404 16643 32456 16652
rect 32404 16609 32413 16643
rect 32413 16609 32447 16643
rect 32447 16609 32456 16643
rect 32404 16600 32456 16609
rect 32956 16532 33008 16584
rect 34336 16668 34388 16720
rect 25688 16396 25740 16448
rect 30656 16396 30708 16448
rect 32496 16396 32548 16448
rect 32956 16396 33008 16448
rect 34612 16532 34664 16584
rect 33232 16464 33284 16516
rect 34152 16464 34204 16516
rect 35164 16507 35216 16516
rect 35164 16473 35173 16507
rect 35173 16473 35207 16507
rect 35207 16473 35216 16507
rect 35164 16464 35216 16473
rect 35256 16507 35308 16516
rect 35256 16473 35265 16507
rect 35265 16473 35299 16507
rect 35299 16473 35308 16507
rect 35256 16464 35308 16473
rect 35348 16396 35400 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 2596 16192 2648 16244
rect 3608 16192 3660 16244
rect 1676 16167 1728 16176
rect 1676 16133 1685 16167
rect 1685 16133 1719 16167
rect 1719 16133 1728 16167
rect 1676 16124 1728 16133
rect 3056 16124 3108 16176
rect 4620 16124 4672 16176
rect 5356 16124 5408 16176
rect 6276 16192 6328 16244
rect 7472 16192 7524 16244
rect 7564 16192 7616 16244
rect 11980 16192 12032 16244
rect 12808 16192 12860 16244
rect 13820 16192 13872 16244
rect 14372 16192 14424 16244
rect 16120 16192 16172 16244
rect 17500 16192 17552 16244
rect 17684 16192 17736 16244
rect 3792 16099 3844 16108
rect 3792 16065 3801 16099
rect 3801 16065 3835 16099
rect 3835 16065 3844 16099
rect 3792 16056 3844 16065
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 3884 16056 3936 16065
rect 7012 16124 7064 16176
rect 7104 16056 7156 16108
rect 8024 16056 8076 16108
rect 8484 16056 8536 16108
rect 9588 16056 9640 16108
rect 4068 16031 4120 16040
rect 4068 15997 4077 16031
rect 4077 15997 4111 16031
rect 4111 15997 4120 16031
rect 4068 15988 4120 15997
rect 5908 16031 5960 16040
rect 5908 15997 5917 16031
rect 5917 15997 5951 16031
rect 5951 15997 5960 16031
rect 5908 15988 5960 15997
rect 6460 15988 6512 16040
rect 6920 16031 6972 16040
rect 6920 15997 6929 16031
rect 6929 15997 6963 16031
rect 6963 15997 6972 16031
rect 6920 15988 6972 15997
rect 3424 15963 3476 15972
rect 3424 15929 3433 15963
rect 3433 15929 3467 15963
rect 3467 15929 3476 15963
rect 3424 15920 3476 15929
rect 9680 15988 9732 16040
rect 10600 15988 10652 16040
rect 11060 16099 11112 16108
rect 11060 16065 11069 16099
rect 11069 16065 11103 16099
rect 11103 16065 11112 16099
rect 11060 16056 11112 16065
rect 11520 16056 11572 16108
rect 12440 16056 12492 16108
rect 13544 16124 13596 16176
rect 12716 16056 12768 16108
rect 13176 16056 13228 16108
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 14004 16124 14056 16176
rect 16764 16124 16816 16176
rect 16948 16124 17000 16176
rect 13912 16056 13964 16108
rect 13268 15988 13320 16040
rect 12348 15920 12400 15972
rect 12808 15920 12860 15972
rect 14832 15920 14884 15972
rect 15568 16056 15620 16108
rect 16212 16056 16264 16108
rect 16672 15988 16724 16040
rect 17408 16099 17460 16108
rect 17408 16065 17417 16099
rect 17417 16065 17451 16099
rect 17451 16065 17460 16099
rect 17408 16056 17460 16065
rect 17868 16124 17920 16176
rect 18696 16167 18748 16176
rect 18696 16133 18705 16167
rect 18705 16133 18739 16167
rect 18739 16133 18748 16167
rect 18696 16124 18748 16133
rect 19156 16235 19208 16244
rect 19156 16201 19165 16235
rect 19165 16201 19199 16235
rect 19199 16201 19208 16235
rect 19156 16192 19208 16201
rect 19248 16192 19300 16244
rect 20536 16192 20588 16244
rect 23388 16192 23440 16244
rect 24768 16192 24820 16244
rect 25136 16192 25188 16244
rect 17960 16056 18012 16108
rect 18512 16056 18564 16108
rect 18972 16099 19024 16108
rect 18972 16065 18981 16099
rect 18981 16065 19015 16099
rect 19015 16065 19024 16099
rect 18972 16056 19024 16065
rect 19432 16099 19484 16108
rect 19432 16065 19439 16099
rect 19439 16065 19484 16099
rect 18788 16031 18840 16040
rect 18788 15997 18797 16031
rect 18797 15997 18831 16031
rect 18831 15997 18840 16031
rect 18788 15988 18840 15997
rect 19156 15988 19208 16040
rect 19432 16056 19484 16065
rect 20076 16124 20128 16176
rect 19708 16099 19760 16108
rect 19708 16065 19722 16099
rect 19722 16065 19756 16099
rect 19756 16065 19760 16099
rect 22836 16124 22888 16176
rect 25044 16167 25096 16176
rect 25044 16133 25071 16167
rect 25071 16133 25096 16167
rect 25044 16124 25096 16133
rect 25780 16235 25832 16244
rect 25780 16201 25789 16235
rect 25789 16201 25823 16235
rect 25823 16201 25832 16235
rect 25780 16192 25832 16201
rect 27620 16235 27672 16244
rect 27620 16201 27629 16235
rect 27629 16201 27663 16235
rect 27663 16201 27672 16235
rect 27620 16192 27672 16201
rect 19708 16056 19760 16065
rect 20996 16056 21048 16108
rect 6460 15852 6512 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 10692 15852 10744 15904
rect 12992 15852 13044 15904
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 19800 15920 19852 15972
rect 19892 15963 19944 15972
rect 19892 15929 19901 15963
rect 19901 15929 19935 15963
rect 19935 15929 19944 15963
rect 19892 15920 19944 15929
rect 19340 15852 19392 15904
rect 19708 15852 19760 15904
rect 20168 15988 20220 16040
rect 21824 16031 21876 16040
rect 21824 15997 21833 16031
rect 21833 15997 21867 16031
rect 21867 15997 21876 16031
rect 21824 15988 21876 15997
rect 22284 16099 22336 16108
rect 22284 16065 22293 16099
rect 22293 16065 22327 16099
rect 22327 16065 22336 16099
rect 22284 16056 22336 16065
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 24124 16056 24176 16108
rect 23296 15988 23348 16040
rect 23480 15988 23532 16040
rect 22284 15920 22336 15972
rect 20076 15852 20128 15904
rect 24308 15920 24360 15972
rect 24492 16099 24544 16108
rect 24492 16065 24501 16099
rect 24501 16065 24535 16099
rect 24535 16065 24544 16099
rect 24492 16056 24544 16065
rect 24584 16099 24636 16108
rect 26332 16124 26384 16176
rect 24584 16065 24619 16099
rect 24619 16065 24636 16099
rect 24584 16056 24636 16065
rect 25688 16056 25740 16108
rect 25320 15852 25372 15904
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 26608 16056 26660 16108
rect 26700 16099 26752 16108
rect 26700 16065 26709 16099
rect 26709 16065 26743 16099
rect 26743 16065 26752 16099
rect 26700 16056 26752 16065
rect 26792 16099 26844 16108
rect 26792 16065 26801 16099
rect 26801 16065 26835 16099
rect 26835 16065 26844 16099
rect 26792 16056 26844 16065
rect 27620 15988 27672 16040
rect 27896 16192 27948 16244
rect 28080 16124 28132 16176
rect 29828 16192 29880 16244
rect 30564 16124 30616 16176
rect 30748 16124 30800 16176
rect 27896 16099 27948 16108
rect 27896 16065 27905 16099
rect 27905 16065 27939 16099
rect 27939 16065 27948 16099
rect 27896 16056 27948 16065
rect 28448 16056 28500 16108
rect 28632 16056 28684 16108
rect 29184 16099 29236 16108
rect 29184 16065 29193 16099
rect 29193 16065 29227 16099
rect 29227 16065 29236 16099
rect 29184 16056 29236 16065
rect 29368 16056 29420 16108
rect 30380 16056 30432 16108
rect 30932 16056 30984 16108
rect 29920 15988 29972 16040
rect 30196 15988 30248 16040
rect 30564 15988 30616 16040
rect 31208 16056 31260 16108
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 31576 16056 31628 16108
rect 25964 15920 26016 15972
rect 30104 15920 30156 15972
rect 31944 16192 31996 16244
rect 32772 16192 32824 16244
rect 34520 16192 34572 16244
rect 34704 16192 34756 16244
rect 33324 15988 33376 16040
rect 34428 15988 34480 16040
rect 35164 15920 35216 15972
rect 28356 15852 28408 15904
rect 30656 15895 30708 15904
rect 30656 15861 30665 15895
rect 30665 15861 30699 15895
rect 30699 15861 30708 15895
rect 30656 15852 30708 15861
rect 31576 15852 31628 15904
rect 31852 15852 31904 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3792 15691 3844 15700
rect 3792 15657 3801 15691
rect 3801 15657 3835 15691
rect 3835 15657 3844 15691
rect 3792 15648 3844 15657
rect 5908 15648 5960 15700
rect 4712 15512 4764 15564
rect 6920 15512 6972 15564
rect 8576 15648 8628 15700
rect 8208 15580 8260 15632
rect 8392 15580 8444 15632
rect 7748 15555 7800 15564
rect 7748 15521 7757 15555
rect 7757 15521 7791 15555
rect 7791 15521 7800 15555
rect 7748 15512 7800 15521
rect 8760 15512 8812 15564
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 8300 15444 8352 15496
rect 8852 15444 8904 15496
rect 8944 15444 8996 15496
rect 9404 15555 9456 15564
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 10140 15580 10192 15632
rect 12716 15648 12768 15700
rect 12900 15691 12952 15700
rect 12900 15657 12909 15691
rect 12909 15657 12943 15691
rect 12943 15657 12952 15691
rect 12900 15648 12952 15657
rect 14648 15648 14700 15700
rect 15016 15691 15068 15700
rect 15016 15657 15025 15691
rect 15025 15657 15059 15691
rect 15059 15657 15068 15691
rect 15016 15648 15068 15657
rect 15476 15691 15528 15700
rect 15476 15657 15485 15691
rect 15485 15657 15519 15691
rect 15519 15657 15528 15691
rect 15476 15648 15528 15657
rect 12624 15580 12676 15632
rect 13084 15580 13136 15632
rect 14740 15580 14792 15632
rect 16396 15648 16448 15700
rect 17132 15648 17184 15700
rect 18788 15648 18840 15700
rect 20904 15648 20956 15700
rect 21916 15648 21968 15700
rect 22376 15648 22428 15700
rect 23112 15648 23164 15700
rect 25412 15648 25464 15700
rect 26148 15648 26200 15700
rect 16488 15580 16540 15632
rect 17040 15580 17092 15632
rect 19524 15580 19576 15632
rect 19800 15580 19852 15632
rect 22284 15580 22336 15632
rect 27896 15648 27948 15700
rect 30104 15648 30156 15700
rect 31392 15648 31444 15700
rect 31484 15691 31536 15700
rect 31484 15657 31493 15691
rect 31493 15657 31527 15691
rect 31527 15657 31536 15691
rect 31484 15648 31536 15657
rect 33324 15648 33376 15700
rect 9956 15487 10008 15496
rect 9956 15453 9965 15487
rect 9965 15453 9999 15487
rect 9999 15453 10008 15487
rect 9956 15444 10008 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 10968 15512 11020 15564
rect 10416 15444 10468 15496
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 10692 15487 10744 15496
rect 10692 15453 10705 15487
rect 10705 15453 10744 15487
rect 10692 15444 10744 15453
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 12808 15512 12860 15564
rect 16672 15512 16724 15564
rect 18144 15512 18196 15564
rect 18512 15512 18564 15564
rect 19432 15512 19484 15564
rect 7656 15308 7708 15360
rect 8392 15308 8444 15360
rect 8484 15308 8536 15360
rect 9404 15308 9456 15360
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 15844 15444 15896 15496
rect 16212 15444 16264 15496
rect 17408 15444 17460 15496
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 13360 15376 13412 15428
rect 16304 15419 16356 15428
rect 16304 15385 16313 15419
rect 16313 15385 16347 15419
rect 16347 15385 16356 15419
rect 16304 15376 16356 15385
rect 17960 15376 18012 15428
rect 19432 15376 19484 15428
rect 20260 15444 20312 15496
rect 23848 15512 23900 15564
rect 25044 15512 25096 15564
rect 31668 15580 31720 15632
rect 36176 15580 36228 15632
rect 20812 15444 20864 15496
rect 21364 15444 21416 15496
rect 21824 15444 21876 15496
rect 22100 15487 22152 15496
rect 22100 15453 22109 15487
rect 22109 15453 22143 15487
rect 22143 15453 22152 15487
rect 22100 15444 22152 15453
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 22652 15444 22704 15496
rect 22836 15444 22888 15496
rect 24768 15444 24820 15496
rect 25688 15444 25740 15496
rect 26424 15487 26476 15496
rect 26424 15453 26433 15487
rect 26433 15453 26467 15487
rect 26467 15453 26476 15487
rect 26424 15444 26476 15453
rect 22744 15419 22796 15428
rect 22744 15385 22753 15419
rect 22753 15385 22787 15419
rect 22787 15385 22796 15419
rect 22744 15376 22796 15385
rect 24492 15376 24544 15428
rect 26792 15444 26844 15496
rect 14372 15308 14424 15360
rect 15476 15308 15528 15360
rect 15660 15351 15712 15360
rect 15660 15317 15669 15351
rect 15669 15317 15703 15351
rect 15703 15317 15712 15351
rect 15660 15308 15712 15317
rect 15752 15308 15804 15360
rect 16120 15308 16172 15360
rect 16212 15308 16264 15360
rect 19708 15308 19760 15360
rect 19800 15308 19852 15360
rect 22928 15308 22980 15360
rect 23296 15308 23348 15360
rect 25964 15308 26016 15360
rect 26148 15308 26200 15360
rect 26608 15308 26660 15360
rect 27160 15444 27212 15496
rect 27436 15444 27488 15496
rect 29000 15512 29052 15564
rect 29368 15512 29420 15564
rect 31024 15512 31076 15564
rect 28632 15487 28684 15496
rect 28632 15453 28641 15487
rect 28641 15453 28675 15487
rect 28675 15453 28684 15487
rect 28632 15444 28684 15453
rect 28816 15444 28868 15496
rect 29736 15444 29788 15496
rect 30748 15444 30800 15496
rect 31392 15444 31444 15496
rect 31484 15487 31536 15496
rect 31484 15453 31493 15487
rect 31493 15453 31527 15487
rect 31527 15453 31536 15487
rect 31484 15444 31536 15453
rect 31576 15487 31628 15496
rect 31576 15453 31585 15487
rect 31585 15453 31619 15487
rect 31619 15453 31628 15487
rect 31576 15444 31628 15453
rect 28724 15419 28776 15428
rect 28724 15385 28733 15419
rect 28733 15385 28767 15419
rect 28767 15385 28776 15419
rect 28724 15376 28776 15385
rect 33048 15444 33100 15496
rect 33232 15487 33284 15496
rect 33232 15453 33236 15487
rect 33236 15453 33270 15487
rect 33270 15453 33284 15487
rect 33232 15444 33284 15453
rect 33784 15512 33836 15564
rect 33692 15487 33744 15496
rect 33692 15453 33701 15487
rect 33701 15453 33735 15487
rect 33735 15453 33744 15487
rect 33692 15444 33744 15453
rect 32864 15376 32916 15428
rect 27160 15308 27212 15360
rect 27712 15308 27764 15360
rect 28264 15308 28316 15360
rect 28356 15351 28408 15360
rect 28356 15317 28365 15351
rect 28365 15317 28399 15351
rect 28399 15317 28408 15351
rect 28356 15308 28408 15317
rect 31300 15351 31352 15360
rect 31300 15317 31309 15351
rect 31309 15317 31343 15351
rect 31343 15317 31352 15351
rect 31300 15308 31352 15317
rect 33048 15351 33100 15360
rect 33048 15317 33057 15351
rect 33057 15317 33091 15351
rect 33091 15317 33100 15351
rect 33048 15308 33100 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 4620 15104 4672 15156
rect 5264 15104 5316 15156
rect 7196 15104 7248 15156
rect 7472 15104 7524 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 8392 15104 8444 15156
rect 8760 15104 8812 15156
rect 12532 15104 12584 15156
rect 12716 15104 12768 15156
rect 13912 15104 13964 15156
rect 15660 15104 15712 15156
rect 16212 15104 16264 15156
rect 16304 15104 16356 15156
rect 18236 15104 18288 15156
rect 18328 15104 18380 15156
rect 19064 15147 19116 15156
rect 19064 15113 19091 15147
rect 19091 15113 19116 15147
rect 2596 14968 2648 15020
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 3976 14900 4028 14952
rect 6736 14968 6788 15020
rect 5540 14900 5592 14952
rect 7196 14968 7248 15020
rect 9680 15036 9732 15088
rect 10324 15036 10376 15088
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 8024 14943 8076 14952
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 7932 14832 7984 14884
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 9496 14968 9548 15020
rect 11704 15036 11756 15088
rect 10416 15011 10468 15020
rect 10416 14977 10425 15011
rect 10425 14977 10459 15011
rect 10459 14977 10468 15011
rect 10416 14968 10468 14977
rect 10692 14968 10744 15020
rect 11612 14968 11664 15020
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 14832 15036 14884 15088
rect 15200 15079 15252 15088
rect 15200 15045 15209 15079
rect 15209 15045 15243 15079
rect 15243 15045 15252 15079
rect 15200 15036 15252 15045
rect 9588 14900 9640 14952
rect 12992 14968 13044 15020
rect 4804 14764 4856 14816
rect 5264 14764 5316 14816
rect 8024 14764 8076 14816
rect 8852 14764 8904 14816
rect 9588 14764 9640 14816
rect 10232 14764 10284 14816
rect 10784 14764 10836 14816
rect 12072 14764 12124 14816
rect 12900 14900 12952 14952
rect 13452 14900 13504 14952
rect 13820 14900 13872 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 14648 14968 14700 15020
rect 15660 14968 15712 15020
rect 16396 15036 16448 15088
rect 19064 15104 19116 15113
rect 19156 15104 19208 15156
rect 20904 15104 20956 15156
rect 21456 15104 21508 15156
rect 22560 15104 22612 15156
rect 23020 15104 23072 15156
rect 23572 15104 23624 15156
rect 16120 14968 16172 15020
rect 16764 14968 16816 15020
rect 17960 14968 18012 15020
rect 15108 14900 15160 14952
rect 15568 14900 15620 14952
rect 17592 14900 17644 14952
rect 18236 14968 18288 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 18788 14968 18840 15020
rect 19156 14968 19208 15020
rect 19524 14968 19576 15020
rect 12256 14832 12308 14884
rect 13268 14832 13320 14884
rect 15384 14832 15436 14884
rect 14004 14764 14056 14816
rect 14648 14764 14700 14816
rect 14740 14807 14792 14816
rect 14740 14773 14749 14807
rect 14749 14773 14783 14807
rect 14783 14773 14792 14807
rect 14740 14764 14792 14773
rect 14832 14764 14884 14816
rect 15844 14832 15896 14884
rect 17500 14832 17552 14884
rect 18144 14832 18196 14884
rect 16580 14764 16632 14816
rect 17776 14764 17828 14816
rect 19340 14900 19392 14952
rect 19892 14968 19944 15020
rect 20720 15036 20772 15088
rect 20168 14968 20220 15020
rect 20996 14968 21048 15020
rect 21456 15011 21508 15020
rect 21456 14977 21465 15011
rect 21465 14977 21499 15011
rect 21499 14977 21508 15011
rect 21456 14968 21508 14977
rect 22100 15011 22152 15020
rect 22100 14977 22109 15011
rect 22109 14977 22143 15011
rect 22143 14977 22152 15011
rect 22100 14968 22152 14977
rect 22284 14968 22336 15020
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 22928 14968 22980 15020
rect 23204 15036 23256 15088
rect 24032 15104 24084 15156
rect 26332 15147 26384 15156
rect 26332 15113 26341 15147
rect 26341 15113 26375 15147
rect 26375 15113 26384 15147
rect 26332 15104 26384 15113
rect 20260 14900 20312 14952
rect 19248 14832 19300 14884
rect 20076 14875 20128 14884
rect 20076 14841 20085 14875
rect 20085 14841 20119 14875
rect 20119 14841 20128 14875
rect 20076 14832 20128 14841
rect 21640 14900 21692 14952
rect 22008 14832 22060 14884
rect 18972 14764 19024 14816
rect 19984 14764 20036 14816
rect 20168 14764 20220 14816
rect 21180 14764 21232 14816
rect 21456 14764 21508 14816
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 22376 14764 22428 14816
rect 23388 14968 23440 15020
rect 24216 15036 24268 15088
rect 23480 14943 23532 14952
rect 23480 14909 23489 14943
rect 23489 14909 23523 14943
rect 23523 14909 23532 14943
rect 23480 14900 23532 14909
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 25320 14968 25372 15020
rect 26976 15104 27028 15156
rect 27436 15104 27488 15156
rect 27620 15104 27672 15156
rect 28908 15104 28960 15156
rect 24400 14943 24452 14952
rect 24400 14909 24409 14943
rect 24409 14909 24443 14943
rect 24443 14909 24452 14943
rect 24400 14900 24452 14909
rect 25044 14900 25096 14952
rect 25688 14900 25740 14952
rect 23020 14764 23072 14816
rect 23480 14764 23532 14816
rect 25228 14832 25280 14884
rect 25872 14832 25924 14884
rect 27344 15011 27396 15020
rect 27344 14977 27353 15011
rect 27353 14977 27387 15011
rect 27387 14977 27396 15011
rect 27344 14968 27396 14977
rect 27528 14968 27580 15020
rect 27804 15036 27856 15088
rect 28356 14968 28408 15020
rect 28816 15079 28868 15088
rect 28816 15045 28825 15079
rect 28825 15045 28859 15079
rect 28859 15045 28868 15079
rect 28816 15036 28868 15045
rect 29276 15079 29328 15088
rect 29276 15045 29285 15079
rect 29285 15045 29319 15079
rect 29319 15045 29328 15079
rect 29276 15036 29328 15045
rect 28908 15011 28960 15020
rect 28908 14977 28917 15011
rect 28917 14977 28951 15011
rect 28951 14977 28960 15011
rect 28908 14968 28960 14977
rect 29000 15011 29052 15020
rect 29000 14977 29014 15011
rect 29014 14977 29048 15011
rect 29048 14977 29052 15011
rect 29000 14968 29052 14977
rect 28816 14900 28868 14952
rect 29276 14900 29328 14952
rect 29644 15036 29696 15088
rect 29828 15011 29880 15020
rect 29828 14977 29837 15011
rect 29837 14977 29871 15011
rect 29871 14977 29880 15011
rect 29828 14968 29880 14977
rect 30748 15104 30800 15156
rect 32956 15104 33008 15156
rect 33416 15104 33468 15156
rect 31760 15036 31812 15088
rect 33232 15036 33284 15088
rect 29460 14943 29512 14952
rect 29460 14909 29469 14943
rect 29469 14909 29503 14943
rect 29503 14909 29512 14943
rect 29460 14900 29512 14909
rect 29644 14900 29696 14952
rect 30288 14900 30340 14952
rect 32220 14900 32272 14952
rect 32496 15011 32548 15020
rect 32496 14977 32505 15011
rect 32505 14977 32539 15011
rect 32539 14977 32548 15011
rect 32496 14968 32548 14977
rect 32588 15011 32640 15020
rect 32588 14977 32597 15011
rect 32597 14977 32631 15011
rect 32631 14977 32640 15011
rect 32588 14968 32640 14977
rect 33784 14968 33836 15020
rect 24032 14764 24084 14816
rect 24216 14807 24268 14816
rect 24216 14773 24225 14807
rect 24225 14773 24259 14807
rect 24259 14773 24268 14807
rect 24216 14764 24268 14773
rect 24768 14764 24820 14816
rect 26792 14764 26844 14816
rect 28540 14764 28592 14816
rect 28816 14764 28868 14816
rect 30656 14764 30708 14816
rect 31484 14807 31536 14816
rect 31484 14773 31493 14807
rect 31493 14773 31527 14807
rect 31527 14773 31536 14807
rect 31484 14764 31536 14773
rect 31576 14764 31628 14816
rect 31944 14764 31996 14816
rect 32404 14764 32456 14816
rect 33508 14764 33560 14816
rect 35072 15011 35124 15020
rect 35072 14977 35081 15011
rect 35081 14977 35115 15011
rect 35115 14977 35124 15011
rect 35072 14968 35124 14977
rect 34796 14900 34848 14952
rect 36176 14968 36228 15020
rect 34796 14807 34848 14816
rect 34796 14773 34805 14807
rect 34805 14773 34839 14807
rect 34839 14773 34848 14807
rect 34796 14764 34848 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3240 14560 3292 14612
rect 7104 14603 7156 14612
rect 7104 14569 7113 14603
rect 7113 14569 7147 14603
rect 7147 14569 7156 14603
rect 7104 14560 7156 14569
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 11060 14560 11112 14612
rect 12440 14560 12492 14612
rect 12900 14603 12952 14612
rect 12900 14569 12909 14603
rect 12909 14569 12943 14603
rect 12943 14569 12952 14603
rect 12900 14560 12952 14569
rect 13452 14560 13504 14612
rect 14832 14560 14884 14612
rect 15476 14560 15528 14612
rect 16212 14560 16264 14612
rect 4620 14356 4672 14408
rect 4804 14356 4856 14408
rect 5540 14492 5592 14544
rect 5356 14424 5408 14476
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 9312 14492 9364 14544
rect 6828 14424 6880 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 4436 14331 4488 14340
rect 4436 14297 4445 14331
rect 4445 14297 4479 14331
rect 4479 14297 4488 14331
rect 4436 14288 4488 14297
rect 4528 14331 4580 14340
rect 4528 14297 4537 14331
rect 4537 14297 4571 14331
rect 4571 14297 4580 14331
rect 4528 14288 4580 14297
rect 4620 14220 4672 14272
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 5264 14356 5316 14365
rect 5540 14356 5592 14408
rect 6368 14356 6420 14408
rect 8484 14424 8536 14476
rect 8852 14424 8904 14476
rect 5264 14220 5316 14272
rect 7472 14288 7524 14340
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 8392 14356 8444 14408
rect 8484 14288 8536 14340
rect 9680 14356 9732 14408
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 9956 14356 10008 14408
rect 10508 14424 10560 14476
rect 11336 14467 11388 14476
rect 11336 14433 11345 14467
rect 11345 14433 11379 14467
rect 11379 14433 11388 14467
rect 11336 14424 11388 14433
rect 12624 14492 12676 14544
rect 14096 14492 14148 14544
rect 14740 14492 14792 14544
rect 15936 14492 15988 14544
rect 17592 14535 17644 14544
rect 17592 14501 17601 14535
rect 17601 14501 17635 14535
rect 17635 14501 17644 14535
rect 17592 14492 17644 14501
rect 17684 14535 17736 14544
rect 17684 14501 17693 14535
rect 17693 14501 17727 14535
rect 17727 14501 17736 14535
rect 17684 14492 17736 14501
rect 18328 14560 18380 14612
rect 19064 14560 19116 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 21364 14603 21416 14612
rect 21364 14569 21373 14603
rect 21373 14569 21407 14603
rect 21407 14569 21416 14603
rect 21364 14560 21416 14569
rect 21456 14603 21508 14612
rect 21456 14569 21465 14603
rect 21465 14569 21499 14603
rect 21499 14569 21508 14603
rect 21456 14560 21508 14569
rect 21824 14560 21876 14612
rect 22192 14560 22244 14612
rect 23664 14560 23716 14612
rect 23848 14560 23900 14612
rect 24400 14560 24452 14612
rect 18420 14492 18472 14544
rect 10876 14356 10928 14408
rect 9404 14288 9456 14340
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 12900 14356 12952 14408
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 14464 14424 14516 14476
rect 17040 14424 17092 14476
rect 19248 14492 19300 14544
rect 8208 14220 8260 14272
rect 8392 14220 8444 14272
rect 12624 14288 12676 14340
rect 11244 14220 11296 14272
rect 11612 14220 11664 14272
rect 11888 14220 11940 14272
rect 12440 14220 12492 14272
rect 12808 14220 12860 14272
rect 13636 14399 13688 14408
rect 13636 14365 13645 14399
rect 13645 14365 13679 14399
rect 13679 14365 13688 14399
rect 13636 14356 13688 14365
rect 13820 14399 13872 14408
rect 13820 14365 13829 14399
rect 13829 14365 13863 14399
rect 13863 14365 13872 14399
rect 13820 14356 13872 14365
rect 15016 14356 15068 14408
rect 15200 14399 15252 14408
rect 15200 14365 15209 14399
rect 15209 14365 15243 14399
rect 15243 14365 15252 14399
rect 15200 14356 15252 14365
rect 14740 14331 14792 14340
rect 14740 14297 14749 14331
rect 14749 14297 14783 14331
rect 14783 14297 14792 14331
rect 14740 14288 14792 14297
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 15936 14288 15988 14340
rect 16580 14331 16632 14340
rect 16580 14297 16589 14331
rect 16589 14297 16623 14331
rect 16623 14297 16632 14331
rect 16580 14288 16632 14297
rect 17592 14356 17644 14408
rect 17868 14288 17920 14340
rect 17960 14288 18012 14340
rect 13452 14220 13504 14272
rect 15016 14220 15068 14272
rect 16120 14220 16172 14272
rect 17224 14220 17276 14272
rect 18144 14356 18196 14408
rect 18328 14356 18380 14408
rect 20536 14424 20588 14476
rect 21364 14424 21416 14476
rect 23112 14424 23164 14476
rect 26056 14424 26108 14476
rect 18788 14356 18840 14408
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 18972 14356 19024 14408
rect 19800 14288 19852 14340
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20260 14356 20312 14365
rect 20444 14356 20496 14408
rect 20904 14356 20956 14408
rect 22008 14356 22060 14408
rect 22284 14356 22336 14408
rect 22468 14356 22520 14408
rect 23204 14356 23256 14408
rect 23480 14356 23532 14408
rect 24860 14399 24912 14408
rect 24860 14365 24869 14399
rect 24869 14365 24903 14399
rect 24903 14365 24912 14399
rect 24860 14356 24912 14365
rect 24952 14356 25004 14408
rect 25596 14399 25648 14408
rect 25596 14365 25605 14399
rect 25605 14365 25639 14399
rect 25639 14365 25648 14399
rect 25596 14356 25648 14365
rect 25688 14356 25740 14408
rect 27436 14492 27488 14544
rect 18328 14220 18380 14272
rect 18512 14220 18564 14272
rect 18788 14220 18840 14272
rect 19156 14220 19208 14272
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 21364 14220 21416 14272
rect 22560 14220 22612 14272
rect 23940 14288 23992 14340
rect 26056 14220 26108 14272
rect 27344 14399 27396 14408
rect 27344 14365 27353 14399
rect 27353 14365 27387 14399
rect 27387 14365 27396 14399
rect 27344 14356 27396 14365
rect 27620 14560 27672 14612
rect 29460 14560 29512 14612
rect 29736 14560 29788 14612
rect 32496 14560 32548 14612
rect 28172 14492 28224 14544
rect 28632 14492 28684 14544
rect 28724 14492 28776 14544
rect 29828 14492 29880 14544
rect 31576 14492 31628 14544
rect 31944 14492 31996 14544
rect 34520 14492 34572 14544
rect 29276 14424 29328 14476
rect 29460 14424 29512 14476
rect 26976 14288 27028 14340
rect 27804 14399 27856 14408
rect 27804 14365 27813 14399
rect 27813 14365 27847 14399
rect 27847 14365 27856 14399
rect 27804 14356 27856 14365
rect 27988 14399 28040 14408
rect 27988 14365 27997 14399
rect 27997 14365 28031 14399
rect 28031 14365 28040 14399
rect 27988 14356 28040 14365
rect 28172 14399 28224 14408
rect 28172 14365 28181 14399
rect 28181 14365 28215 14399
rect 28215 14365 28224 14399
rect 28172 14356 28224 14365
rect 30288 14356 30340 14408
rect 30564 14399 30616 14408
rect 30564 14365 30574 14399
rect 30574 14365 30608 14399
rect 30608 14365 30616 14399
rect 31116 14424 31168 14476
rect 30564 14356 30616 14365
rect 31024 14356 31076 14408
rect 31484 14356 31536 14408
rect 27896 14288 27948 14340
rect 27712 14220 27764 14272
rect 29460 14288 29512 14340
rect 29644 14288 29696 14340
rect 28908 14220 28960 14272
rect 30104 14220 30156 14272
rect 30564 14220 30616 14272
rect 32128 14220 32180 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 5264 14016 5316 14068
rect 5724 14016 5776 14068
rect 6368 14016 6420 14068
rect 4804 13991 4856 14000
rect 4804 13957 4813 13991
rect 4813 13957 4847 13991
rect 4847 13957 4856 13991
rect 4804 13948 4856 13957
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 3976 13880 4028 13932
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 8392 14016 8444 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 11336 14016 11388 14068
rect 12716 14059 12768 14068
rect 12716 14025 12725 14059
rect 12725 14025 12759 14059
rect 12759 14025 12768 14059
rect 12716 14016 12768 14025
rect 14648 14016 14700 14068
rect 8024 13991 8076 14000
rect 8024 13957 8033 13991
rect 8033 13957 8067 13991
rect 8067 13957 8076 13991
rect 8024 13948 8076 13957
rect 4712 13812 4764 13864
rect 5448 13880 5500 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 6092 13923 6144 13932
rect 6092 13889 6101 13923
rect 6101 13889 6135 13923
rect 6135 13889 6144 13923
rect 6092 13880 6144 13889
rect 7380 13880 7432 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 7656 13880 7708 13932
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 7932 13880 7984 13889
rect 5540 13744 5592 13796
rect 5356 13676 5408 13728
rect 5908 13812 5960 13864
rect 8484 13923 8536 13932
rect 8484 13889 8493 13923
rect 8493 13889 8527 13923
rect 8527 13889 8536 13923
rect 8484 13880 8536 13889
rect 8852 13880 8904 13932
rect 9404 13880 9456 13932
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 9772 13880 9824 13932
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10140 13880 10192 13932
rect 10692 13948 10744 14000
rect 9588 13812 9640 13864
rect 8208 13787 8260 13796
rect 8208 13753 8217 13787
rect 8217 13753 8251 13787
rect 8251 13753 8260 13787
rect 8208 13744 8260 13753
rect 10324 13744 10376 13796
rect 11060 13948 11112 14000
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 13912 13948 13964 14000
rect 15108 13991 15160 14000
rect 15108 13957 15117 13991
rect 15117 13957 15151 13991
rect 15151 13957 15160 13991
rect 15108 13948 15160 13957
rect 11888 13744 11940 13796
rect 12624 13880 12676 13932
rect 13176 13923 13228 13932
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 13452 13880 13504 13932
rect 13820 13880 13872 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 13636 13812 13688 13864
rect 14464 13880 14516 13932
rect 14832 13880 14884 13932
rect 15476 14059 15528 14068
rect 15476 14025 15485 14059
rect 15485 14025 15519 14059
rect 15519 14025 15528 14059
rect 15476 14016 15528 14025
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 17776 14016 17828 14068
rect 18328 14016 18380 14068
rect 19156 14016 19208 14068
rect 20260 14016 20312 14068
rect 20444 14016 20496 14068
rect 21180 14016 21232 14068
rect 23388 14016 23440 14068
rect 26608 14059 26660 14068
rect 26608 14025 26617 14059
rect 26617 14025 26651 14059
rect 26651 14025 26660 14059
rect 26608 14016 26660 14025
rect 26976 14016 27028 14068
rect 27988 14016 28040 14068
rect 16580 13948 16632 14000
rect 15384 13880 15436 13932
rect 16396 13880 16448 13932
rect 17684 13948 17736 14000
rect 17868 13948 17920 14000
rect 18880 13948 18932 14000
rect 19432 13948 19484 14000
rect 19708 13991 19760 14000
rect 19708 13957 19717 13991
rect 19717 13957 19751 13991
rect 19751 13957 19760 13991
rect 19708 13948 19760 13957
rect 19892 13991 19944 14000
rect 19892 13957 19927 13991
rect 19927 13957 19944 13991
rect 19892 13948 19944 13957
rect 19800 13880 19852 13932
rect 15476 13812 15528 13864
rect 18972 13812 19024 13864
rect 19708 13812 19760 13864
rect 20536 13812 20588 13864
rect 20720 13812 20772 13864
rect 15568 13744 15620 13796
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 12992 13676 13044 13728
rect 16764 13744 16816 13796
rect 17868 13744 17920 13796
rect 23204 13744 23256 13796
rect 24952 13855 25004 13864
rect 24952 13821 24961 13855
rect 24961 13821 24995 13855
rect 24995 13821 25004 13855
rect 24952 13812 25004 13821
rect 25688 13880 25740 13932
rect 27436 13948 27488 14000
rect 29920 14016 29972 14068
rect 32956 14016 33008 14068
rect 25596 13812 25648 13864
rect 26608 13812 26660 13864
rect 26976 13744 27028 13796
rect 27620 13880 27672 13932
rect 28172 13923 28224 13932
rect 28172 13889 28181 13923
rect 28181 13889 28215 13923
rect 28215 13889 28224 13923
rect 28172 13880 28224 13889
rect 28264 13923 28316 13932
rect 28264 13889 28273 13923
rect 28273 13889 28307 13923
rect 28307 13889 28316 13923
rect 28264 13880 28316 13889
rect 28356 13923 28408 13932
rect 28356 13889 28365 13923
rect 28365 13889 28399 13923
rect 28399 13889 28408 13923
rect 28356 13880 28408 13889
rect 28724 13880 28776 13932
rect 28908 13923 28960 13932
rect 28908 13889 28912 13923
rect 28912 13889 28946 13923
rect 28946 13889 28960 13923
rect 28908 13880 28960 13889
rect 29092 13923 29144 13932
rect 29092 13889 29101 13923
rect 29101 13889 29135 13923
rect 29135 13889 29144 13923
rect 29092 13880 29144 13889
rect 29368 13889 29388 13922
rect 29388 13889 29420 13922
rect 29368 13870 29420 13889
rect 17316 13676 17368 13728
rect 19340 13676 19392 13728
rect 19883 13719 19935 13728
rect 19883 13685 19892 13719
rect 19892 13685 19926 13719
rect 19926 13685 19935 13719
rect 19883 13676 19935 13685
rect 21640 13676 21692 13728
rect 23940 13676 23992 13728
rect 26240 13676 26292 13728
rect 27160 13676 27212 13728
rect 27988 13855 28040 13864
rect 27988 13821 27997 13855
rect 27997 13821 28031 13855
rect 28031 13821 28040 13855
rect 27988 13812 28040 13821
rect 28632 13855 28684 13864
rect 28632 13821 28641 13855
rect 28641 13821 28675 13855
rect 28675 13821 28684 13855
rect 28632 13812 28684 13821
rect 32128 13991 32180 14000
rect 32128 13957 32137 13991
rect 32137 13957 32171 13991
rect 32171 13957 32180 13991
rect 32128 13948 32180 13957
rect 27988 13676 28040 13728
rect 28264 13676 28316 13728
rect 28816 13744 28868 13796
rect 28908 13744 28960 13796
rect 29460 13744 29512 13796
rect 30104 13880 30156 13932
rect 30656 13923 30708 13932
rect 30656 13889 30665 13923
rect 30665 13889 30699 13923
rect 30699 13889 30708 13923
rect 30656 13880 30708 13889
rect 33600 13880 33652 13932
rect 29920 13744 29972 13796
rect 30196 13812 30248 13864
rect 31944 13812 31996 13864
rect 31760 13676 31812 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4620 13472 4672 13524
rect 6092 13472 6144 13524
rect 9496 13472 9548 13524
rect 10140 13472 10192 13524
rect 6736 13404 6788 13456
rect 15660 13472 15712 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 17500 13472 17552 13524
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 18696 13515 18748 13524
rect 18696 13481 18705 13515
rect 18705 13481 18739 13515
rect 18739 13481 18748 13515
rect 18696 13472 18748 13481
rect 19340 13472 19392 13524
rect 5356 13336 5408 13388
rect 5540 13336 5592 13388
rect 13360 13404 13412 13456
rect 4712 13200 4764 13252
rect 5724 13268 5776 13320
rect 6092 13268 6144 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 9404 13268 9456 13320
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 12072 13336 12124 13388
rect 5540 13200 5592 13252
rect 9680 13200 9732 13252
rect 10232 13200 10284 13252
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11060 13268 11112 13320
rect 13728 13336 13780 13388
rect 14096 13336 14148 13388
rect 17592 13404 17644 13456
rect 20352 13472 20404 13524
rect 21088 13472 21140 13524
rect 11244 13200 11296 13252
rect 6920 13132 6972 13184
rect 8944 13132 8996 13184
rect 13176 13268 13228 13320
rect 15016 13200 15068 13252
rect 16028 13268 16080 13320
rect 16212 13311 16264 13320
rect 16212 13277 16221 13311
rect 16221 13277 16255 13311
rect 16255 13277 16264 13311
rect 16212 13268 16264 13277
rect 18052 13336 18104 13388
rect 17868 13268 17920 13320
rect 18328 13268 18380 13320
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 15660 13132 15712 13184
rect 18144 13200 18196 13252
rect 19156 13200 19208 13252
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 20168 13336 20220 13388
rect 20444 13336 20496 13388
rect 20260 13311 20312 13320
rect 20260 13277 20269 13311
rect 20269 13277 20303 13311
rect 20303 13277 20312 13311
rect 20260 13268 20312 13277
rect 20352 13311 20404 13320
rect 20352 13277 20362 13311
rect 20362 13277 20396 13311
rect 20396 13277 20404 13311
rect 20352 13268 20404 13277
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 20076 13200 20128 13252
rect 20168 13200 20220 13252
rect 17500 13175 17552 13184
rect 17500 13141 17509 13175
rect 17509 13141 17543 13175
rect 17543 13141 17552 13175
rect 17500 13132 17552 13141
rect 17592 13132 17644 13184
rect 18420 13132 18472 13184
rect 19524 13132 19576 13184
rect 20260 13132 20312 13184
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 22100 13472 22152 13524
rect 26424 13472 26476 13524
rect 26700 13472 26752 13524
rect 28172 13472 28224 13524
rect 28724 13472 28776 13524
rect 28908 13472 28960 13524
rect 31576 13472 31628 13524
rect 21548 13404 21600 13456
rect 23112 13404 23164 13456
rect 27344 13404 27396 13456
rect 31760 13472 31812 13524
rect 34796 13472 34848 13524
rect 33048 13404 33100 13456
rect 33140 13447 33192 13456
rect 33140 13413 33149 13447
rect 33149 13413 33183 13447
rect 33183 13413 33192 13447
rect 33140 13404 33192 13413
rect 25688 13379 25740 13388
rect 25688 13345 25697 13379
rect 25697 13345 25731 13379
rect 25731 13345 25740 13379
rect 25688 13336 25740 13345
rect 21640 13311 21692 13320
rect 21640 13277 21649 13311
rect 21649 13277 21683 13311
rect 21683 13277 21692 13311
rect 21640 13268 21692 13277
rect 21088 13200 21140 13252
rect 21916 13268 21968 13320
rect 24768 13268 24820 13320
rect 23664 13200 23716 13252
rect 25596 13311 25648 13320
rect 25596 13277 25605 13311
rect 25605 13277 25639 13311
rect 25639 13277 25648 13311
rect 25596 13268 25648 13277
rect 26056 13268 26108 13320
rect 26608 13268 26660 13320
rect 28080 13336 28132 13388
rect 29000 13336 29052 13388
rect 31852 13379 31904 13388
rect 31852 13345 31861 13379
rect 31861 13345 31895 13379
rect 31895 13345 31904 13379
rect 31852 13336 31904 13345
rect 35440 13404 35492 13456
rect 35348 13336 35400 13388
rect 26884 13268 26936 13320
rect 26976 13311 27028 13320
rect 26976 13277 26985 13311
rect 26985 13277 27019 13311
rect 27019 13277 27028 13311
rect 26976 13268 27028 13277
rect 28448 13268 28500 13320
rect 28632 13268 28684 13320
rect 29276 13268 29328 13320
rect 29920 13268 29972 13320
rect 31944 13311 31996 13320
rect 31944 13277 31953 13311
rect 31953 13277 31987 13311
rect 31987 13277 31996 13311
rect 31944 13268 31996 13277
rect 32496 13268 32548 13320
rect 33876 13268 33928 13320
rect 34336 13311 34388 13320
rect 34336 13277 34345 13311
rect 34345 13277 34379 13311
rect 34379 13277 34388 13311
rect 34336 13268 34388 13277
rect 27160 13200 27212 13252
rect 29000 13200 29052 13252
rect 31668 13243 31720 13252
rect 31668 13209 31677 13243
rect 31677 13209 31711 13243
rect 31711 13209 31720 13243
rect 31668 13200 31720 13209
rect 33048 13200 33100 13252
rect 22284 13132 22336 13184
rect 23572 13132 23624 13184
rect 26792 13132 26844 13184
rect 27620 13132 27672 13184
rect 32128 13175 32180 13184
rect 32128 13141 32137 13175
rect 32137 13141 32171 13175
rect 32171 13141 32180 13175
rect 32128 13132 32180 13141
rect 34520 13175 34572 13184
rect 34520 13141 34529 13175
rect 34529 13141 34563 13175
rect 34563 13141 34572 13175
rect 34520 13132 34572 13141
rect 34796 13175 34848 13184
rect 34796 13141 34805 13175
rect 34805 13141 34839 13175
rect 34839 13141 34848 13175
rect 34796 13132 34848 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 8484 12928 8536 12980
rect 9036 12928 9088 12980
rect 5724 12903 5776 12912
rect 5724 12869 5733 12903
rect 5733 12869 5767 12903
rect 5767 12869 5776 12903
rect 5724 12860 5776 12869
rect 5908 12792 5960 12844
rect 7196 12860 7248 12912
rect 7656 12860 7708 12912
rect 10416 12928 10468 12980
rect 10968 12928 11020 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 15752 12971 15804 12980
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 17316 12928 17368 12980
rect 18604 12928 18656 12980
rect 19708 12928 19760 12980
rect 19984 12928 20036 12980
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 6920 12724 6972 12776
rect 7472 12724 7524 12776
rect 7564 12767 7616 12776
rect 7564 12733 7573 12767
rect 7573 12733 7607 12767
rect 7607 12733 7616 12767
rect 7564 12724 7616 12733
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 8300 12835 8352 12844
rect 8300 12801 8309 12835
rect 8309 12801 8343 12835
rect 8343 12801 8352 12835
rect 8300 12792 8352 12801
rect 8208 12724 8260 12776
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9680 12860 9732 12912
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 9220 12792 9272 12844
rect 10140 12792 10192 12844
rect 12072 12860 12124 12912
rect 14188 12860 14240 12912
rect 10324 12724 10376 12776
rect 10600 12724 10652 12776
rect 8668 12656 8720 12708
rect 9220 12656 9272 12708
rect 9312 12656 9364 12708
rect 9588 12656 9640 12708
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 11336 12792 11388 12844
rect 11796 12792 11848 12844
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 15476 12792 15528 12844
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 15568 12792 15620 12801
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 16028 12792 16080 12844
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 14556 12724 14608 12776
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 17776 12792 17828 12844
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 19248 12792 19300 12844
rect 19800 12792 19852 12844
rect 19892 12792 19944 12844
rect 21180 12928 21232 12980
rect 25228 12928 25280 12980
rect 26240 12928 26292 12980
rect 26700 12928 26752 12980
rect 20628 12860 20680 12912
rect 20996 12860 21048 12912
rect 21732 12860 21784 12912
rect 24584 12860 24636 12912
rect 25872 12860 25924 12912
rect 21364 12792 21416 12844
rect 22100 12792 22152 12844
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 22560 12792 22612 12801
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 23664 12835 23716 12844
rect 23664 12801 23673 12835
rect 23673 12801 23707 12835
rect 23707 12801 23716 12835
rect 23664 12792 23716 12801
rect 24216 12835 24268 12844
rect 24216 12801 24225 12835
rect 24225 12801 24259 12835
rect 24259 12801 24268 12835
rect 24216 12792 24268 12801
rect 25596 12792 25648 12844
rect 26608 12860 26660 12912
rect 27252 12860 27304 12912
rect 27344 12860 27396 12912
rect 28172 12860 28224 12912
rect 19524 12724 19576 12776
rect 23020 12724 23072 12776
rect 24400 12767 24452 12776
rect 24400 12733 24409 12767
rect 24409 12733 24443 12767
rect 24443 12733 24452 12767
rect 24400 12724 24452 12733
rect 11428 12656 11480 12708
rect 12532 12656 12584 12708
rect 13176 12656 13228 12708
rect 13360 12656 13412 12708
rect 15200 12656 15252 12708
rect 15752 12656 15804 12708
rect 17316 12656 17368 12708
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 8576 12588 8628 12640
rect 8760 12588 8812 12640
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 10324 12588 10376 12640
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 12072 12588 12124 12640
rect 13084 12588 13136 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 16304 12588 16356 12640
rect 16948 12588 17000 12640
rect 18144 12656 18196 12708
rect 24216 12656 24268 12708
rect 24768 12724 24820 12776
rect 25504 12767 25556 12776
rect 25504 12733 25513 12767
rect 25513 12733 25547 12767
rect 25547 12733 25556 12767
rect 25504 12724 25556 12733
rect 25688 12724 25740 12776
rect 26700 12835 26752 12844
rect 26700 12801 26709 12835
rect 26709 12801 26743 12835
rect 26743 12801 26752 12835
rect 26700 12792 26752 12801
rect 27068 12835 27120 12844
rect 27068 12801 27077 12835
rect 27077 12801 27111 12835
rect 27111 12801 27120 12835
rect 27068 12792 27120 12801
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 24676 12699 24728 12708
rect 24676 12665 24685 12699
rect 24685 12665 24719 12699
rect 24719 12665 24728 12699
rect 24676 12656 24728 12665
rect 24952 12656 25004 12708
rect 25872 12699 25924 12708
rect 25872 12665 25881 12699
rect 25881 12665 25915 12699
rect 25915 12665 25924 12699
rect 25872 12656 25924 12665
rect 26792 12724 26844 12776
rect 27160 12724 27212 12776
rect 27896 12792 27948 12844
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 28724 12792 28776 12844
rect 29000 12835 29052 12844
rect 29000 12801 29009 12835
rect 29009 12801 29043 12835
rect 29043 12801 29052 12835
rect 29000 12792 29052 12801
rect 29460 12792 29512 12844
rect 27620 12724 27672 12776
rect 30472 12792 30524 12844
rect 30748 12835 30800 12844
rect 30748 12801 30755 12835
rect 30755 12801 30800 12835
rect 30748 12792 30800 12801
rect 32312 12928 32364 12980
rect 32496 12928 32548 12980
rect 33416 12928 33468 12980
rect 33692 12928 33744 12980
rect 31024 12835 31076 12844
rect 31024 12801 31038 12835
rect 31038 12801 31072 12835
rect 31072 12801 31076 12835
rect 31024 12792 31076 12801
rect 31760 12792 31812 12844
rect 26884 12656 26936 12708
rect 28080 12656 28132 12708
rect 20536 12631 20588 12640
rect 20536 12597 20545 12631
rect 20545 12597 20579 12631
rect 20579 12597 20588 12631
rect 20536 12588 20588 12597
rect 22744 12588 22796 12640
rect 28264 12588 28316 12640
rect 30748 12656 30800 12708
rect 30932 12656 30984 12708
rect 28724 12588 28776 12640
rect 28816 12631 28868 12640
rect 28816 12597 28825 12631
rect 28825 12597 28859 12631
rect 28859 12597 28868 12631
rect 28816 12588 28868 12597
rect 29092 12588 29144 12640
rect 32864 12588 32916 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3976 12427 4028 12436
rect 3976 12393 3985 12427
rect 3985 12393 4019 12427
rect 4019 12393 4028 12427
rect 3976 12384 4028 12393
rect 4712 12384 4764 12436
rect 5448 12384 5500 12436
rect 8208 12384 8260 12436
rect 5540 12316 5592 12368
rect 8392 12316 8444 12368
rect 2412 12248 2464 12300
rect 5724 12248 5776 12300
rect 7012 12248 7064 12300
rect 7564 12248 7616 12300
rect 4344 12180 4396 12232
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 5264 12180 5316 12232
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 8300 12248 8352 12300
rect 4712 12112 4764 12164
rect 4160 12044 4212 12096
rect 4436 12044 4488 12096
rect 4804 12044 4856 12096
rect 6920 12112 6972 12164
rect 7564 12155 7616 12164
rect 7564 12121 7573 12155
rect 7573 12121 7607 12155
rect 7607 12121 7616 12155
rect 7564 12112 7616 12121
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 9036 12384 9088 12436
rect 9404 12384 9456 12436
rect 8944 12316 8996 12368
rect 9864 12384 9916 12436
rect 9772 12316 9824 12368
rect 10232 12316 10284 12368
rect 10876 12316 10928 12368
rect 10968 12316 11020 12368
rect 11152 12316 11204 12368
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 9312 12248 9364 12300
rect 9404 12248 9456 12300
rect 10600 12248 10652 12300
rect 11336 12291 11388 12300
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 9680 12180 9732 12232
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 10048 12180 10100 12232
rect 11336 12257 11345 12291
rect 11345 12257 11379 12291
rect 11379 12257 11388 12291
rect 11336 12248 11388 12257
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 8116 12044 8168 12096
rect 9312 12112 9364 12164
rect 9496 12155 9548 12164
rect 9496 12121 9505 12155
rect 9505 12121 9539 12155
rect 9539 12121 9548 12155
rect 9496 12112 9548 12121
rect 10968 12155 11020 12164
rect 10968 12121 10977 12155
rect 10977 12121 11011 12155
rect 11011 12121 11020 12155
rect 10968 12112 11020 12121
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11244 12223 11296 12232
rect 11244 12189 11253 12223
rect 11253 12189 11287 12223
rect 11287 12189 11296 12223
rect 11244 12180 11296 12189
rect 12900 12316 12952 12368
rect 12072 12291 12124 12300
rect 12072 12257 12081 12291
rect 12081 12257 12115 12291
rect 12115 12257 12124 12291
rect 12072 12248 12124 12257
rect 12164 12291 12216 12300
rect 12164 12257 12173 12291
rect 12173 12257 12207 12291
rect 12207 12257 12216 12291
rect 12164 12248 12216 12257
rect 13452 12316 13504 12368
rect 14648 12384 14700 12436
rect 14740 12427 14792 12436
rect 14740 12393 14749 12427
rect 14749 12393 14783 12427
rect 14783 12393 14792 12427
rect 14740 12384 14792 12393
rect 15200 12427 15252 12436
rect 15200 12393 15209 12427
rect 15209 12393 15243 12427
rect 15243 12393 15252 12427
rect 15200 12384 15252 12393
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 18052 12427 18104 12436
rect 18052 12393 18061 12427
rect 18061 12393 18095 12427
rect 18095 12393 18104 12427
rect 18052 12384 18104 12393
rect 18696 12384 18748 12436
rect 18972 12384 19024 12436
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 20168 12384 20220 12436
rect 20812 12384 20864 12436
rect 21364 12427 21416 12436
rect 21364 12393 21373 12427
rect 21373 12393 21407 12427
rect 21407 12393 21416 12427
rect 21364 12384 21416 12393
rect 22468 12384 22520 12436
rect 23020 12384 23072 12436
rect 23204 12384 23256 12436
rect 23388 12384 23440 12436
rect 23664 12384 23716 12436
rect 23756 12384 23808 12436
rect 24308 12384 24360 12436
rect 24400 12427 24452 12436
rect 24400 12393 24409 12427
rect 24409 12393 24443 12427
rect 24443 12393 24452 12427
rect 24400 12384 24452 12393
rect 26148 12384 26200 12436
rect 28448 12384 28500 12436
rect 28724 12384 28776 12436
rect 32220 12384 32272 12436
rect 11704 12180 11756 12232
rect 11888 12180 11940 12232
rect 11980 12223 12032 12232
rect 11980 12189 11989 12223
rect 11989 12189 12023 12223
rect 12023 12189 12032 12223
rect 11980 12180 12032 12189
rect 12440 12180 12492 12232
rect 9772 12044 9824 12096
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 10324 12044 10376 12053
rect 10508 12044 10560 12096
rect 10692 12044 10744 12096
rect 13820 12180 13872 12232
rect 14004 12180 14056 12232
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 12716 12044 12768 12096
rect 13544 12087 13596 12096
rect 13544 12053 13553 12087
rect 13553 12053 13587 12087
rect 13587 12053 13596 12087
rect 13544 12044 13596 12053
rect 13728 12087 13780 12096
rect 13728 12053 13755 12087
rect 13755 12053 13780 12087
rect 13728 12044 13780 12053
rect 14556 12180 14608 12232
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 16120 12223 16172 12232
rect 16120 12189 16129 12223
rect 16129 12189 16163 12223
rect 16163 12189 16172 12223
rect 16120 12180 16172 12189
rect 16212 12223 16264 12232
rect 16212 12189 16222 12223
rect 16222 12189 16256 12223
rect 16256 12189 16264 12223
rect 16212 12180 16264 12189
rect 14648 12155 14700 12164
rect 14648 12121 14657 12155
rect 14657 12121 14691 12155
rect 14691 12121 14700 12155
rect 14648 12112 14700 12121
rect 19708 12316 19760 12368
rect 19800 12316 19852 12368
rect 21088 12316 21140 12368
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 18604 12248 18656 12300
rect 18972 12248 19024 12300
rect 19340 12248 19392 12300
rect 16488 12223 16540 12232
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 16580 12223 16632 12232
rect 16580 12189 16594 12223
rect 16594 12189 16628 12223
rect 16628 12189 16632 12223
rect 16580 12180 16632 12189
rect 16396 12155 16448 12164
rect 16396 12121 16405 12155
rect 16405 12121 16439 12155
rect 16439 12121 16448 12155
rect 17040 12180 17092 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 18144 12180 18196 12232
rect 16396 12112 16448 12121
rect 16948 12112 17000 12164
rect 18420 12112 18472 12164
rect 17868 12044 17920 12096
rect 21548 12248 21600 12300
rect 18880 12155 18932 12164
rect 18880 12121 18907 12155
rect 18907 12121 18932 12155
rect 18880 12112 18932 12121
rect 19156 12112 19208 12164
rect 19800 12112 19852 12164
rect 19892 12112 19944 12164
rect 20076 12112 20128 12164
rect 21272 12180 21324 12232
rect 29736 12316 29788 12368
rect 22560 12291 22612 12300
rect 22560 12257 22569 12291
rect 22569 12257 22603 12291
rect 22603 12257 22612 12291
rect 22560 12248 22612 12257
rect 26516 12248 26568 12300
rect 26884 12248 26936 12300
rect 27620 12248 27672 12300
rect 28264 12248 28316 12300
rect 28448 12248 28500 12300
rect 28816 12248 28868 12300
rect 33140 12427 33192 12436
rect 33140 12393 33149 12427
rect 33149 12393 33183 12427
rect 33183 12393 33192 12427
rect 33140 12384 33192 12393
rect 24032 12223 24084 12232
rect 24032 12189 24041 12223
rect 24041 12189 24075 12223
rect 24075 12189 24084 12223
rect 24032 12180 24084 12189
rect 24308 12180 24360 12232
rect 20628 12112 20680 12164
rect 21088 12155 21140 12164
rect 21088 12121 21097 12155
rect 21097 12121 21131 12155
rect 21131 12121 21140 12155
rect 21088 12112 21140 12121
rect 21456 12112 21508 12164
rect 21916 12112 21968 12164
rect 19432 12044 19484 12096
rect 20720 12044 20772 12096
rect 21180 12044 21232 12096
rect 22560 12112 22612 12164
rect 23388 12155 23440 12164
rect 23388 12121 23397 12155
rect 23397 12121 23431 12155
rect 23431 12121 23440 12155
rect 23388 12112 23440 12121
rect 23572 12112 23624 12164
rect 23940 12112 23992 12164
rect 24400 12112 24452 12164
rect 25872 12180 25924 12232
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 26608 12180 26660 12189
rect 26792 12180 26844 12232
rect 27160 12223 27212 12232
rect 27160 12189 27169 12223
rect 27169 12189 27203 12223
rect 27203 12189 27212 12223
rect 27160 12180 27212 12189
rect 27344 12223 27396 12232
rect 27344 12189 27353 12223
rect 27353 12189 27387 12223
rect 27387 12189 27396 12223
rect 27344 12180 27396 12189
rect 28908 12223 28960 12232
rect 28908 12189 28917 12223
rect 28917 12189 28951 12223
rect 28951 12189 28960 12223
rect 28908 12180 28960 12189
rect 32128 12180 32180 12232
rect 26332 12112 26384 12164
rect 27620 12155 27672 12164
rect 27620 12121 27629 12155
rect 27629 12121 27663 12155
rect 27663 12121 27672 12155
rect 27620 12112 27672 12121
rect 28080 12112 28132 12164
rect 28264 12112 28316 12164
rect 32496 12223 32548 12232
rect 32496 12189 32505 12223
rect 32505 12189 32539 12223
rect 32539 12189 32548 12223
rect 32496 12180 32548 12189
rect 32680 12180 32732 12232
rect 32956 12223 33008 12232
rect 32956 12189 32965 12223
rect 32965 12189 32999 12223
rect 32999 12189 33008 12223
rect 32956 12180 33008 12189
rect 34520 12180 34572 12232
rect 35256 12112 35308 12164
rect 23020 12044 23072 12096
rect 24860 12044 24912 12096
rect 25044 12044 25096 12096
rect 25228 12044 25280 12096
rect 26240 12044 26292 12096
rect 27160 12044 27212 12096
rect 27988 12044 28040 12096
rect 28724 12087 28776 12096
rect 28724 12053 28733 12087
rect 28733 12053 28767 12087
rect 28767 12053 28776 12087
rect 28724 12044 28776 12053
rect 31484 12044 31536 12096
rect 32036 12044 32088 12096
rect 32588 12044 32640 12096
rect 32772 12087 32824 12096
rect 32772 12053 32781 12087
rect 32781 12053 32815 12087
rect 32815 12053 32824 12087
rect 32772 12044 32824 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 4160 11840 4212 11892
rect 4528 11840 4580 11892
rect 4712 11883 4764 11892
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 5264 11840 5316 11892
rect 3884 11772 3936 11824
rect 7564 11840 7616 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 7840 11840 7892 11892
rect 8208 11840 8260 11892
rect 8392 11840 8444 11892
rect 9496 11840 9548 11892
rect 9956 11840 10008 11892
rect 10784 11840 10836 11892
rect 11244 11840 11296 11892
rect 12900 11840 12952 11892
rect 13176 11840 13228 11892
rect 14648 11840 14700 11892
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 4804 11704 4856 11756
rect 4344 11568 4396 11620
rect 4804 11568 4856 11620
rect 5356 11704 5408 11756
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 7472 11704 7524 11756
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 8668 11704 8720 11756
rect 9220 11704 9272 11756
rect 12808 11772 12860 11824
rect 13728 11772 13780 11824
rect 9680 11704 9732 11756
rect 10416 11704 10468 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 10968 11704 11020 11713
rect 11244 11704 11296 11756
rect 12072 11704 12124 11756
rect 12256 11704 12308 11756
rect 12992 11704 13044 11756
rect 5816 11568 5868 11620
rect 6460 11679 6512 11688
rect 6460 11645 6469 11679
rect 6469 11645 6503 11679
rect 6503 11645 6512 11679
rect 6460 11636 6512 11645
rect 8208 11568 8260 11620
rect 5540 11500 5592 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 6184 11500 6236 11552
rect 7288 11500 7340 11552
rect 7748 11500 7800 11552
rect 8484 11500 8536 11552
rect 8576 11500 8628 11552
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 9772 11636 9824 11688
rect 9864 11636 9916 11688
rect 11060 11636 11112 11688
rect 9312 11568 9364 11620
rect 11888 11636 11940 11688
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 10232 11500 10284 11552
rect 13268 11704 13320 11756
rect 16120 11840 16172 11892
rect 25136 11840 25188 11892
rect 26792 11840 26844 11892
rect 26976 11840 27028 11892
rect 27988 11840 28040 11892
rect 28172 11840 28224 11892
rect 15384 11772 15436 11824
rect 16672 11772 16724 11824
rect 17868 11772 17920 11824
rect 18420 11815 18472 11824
rect 18420 11781 18429 11815
rect 18429 11781 18463 11815
rect 18463 11781 18472 11815
rect 18420 11772 18472 11781
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 13820 11636 13872 11688
rect 14740 11636 14792 11688
rect 14832 11636 14884 11688
rect 16948 11636 17000 11688
rect 12256 11568 12308 11620
rect 13084 11568 13136 11620
rect 15660 11500 15712 11552
rect 17132 11568 17184 11620
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 19064 11772 19116 11824
rect 18144 11704 18196 11713
rect 18052 11636 18104 11688
rect 18512 11636 18564 11688
rect 19432 11704 19484 11756
rect 20352 11772 20404 11824
rect 20628 11772 20680 11824
rect 20720 11815 20772 11824
rect 20720 11781 20761 11815
rect 20761 11781 20772 11815
rect 20720 11772 20772 11781
rect 23388 11772 23440 11824
rect 23664 11772 23716 11824
rect 19616 11636 19668 11688
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 21364 11704 21416 11756
rect 22008 11704 22060 11756
rect 22284 11636 22336 11688
rect 23296 11704 23348 11756
rect 24860 11772 24912 11824
rect 25412 11772 25464 11824
rect 26516 11772 26568 11824
rect 28540 11815 28592 11824
rect 24768 11704 24820 11756
rect 25044 11704 25096 11756
rect 25228 11747 25280 11756
rect 25228 11713 25237 11747
rect 25237 11713 25271 11747
rect 25271 11713 25280 11747
rect 25228 11704 25280 11713
rect 26148 11704 26200 11756
rect 27344 11704 27396 11756
rect 28264 11747 28316 11756
rect 28264 11713 28273 11747
rect 28273 11713 28307 11747
rect 28307 11713 28316 11747
rect 28264 11704 28316 11713
rect 28540 11781 28557 11815
rect 28557 11781 28592 11815
rect 28540 11772 28592 11781
rect 28908 11772 28960 11824
rect 30932 11772 30984 11824
rect 31484 11840 31536 11892
rect 23848 11636 23900 11688
rect 25412 11636 25464 11688
rect 25504 11679 25556 11688
rect 25504 11645 25513 11679
rect 25513 11645 25547 11679
rect 25547 11645 25556 11679
rect 25504 11636 25556 11645
rect 27068 11636 27120 11688
rect 27160 11679 27212 11688
rect 27160 11645 27169 11679
rect 27169 11645 27203 11679
rect 27203 11645 27212 11679
rect 27160 11636 27212 11645
rect 27252 11679 27304 11688
rect 27252 11645 27261 11679
rect 27261 11645 27295 11679
rect 27295 11645 27304 11679
rect 27252 11636 27304 11645
rect 27528 11679 27580 11688
rect 27528 11645 27537 11679
rect 27537 11645 27571 11679
rect 27571 11645 27580 11679
rect 27528 11636 27580 11645
rect 27804 11636 27856 11688
rect 28816 11747 28868 11756
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 30288 11704 30340 11756
rect 30564 11704 30616 11756
rect 32036 11840 32088 11892
rect 33692 11840 33744 11892
rect 35256 11840 35308 11892
rect 31208 11704 31260 11756
rect 31760 11704 31812 11756
rect 34428 11772 34480 11824
rect 34888 11815 34940 11824
rect 34888 11781 34897 11815
rect 34897 11781 34931 11815
rect 34931 11781 34940 11815
rect 34888 11772 34940 11781
rect 29552 11636 29604 11688
rect 32404 11679 32456 11688
rect 32404 11645 32413 11679
rect 32413 11645 32447 11679
rect 32447 11645 32456 11679
rect 32404 11636 32456 11645
rect 33324 11747 33376 11756
rect 33324 11713 33341 11747
rect 33341 11713 33376 11747
rect 33324 11704 33376 11713
rect 33416 11747 33468 11756
rect 33416 11713 33425 11747
rect 33425 11713 33459 11747
rect 33459 11713 33468 11747
rect 33416 11704 33468 11713
rect 33508 11747 33560 11756
rect 33508 11713 33517 11747
rect 33517 11713 33551 11747
rect 33551 11713 33560 11747
rect 33508 11704 33560 11713
rect 33600 11747 33652 11756
rect 33600 11713 33609 11747
rect 33609 11713 33643 11747
rect 33643 11713 33652 11747
rect 33600 11704 33652 11713
rect 33692 11704 33744 11756
rect 33968 11747 34020 11756
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 33968 11704 34020 11713
rect 34612 11704 34664 11756
rect 16672 11500 16724 11552
rect 16948 11500 17000 11552
rect 18512 11500 18564 11552
rect 19340 11500 19392 11552
rect 20536 11500 20588 11552
rect 20720 11543 20772 11552
rect 20720 11509 20729 11543
rect 20729 11509 20763 11543
rect 20763 11509 20772 11543
rect 20720 11500 20772 11509
rect 25780 11568 25832 11620
rect 27620 11568 27672 11620
rect 29276 11568 29328 11620
rect 34336 11568 34388 11620
rect 34612 11568 34664 11620
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 22468 11500 22520 11552
rect 23848 11500 23900 11552
rect 24492 11500 24544 11552
rect 24584 11500 24636 11552
rect 28448 11500 28500 11552
rect 29184 11543 29236 11552
rect 29184 11509 29193 11543
rect 29193 11509 29227 11543
rect 29227 11509 29236 11543
rect 29184 11500 29236 11509
rect 32496 11543 32548 11552
rect 32496 11509 32505 11543
rect 32505 11509 32539 11543
rect 32539 11509 32548 11543
rect 32496 11500 32548 11509
rect 32680 11500 32732 11552
rect 33784 11543 33836 11552
rect 33784 11509 33793 11543
rect 33793 11509 33827 11543
rect 33827 11509 33836 11543
rect 33784 11500 33836 11509
rect 33876 11543 33928 11552
rect 33876 11509 33885 11543
rect 33885 11509 33919 11543
rect 33919 11509 33928 11543
rect 33876 11500 33928 11509
rect 33968 11500 34020 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 5356 11296 5408 11348
rect 5816 11339 5868 11348
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 5448 11228 5500 11280
rect 6276 11296 6328 11348
rect 6644 11228 6696 11280
rect 7656 11296 7708 11348
rect 11152 11296 11204 11348
rect 13452 11296 13504 11348
rect 17960 11296 18012 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18236 11296 18288 11348
rect 19064 11296 19116 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 6920 11160 6972 11212
rect 6092 11092 6144 11144
rect 4068 11024 4120 11076
rect 5632 11024 5684 11076
rect 6460 11092 6512 11144
rect 7472 11067 7524 11076
rect 7472 11033 7499 11067
rect 7499 11033 7524 11067
rect 7472 11024 7524 11033
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 9128 11228 9180 11280
rect 9404 11228 9456 11280
rect 13544 11228 13596 11280
rect 15476 11228 15528 11280
rect 15844 11228 15896 11280
rect 19892 11296 19944 11348
rect 19984 11296 20036 11348
rect 19708 11228 19760 11280
rect 20168 11228 20220 11280
rect 20352 11271 20404 11280
rect 20352 11237 20361 11271
rect 20361 11237 20395 11271
rect 20395 11237 20404 11271
rect 20352 11228 20404 11237
rect 10140 11160 10192 11212
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 9312 11092 9364 11144
rect 12256 11092 12308 11144
rect 13084 11160 13136 11212
rect 13452 11160 13504 11212
rect 7840 11024 7892 11076
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 9404 11024 9456 11076
rect 12900 11092 12952 11144
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 16212 11092 16264 11144
rect 16856 11160 16908 11212
rect 19340 11160 19392 11212
rect 20720 11296 20772 11348
rect 21272 11296 21324 11348
rect 21456 11339 21508 11348
rect 21456 11305 21465 11339
rect 21465 11305 21499 11339
rect 21499 11305 21508 11339
rect 21456 11296 21508 11305
rect 21548 11296 21600 11348
rect 22284 11296 22336 11348
rect 20812 11228 20864 11280
rect 21180 11228 21232 11280
rect 22008 11228 22060 11280
rect 22836 11296 22888 11348
rect 23020 11339 23072 11348
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 23664 11296 23716 11348
rect 24216 11296 24268 11348
rect 24860 11296 24912 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 23388 11228 23440 11280
rect 25412 11296 25464 11348
rect 27160 11296 27212 11348
rect 27896 11296 27948 11348
rect 28540 11296 28592 11348
rect 29000 11296 29052 11348
rect 29184 11296 29236 11348
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 16764 11092 16816 11144
rect 17040 11092 17092 11144
rect 5908 10956 5960 11008
rect 9680 10956 9732 11008
rect 10968 10956 11020 11008
rect 12624 10956 12676 11008
rect 15384 11024 15436 11076
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20536 11160 20588 11212
rect 19892 11135 19944 11144
rect 13268 10956 13320 11008
rect 14924 10956 14976 11008
rect 17776 10956 17828 11008
rect 17868 10999 17920 11008
rect 17868 10965 17877 10999
rect 17877 10965 17911 10999
rect 17911 10965 17920 10999
rect 17868 10956 17920 10965
rect 18788 11024 18840 11076
rect 19616 11024 19668 11076
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 20076 11092 20128 11144
rect 20628 11092 20680 11144
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 20904 11160 20956 11212
rect 22836 11160 22888 11212
rect 20904 11024 20956 11076
rect 21364 11092 21416 11144
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 22468 11135 22520 11144
rect 22468 11101 22477 11135
rect 22477 11101 22511 11135
rect 22511 11101 22520 11135
rect 22468 11092 22520 11101
rect 23572 11160 23624 11212
rect 25044 11160 25096 11212
rect 25596 11160 25648 11212
rect 21548 10956 21600 11008
rect 21640 10956 21692 11008
rect 22284 11024 22336 11076
rect 22744 11067 22796 11076
rect 22744 11033 22753 11067
rect 22753 11033 22787 11067
rect 22787 11033 22796 11067
rect 22744 11024 22796 11033
rect 22652 10956 22704 11008
rect 22928 11024 22980 11076
rect 24492 11135 24544 11144
rect 24492 11101 24501 11135
rect 24501 11101 24535 11135
rect 24535 11101 24544 11135
rect 24492 11092 24544 11101
rect 25872 11228 25924 11280
rect 23572 11024 23624 11076
rect 24584 11024 24636 11076
rect 25596 11024 25648 11076
rect 23112 10956 23164 11008
rect 23848 10956 23900 11008
rect 25228 10956 25280 11008
rect 26884 11135 26936 11144
rect 26884 11101 26893 11135
rect 26893 11101 26927 11135
rect 26927 11101 26936 11135
rect 26884 11092 26936 11101
rect 28080 11135 28132 11144
rect 28080 11101 28089 11135
rect 28089 11101 28123 11135
rect 28123 11101 28132 11135
rect 28080 11092 28132 11101
rect 28172 11135 28224 11144
rect 28172 11101 28181 11135
rect 28181 11101 28215 11135
rect 28215 11101 28224 11135
rect 28172 11092 28224 11101
rect 28356 11135 28408 11144
rect 28356 11101 28365 11135
rect 28365 11101 28399 11135
rect 28399 11101 28408 11135
rect 28356 11092 28408 11101
rect 28448 11135 28500 11144
rect 28448 11101 28457 11135
rect 28457 11101 28491 11135
rect 28491 11101 28500 11135
rect 28448 11092 28500 11101
rect 28816 11228 28868 11280
rect 28632 11092 28684 11144
rect 29000 11135 29052 11144
rect 29000 11101 29009 11135
rect 29009 11101 29043 11135
rect 29043 11101 29052 11135
rect 29000 11092 29052 11101
rect 30380 11339 30432 11348
rect 30380 11305 30389 11339
rect 30389 11305 30423 11339
rect 30423 11305 30432 11339
rect 30380 11296 30432 11305
rect 33692 11296 33744 11348
rect 33784 11339 33836 11348
rect 33784 11305 33793 11339
rect 33793 11305 33827 11339
rect 33827 11305 33836 11339
rect 33784 11296 33836 11305
rect 29184 11135 29236 11144
rect 29184 11101 29193 11135
rect 29193 11101 29227 11135
rect 29227 11101 29236 11135
rect 29184 11092 29236 11101
rect 30380 11160 30432 11212
rect 30564 11135 30616 11144
rect 30564 11101 30573 11135
rect 30573 11101 30607 11135
rect 30607 11101 30616 11135
rect 30564 11092 30616 11101
rect 34336 11228 34388 11280
rect 34612 11160 34664 11212
rect 32680 11135 32732 11144
rect 32680 11101 32689 11135
rect 32689 11101 32723 11135
rect 32723 11101 32732 11135
rect 32680 11092 32732 11101
rect 33692 11135 33744 11144
rect 33692 11101 33701 11135
rect 33701 11101 33735 11135
rect 33735 11101 33744 11135
rect 33692 11092 33744 11101
rect 34796 11092 34848 11144
rect 28448 10956 28500 11008
rect 28632 10956 28684 11008
rect 30656 11024 30708 11076
rect 32404 11024 32456 11076
rect 32956 11024 33008 11076
rect 29184 10956 29236 11008
rect 30104 10956 30156 11008
rect 30840 10956 30892 11008
rect 33232 10956 33284 11008
rect 33508 10956 33560 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 4804 10752 4856 10804
rect 6000 10752 6052 10804
rect 5908 10727 5960 10736
rect 5908 10693 5917 10727
rect 5917 10693 5951 10727
rect 5951 10693 5960 10727
rect 5908 10684 5960 10693
rect 7012 10752 7064 10804
rect 8208 10752 8260 10804
rect 11520 10752 11572 10804
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 6920 10548 6972 10600
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 8024 10480 8076 10532
rect 7196 10412 7248 10464
rect 7380 10412 7432 10464
rect 7656 10412 7708 10464
rect 8484 10548 8536 10600
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 10140 10616 10192 10668
rect 10232 10659 10284 10668
rect 10232 10625 10241 10659
rect 10241 10625 10275 10659
rect 10275 10625 10284 10659
rect 10232 10616 10284 10625
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 11336 10684 11388 10736
rect 11152 10616 11204 10668
rect 11704 10616 11756 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 11704 10480 11756 10532
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13452 10659 13504 10668
rect 13452 10625 13461 10659
rect 13461 10625 13495 10659
rect 13495 10625 13504 10659
rect 13452 10616 13504 10625
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 13360 10480 13412 10532
rect 14188 10548 14240 10600
rect 14648 10480 14700 10532
rect 18512 10752 18564 10804
rect 19432 10752 19484 10804
rect 16580 10684 16632 10736
rect 17868 10684 17920 10736
rect 17960 10684 18012 10736
rect 25596 10752 25648 10804
rect 21364 10684 21416 10736
rect 21548 10684 21600 10736
rect 23848 10727 23900 10736
rect 23848 10693 23857 10727
rect 23857 10693 23891 10727
rect 23891 10693 23900 10727
rect 23848 10684 23900 10693
rect 24492 10684 24544 10736
rect 27344 10752 27396 10804
rect 27804 10752 27856 10804
rect 28540 10752 28592 10804
rect 17316 10616 17368 10668
rect 19432 10616 19484 10668
rect 16212 10548 16264 10600
rect 18696 10548 18748 10600
rect 19984 10659 20036 10668
rect 19984 10625 19993 10659
rect 19993 10625 20027 10659
rect 20027 10625 20036 10659
rect 19984 10616 20036 10625
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 22008 10616 22060 10668
rect 23572 10659 23624 10668
rect 23572 10625 23581 10659
rect 23581 10625 23615 10659
rect 23615 10625 23624 10659
rect 23572 10616 23624 10625
rect 23664 10616 23716 10668
rect 22468 10548 22520 10600
rect 22928 10548 22980 10600
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 24768 10616 24820 10668
rect 25228 10659 25280 10668
rect 25228 10625 25237 10659
rect 25237 10625 25271 10659
rect 25271 10625 25280 10659
rect 25228 10616 25280 10625
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 25596 10616 25648 10668
rect 27252 10684 27304 10736
rect 28172 10684 28224 10736
rect 25320 10548 25372 10600
rect 26148 10616 26200 10668
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 26424 10616 26476 10668
rect 26700 10659 26752 10668
rect 26700 10625 26709 10659
rect 26709 10625 26743 10659
rect 26743 10625 26752 10659
rect 26700 10616 26752 10625
rect 27068 10616 27120 10668
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 27988 10616 28040 10668
rect 27344 10548 27396 10600
rect 27896 10548 27948 10600
rect 28540 10659 28592 10668
rect 28540 10625 28549 10659
rect 28549 10625 28583 10659
rect 28583 10625 28592 10659
rect 28540 10616 28592 10625
rect 28724 10684 28776 10736
rect 29184 10752 29236 10804
rect 29276 10795 29328 10804
rect 29276 10761 29285 10795
rect 29285 10761 29319 10795
rect 29319 10761 29328 10795
rect 29276 10752 29328 10761
rect 33140 10752 33192 10804
rect 34704 10752 34756 10804
rect 28724 10548 28776 10600
rect 29736 10616 29788 10668
rect 29920 10616 29972 10668
rect 31300 10684 31352 10736
rect 34336 10727 34388 10736
rect 34336 10693 34345 10727
rect 34345 10693 34379 10727
rect 34379 10693 34388 10727
rect 34336 10684 34388 10693
rect 34796 10684 34848 10736
rect 31024 10616 31076 10668
rect 33692 10616 33744 10668
rect 34612 10616 34664 10668
rect 21456 10480 21508 10532
rect 25412 10480 25464 10532
rect 26240 10480 26292 10532
rect 27804 10480 27856 10532
rect 28080 10480 28132 10532
rect 8300 10412 8352 10464
rect 9680 10412 9732 10464
rect 9772 10412 9824 10464
rect 12348 10412 12400 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 16764 10412 16816 10464
rect 17224 10412 17276 10464
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 22192 10412 22244 10464
rect 23940 10412 23992 10464
rect 24400 10412 24452 10464
rect 24584 10412 24636 10464
rect 27160 10412 27212 10464
rect 27344 10412 27396 10464
rect 28172 10412 28224 10464
rect 28356 10480 28408 10532
rect 30656 10548 30708 10600
rect 30288 10480 30340 10532
rect 35440 10659 35492 10668
rect 35440 10625 35449 10659
rect 35449 10625 35483 10659
rect 35483 10625 35492 10659
rect 35440 10616 35492 10625
rect 32312 10455 32364 10464
rect 32312 10421 32321 10455
rect 32321 10421 32355 10455
rect 32355 10421 32364 10455
rect 32312 10412 32364 10421
rect 36176 10412 36228 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6276 10251 6328 10260
rect 6276 10217 6285 10251
rect 6285 10217 6319 10251
rect 6319 10217 6328 10251
rect 6276 10208 6328 10217
rect 6552 10208 6604 10260
rect 6920 10208 6972 10260
rect 7932 10208 7984 10260
rect 8760 10208 8812 10260
rect 9956 10208 10008 10260
rect 10692 10208 10744 10260
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 16212 10208 16264 10260
rect 16580 10251 16632 10260
rect 16580 10217 16589 10251
rect 16589 10217 16623 10251
rect 16623 10217 16632 10251
rect 16580 10208 16632 10217
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 17776 10208 17828 10260
rect 20168 10208 20220 10260
rect 20720 10208 20772 10260
rect 21916 10208 21968 10260
rect 22192 10251 22244 10260
rect 22192 10217 22201 10251
rect 22201 10217 22235 10251
rect 22235 10217 22244 10251
rect 22192 10208 22244 10217
rect 22836 10208 22888 10260
rect 25412 10208 25464 10260
rect 6092 10140 6144 10192
rect 2872 10072 2924 10124
rect 4068 10072 4120 10124
rect 4620 10072 4672 10124
rect 9772 10140 9824 10192
rect 7012 10072 7064 10124
rect 7104 10072 7156 10124
rect 5724 10004 5776 10056
rect 5908 10047 5960 10056
rect 5908 10013 5914 10047
rect 5914 10013 5948 10047
rect 5948 10013 5960 10047
rect 5908 10004 5960 10013
rect 6828 10004 6880 10056
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 8668 10115 8720 10124
rect 8668 10081 8677 10115
rect 8677 10081 8711 10115
rect 8711 10081 8720 10115
rect 8668 10072 8720 10081
rect 9404 10072 9456 10124
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 8392 10004 8444 10056
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 9128 9979 9180 9988
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6000 9868 6052 9920
rect 7472 9911 7524 9920
rect 7472 9877 7481 9911
rect 7481 9877 7515 9911
rect 7515 9877 7524 9911
rect 7472 9868 7524 9877
rect 9128 9945 9137 9979
rect 9137 9945 9171 9979
rect 9171 9945 9180 9979
rect 9128 9936 9180 9945
rect 9588 10004 9640 10056
rect 10324 10140 10376 10192
rect 10232 10072 10284 10124
rect 9956 10004 10008 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 16396 10183 16448 10192
rect 16396 10149 16405 10183
rect 16405 10149 16439 10183
rect 16439 10149 16448 10183
rect 16396 10140 16448 10149
rect 13268 10072 13320 10124
rect 13912 10072 13964 10124
rect 10968 10004 11020 10056
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11244 10004 11296 10056
rect 11520 10004 11572 10056
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 16488 10115 16540 10124
rect 16488 10081 16497 10115
rect 16497 10081 16531 10115
rect 16531 10081 16540 10115
rect 16488 10072 16540 10081
rect 16672 10072 16724 10124
rect 14832 10004 14884 10056
rect 13544 9936 13596 9988
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 17224 10072 17276 10124
rect 18420 10072 18472 10124
rect 18696 10140 18748 10192
rect 18880 10183 18932 10192
rect 18880 10149 18889 10183
rect 18889 10149 18923 10183
rect 18923 10149 18932 10183
rect 18880 10140 18932 10149
rect 19616 10140 19668 10192
rect 19708 10072 19760 10124
rect 22928 10072 22980 10124
rect 25688 10072 25740 10124
rect 26240 10072 26292 10124
rect 27896 10140 27948 10192
rect 28724 10183 28776 10192
rect 28724 10149 28733 10183
rect 28733 10149 28767 10183
rect 28767 10149 28776 10183
rect 28724 10140 28776 10149
rect 29460 10208 29512 10260
rect 31024 10251 31076 10260
rect 31024 10217 31033 10251
rect 31033 10217 31067 10251
rect 31067 10217 31076 10251
rect 31024 10208 31076 10217
rect 31208 10140 31260 10192
rect 26424 10115 26476 10124
rect 26424 10081 26433 10115
rect 26433 10081 26467 10115
rect 26467 10081 26476 10115
rect 26424 10072 26476 10081
rect 26700 10072 26752 10124
rect 28356 10072 28408 10124
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17960 9936 18012 9988
rect 18144 9936 18196 9988
rect 19432 10004 19484 10056
rect 19984 10004 20036 10056
rect 19340 9936 19392 9988
rect 19892 9936 19944 9988
rect 20260 10047 20312 10056
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 12900 9868 12952 9920
rect 13360 9868 13412 9920
rect 13820 9868 13872 9920
rect 14740 9868 14792 9920
rect 14924 9868 14976 9920
rect 19708 9868 19760 9920
rect 20168 9936 20220 9988
rect 20628 10004 20680 10056
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 21272 9979 21324 9988
rect 21272 9945 21281 9979
rect 21281 9945 21315 9979
rect 21315 9945 21324 9979
rect 21272 9936 21324 9945
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 23940 10004 23992 10056
rect 22928 9936 22980 9988
rect 24308 9936 24360 9988
rect 25228 10004 25280 10056
rect 25596 9936 25648 9988
rect 26056 9936 26108 9988
rect 21364 9868 21416 9920
rect 21824 9868 21876 9920
rect 26516 9936 26568 9988
rect 27068 9868 27120 9920
rect 27344 10004 27396 10056
rect 27896 10047 27948 10056
rect 27896 10013 27905 10047
rect 27905 10013 27939 10047
rect 27939 10013 27948 10047
rect 27896 10004 27948 10013
rect 28172 10004 28224 10056
rect 28080 9936 28132 9988
rect 28908 10013 28929 10034
rect 28929 10013 28960 10034
rect 28908 9982 28960 10013
rect 29184 10004 29236 10056
rect 29552 10004 29604 10056
rect 29828 10047 29880 10056
rect 29828 10013 29845 10047
rect 29845 10013 29880 10047
rect 29828 10004 29880 10013
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 30196 10004 30248 10056
rect 30748 10047 30800 10056
rect 30748 10013 30757 10047
rect 30757 10013 30791 10047
rect 30791 10013 30800 10047
rect 30748 10004 30800 10013
rect 31208 10047 31260 10056
rect 29920 9979 29972 9988
rect 29920 9945 29929 9979
rect 29929 9945 29963 9979
rect 29963 9945 29972 9979
rect 29920 9936 29972 9945
rect 31208 10013 31212 10047
rect 31212 10013 31246 10047
rect 31246 10013 31260 10047
rect 31208 10004 31260 10013
rect 31392 10072 31444 10124
rect 31668 10047 31720 10056
rect 31668 10013 31677 10047
rect 31677 10013 31711 10047
rect 31711 10013 31720 10047
rect 31668 10004 31720 10013
rect 29736 9868 29788 9920
rect 29828 9868 29880 9920
rect 30932 9936 30984 9988
rect 34336 9936 34388 9988
rect 30196 9868 30248 9920
rect 30380 9868 30432 9920
rect 31116 9868 31168 9920
rect 31484 9868 31536 9920
rect 36268 9868 36320 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 10600 9664 10652 9716
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 6184 9596 6236 9648
rect 5816 9528 5868 9580
rect 6000 9528 6052 9580
rect 4068 9460 4120 9512
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7104 9571 7156 9580
rect 7104 9537 7112 9571
rect 7112 9537 7146 9571
rect 7146 9537 7156 9571
rect 7104 9528 7156 9537
rect 7472 9528 7524 9580
rect 11060 9596 11112 9648
rect 14188 9596 14240 9648
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 6184 9435 6236 9444
rect 6184 9401 6193 9435
rect 6193 9401 6227 9435
rect 6227 9401 6236 9435
rect 6184 9392 6236 9401
rect 8944 9460 8996 9512
rect 10324 9460 10376 9512
rect 11152 9528 11204 9580
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 12532 9528 12584 9580
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 14924 9596 14976 9648
rect 16028 9664 16080 9716
rect 17960 9664 18012 9716
rect 18144 9664 18196 9716
rect 18236 9664 18288 9716
rect 18696 9664 18748 9716
rect 11336 9460 11388 9512
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 12624 9392 12676 9444
rect 14740 9571 14792 9580
rect 14740 9537 14749 9571
rect 14749 9537 14783 9571
rect 14783 9537 14792 9571
rect 14740 9528 14792 9537
rect 17316 9596 17368 9648
rect 24584 9664 24636 9716
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16396 9528 16448 9580
rect 15108 9460 15160 9512
rect 15660 9503 15712 9512
rect 15660 9469 15669 9503
rect 15669 9469 15703 9503
rect 15703 9469 15712 9503
rect 15660 9460 15712 9469
rect 17040 9460 17092 9512
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 18512 9528 18564 9580
rect 18696 9528 18748 9580
rect 18972 9528 19024 9580
rect 19432 9528 19484 9580
rect 19616 9571 19668 9580
rect 19616 9537 19625 9571
rect 19625 9537 19659 9571
rect 19659 9537 19668 9571
rect 19616 9528 19668 9537
rect 21272 9596 21324 9648
rect 20628 9528 20680 9580
rect 19800 9460 19852 9512
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 22928 9571 22980 9580
rect 22928 9537 22937 9571
rect 22937 9537 22971 9571
rect 22971 9537 22980 9571
rect 22928 9528 22980 9537
rect 23204 9528 23256 9580
rect 23848 9596 23900 9648
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 24584 9571 24636 9580
rect 24584 9537 24593 9571
rect 24593 9537 24627 9571
rect 24627 9537 24636 9571
rect 24584 9528 24636 9537
rect 25504 9528 25556 9580
rect 26056 9571 26108 9580
rect 26056 9537 26065 9571
rect 26065 9537 26099 9571
rect 26099 9537 26108 9571
rect 26056 9528 26108 9537
rect 26976 9596 27028 9648
rect 26700 9528 26752 9580
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 28540 9664 28592 9716
rect 28724 9596 28776 9648
rect 29460 9596 29512 9648
rect 29552 9596 29604 9648
rect 32036 9664 32088 9716
rect 33692 9664 33744 9716
rect 34336 9664 34388 9716
rect 34796 9664 34848 9716
rect 30380 9596 30432 9648
rect 16764 9392 16816 9444
rect 18880 9392 18932 9444
rect 15292 9324 15344 9376
rect 17500 9324 17552 9376
rect 18144 9324 18196 9376
rect 18604 9324 18656 9376
rect 19064 9324 19116 9376
rect 22560 9392 22612 9444
rect 23020 9392 23072 9444
rect 23572 9435 23624 9444
rect 23572 9401 23581 9435
rect 23581 9401 23615 9435
rect 23615 9401 23624 9435
rect 23572 9392 23624 9401
rect 25044 9460 25096 9512
rect 25136 9460 25188 9512
rect 25964 9460 26016 9512
rect 22468 9324 22520 9376
rect 22836 9324 22888 9376
rect 23388 9324 23440 9376
rect 25412 9324 25464 9376
rect 25872 9392 25924 9444
rect 27436 9460 27488 9512
rect 29276 9528 29328 9580
rect 29828 9528 29880 9580
rect 30012 9528 30064 9580
rect 32864 9571 32916 9580
rect 32864 9537 32873 9571
rect 32873 9537 32907 9571
rect 32907 9537 32916 9571
rect 32864 9528 32916 9537
rect 33048 9571 33100 9580
rect 33048 9537 33065 9571
rect 33065 9537 33100 9571
rect 33048 9528 33100 9537
rect 33140 9571 33192 9580
rect 33140 9537 33149 9571
rect 33149 9537 33183 9571
rect 33183 9537 33192 9571
rect 33140 9528 33192 9537
rect 33232 9571 33284 9580
rect 33232 9537 33241 9571
rect 33241 9537 33275 9571
rect 33275 9537 33284 9571
rect 33232 9528 33284 9537
rect 33324 9571 33376 9580
rect 33324 9537 33333 9571
rect 33333 9537 33367 9571
rect 33367 9537 33376 9571
rect 33324 9528 33376 9537
rect 33508 9528 33560 9580
rect 33600 9571 33652 9580
rect 33600 9537 33609 9571
rect 33609 9537 33643 9571
rect 33643 9537 33652 9571
rect 33600 9528 33652 9537
rect 34336 9571 34388 9580
rect 34336 9537 34346 9571
rect 34346 9537 34380 9571
rect 34380 9537 34388 9571
rect 34336 9528 34388 9537
rect 27804 9460 27856 9512
rect 28448 9460 28500 9512
rect 28908 9460 28960 9512
rect 26332 9435 26384 9444
rect 26332 9401 26341 9435
rect 26341 9401 26375 9435
rect 26375 9401 26384 9435
rect 26332 9392 26384 9401
rect 27712 9392 27764 9444
rect 33232 9392 33284 9444
rect 28724 9324 28776 9376
rect 28908 9324 28960 9376
rect 29920 9324 29972 9376
rect 30104 9324 30156 9376
rect 33324 9324 33376 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 5908 9120 5960 9172
rect 6920 9120 6972 9172
rect 7104 9120 7156 9172
rect 5816 8984 5868 9036
rect 15200 9120 15252 9172
rect 16120 9120 16172 9172
rect 17408 9120 17460 9172
rect 18604 9163 18656 9172
rect 18604 9129 18613 9163
rect 18613 9129 18647 9163
rect 18647 9129 18656 9163
rect 18604 9120 18656 9129
rect 19340 9120 19392 9172
rect 21364 9120 21416 9172
rect 21456 9163 21508 9172
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 22008 9120 22060 9172
rect 22652 9163 22704 9172
rect 22652 9129 22661 9163
rect 22661 9129 22695 9163
rect 22695 9129 22704 9163
rect 22652 9120 22704 9129
rect 22744 9120 22796 9172
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 25044 9163 25096 9172
rect 25044 9129 25053 9163
rect 25053 9129 25087 9163
rect 25087 9129 25096 9163
rect 25044 9120 25096 9129
rect 25964 9120 26016 9172
rect 8300 9052 8352 9104
rect 4068 8916 4120 8968
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 6828 8916 6880 8968
rect 4804 8891 4856 8900
rect 4804 8857 4813 8891
rect 4813 8857 4847 8891
rect 4847 8857 4856 8891
rect 4804 8848 4856 8857
rect 6644 8780 6696 8832
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 9036 8916 9088 8968
rect 17500 9095 17552 9104
rect 17500 9061 17509 9095
rect 17509 9061 17543 9095
rect 17543 9061 17552 9095
rect 17500 9052 17552 9061
rect 17868 9052 17920 9104
rect 20536 9052 20588 9104
rect 22560 9052 22612 9104
rect 25596 9052 25648 9104
rect 26240 9052 26292 9104
rect 26792 9095 26844 9104
rect 26792 9061 26801 9095
rect 26801 9061 26835 9095
rect 26835 9061 26844 9095
rect 26792 9052 26844 9061
rect 26976 9095 27028 9104
rect 26976 9061 26985 9095
rect 26985 9061 27019 9095
rect 27019 9061 27028 9095
rect 26976 9052 27028 9061
rect 10048 8984 10100 9036
rect 12716 8984 12768 9036
rect 18972 8984 19024 9036
rect 20628 8984 20680 9036
rect 25688 9027 25740 9036
rect 25688 8993 25697 9027
rect 25697 8993 25731 9027
rect 25731 8993 25740 9027
rect 25688 8984 25740 8993
rect 26700 8984 26752 9036
rect 9864 8916 9916 8968
rect 11060 8916 11112 8968
rect 11520 8916 11572 8968
rect 7380 8848 7432 8900
rect 8116 8848 8168 8900
rect 8392 8848 8444 8900
rect 8668 8780 8720 8832
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 15936 8916 15988 8968
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 17592 8916 17644 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 18328 8916 18380 8968
rect 18420 8959 18472 8968
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 18604 8916 18656 8968
rect 19432 8916 19484 8968
rect 19984 8916 20036 8968
rect 20260 8916 20312 8968
rect 21456 8916 21508 8968
rect 21548 8959 21600 8968
rect 21548 8925 21557 8959
rect 21557 8925 21591 8959
rect 21591 8925 21600 8959
rect 21548 8916 21600 8925
rect 23112 8916 23164 8968
rect 24676 8959 24728 8968
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24676 8916 24728 8925
rect 12072 8891 12124 8900
rect 12072 8857 12081 8891
rect 12081 8857 12115 8891
rect 12115 8857 12124 8891
rect 12072 8848 12124 8857
rect 14832 8848 14884 8900
rect 16212 8848 16264 8900
rect 10416 8780 10468 8832
rect 10876 8780 10928 8832
rect 13360 8780 13412 8832
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 17040 8780 17092 8832
rect 17316 8848 17368 8900
rect 18512 8848 18564 8900
rect 18788 8848 18840 8900
rect 19064 8891 19116 8900
rect 19064 8857 19073 8891
rect 19073 8857 19107 8891
rect 19107 8857 19116 8891
rect 19064 8848 19116 8857
rect 22836 8891 22888 8900
rect 22836 8857 22863 8891
rect 22863 8857 22888 8891
rect 22836 8848 22888 8857
rect 21272 8780 21324 8832
rect 21916 8780 21968 8832
rect 22928 8780 22980 8832
rect 23940 8848 23992 8900
rect 24584 8780 24636 8832
rect 26240 8916 26292 8968
rect 27988 8984 28040 9036
rect 26516 8848 26568 8900
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 28172 8916 28224 8968
rect 28356 8916 28408 8968
rect 29368 9052 29420 9104
rect 29736 9052 29788 9104
rect 29184 8984 29236 9036
rect 27804 8848 27856 8900
rect 28816 8848 28868 8900
rect 29552 8959 29604 8968
rect 29552 8925 29561 8959
rect 29561 8925 29595 8959
rect 29595 8925 29604 8959
rect 29552 8916 29604 8925
rect 29644 8916 29696 8968
rect 28632 8780 28684 8832
rect 29000 8780 29052 8832
rect 30196 8848 30248 8900
rect 29920 8780 29972 8832
rect 31576 9120 31628 9172
rect 32680 9120 32732 9172
rect 33600 9120 33652 9172
rect 31392 8984 31444 9036
rect 32496 8984 32548 9036
rect 31208 8916 31260 8968
rect 31668 8959 31720 8968
rect 31668 8925 31677 8959
rect 31677 8925 31711 8959
rect 31711 8925 31720 8959
rect 31668 8916 31720 8925
rect 33140 8916 33192 8968
rect 33876 9052 33928 9104
rect 35992 8916 36044 8968
rect 32864 8848 32916 8900
rect 32496 8780 32548 8832
rect 32680 8780 32732 8832
rect 33048 8823 33100 8832
rect 33048 8789 33057 8823
rect 33057 8789 33091 8823
rect 33091 8789 33100 8823
rect 33048 8780 33100 8789
rect 33508 8891 33560 8900
rect 33508 8857 33517 8891
rect 33517 8857 33551 8891
rect 33551 8857 33560 8891
rect 33508 8848 33560 8857
rect 34980 8780 35032 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 4804 8576 4856 8628
rect 9036 8619 9088 8628
rect 9036 8585 9045 8619
rect 9045 8585 9079 8619
rect 9079 8585 9088 8619
rect 9036 8576 9088 8585
rect 12072 8576 12124 8628
rect 9128 8508 9180 8560
rect 6736 8440 6788 8492
rect 7104 8440 7156 8492
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 10508 8508 10560 8560
rect 12808 8508 12860 8560
rect 5724 8372 5776 8424
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 7196 8372 7248 8424
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 11336 8440 11388 8492
rect 15200 8576 15252 8628
rect 13360 8551 13412 8560
rect 13360 8517 13369 8551
rect 13369 8517 13403 8551
rect 13403 8517 13412 8551
rect 13360 8508 13412 8517
rect 14464 8440 14516 8492
rect 14648 8440 14700 8492
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 17684 8576 17736 8628
rect 18696 8619 18748 8628
rect 18696 8585 18705 8619
rect 18705 8585 18739 8619
rect 18739 8585 18748 8619
rect 18696 8576 18748 8585
rect 19432 8576 19484 8628
rect 21180 8576 21232 8628
rect 21640 8576 21692 8628
rect 7288 8236 7340 8288
rect 9312 8304 9364 8356
rect 10876 8415 10928 8424
rect 10876 8381 10885 8415
rect 10885 8381 10919 8415
rect 10919 8381 10928 8415
rect 10876 8372 10928 8381
rect 11520 8372 11572 8424
rect 10140 8347 10192 8356
rect 10140 8313 10149 8347
rect 10149 8313 10183 8347
rect 10183 8313 10192 8347
rect 10140 8304 10192 8313
rect 10232 8347 10284 8356
rect 10232 8313 10241 8347
rect 10241 8313 10275 8347
rect 10275 8313 10284 8347
rect 10232 8304 10284 8313
rect 14740 8372 14792 8424
rect 14832 8415 14884 8424
rect 14832 8381 14841 8415
rect 14841 8381 14875 8415
rect 14875 8381 14884 8415
rect 14832 8372 14884 8381
rect 14924 8372 14976 8424
rect 17500 8440 17552 8492
rect 18420 8508 18472 8560
rect 19156 8508 19208 8560
rect 18052 8440 18104 8492
rect 18328 8483 18380 8492
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 18328 8440 18380 8449
rect 18604 8440 18656 8492
rect 17960 8372 18012 8424
rect 10692 8279 10744 8288
rect 10692 8245 10701 8279
rect 10701 8245 10735 8279
rect 10735 8245 10744 8279
rect 10692 8236 10744 8245
rect 13912 8236 13964 8288
rect 17408 8304 17460 8356
rect 17500 8347 17552 8356
rect 17500 8313 17509 8347
rect 17509 8313 17543 8347
rect 17543 8313 17552 8347
rect 17500 8304 17552 8313
rect 14740 8236 14792 8288
rect 15108 8236 15160 8288
rect 16028 8236 16080 8288
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 17684 8304 17736 8356
rect 19340 8483 19392 8492
rect 19340 8449 19349 8483
rect 19349 8449 19383 8483
rect 19383 8449 19392 8483
rect 19340 8440 19392 8449
rect 19524 8508 19576 8560
rect 20444 8440 20496 8492
rect 20720 8508 20772 8560
rect 21456 8508 21508 8560
rect 22560 8576 22612 8628
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 20628 8440 20680 8492
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 23848 8508 23900 8560
rect 20720 8372 20772 8424
rect 21548 8372 21600 8424
rect 22008 8372 22060 8424
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 24400 8576 24452 8628
rect 24676 8576 24728 8628
rect 27252 8576 27304 8628
rect 28540 8576 28592 8628
rect 28632 8576 28684 8628
rect 25504 8508 25556 8560
rect 30472 8576 30524 8628
rect 31208 8576 31260 8628
rect 31760 8576 31812 8628
rect 24400 8440 24452 8492
rect 24584 8483 24636 8492
rect 24584 8449 24593 8483
rect 24593 8449 24627 8483
rect 24627 8449 24636 8483
rect 24584 8440 24636 8449
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 24768 8440 24820 8492
rect 25872 8440 25924 8492
rect 24124 8372 24176 8424
rect 26792 8440 26844 8492
rect 26976 8440 27028 8492
rect 26240 8372 26292 8424
rect 26700 8415 26752 8424
rect 26700 8381 26709 8415
rect 26709 8381 26743 8415
rect 26743 8381 26752 8415
rect 26700 8372 26752 8381
rect 28632 8440 28684 8492
rect 28816 8440 28868 8492
rect 29828 8508 29880 8560
rect 30288 8551 30340 8560
rect 30288 8517 30297 8551
rect 30297 8517 30331 8551
rect 30331 8517 30340 8551
rect 30288 8508 30340 8517
rect 30104 8440 30156 8492
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30932 8483 30984 8492
rect 30196 8440 30248 8449
rect 30932 8449 30941 8483
rect 30941 8449 30975 8483
rect 30975 8449 30984 8483
rect 30932 8440 30984 8449
rect 33416 8576 33468 8628
rect 33876 8576 33928 8628
rect 34980 8619 35032 8628
rect 34980 8585 34989 8619
rect 34989 8585 35023 8619
rect 35023 8585 35032 8619
rect 34980 8576 35032 8585
rect 34520 8508 34572 8560
rect 28540 8372 28592 8424
rect 28908 8372 28960 8424
rect 29092 8372 29144 8424
rect 29828 8415 29880 8424
rect 29828 8381 29837 8415
rect 29837 8381 29871 8415
rect 29871 8381 29880 8415
rect 29828 8372 29880 8381
rect 31392 8440 31444 8492
rect 19524 8304 19576 8356
rect 20536 8304 20588 8356
rect 20904 8304 20956 8356
rect 19616 8236 19668 8288
rect 20076 8236 20128 8288
rect 22008 8279 22060 8288
rect 22008 8245 22017 8279
rect 22017 8245 22051 8279
rect 22051 8245 22060 8279
rect 22008 8236 22060 8245
rect 24400 8347 24452 8356
rect 24400 8313 24409 8347
rect 24409 8313 24443 8347
rect 24443 8313 24452 8347
rect 24400 8304 24452 8313
rect 25504 8304 25556 8356
rect 27712 8304 27764 8356
rect 31208 8304 31260 8356
rect 31484 8415 31536 8424
rect 31484 8381 31493 8415
rect 31493 8381 31527 8415
rect 31527 8381 31536 8415
rect 31484 8372 31536 8381
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 33508 8440 33560 8492
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 34796 8483 34848 8492
rect 34796 8449 34805 8483
rect 34805 8449 34839 8483
rect 34839 8449 34848 8483
rect 34796 8440 34848 8449
rect 31576 8304 31628 8356
rect 26516 8236 26568 8288
rect 27988 8236 28040 8288
rect 28540 8279 28592 8288
rect 28540 8245 28549 8279
rect 28549 8245 28583 8279
rect 28583 8245 28592 8279
rect 28540 8236 28592 8245
rect 28632 8279 28684 8288
rect 28632 8245 28641 8279
rect 28641 8245 28675 8279
rect 28675 8245 28684 8279
rect 28632 8236 28684 8245
rect 31024 8236 31076 8288
rect 32864 8347 32916 8356
rect 32864 8313 32873 8347
rect 32873 8313 32907 8347
rect 32907 8313 32916 8347
rect 32864 8304 32916 8313
rect 33048 8304 33100 8356
rect 34244 8304 34296 8356
rect 33508 8236 33560 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 8484 8032 8536 8084
rect 9496 8032 9548 8084
rect 9404 7964 9456 8016
rect 9864 8032 9916 8084
rect 10140 8032 10192 8084
rect 10232 8032 10284 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 6920 7760 6972 7812
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 9128 7828 9180 7880
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 10324 7828 10376 7880
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 13636 8032 13688 8084
rect 14740 8032 14792 8084
rect 16856 8032 16908 8084
rect 17316 8075 17368 8084
rect 17316 8041 17325 8075
rect 17325 8041 17359 8075
rect 17359 8041 17368 8075
rect 17316 8032 17368 8041
rect 11520 7828 11572 7880
rect 19064 8032 19116 8084
rect 19432 8032 19484 8084
rect 20996 8075 21048 8084
rect 20996 8041 21005 8075
rect 21005 8041 21039 8075
rect 21039 8041 21048 8075
rect 20996 8032 21048 8041
rect 21548 8032 21600 8084
rect 16028 7939 16080 7948
rect 16028 7905 16037 7939
rect 16037 7905 16071 7939
rect 16071 7905 16080 7939
rect 16028 7896 16080 7905
rect 11980 7803 12032 7812
rect 11980 7769 11989 7803
rect 11989 7769 12023 7803
rect 12023 7769 12032 7803
rect 11980 7760 12032 7769
rect 14464 7760 14516 7812
rect 15108 7871 15160 7880
rect 15108 7837 15122 7871
rect 15122 7837 15156 7871
rect 15156 7837 15160 7871
rect 15108 7828 15160 7837
rect 15292 7828 15344 7880
rect 16580 7828 16632 7880
rect 17132 7828 17184 7880
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 14832 7760 14884 7812
rect 14924 7803 14976 7812
rect 14924 7769 14933 7803
rect 14933 7769 14967 7803
rect 14967 7769 14976 7803
rect 14924 7760 14976 7769
rect 8208 7692 8260 7744
rect 10968 7692 11020 7744
rect 11520 7692 11572 7744
rect 11796 7692 11848 7744
rect 11888 7692 11940 7744
rect 14556 7692 14608 7744
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 15752 7735 15804 7744
rect 15752 7701 15761 7735
rect 15761 7701 15795 7735
rect 15795 7701 15804 7735
rect 15752 7692 15804 7701
rect 16580 7735 16632 7744
rect 16580 7701 16589 7735
rect 16589 7701 16623 7735
rect 16623 7701 16632 7735
rect 16580 7692 16632 7701
rect 16948 7760 17000 7812
rect 19340 7896 19392 7948
rect 24032 8032 24084 8084
rect 26792 8075 26844 8084
rect 26792 8041 26801 8075
rect 26801 8041 26835 8075
rect 26835 8041 26844 8075
rect 26792 8032 26844 8041
rect 27068 8032 27120 8084
rect 28816 8032 28868 8084
rect 29184 8032 29236 8084
rect 29276 8032 29328 8084
rect 36544 8032 36596 8084
rect 21732 7964 21784 8016
rect 22100 7964 22152 8016
rect 25504 7964 25556 8016
rect 26240 7964 26292 8016
rect 26516 7964 26568 8016
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 19984 7828 20036 7880
rect 21088 7828 21140 7880
rect 21456 7828 21508 7880
rect 24124 7896 24176 7948
rect 27804 7964 27856 8016
rect 29368 7964 29420 8016
rect 29736 7964 29788 8016
rect 30380 7964 30432 8016
rect 30932 7964 30984 8016
rect 31944 7964 31996 8016
rect 33048 7964 33100 8016
rect 23756 7828 23808 7880
rect 24584 7828 24636 7880
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 25688 7828 25740 7880
rect 28632 7896 28684 7948
rect 27712 7828 27764 7880
rect 27896 7871 27948 7880
rect 27896 7837 27905 7871
rect 27905 7837 27939 7871
rect 27939 7837 27948 7871
rect 27896 7828 27948 7837
rect 27988 7828 28040 7880
rect 28908 7828 28960 7880
rect 29920 7896 29972 7948
rect 30472 7896 30524 7948
rect 31392 7896 31444 7948
rect 32680 7896 32732 7948
rect 19156 7760 19208 7812
rect 19340 7692 19392 7744
rect 24676 7760 24728 7812
rect 25596 7760 25648 7812
rect 19616 7692 19668 7744
rect 21916 7692 21968 7744
rect 22928 7692 22980 7744
rect 26056 7692 26108 7744
rect 26700 7692 26752 7744
rect 27436 7735 27488 7744
rect 27436 7701 27445 7735
rect 27445 7701 27479 7735
rect 27479 7701 27488 7735
rect 27436 7692 27488 7701
rect 28816 7760 28868 7812
rect 29184 7760 29236 7812
rect 29460 7760 29512 7812
rect 30196 7760 30248 7812
rect 31024 7871 31076 7880
rect 31024 7837 31033 7871
rect 31033 7837 31067 7871
rect 31067 7837 31076 7871
rect 31024 7828 31076 7837
rect 31944 7828 31996 7880
rect 29276 7692 29328 7744
rect 30104 7692 30156 7744
rect 30840 7760 30892 7812
rect 32864 7828 32916 7880
rect 33508 7871 33560 7880
rect 33508 7837 33517 7871
rect 33517 7837 33551 7871
rect 33551 7837 33560 7871
rect 33508 7828 33560 7837
rect 33876 7896 33928 7948
rect 34244 7964 34296 8016
rect 34336 7828 34388 7880
rect 36084 7828 36136 7880
rect 34060 7760 34112 7812
rect 34428 7803 34480 7812
rect 34428 7769 34437 7803
rect 34437 7769 34471 7803
rect 34471 7769 34480 7803
rect 34428 7760 34480 7769
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 31668 7692 31720 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 11612 7531 11664 7540
rect 11612 7497 11621 7531
rect 11621 7497 11655 7531
rect 11655 7497 11664 7531
rect 11612 7488 11664 7497
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 12072 7488 12124 7540
rect 11520 7463 11572 7472
rect 11520 7429 11529 7463
rect 11529 7429 11563 7463
rect 11563 7429 11572 7463
rect 11520 7420 11572 7429
rect 11888 7463 11940 7472
rect 11888 7429 11897 7463
rect 11897 7429 11931 7463
rect 11931 7429 11940 7463
rect 11888 7420 11940 7429
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 14924 7488 14976 7540
rect 15752 7488 15804 7540
rect 12072 7352 12124 7404
rect 12532 7395 12584 7404
rect 12532 7361 12541 7395
rect 12541 7361 12575 7395
rect 12575 7361 12584 7395
rect 12532 7352 12584 7361
rect 12716 7352 12768 7404
rect 13912 7352 13964 7404
rect 15108 7420 15160 7472
rect 21916 7488 21968 7540
rect 22192 7531 22244 7540
rect 22192 7497 22201 7531
rect 22201 7497 22235 7531
rect 22235 7497 22244 7531
rect 22192 7488 22244 7497
rect 23664 7488 23716 7540
rect 18788 7420 18840 7472
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 13268 7284 13320 7336
rect 14188 7327 14240 7336
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 15108 7327 15160 7336
rect 15108 7293 15117 7327
rect 15117 7293 15151 7327
rect 15151 7293 15160 7327
rect 15108 7284 15160 7293
rect 16948 7352 17000 7404
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 17776 7352 17828 7404
rect 19524 7420 19576 7472
rect 19248 7395 19300 7404
rect 19248 7361 19257 7395
rect 19257 7361 19291 7395
rect 19291 7361 19300 7395
rect 19248 7352 19300 7361
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19800 7352 19852 7404
rect 20904 7420 20956 7472
rect 21640 7420 21692 7472
rect 22008 7463 22060 7472
rect 22008 7429 22017 7463
rect 22017 7429 22051 7463
rect 22051 7429 22060 7463
rect 22008 7420 22060 7429
rect 22100 7463 22152 7472
rect 22100 7429 22109 7463
rect 22109 7429 22143 7463
rect 22143 7429 22152 7463
rect 22100 7420 22152 7429
rect 22652 7420 22704 7472
rect 23388 7420 23440 7472
rect 23940 7420 23992 7472
rect 21272 7352 21324 7404
rect 21548 7352 21600 7404
rect 22928 7352 22980 7404
rect 24124 7395 24176 7404
rect 15752 7284 15804 7336
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 16856 7216 16908 7268
rect 15108 7148 15160 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 17040 7259 17092 7268
rect 17040 7225 17049 7259
rect 17049 7225 17083 7259
rect 17083 7225 17092 7259
rect 17040 7216 17092 7225
rect 19616 7216 19668 7268
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 20168 7327 20220 7336
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 20352 7259 20404 7268
rect 20352 7225 20361 7259
rect 20361 7225 20395 7259
rect 20395 7225 20404 7259
rect 20352 7216 20404 7225
rect 20904 7216 20956 7268
rect 21824 7216 21876 7268
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24492 7488 24544 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 25596 7531 25648 7540
rect 25596 7497 25605 7531
rect 25605 7497 25639 7531
rect 25639 7497 25648 7531
rect 25596 7488 25648 7497
rect 26424 7488 26476 7540
rect 24400 7395 24452 7404
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 23848 7284 23900 7336
rect 24768 7284 24820 7336
rect 25320 7352 25372 7404
rect 25504 7395 25556 7404
rect 25504 7361 25513 7395
rect 25513 7361 25547 7395
rect 25547 7361 25556 7395
rect 25504 7352 25556 7361
rect 26516 7352 26568 7404
rect 26792 7352 26844 7404
rect 29000 7531 29052 7540
rect 29000 7497 29009 7531
rect 29009 7497 29043 7531
rect 29043 7497 29052 7531
rect 29000 7488 29052 7497
rect 30380 7488 30432 7540
rect 30748 7488 30800 7540
rect 27896 7420 27948 7472
rect 28816 7420 28868 7472
rect 27436 7352 27488 7404
rect 28080 7352 28132 7404
rect 28724 7352 28776 7404
rect 25780 7284 25832 7336
rect 26056 7284 26108 7336
rect 26240 7284 26292 7336
rect 28172 7284 28224 7336
rect 28908 7284 28960 7336
rect 29920 7352 29972 7404
rect 30104 7352 30156 7404
rect 30288 7352 30340 7404
rect 30932 7463 30984 7472
rect 30932 7429 30941 7463
rect 30941 7429 30975 7463
rect 30975 7429 30984 7463
rect 30932 7420 30984 7429
rect 31300 7420 31352 7472
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 31024 7284 31076 7336
rect 31300 7284 31352 7336
rect 31576 7352 31628 7404
rect 34152 7488 34204 7540
rect 34796 7488 34848 7540
rect 33968 7420 34020 7472
rect 34336 7420 34388 7472
rect 33140 7284 33192 7336
rect 19156 7148 19208 7200
rect 20444 7148 20496 7200
rect 20812 7148 20864 7200
rect 26792 7216 26844 7268
rect 27620 7216 27672 7268
rect 28540 7216 28592 7268
rect 22652 7148 22704 7200
rect 23848 7148 23900 7200
rect 26424 7148 26476 7200
rect 26608 7148 26660 7200
rect 27436 7148 27488 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 15292 6944 15344 6996
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 22008 6944 22060 6996
rect 22284 6944 22336 6996
rect 22652 6987 22704 6996
rect 22652 6953 22661 6987
rect 22661 6953 22695 6987
rect 22695 6953 22704 6987
rect 22652 6944 22704 6953
rect 23388 6987 23440 6996
rect 23388 6953 23397 6987
rect 23397 6953 23431 6987
rect 23431 6953 23440 6987
rect 23388 6944 23440 6953
rect 12992 6808 13044 6860
rect 14188 6876 14240 6928
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 11704 6715 11756 6724
rect 11704 6681 11713 6715
rect 11713 6681 11747 6715
rect 11747 6681 11756 6715
rect 11704 6672 11756 6681
rect 13636 6783 13688 6792
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 20168 6876 20220 6928
rect 25872 6944 25924 6996
rect 17132 6808 17184 6860
rect 24768 6876 24820 6928
rect 16764 6740 16816 6792
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 14004 6604 14056 6656
rect 14464 6604 14516 6656
rect 17040 6672 17092 6724
rect 17684 6740 17736 6792
rect 17776 6783 17828 6792
rect 17776 6749 17785 6783
rect 17785 6749 17819 6783
rect 17819 6749 17828 6783
rect 17776 6740 17828 6749
rect 19524 6740 19576 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 17592 6604 17644 6656
rect 19340 6672 19392 6724
rect 20076 6672 20128 6724
rect 20720 6672 20772 6724
rect 22100 6740 22152 6792
rect 21548 6715 21600 6724
rect 21548 6681 21557 6715
rect 21557 6681 21591 6715
rect 21591 6681 21600 6715
rect 21548 6672 21600 6681
rect 19708 6604 19760 6656
rect 23112 6783 23164 6792
rect 23112 6749 23121 6783
rect 23121 6749 23155 6783
rect 23155 6749 23164 6783
rect 23112 6740 23164 6749
rect 23480 6740 23532 6792
rect 24676 6740 24728 6792
rect 24768 6783 24820 6792
rect 24768 6749 24777 6783
rect 24777 6749 24811 6783
rect 24811 6749 24820 6783
rect 24768 6740 24820 6749
rect 26332 6944 26384 6996
rect 27528 6944 27580 6996
rect 26056 6851 26108 6860
rect 26056 6817 26065 6851
rect 26065 6817 26099 6851
rect 26099 6817 26108 6851
rect 26056 6808 26108 6817
rect 27252 6876 27304 6928
rect 28816 6876 28868 6928
rect 29184 6944 29236 6996
rect 26332 6808 26384 6860
rect 29368 6808 29420 6860
rect 29920 6808 29972 6860
rect 23480 6604 23532 6656
rect 23664 6715 23716 6724
rect 23664 6681 23673 6715
rect 23673 6681 23707 6715
rect 23707 6681 23716 6715
rect 23664 6672 23716 6681
rect 23848 6715 23900 6724
rect 23848 6681 23857 6715
rect 23857 6681 23891 6715
rect 23891 6681 23900 6715
rect 23848 6672 23900 6681
rect 26424 6740 26476 6792
rect 26516 6740 26568 6792
rect 25228 6672 25280 6724
rect 26792 6740 26844 6792
rect 27344 6783 27396 6792
rect 27344 6749 27353 6783
rect 27353 6749 27387 6783
rect 27387 6749 27396 6783
rect 27344 6740 27396 6749
rect 27528 6740 27580 6792
rect 28632 6740 28684 6792
rect 30656 6944 30708 6996
rect 32588 6944 32640 6996
rect 34428 6944 34480 6996
rect 30840 6851 30892 6860
rect 30840 6817 30858 6851
rect 30858 6817 30892 6851
rect 30840 6808 30892 6817
rect 30932 6808 30984 6860
rect 31300 6851 31352 6860
rect 31300 6817 31309 6851
rect 31309 6817 31343 6851
rect 31343 6817 31352 6851
rect 31300 6808 31352 6817
rect 33140 6808 33192 6860
rect 28448 6715 28500 6724
rect 28448 6681 28457 6715
rect 28457 6681 28491 6715
rect 28491 6681 28500 6715
rect 28448 6672 28500 6681
rect 28724 6672 28776 6724
rect 29552 6672 29604 6724
rect 33784 6672 33836 6724
rect 34336 6672 34388 6724
rect 23940 6604 23992 6656
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 26608 6604 26660 6656
rect 28080 6604 28132 6656
rect 28356 6604 28408 6656
rect 30564 6604 30616 6656
rect 31760 6604 31812 6656
rect 32128 6604 32180 6656
rect 36360 6604 36412 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 11704 6400 11756 6452
rect 13268 6332 13320 6384
rect 13360 6375 13412 6384
rect 13360 6341 13369 6375
rect 13369 6341 13403 6375
rect 13403 6341 13412 6375
rect 13360 6332 13412 6341
rect 15016 6332 15068 6384
rect 17684 6400 17736 6452
rect 23112 6400 23164 6452
rect 25044 6400 25096 6452
rect 11980 6307 12032 6316
rect 11980 6273 11989 6307
rect 11989 6273 12023 6307
rect 12023 6273 12032 6307
rect 11980 6264 12032 6273
rect 12072 6307 12124 6316
rect 12072 6273 12081 6307
rect 12081 6273 12115 6307
rect 12115 6273 12124 6307
rect 12072 6264 12124 6273
rect 11888 6196 11940 6248
rect 13084 6239 13136 6248
rect 13084 6205 13093 6239
rect 13093 6205 13127 6239
rect 13127 6205 13136 6239
rect 13084 6196 13136 6205
rect 14004 6196 14056 6248
rect 14924 6264 14976 6316
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 17592 6375 17644 6384
rect 17592 6341 17601 6375
rect 17601 6341 17635 6375
rect 17635 6341 17644 6375
rect 17592 6332 17644 6341
rect 18880 6332 18932 6384
rect 20444 6332 20496 6384
rect 20536 6375 20588 6384
rect 20536 6341 20545 6375
rect 20545 6341 20579 6375
rect 20579 6341 20588 6375
rect 20536 6332 20588 6341
rect 24400 6332 24452 6384
rect 26608 6400 26660 6452
rect 26700 6332 26752 6384
rect 27528 6400 27580 6452
rect 27344 6332 27396 6384
rect 28448 6400 28500 6452
rect 30196 6443 30248 6452
rect 30196 6409 30205 6443
rect 30205 6409 30239 6443
rect 30239 6409 30248 6443
rect 30196 6400 30248 6409
rect 28632 6332 28684 6384
rect 28724 6375 28776 6384
rect 28724 6341 28733 6375
rect 28733 6341 28767 6375
rect 28767 6341 28776 6375
rect 28724 6332 28776 6341
rect 16672 6264 16724 6316
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 17224 6264 17276 6316
rect 18972 6264 19024 6316
rect 19156 6196 19208 6248
rect 19340 6239 19392 6248
rect 19340 6205 19349 6239
rect 19349 6205 19383 6239
rect 19383 6205 19392 6239
rect 19340 6196 19392 6205
rect 19524 6196 19576 6248
rect 19800 6128 19852 6180
rect 21640 6264 21692 6316
rect 21916 6264 21968 6316
rect 23664 6264 23716 6316
rect 25780 6307 25832 6316
rect 25780 6273 25789 6307
rect 25789 6273 25823 6307
rect 25823 6273 25832 6307
rect 25780 6264 25832 6273
rect 25872 6264 25924 6316
rect 27252 6264 27304 6316
rect 27528 6264 27580 6316
rect 28264 6264 28316 6316
rect 33140 6400 33192 6452
rect 34520 6400 34572 6452
rect 33784 6332 33836 6384
rect 24584 6196 24636 6248
rect 26792 6196 26844 6248
rect 27068 6239 27120 6248
rect 27068 6205 27077 6239
rect 27077 6205 27111 6239
rect 27111 6205 27120 6239
rect 27068 6196 27120 6205
rect 29368 6196 29420 6248
rect 29920 6196 29972 6248
rect 23020 6128 23072 6180
rect 23940 6128 23992 6180
rect 24768 6128 24820 6180
rect 32772 6196 32824 6248
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 15476 6060 15528 6112
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 17224 6060 17276 6112
rect 17776 6060 17828 6112
rect 19432 6103 19484 6112
rect 19432 6069 19441 6103
rect 19441 6069 19475 6103
rect 19475 6069 19484 6103
rect 19432 6060 19484 6069
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 22008 6060 22060 6112
rect 25136 6060 25188 6112
rect 25688 6103 25740 6112
rect 25688 6069 25697 6103
rect 25697 6069 25731 6103
rect 25731 6069 25740 6103
rect 25688 6060 25740 6069
rect 26516 6103 26568 6112
rect 26516 6069 26525 6103
rect 26525 6069 26559 6103
rect 26559 6069 26568 6103
rect 26516 6060 26568 6069
rect 27344 6060 27396 6112
rect 32128 6060 32180 6112
rect 33784 6060 33836 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 13728 5856 13780 5908
rect 14280 5856 14332 5908
rect 11428 5720 11480 5772
rect 12624 5788 12676 5840
rect 17316 5856 17368 5908
rect 18880 5856 18932 5908
rect 19064 5856 19116 5908
rect 12256 5652 12308 5704
rect 13636 5720 13688 5772
rect 11888 5559 11940 5568
rect 11888 5525 11897 5559
rect 11897 5525 11931 5559
rect 11931 5525 11940 5559
rect 11888 5516 11940 5525
rect 12808 5584 12860 5636
rect 13820 5695 13872 5704
rect 13820 5661 13829 5695
rect 13829 5661 13863 5695
rect 13863 5661 13872 5695
rect 13820 5652 13872 5661
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 15476 5720 15528 5729
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 19616 5788 19668 5840
rect 20628 5788 20680 5840
rect 21732 5788 21784 5840
rect 21824 5788 21876 5840
rect 18420 5652 18472 5661
rect 18972 5695 19024 5704
rect 18972 5661 18981 5695
rect 18981 5661 19015 5695
rect 19015 5661 19024 5695
rect 18972 5652 19024 5661
rect 19156 5652 19208 5704
rect 19524 5652 19576 5704
rect 21088 5720 21140 5772
rect 20996 5652 21048 5704
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 21732 5695 21784 5704
rect 21732 5661 21741 5695
rect 21741 5661 21775 5695
rect 21775 5661 21784 5695
rect 21732 5652 21784 5661
rect 22008 5695 22060 5704
rect 22008 5661 22017 5695
rect 22017 5661 22051 5695
rect 22051 5661 22060 5695
rect 22008 5652 22060 5661
rect 22100 5695 22152 5704
rect 22100 5661 22109 5695
rect 22109 5661 22143 5695
rect 22143 5661 22152 5695
rect 22100 5652 22152 5661
rect 14004 5516 14056 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14832 5516 14884 5568
rect 16764 5584 16816 5636
rect 17316 5584 17368 5636
rect 20812 5584 20864 5636
rect 21824 5584 21876 5636
rect 22928 5652 22980 5704
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 23848 5856 23900 5908
rect 29644 5856 29696 5908
rect 34152 5856 34204 5908
rect 23940 5788 23992 5840
rect 24492 5720 24544 5772
rect 23388 5695 23440 5704
rect 23388 5661 23397 5695
rect 23397 5661 23431 5695
rect 23431 5661 23440 5695
rect 23388 5652 23440 5661
rect 23940 5695 23992 5704
rect 23940 5661 23949 5695
rect 23949 5661 23983 5695
rect 23983 5661 23992 5695
rect 23940 5652 23992 5661
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 24676 5652 24728 5661
rect 24768 5652 24820 5704
rect 28264 5720 28316 5772
rect 33140 5720 33192 5772
rect 16856 5516 16908 5568
rect 17500 5516 17552 5568
rect 17960 5516 18012 5568
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 20720 5516 20772 5525
rect 22100 5516 22152 5568
rect 22284 5559 22336 5568
rect 22284 5525 22293 5559
rect 22293 5525 22327 5559
rect 22327 5525 22336 5559
rect 22284 5516 22336 5525
rect 25688 5652 25740 5704
rect 29920 5652 29972 5704
rect 23572 5559 23624 5568
rect 23572 5525 23581 5559
rect 23581 5525 23615 5559
rect 23615 5525 23624 5559
rect 23572 5516 23624 5525
rect 24492 5516 24544 5568
rect 31024 5627 31076 5636
rect 31024 5593 31033 5627
rect 31033 5593 31067 5627
rect 31067 5593 31076 5627
rect 31024 5584 31076 5593
rect 32404 5627 32456 5636
rect 32404 5593 32413 5627
rect 32413 5593 32447 5627
rect 32447 5593 32456 5627
rect 32404 5584 32456 5593
rect 33784 5584 33836 5636
rect 25320 5516 25372 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 12164 5312 12216 5364
rect 13820 5312 13872 5364
rect 14004 5244 14056 5296
rect 14096 5287 14148 5296
rect 14096 5253 14105 5287
rect 14105 5253 14139 5287
rect 14139 5253 14148 5287
rect 14096 5244 14148 5253
rect 12164 5219 12216 5228
rect 12164 5185 12173 5219
rect 12173 5185 12207 5219
rect 12207 5185 12216 5219
rect 12164 5176 12216 5185
rect 15292 5244 15344 5296
rect 17592 5312 17644 5364
rect 17868 5312 17920 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 19616 5312 19668 5364
rect 17960 5244 18012 5296
rect 19340 5244 19392 5296
rect 20352 5244 20404 5296
rect 17500 5219 17552 5228
rect 17500 5185 17509 5219
rect 17509 5185 17543 5219
rect 17543 5185 17552 5219
rect 17500 5176 17552 5185
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 19616 5219 19668 5228
rect 19616 5185 19625 5219
rect 19625 5185 19659 5219
rect 19659 5185 19668 5219
rect 19616 5176 19668 5185
rect 22376 5244 22428 5296
rect 22560 5244 22612 5296
rect 24768 5244 24820 5296
rect 26424 5312 26476 5364
rect 26884 5312 26936 5364
rect 25136 5244 25188 5296
rect 12256 5108 12308 5160
rect 14924 5108 14976 5160
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 16212 5108 16264 5160
rect 16856 5108 16908 5160
rect 17776 5151 17828 5160
rect 17776 5117 17785 5151
rect 17785 5117 17819 5151
rect 17819 5117 17828 5151
rect 17776 5108 17828 5117
rect 19248 5108 19300 5160
rect 20352 5108 20404 5160
rect 11520 4972 11572 5024
rect 14648 4972 14700 5024
rect 16304 4972 16356 5024
rect 16488 4972 16540 5024
rect 21088 5040 21140 5092
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 22100 5108 22152 5117
rect 24400 5219 24452 5228
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 24400 5176 24452 5185
rect 24492 5219 24544 5228
rect 24492 5185 24501 5219
rect 24501 5185 24535 5219
rect 24535 5185 24544 5219
rect 24492 5176 24544 5185
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 20996 4972 21048 5024
rect 24400 4972 24452 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 16120 4768 16172 4820
rect 19616 4768 19668 4820
rect 20352 4811 20404 4820
rect 20352 4777 20361 4811
rect 20361 4777 20395 4811
rect 20395 4777 20404 4811
rect 20352 4768 20404 4777
rect 22928 4768 22980 4820
rect 26700 4768 26752 4820
rect 18420 4700 18472 4752
rect 20260 4700 20312 4752
rect 13084 4632 13136 4684
rect 15200 4632 15252 4684
rect 15292 4632 15344 4684
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 16856 4632 16908 4684
rect 13820 4564 13872 4616
rect 18696 4607 18748 4616
rect 18696 4573 18705 4607
rect 18705 4573 18739 4607
rect 18739 4573 18748 4607
rect 18696 4564 18748 4573
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 19892 4607 19944 4616
rect 19892 4573 19901 4607
rect 19901 4573 19935 4607
rect 19935 4573 19944 4607
rect 19892 4564 19944 4573
rect 21272 4632 21324 4684
rect 22100 4675 22152 4684
rect 22100 4641 22109 4675
rect 22109 4641 22143 4675
rect 22143 4641 22152 4675
rect 22100 4632 22152 4641
rect 23112 4632 23164 4684
rect 24860 4632 24912 4684
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 11428 4496 11480 4548
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 13176 4496 13228 4548
rect 14004 4496 14056 4548
rect 14648 4539 14700 4548
rect 14648 4505 14657 4539
rect 14657 4505 14691 4539
rect 14691 4505 14700 4539
rect 14648 4496 14700 4505
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 14924 4428 14976 4480
rect 16212 4428 16264 4480
rect 18236 4496 18288 4548
rect 19064 4496 19116 4548
rect 18144 4471 18196 4480
rect 18144 4437 18153 4471
rect 18153 4437 18187 4471
rect 18187 4437 18196 4471
rect 18144 4428 18196 4437
rect 20812 4564 20864 4616
rect 21916 4564 21968 4616
rect 21088 4496 21140 4548
rect 22284 4496 22336 4548
rect 22652 4496 22704 4548
rect 25228 4496 25280 4548
rect 27344 4428 27396 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 12164 4224 12216 4276
rect 14924 4267 14976 4276
rect 14924 4233 14933 4267
rect 14933 4233 14967 4267
rect 14967 4233 14976 4267
rect 14924 4224 14976 4233
rect 13176 4156 13228 4208
rect 4068 4088 4120 4140
rect 15292 4156 15344 4208
rect 14740 4088 14792 4140
rect 15844 4088 15896 4140
rect 17684 4224 17736 4276
rect 17592 4156 17644 4208
rect 18144 4156 18196 4208
rect 19064 4156 19116 4208
rect 17684 4131 17736 4140
rect 17684 4097 17693 4131
rect 17693 4097 17727 4131
rect 17727 4097 17736 4131
rect 17684 4088 17736 4097
rect 11336 4063 11388 4072
rect 11336 4029 11345 4063
rect 11345 4029 11379 4063
rect 11379 4029 11388 4063
rect 11336 4020 11388 4029
rect 12992 4020 13044 4072
rect 940 3952 992 4004
rect 15384 4020 15436 4072
rect 16948 3952 17000 4004
rect 17776 4063 17828 4072
rect 17776 4029 17785 4063
rect 17785 4029 17819 4063
rect 17819 4029 17828 4063
rect 17776 4020 17828 4029
rect 18512 4020 18564 4072
rect 19892 4267 19944 4276
rect 19892 4233 19901 4267
rect 19901 4233 19935 4267
rect 19935 4233 19944 4267
rect 19892 4224 19944 4233
rect 22652 4156 22704 4208
rect 24032 4156 24084 4208
rect 19432 4088 19484 4140
rect 19524 4020 19576 4072
rect 19800 4063 19852 4072
rect 19800 4029 19809 4063
rect 19809 4029 19843 4063
rect 19843 4029 19852 4063
rect 19800 4020 19852 4029
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 23296 4131 23348 4140
rect 23296 4097 23305 4131
rect 23305 4097 23339 4131
rect 23339 4097 23348 4131
rect 23296 4088 23348 4097
rect 24860 4088 24912 4140
rect 20720 4020 20772 4072
rect 23572 4063 23624 4072
rect 23572 4029 23581 4063
rect 23581 4029 23615 4063
rect 23615 4029 23624 4063
rect 23572 4020 23624 4029
rect 23940 4020 23992 4072
rect 26332 4020 26384 4072
rect 36452 4088 36504 4140
rect 19708 3952 19760 4004
rect 10968 3884 11020 3936
rect 13820 3884 13872 3936
rect 15568 3884 15620 3936
rect 18696 3884 18748 3936
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 26608 3884 26660 3936
rect 26700 3927 26752 3936
rect 26700 3893 26709 3927
rect 26709 3893 26743 3927
rect 26743 3893 26752 3927
rect 26700 3884 26752 3893
rect 36728 3884 36780 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 12256 3680 12308 3732
rect 12256 3544 12308 3596
rect 13636 3544 13688 3596
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 16948 3723 17000 3732
rect 16948 3689 16957 3723
rect 16957 3689 16991 3723
rect 16991 3689 17000 3723
rect 16948 3680 17000 3689
rect 17684 3680 17736 3732
rect 26332 3680 26384 3732
rect 27344 3680 27396 3732
rect 36084 3680 36136 3732
rect 17592 3612 17644 3664
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11244 3476 11296 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 12808 3476 12860 3528
rect 13084 3476 13136 3528
rect 13728 3476 13780 3528
rect 11704 3451 11756 3460
rect 11704 3417 11713 3451
rect 11713 3417 11747 3451
rect 11747 3417 11756 3451
rect 11704 3408 11756 3417
rect 9864 3340 9916 3392
rect 12716 3340 12768 3392
rect 14648 3408 14700 3460
rect 15200 3587 15252 3596
rect 15200 3553 15209 3587
rect 15209 3553 15243 3587
rect 15243 3553 15252 3587
rect 15200 3544 15252 3553
rect 15476 3544 15528 3596
rect 16764 3476 16816 3528
rect 15384 3408 15436 3460
rect 15568 3408 15620 3460
rect 16120 3408 16172 3460
rect 20352 3612 20404 3664
rect 23940 3612 23992 3664
rect 18604 3544 18656 3596
rect 18420 3476 18472 3528
rect 18788 3476 18840 3528
rect 19156 3476 19208 3528
rect 19524 3476 19576 3528
rect 23296 3544 23348 3596
rect 26700 3612 26752 3664
rect 26608 3544 26660 3596
rect 27344 3519 27396 3528
rect 27344 3485 27353 3519
rect 27353 3485 27387 3519
rect 27387 3485 27396 3519
rect 27344 3476 27396 3485
rect 13452 3340 13504 3392
rect 17040 3383 17092 3392
rect 17040 3349 17049 3383
rect 17049 3349 17083 3383
rect 17083 3349 17092 3383
rect 17040 3340 17092 3349
rect 17132 3340 17184 3392
rect 24032 3408 24084 3460
rect 18144 3340 18196 3392
rect 25136 3408 25188 3460
rect 36084 3451 36136 3460
rect 36084 3417 36093 3451
rect 36093 3417 36127 3451
rect 36127 3417 36136 3451
rect 36084 3408 36136 3417
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 26240 3340 26292 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 11428 3136 11480 3188
rect 11704 3136 11756 3188
rect 12716 3136 12768 3188
rect 9864 3111 9916 3120
rect 9864 3077 9873 3111
rect 9873 3077 9907 3111
rect 9907 3077 9916 3111
rect 9864 3068 9916 3077
rect 11980 3000 12032 3052
rect 13452 3068 13504 3120
rect 13728 3068 13780 3120
rect 15292 3068 15344 3120
rect 16120 3000 16172 3052
rect 17776 3136 17828 3188
rect 17132 3111 17184 3120
rect 17132 3077 17141 3111
rect 17141 3077 17175 3111
rect 17175 3077 17184 3111
rect 17132 3068 17184 3077
rect 18236 3000 18288 3052
rect 22100 3136 22152 3188
rect 24032 3136 24084 3188
rect 19432 3068 19484 3120
rect 23296 3068 23348 3120
rect 24860 3136 24912 3188
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 26240 3068 26292 3120
rect 26424 3000 26476 3052
rect 11336 2975 11388 2984
rect 11336 2941 11345 2975
rect 11345 2941 11379 2975
rect 11379 2941 11388 2975
rect 11336 2932 11388 2941
rect 12256 2932 12308 2984
rect 12808 2864 12860 2916
rect 15200 2796 15252 2848
rect 16764 2932 16816 2984
rect 18972 2975 19024 2984
rect 18972 2941 18981 2975
rect 18981 2941 19015 2975
rect 19015 2941 19024 2975
rect 18972 2932 19024 2941
rect 20444 2975 20496 2984
rect 20444 2941 20453 2975
rect 20453 2941 20487 2975
rect 20487 2941 20496 2975
rect 20444 2932 20496 2941
rect 18144 2796 18196 2848
rect 19708 2796 19760 2848
rect 23848 2796 23900 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 14648 2635 14700 2644
rect 14648 2601 14657 2635
rect 14657 2601 14691 2635
rect 14691 2601 14700 2635
rect 14648 2592 14700 2601
rect 17500 2592 17552 2644
rect 18972 2592 19024 2644
rect 18420 2567 18472 2576
rect 18420 2533 18429 2567
rect 18429 2533 18463 2567
rect 18463 2533 18472 2567
rect 18420 2524 18472 2533
rect 11336 2456 11388 2508
rect 11888 2388 11940 2440
rect 15200 2499 15252 2508
rect 15200 2465 15209 2499
rect 15209 2465 15243 2499
rect 15243 2465 15252 2499
rect 15200 2456 15252 2465
rect 15476 2456 15528 2508
rect 17040 2456 17092 2508
rect 19708 2456 19760 2508
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 13820 2388 13872 2440
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 24492 2388 24544 2440
rect 24952 2388 25004 2440
rect 18236 2320 18288 2372
rect 11612 2252 11664 2304
rect 12256 2252 12308 2304
rect 12900 2252 12952 2304
rect 13544 2252 13596 2304
rect 14188 2252 14240 2304
rect 15476 2252 15528 2304
rect 16120 2252 16172 2304
rect 25136 2252 25188 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 5814 39039 5870 39839
rect 6458 39039 6514 39839
rect 7102 39039 7158 39839
rect 7746 39039 7802 39839
rect 8390 39039 8446 39839
rect 9034 39039 9090 39839
rect 9678 39039 9734 39839
rect 10322 39039 10378 39839
rect 10966 39039 11022 39839
rect 11610 39039 11666 39839
rect 12254 39039 12310 39839
rect 12898 39039 12954 39839
rect 13004 39086 13400 39114
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 5828 37262 5856 39039
rect 6472 37482 6500 39039
rect 6472 37454 6592 37482
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 4436 37120 4488 37126
rect 4436 37062 4488 37068
rect 4448 36854 4476 37062
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4436 36848 4488 36854
rect 4436 36790 4488 36796
rect 5828 36786 5856 37198
rect 5816 36780 5868 36786
rect 5816 36722 5868 36728
rect 5540 36576 5592 36582
rect 5540 36518 5592 36524
rect 6460 36576 6512 36582
rect 6460 36518 6512 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5552 35630 5580 36518
rect 6472 36242 6500 36518
rect 6460 36236 6512 36242
rect 6460 36178 6512 36184
rect 5540 35624 5592 35630
rect 5540 35566 5592 35572
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 5552 35154 5580 35566
rect 6564 35154 6592 37454
rect 6920 36712 6972 36718
rect 6920 36654 6972 36660
rect 6932 36378 6960 36654
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 7116 35630 7144 39039
rect 7564 37324 7616 37330
rect 7564 37266 7616 37272
rect 7472 37120 7524 37126
rect 7472 37062 7524 37068
rect 7380 36848 7432 36854
rect 7380 36790 7432 36796
rect 7392 36038 7420 36790
rect 7484 36242 7512 37062
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 7380 36032 7432 36038
rect 7380 35974 7432 35980
rect 7392 35834 7420 35974
rect 7380 35828 7432 35834
rect 7380 35770 7432 35776
rect 7012 35624 7064 35630
rect 7012 35566 7064 35572
rect 7104 35624 7156 35630
rect 7104 35566 7156 35572
rect 7024 35290 7052 35566
rect 7012 35284 7064 35290
rect 7012 35226 7064 35232
rect 7116 35154 7144 35566
rect 7576 35154 7604 37266
rect 7760 35894 7788 39039
rect 8404 37262 8432 39039
rect 9048 37346 9076 39039
rect 8956 37318 9076 37346
rect 9588 37324 9640 37330
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 8300 37188 8352 37194
rect 8300 37130 8352 37136
rect 8024 36780 8076 36786
rect 8024 36722 8076 36728
rect 8036 36106 8064 36722
rect 8312 36582 8340 37130
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 8404 36242 8432 37198
rect 8760 36712 8812 36718
rect 8760 36654 8812 36660
rect 8772 36310 8800 36654
rect 8760 36304 8812 36310
rect 8760 36246 8812 36252
rect 8392 36236 8444 36242
rect 8392 36178 8444 36184
rect 8024 36100 8076 36106
rect 8024 36042 8076 36048
rect 7760 35866 7880 35894
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 6552 35148 6604 35154
rect 6552 35090 6604 35096
rect 7104 35148 7156 35154
rect 7104 35090 7156 35096
rect 7564 35148 7616 35154
rect 7564 35090 7616 35096
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 5460 34746 5488 34954
rect 5448 34740 5500 34746
rect 5448 34682 5500 34688
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5552 34066 5580 35090
rect 6564 34746 6592 35090
rect 6552 34740 6604 34746
rect 6552 34682 6604 34688
rect 7576 34542 7604 35090
rect 7564 34536 7616 34542
rect 7564 34478 7616 34484
rect 5540 34060 5592 34066
rect 5540 34002 5592 34008
rect 6368 34060 6420 34066
rect 6368 34002 6420 34008
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 6380 33522 6408 34002
rect 7012 33924 7064 33930
rect 7012 33866 7064 33872
rect 7024 33658 7052 33866
rect 7012 33652 7064 33658
rect 7012 33594 7064 33600
rect 6368 33516 6420 33522
rect 6368 33458 6420 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 2688 32496 2740 32502
rect 2688 32438 2740 32444
rect 2700 31822 2728 32438
rect 4896 32428 4948 32434
rect 4896 32370 4948 32376
rect 5356 32428 5408 32434
rect 5356 32370 5408 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4908 32026 4936 32370
rect 4896 32020 4948 32026
rect 4896 31962 4948 31968
rect 2688 31816 2740 31822
rect 2688 31758 2740 31764
rect 2700 31385 2728 31758
rect 4068 31748 4120 31754
rect 4068 31690 4120 31696
rect 5264 31748 5316 31754
rect 5264 31690 5316 31696
rect 2686 31376 2742 31385
rect 2686 31311 2742 31320
rect 3700 31204 3752 31210
rect 3700 31146 3752 31152
rect 3712 30326 3740 31146
rect 4080 30666 4108 31690
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5276 31362 5304 31690
rect 5368 31686 5396 32370
rect 5540 32224 5592 32230
rect 5540 32166 5592 32172
rect 5552 31890 5580 32166
rect 5540 31884 5592 31890
rect 5540 31826 5592 31832
rect 5356 31680 5408 31686
rect 5356 31622 5408 31628
rect 5368 31414 5396 31622
rect 6380 31414 6408 33458
rect 7852 33454 7880 35866
rect 7932 35760 7984 35766
rect 7932 35702 7984 35708
rect 7944 35018 7972 35702
rect 7932 35012 7984 35018
rect 7932 34954 7984 34960
rect 7944 33862 7972 34954
rect 8298 34640 8354 34649
rect 8298 34575 8300 34584
rect 8352 34575 8354 34584
rect 8300 34546 8352 34552
rect 8666 34504 8722 34513
rect 8666 34439 8668 34448
rect 8720 34439 8722 34448
rect 8668 34410 8720 34416
rect 8956 34134 8984 37318
rect 9588 37266 9640 37272
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 9048 36718 9076 37062
rect 9036 36712 9088 36718
rect 9036 36654 9088 36660
rect 9220 36576 9272 36582
rect 9220 36518 9272 36524
rect 9232 35698 9260 36518
rect 9600 36242 9628 37266
rect 9692 36922 9720 39039
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 9680 36916 9732 36922
rect 9680 36858 9732 36864
rect 9588 36236 9640 36242
rect 9588 36178 9640 36184
rect 9692 36174 9720 36858
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9772 36100 9824 36106
rect 9772 36042 9824 36048
rect 9784 35698 9812 36042
rect 9220 35692 9272 35698
rect 9220 35634 9272 35640
rect 9496 35692 9548 35698
rect 9496 35634 9548 35640
rect 9772 35692 9824 35698
rect 9772 35634 9824 35640
rect 9312 35624 9364 35630
rect 9312 35566 9364 35572
rect 9324 35290 9352 35566
rect 9312 35284 9364 35290
rect 9312 35226 9364 35232
rect 9220 35080 9272 35086
rect 9220 35022 9272 35028
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9232 34746 9260 35022
rect 9220 34740 9272 34746
rect 9220 34682 9272 34688
rect 9416 34678 9444 35022
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 9508 34542 9536 35634
rect 9784 34610 9812 35634
rect 9956 35624 10008 35630
rect 9956 35566 10008 35572
rect 9968 35290 9996 35566
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 10060 35222 10088 37062
rect 10232 35556 10284 35562
rect 10232 35498 10284 35504
rect 10244 35329 10272 35498
rect 10230 35320 10286 35329
rect 10230 35255 10286 35264
rect 10048 35216 10100 35222
rect 10048 35158 10100 35164
rect 9956 35080 10008 35086
rect 9956 35022 10008 35028
rect 9772 34604 9824 34610
rect 9772 34546 9824 34552
rect 9496 34536 9548 34542
rect 9496 34478 9548 34484
rect 8944 34128 8996 34134
rect 8944 34070 8996 34076
rect 9508 34066 9536 34478
rect 9784 34377 9812 34546
rect 9968 34406 9996 35022
rect 10060 35018 10088 35158
rect 10232 35080 10284 35086
rect 10232 35022 10284 35028
rect 10048 35012 10100 35018
rect 10048 34954 10100 34960
rect 10060 34474 10088 34954
rect 10244 34610 10272 35022
rect 10232 34604 10284 34610
rect 10232 34546 10284 34552
rect 10048 34468 10100 34474
rect 10048 34410 10100 34416
rect 9956 34400 10008 34406
rect 9770 34368 9826 34377
rect 9956 34342 10008 34348
rect 9770 34303 9826 34312
rect 8668 34060 8720 34066
rect 8668 34002 8720 34008
rect 9496 34060 9548 34066
rect 9496 34002 9548 34008
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7944 33590 7972 33798
rect 7932 33584 7984 33590
rect 7932 33526 7984 33532
rect 8680 33522 8708 34002
rect 10060 33998 10088 34410
rect 10244 34202 10272 34546
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 8852 33992 8904 33998
rect 8852 33934 8904 33940
rect 10048 33992 10100 33998
rect 10048 33934 10100 33940
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 8484 33516 8536 33522
rect 8484 33458 8536 33464
rect 8668 33516 8720 33522
rect 8668 33458 8720 33464
rect 7012 33448 7064 33454
rect 7012 33390 7064 33396
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7024 33114 7052 33390
rect 7012 33108 7064 33114
rect 7012 33050 7064 33056
rect 7852 32910 7880 33390
rect 8496 33046 8524 33458
rect 8300 33040 8352 33046
rect 8300 32982 8352 32988
rect 8484 33040 8536 33046
rect 8484 32982 8536 32988
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 6552 32564 6604 32570
rect 6552 32506 6604 32512
rect 6564 31822 6592 32506
rect 7288 32496 7340 32502
rect 7288 32438 7340 32444
rect 7932 32496 7984 32502
rect 7932 32438 7984 32444
rect 7104 32360 7156 32366
rect 7104 32302 7156 32308
rect 7116 32026 7144 32302
rect 7196 32224 7248 32230
rect 7196 32166 7248 32172
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 6920 31952 6972 31958
rect 6920 31894 6972 31900
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 5184 31334 5304 31362
rect 5356 31408 5408 31414
rect 5356 31350 5408 31356
rect 6368 31408 6420 31414
rect 6368 31350 6420 31356
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5184 30734 5212 31334
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5172 30728 5224 30734
rect 5170 30696 5172 30705
rect 5224 30696 5226 30705
rect 4068 30660 4120 30666
rect 5170 30631 5226 30640
rect 4068 30602 4120 30608
rect 4080 30326 4108 30602
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5552 30326 5580 31078
rect 6380 30784 6408 31350
rect 6288 30756 6408 30784
rect 5632 30660 5684 30666
rect 5632 30602 5684 30608
rect 5644 30394 5672 30602
rect 5632 30388 5684 30394
rect 5632 30330 5684 30336
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 4068 30320 4120 30326
rect 4068 30262 4120 30268
rect 5540 30320 5592 30326
rect 5540 30262 5592 30268
rect 3056 29708 3108 29714
rect 3056 29650 3108 29656
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 2872 29504 2924 29510
rect 2872 29446 2924 29452
rect 1780 29238 1808 29446
rect 1768 29232 1820 29238
rect 1768 29174 1820 29180
rect 1400 29096 1452 29102
rect 1400 29038 1452 29044
rect 1412 28558 1440 29038
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1412 27470 1440 28494
rect 1676 28484 1728 28490
rect 1676 28426 1728 28432
rect 1688 28218 1716 28426
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 2780 28076 2832 28082
rect 2780 28018 2832 28024
rect 2504 27872 2556 27878
rect 2504 27814 2556 27820
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 26858 1440 27406
rect 1676 27396 1728 27402
rect 1676 27338 1728 27344
rect 1688 27130 1716 27338
rect 1676 27124 1728 27130
rect 1676 27066 1728 27072
rect 1400 26852 1452 26858
rect 1400 26794 1452 26800
rect 1412 25838 1440 26794
rect 1400 25832 1452 25838
rect 1400 25774 1452 25780
rect 2228 25832 2280 25838
rect 2228 25774 2280 25780
rect 2412 25832 2464 25838
rect 2412 25774 2464 25780
rect 1412 25702 1440 25774
rect 1400 25696 1452 25702
rect 1400 25638 1452 25644
rect 1412 24750 1440 25638
rect 2240 25498 2268 25774
rect 2424 25702 2452 25774
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2228 25492 2280 25498
rect 2228 25434 2280 25440
rect 2412 25152 2464 25158
rect 2412 25094 2464 25100
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1412 23186 1440 24686
rect 2320 24064 2372 24070
rect 2320 24006 2372 24012
rect 2332 23866 2360 24006
rect 2320 23860 2372 23866
rect 2320 23802 2372 23808
rect 2320 23656 2372 23662
rect 2424 23644 2452 25094
rect 2372 23616 2452 23644
rect 2320 23598 2372 23604
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23186 1716 23462
rect 1400 23180 1452 23186
rect 1400 23122 1452 23128
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 1688 22234 1716 22374
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1412 21554 1440 22034
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 20466 1440 21490
rect 1676 20800 1728 20806
rect 1676 20742 1728 20748
rect 1400 20460 1452 20466
rect 1400 20402 1452 20408
rect 1412 19922 1440 20402
rect 1688 19922 1716 20742
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1412 18834 1440 19858
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 18290 1440 18770
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17882 1716 18158
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 2332 17746 2360 23598
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16182 1716 16934
rect 1676 16176 1728 16182
rect 1676 16118 1728 16124
rect 2424 12306 2452 21830
rect 2516 20602 2544 27814
rect 2792 27674 2820 28018
rect 2780 27668 2832 27674
rect 2780 27610 2832 27616
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 2700 27130 2728 27474
rect 2688 27124 2740 27130
rect 2688 27066 2740 27072
rect 2780 24676 2832 24682
rect 2780 24618 2832 24624
rect 2792 23730 2820 24618
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2596 23656 2648 23662
rect 2596 23598 2648 23604
rect 2608 22574 2636 23598
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2700 22098 2728 23666
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2792 21944 2820 22102
rect 2700 21916 2820 21944
rect 2504 20596 2556 20602
rect 2504 20538 2556 20544
rect 2700 19514 2728 21916
rect 2884 20942 2912 29446
rect 3068 28014 3096 29650
rect 3712 29345 3740 30262
rect 3698 29336 3754 29345
rect 4080 29306 4108 30262
rect 6288 30258 6316 30756
rect 5816 30252 5868 30258
rect 5816 30194 5868 30200
rect 6276 30252 6328 30258
rect 6276 30194 6328 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4344 29640 4396 29646
rect 4344 29582 4396 29588
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 4160 29504 4212 29510
rect 4160 29446 4212 29452
rect 3698 29271 3754 29280
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4172 29238 4200 29446
rect 4160 29232 4212 29238
rect 4356 29209 4384 29582
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4160 29174 4212 29180
rect 4342 29200 4398 29209
rect 4342 29135 4398 29144
rect 4356 29102 4384 29135
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4252 28756 4304 28762
rect 4252 28698 4304 28704
rect 3148 28416 3200 28422
rect 3148 28358 3200 28364
rect 3160 28082 3188 28358
rect 4264 28150 4292 28698
rect 4528 28620 4580 28626
rect 4528 28562 4580 28568
rect 4252 28144 4304 28150
rect 4158 28112 4214 28121
rect 3148 28076 3200 28082
rect 4252 28086 4304 28092
rect 4158 28047 4160 28056
rect 3148 28018 3200 28024
rect 4212 28047 4214 28056
rect 4436 28076 4488 28082
rect 4160 28018 4212 28024
rect 4540 28064 4568 28562
rect 4632 28234 4660 29446
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4804 29300 4856 29306
rect 4804 29242 4856 29248
rect 4710 29200 4766 29209
rect 4710 29135 4766 29144
rect 4724 28626 4752 29135
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 4816 28490 4844 29242
rect 5276 29186 5304 29582
rect 5448 29572 5500 29578
rect 5448 29514 5500 29520
rect 5184 29170 5304 29186
rect 5184 29164 5316 29170
rect 5184 29158 5264 29164
rect 5184 28762 5212 29158
rect 5264 29106 5316 29112
rect 5264 29028 5316 29034
rect 5264 28970 5316 28976
rect 5172 28756 5224 28762
rect 5172 28698 5224 28704
rect 5276 28626 5304 28970
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 5264 28620 5316 28626
rect 5264 28562 5316 28568
rect 4804 28484 4856 28490
rect 4804 28426 4856 28432
rect 5368 28404 5396 28902
rect 5460 28762 5488 29514
rect 5724 29504 5776 29510
rect 5724 29446 5776 29452
rect 5736 29306 5764 29446
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5448 28756 5500 28762
rect 5448 28698 5500 28704
rect 5828 28626 5856 30194
rect 6748 30190 6776 31418
rect 6932 30802 6960 31894
rect 7208 31890 7236 32166
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 7208 31414 7236 31826
rect 7196 31408 7248 31414
rect 7196 31350 7248 31356
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 7208 30734 7236 31350
rect 7196 30728 7248 30734
rect 7196 30670 7248 30676
rect 7104 30592 7156 30598
rect 7104 30534 7156 30540
rect 7116 30326 7144 30534
rect 7104 30320 7156 30326
rect 7104 30262 7156 30268
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6656 29850 6684 30126
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6276 29708 6328 29714
rect 6276 29650 6328 29656
rect 6288 29102 6316 29650
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 6932 29238 6960 29582
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 7116 29306 7144 29446
rect 7104 29300 7156 29306
rect 7104 29242 7156 29248
rect 6644 29232 6696 29238
rect 6920 29232 6972 29238
rect 6696 29180 6868 29186
rect 6644 29174 6868 29180
rect 6920 29174 6972 29180
rect 6656 29158 6868 29174
rect 6276 29096 6328 29102
rect 6276 29038 6328 29044
rect 6092 28960 6144 28966
rect 6092 28902 6144 28908
rect 6104 28626 6132 28902
rect 5816 28620 5868 28626
rect 5816 28562 5868 28568
rect 6092 28620 6144 28626
rect 6092 28562 6144 28568
rect 5448 28416 5500 28422
rect 5368 28376 5448 28404
rect 5448 28358 5500 28364
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4632 28218 4844 28234
rect 4632 28212 4856 28218
rect 4632 28206 4804 28212
rect 4804 28154 4856 28160
rect 4986 28112 5042 28121
rect 4488 28036 4568 28064
rect 4620 28076 4672 28082
rect 4436 28018 4488 28024
rect 5460 28082 5488 28358
rect 4672 28036 4844 28064
rect 4986 28047 4988 28056
rect 4620 28018 4672 28024
rect 3056 28008 3108 28014
rect 3056 27950 3108 27956
rect 3068 26926 3096 27950
rect 4712 27872 4764 27878
rect 4712 27814 4764 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3792 27396 3844 27402
rect 3792 27338 3844 27344
rect 3700 27124 3752 27130
rect 3700 27066 3752 27072
rect 3146 27024 3202 27033
rect 3146 26959 3202 26968
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 2964 25968 3016 25974
rect 2964 25910 3016 25916
rect 2976 24886 3004 25910
rect 3068 25362 3096 26862
rect 3160 26042 3188 26959
rect 3712 26790 3740 27066
rect 3804 27062 3832 27338
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 27062 4108 27270
rect 3792 27056 3844 27062
rect 3792 26998 3844 27004
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 3700 26784 3752 26790
rect 3700 26726 3752 26732
rect 3148 26036 3200 26042
rect 3148 25978 3200 25984
rect 3056 25356 3108 25362
rect 3056 25298 3108 25304
rect 3160 25294 3188 25978
rect 3148 25288 3200 25294
rect 3200 25248 3280 25276
rect 3148 25230 3200 25236
rect 2964 24880 3016 24886
rect 2964 24822 3016 24828
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 3068 23322 3096 23598
rect 3056 23316 3108 23322
rect 3056 23258 3108 23264
rect 3160 23050 3188 23734
rect 3252 23526 3280 25248
rect 3608 24880 3660 24886
rect 3608 24822 3660 24828
rect 3620 24274 3648 24822
rect 3608 24268 3660 24274
rect 3608 24210 3660 24216
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3240 23520 3292 23526
rect 3240 23462 3292 23468
rect 3436 23254 3464 24142
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3148 23044 3200 23050
rect 3148 22986 3200 22992
rect 3424 23044 3476 23050
rect 3424 22986 3476 22992
rect 3160 21978 3188 22986
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 2976 21962 3188 21978
rect 2964 21956 3188 21962
rect 3016 21950 3188 21956
rect 2964 21898 3016 21904
rect 2976 21486 3004 21898
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2884 20058 2912 20742
rect 2976 20466 3004 21422
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2976 19786 3004 20402
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2688 19508 2740 19514
rect 2688 19450 2740 19456
rect 2700 19334 2728 19450
rect 3252 19446 3280 22714
rect 3332 21480 3384 21486
rect 3332 21422 3384 21428
rect 3240 19440 3292 19446
rect 3240 19382 3292 19388
rect 2608 19306 2728 19334
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 2516 16998 2544 17682
rect 2608 17270 2636 19306
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2688 18828 2740 18834
rect 2688 18770 2740 18776
rect 2700 18222 2728 18770
rect 2792 18630 2820 19110
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2976 17814 3004 19246
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17338 2728 17478
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2976 17270 3004 17750
rect 3252 17542 3280 19382
rect 3344 18426 3372 21422
rect 3436 19446 3464 22986
rect 3620 22778 3648 24210
rect 3608 22772 3660 22778
rect 3608 22714 3660 22720
rect 3712 22234 3740 26726
rect 3804 26450 3832 26998
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 3976 25968 4028 25974
rect 4080 25922 4108 26998
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4160 26240 4212 26246
rect 4160 26182 4212 26188
rect 4028 25916 4108 25922
rect 3976 25910 4108 25916
rect 3988 25894 4108 25910
rect 4080 25838 4108 25894
rect 3884 25832 3936 25838
rect 3884 25774 3936 25780
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 3896 25498 3924 25774
rect 4172 25684 4200 26182
rect 4724 25922 4752 27814
rect 4816 27402 4844 28036
rect 5040 28047 5042 28056
rect 5448 28076 5500 28082
rect 4988 28018 5040 28024
rect 5448 28018 5500 28024
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 5000 27470 5028 28018
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 5448 27464 5500 27470
rect 5736 27452 5764 28018
rect 5816 27940 5868 27946
rect 5816 27882 5868 27888
rect 5500 27424 5764 27452
rect 5448 27406 5500 27412
rect 4804 27396 4856 27402
rect 4804 27338 4856 27344
rect 4816 27130 4844 27338
rect 5172 27328 5224 27334
rect 5224 27288 5304 27316
rect 5172 27270 5224 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4804 27124 4856 27130
rect 4804 27066 4856 27072
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4816 26586 4844 26862
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 5184 26314 5212 26726
rect 5172 26308 5224 26314
rect 5172 26250 5224 26256
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4724 25894 4844 25922
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 3988 25656 4200 25684
rect 3884 25492 3936 25498
rect 3884 25434 3936 25440
rect 3792 25356 3844 25362
rect 3792 25298 3844 25304
rect 3804 24750 3832 25298
rect 3988 25158 4016 25656
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3804 22094 3832 24686
rect 3988 23322 4016 25094
rect 4724 24886 4752 25774
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4816 24834 4844 25894
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 4080 24342 4108 24754
rect 4528 24744 4580 24750
rect 4724 24698 4752 24822
rect 4816 24806 4936 24834
rect 4804 24744 4856 24750
rect 4580 24692 4660 24698
rect 4528 24686 4660 24692
rect 4540 24670 4660 24686
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24410 4660 24670
rect 4724 24692 4804 24698
rect 4724 24686 4856 24692
rect 4724 24670 4844 24686
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4068 24336 4120 24342
rect 4068 24278 4120 24284
rect 4080 23866 4108 24278
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4540 23866 4568 24142
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4528 23860 4580 23866
rect 4528 23802 4580 23808
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3988 23050 4016 23258
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 3976 23044 4028 23050
rect 3976 22986 4028 22992
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3712 22066 3832 22094
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3528 18698 3556 20742
rect 3712 19242 3740 22066
rect 3792 21888 3844 21894
rect 3792 21830 3844 21836
rect 3804 21690 3832 21830
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3896 21418 3924 22578
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 3988 22234 4016 22510
rect 4080 22506 4108 23122
rect 4528 23112 4580 23118
rect 4632 23100 4660 24006
rect 4724 23662 4752 24670
rect 4908 24562 4936 24806
rect 4816 24534 4936 24562
rect 4712 23656 4764 23662
rect 4712 23598 4764 23604
rect 4712 23248 4764 23254
rect 4712 23190 4764 23196
rect 4724 23118 4752 23190
rect 4580 23072 4660 23100
rect 4712 23112 4764 23118
rect 4528 23054 4580 23060
rect 4712 23054 4764 23060
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4436 22636 4488 22642
rect 4436 22578 4488 22584
rect 4448 22506 4476 22578
rect 4068 22500 4120 22506
rect 4068 22442 4120 22448
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3988 22098 4016 22170
rect 4080 22137 4108 22442
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4066 22128 4122 22137
rect 3976 22092 4028 22098
rect 4066 22063 4122 22072
rect 4342 22128 4398 22137
rect 4632 22094 4660 22918
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4724 22234 4752 22578
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4342 22063 4344 22072
rect 3976 22034 4028 22040
rect 3884 21412 3936 21418
rect 3884 21354 3936 21360
rect 4080 21010 4108 22063
rect 4396 22063 4398 22072
rect 4540 22066 4660 22094
rect 4344 22034 4396 22040
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4448 21690 4476 21830
rect 4436 21684 4488 21690
rect 4436 21626 4488 21632
rect 4540 21554 4568 22066
rect 4620 21956 4672 21962
rect 4620 21898 4672 21904
rect 4632 21690 4660 21898
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21128 4660 21490
rect 4540 21100 4660 21128
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3804 20602 3832 20742
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 4080 20398 4108 20946
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4356 20602 4384 20878
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 3896 19718 3924 20334
rect 4356 20262 4384 20538
rect 4540 20262 4568 21100
rect 4724 20942 4752 21830
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4712 20936 4764 20942
rect 4712 20878 4764 20884
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 20058 4660 20878
rect 4816 20466 4844 24534
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5172 23860 5224 23866
rect 5172 23802 5224 23808
rect 5184 23730 5212 23802
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 4896 23248 4948 23254
rect 4896 23190 4948 23196
rect 4908 23118 4936 23190
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 5000 23050 5028 23462
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5172 22636 5224 22642
rect 5172 22578 5224 22584
rect 5184 22166 5212 22578
rect 5172 22160 5224 22166
rect 5172 22102 5224 22108
rect 5276 22030 5304 27288
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5460 23866 5488 26454
rect 5736 26314 5764 27424
rect 5828 27130 5856 27882
rect 6184 27396 6236 27402
rect 6184 27338 6236 27344
rect 5816 27124 5868 27130
rect 5816 27066 5868 27072
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5632 25288 5684 25294
rect 5736 25276 5764 26250
rect 5828 26246 5856 27066
rect 6196 26994 6224 27338
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 6184 26988 6236 26994
rect 6184 26930 6236 26936
rect 5920 26382 5948 26930
rect 6288 26858 6316 29038
rect 6840 28914 6868 29158
rect 6840 28886 6960 28914
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6460 27396 6512 27402
rect 6460 27338 6512 27344
rect 6472 27130 6500 27338
rect 6460 27124 6512 27130
rect 6460 27066 6512 27072
rect 6276 26852 6328 26858
rect 6276 26794 6328 26800
rect 6288 26586 6316 26794
rect 6276 26580 6328 26586
rect 6276 26522 6328 26528
rect 6000 26444 6052 26450
rect 6000 26386 6052 26392
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5684 25248 5764 25276
rect 5632 25230 5684 25236
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5356 23724 5408 23730
rect 5356 23666 5408 23672
rect 5368 23254 5396 23666
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5368 22642 5396 23190
rect 5540 22704 5592 22710
rect 5540 22646 5592 22652
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5356 22500 5408 22506
rect 5356 22442 5408 22448
rect 5080 22024 5132 22030
rect 5078 21992 5080 22001
rect 5172 22024 5224 22030
rect 5132 21992 5134 22001
rect 5172 21966 5224 21972
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 5078 21927 5134 21936
rect 5184 21876 5212 21966
rect 5184 21848 5304 21876
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21622 5304 21848
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 4896 21072 4948 21078
rect 4896 21014 4948 21020
rect 5368 21026 5396 22442
rect 5460 21894 5488 22578
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 5552 21554 5580 22646
rect 5644 22642 5672 25094
rect 5736 24886 5764 25248
rect 5828 25226 5856 26182
rect 6012 25974 6040 26386
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6196 26042 6224 26318
rect 6184 26036 6236 26042
rect 6184 25978 6236 25984
rect 6000 25968 6052 25974
rect 5998 25936 6000 25945
rect 6052 25936 6054 25945
rect 5998 25871 6054 25880
rect 6196 25362 6224 25978
rect 6288 25362 6316 26522
rect 6656 25922 6684 28562
rect 6932 27674 6960 28886
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 6828 26920 6880 26926
rect 6826 26888 6828 26897
rect 6880 26888 6882 26897
rect 6826 26823 6882 26832
rect 6736 26308 6788 26314
rect 6736 26250 6788 26256
rect 6748 25974 6776 26250
rect 6564 25894 6684 25922
rect 6736 25968 6788 25974
rect 6736 25910 6788 25916
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 6276 25356 6328 25362
rect 6276 25298 6328 25304
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 5816 25220 5868 25226
rect 5816 25162 5868 25168
rect 5908 25220 5960 25226
rect 5908 25162 5960 25168
rect 5724 24880 5776 24886
rect 5724 24822 5776 24828
rect 5828 23118 5856 25162
rect 5920 24954 5948 25162
rect 6012 24954 6040 25230
rect 5908 24948 5960 24954
rect 5908 24890 5960 24896
rect 6000 24948 6052 24954
rect 6000 24890 6052 24896
rect 5920 24274 5948 24890
rect 6012 24614 6040 24890
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 6196 24206 6224 24550
rect 6288 24342 6316 25298
rect 6460 25152 6512 25158
rect 6380 25112 6460 25140
rect 6276 24336 6328 24342
rect 6276 24278 6328 24284
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 6012 23769 6040 23802
rect 5998 23760 6054 23769
rect 5998 23695 6054 23704
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5632 22636 5684 22642
rect 5632 22578 5684 22584
rect 5816 22636 5868 22642
rect 5816 22578 5868 22584
rect 5724 22568 5776 22574
rect 5724 22510 5776 22516
rect 5632 22500 5684 22506
rect 5632 22442 5684 22448
rect 5644 22098 5672 22442
rect 5632 22092 5684 22098
rect 5632 22034 5684 22040
rect 5644 21554 5672 22034
rect 5736 22030 5764 22510
rect 5724 22024 5776 22030
rect 5722 21992 5724 22001
rect 5776 21992 5778 22001
rect 5722 21927 5778 21936
rect 5736 21604 5764 21927
rect 5828 21672 5856 22578
rect 6012 22030 6040 23462
rect 6288 23186 6316 24006
rect 6276 23180 6328 23186
rect 6276 23122 6328 23128
rect 6380 23066 6408 25112
rect 6460 25094 6512 25100
rect 6460 24880 6512 24886
rect 6460 24822 6512 24828
rect 6472 24206 6500 24822
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6472 23633 6500 24142
rect 6458 23624 6514 23633
rect 6458 23559 6514 23568
rect 6288 23038 6408 23066
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 5828 21644 6040 21672
rect 5736 21576 5948 21604
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 4908 20913 4936 21014
rect 5368 20998 5488 21026
rect 5356 20936 5408 20942
rect 4894 20904 4950 20913
rect 5356 20878 5408 20884
rect 4894 20839 4950 20848
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4526 19952 4582 19961
rect 4526 19887 4582 19896
rect 4540 19854 4568 19887
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3700 19236 3752 19242
rect 3700 19178 3752 19184
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3436 18426 3464 18634
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3344 17746 3372 18362
rect 3712 18358 3740 18566
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 3608 17128 3660 17134
rect 3608 17070 3660 17076
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2700 16658 2728 16730
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 2608 16250 2636 16594
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2608 15026 2636 16186
rect 3068 16182 3096 16390
rect 3056 16176 3108 16182
rect 3056 16118 3108 16124
rect 3436 15978 3464 16594
rect 3620 16250 3648 17070
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3896 16114 3924 19654
rect 4264 19378 4292 19722
rect 4724 19378 4752 20402
rect 5092 20398 5120 20538
rect 5276 20466 5304 20742
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19990 4844 20198
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4908 19854 4936 20266
rect 5368 20058 5396 20878
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4264 19258 4292 19314
rect 4080 19230 4292 19258
rect 4080 18970 4108 19230
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4436 18828 4488 18834
rect 4436 18770 4488 18776
rect 4448 18222 4476 18770
rect 4632 18698 4660 19110
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4436 18216 4488 18222
rect 4436 18158 4488 18164
rect 3976 17264 4028 17270
rect 4080 17252 4108 18158
rect 4540 18068 4568 18566
rect 4540 18040 4660 18068
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18040
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4724 17746 4752 18702
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4028 17224 4108 17252
rect 3976 17206 4028 17212
rect 4080 16726 4108 17224
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16794 4660 17070
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3804 15706 3832 16050
rect 4080 16046 4108 16662
rect 4724 16538 4752 17546
rect 4632 16510 4752 16538
rect 4632 16182 4660 16510
rect 4712 16448 4764 16454
rect 4816 16402 4844 19790
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 5184 18970 5212 19382
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18426 5304 19314
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5368 18358 5396 18566
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5368 17270 5396 18294
rect 5460 17678 5488 20998
rect 5552 20942 5580 21490
rect 5722 21176 5778 21185
rect 5722 21111 5724 21120
rect 5776 21111 5778 21120
rect 5724 21082 5776 21088
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5644 20602 5672 20878
rect 5722 20632 5778 20641
rect 5632 20596 5684 20602
rect 5828 20602 5856 20878
rect 5920 20874 5948 21576
rect 5908 20868 5960 20874
rect 5908 20810 5960 20816
rect 5722 20567 5778 20576
rect 5816 20596 5868 20602
rect 5632 20538 5684 20544
rect 5736 20534 5764 20567
rect 5816 20538 5868 20544
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5920 20466 5948 20810
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 6012 20346 6040 21644
rect 5920 20318 6040 20346
rect 5920 20058 5948 20318
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 6012 19961 6040 20198
rect 6104 19990 6132 21966
rect 6092 19984 6144 19990
rect 5998 19952 6054 19961
rect 6092 19926 6144 19932
rect 5998 19887 6054 19896
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5262 16688 5318 16697
rect 5262 16623 5318 16632
rect 4894 16552 4950 16561
rect 4894 16487 4950 16496
rect 4908 16454 4936 16487
rect 4764 16396 4844 16402
rect 4712 16390 4844 16396
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4724 16374 4844 16390
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 4724 15570 4752 16374
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5276 15162 5304 16623
rect 5368 16522 5396 17206
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16590 5488 16934
rect 5448 16584 5500 16590
rect 5552 16561 5580 18906
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5828 17746 5856 18022
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 6196 17202 6224 21966
rect 6288 21894 6316 23038
rect 6472 22094 6500 23054
rect 6380 22066 6500 22094
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6380 21690 6408 22066
rect 6460 21956 6512 21962
rect 6460 21898 6512 21904
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6288 19718 6316 19926
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 5448 16526 5500 16532
rect 5538 16552 5594 16561
rect 5356 16516 5408 16522
rect 5538 16487 5594 16496
rect 5356 16458 5408 16464
rect 5368 16182 5396 16458
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2608 13938 2636 14962
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3252 14618 3280 14894
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3988 13938 4016 14894
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14600 4660 15098
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4448 14572 4660 14600
rect 4448 14346 4476 14572
rect 4816 14414 4844 14758
rect 5276 14414 5304 14758
rect 5552 14550 5580 14894
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 4620 14408 4672 14414
rect 4804 14408 4856 14414
rect 4672 14368 4752 14396
rect 4620 14350 4672 14356
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3988 12442 4016 13874
rect 4540 13716 4568 14282
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4632 13938 4660 14214
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4724 13870 4752 14368
rect 4804 14350 4856 14356
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 14074 5304 14214
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 4804 14000 4856 14006
rect 4802 13968 4804 13977
rect 4856 13968 4858 13977
rect 4802 13903 4858 13912
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4540 13688 4660 13716
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 13688
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4724 13410 4752 13806
rect 5368 13734 5396 14418
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 13932 5500 13938
rect 5552 13920 5580 14350
rect 5500 13892 5580 13920
rect 5448 13874 5500 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 4632 13382 4752 13410
rect 5368 13394 5396 13670
rect 5552 13394 5580 13738
rect 5356 13388 5408 13394
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3976 12436 4028 12442
rect 4632 12434 4660 13382
rect 5356 13330 5408 13336
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4724 12442 4752 13194
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5368 12986 5396 13330
rect 5552 13258 5580 13330
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 3976 12378 4028 12384
rect 4356 12406 4660 12434
rect 4712 12436 4764 12442
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 3884 11824 3936 11830
rect 3988 11812 4016 12378
rect 4356 12238 4384 12406
rect 4712 12378 4764 12384
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11898 4200 12038
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3936 11784 4016 11812
rect 3884 11766 3936 11772
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2884 10130 2912 11630
rect 4356 11626 4384 12174
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11778 4476 12038
rect 4540 11898 4568 12174
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4724 11898 4752 12106
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4448 11750 4660 11778
rect 4816 11762 4844 12038
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5276 11898 5304 12174
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5368 11762 5396 12038
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 10130 4108 11018
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 11750
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4816 10810 4844 11562
rect 5368 11354 5396 11698
rect 5460 11694 5488 12378
rect 5540 12368 5592 12374
rect 5540 12310 5592 12316
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5460 11286 5488 11630
rect 5552 11558 5580 12310
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5644 11082 5672 16594
rect 6288 16250 6316 16594
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6472 16046 6500 21898
rect 6564 21078 6592 25894
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6656 25498 6684 25774
rect 6644 25492 6696 25498
rect 6644 25434 6696 25440
rect 6932 24313 6960 27610
rect 7208 27538 7236 30670
rect 7300 30598 7328 32438
rect 7944 31958 7972 32438
rect 8208 32428 8260 32434
rect 8208 32370 8260 32376
rect 7932 31952 7984 31958
rect 7932 31894 7984 31900
rect 8220 31822 8248 32370
rect 8312 31890 8340 32982
rect 8864 32570 8892 33934
rect 9680 33856 9732 33862
rect 9680 33798 9732 33804
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9496 33584 9548 33590
rect 9496 33526 9548 33532
rect 9128 32768 9180 32774
rect 9128 32710 9180 32716
rect 8484 32564 8536 32570
rect 8404 32524 8484 32552
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8208 31816 8260 31822
rect 8208 31758 8260 31764
rect 8024 31680 8076 31686
rect 8024 31622 8076 31628
rect 7656 31340 7708 31346
rect 7656 31282 7708 31288
rect 7668 30784 7696 31282
rect 7668 30756 7880 30784
rect 7852 30666 7880 30756
rect 7840 30660 7892 30666
rect 7840 30602 7892 30608
rect 7288 30592 7340 30598
rect 7288 30534 7340 30540
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 7300 29170 7328 29446
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7392 29034 7420 29106
rect 7380 29028 7432 29034
rect 7380 28970 7432 28976
rect 7576 28082 7604 29514
rect 7668 29238 7696 29582
rect 7656 29232 7708 29238
rect 7656 29174 7708 29180
rect 7668 28762 7696 29174
rect 7748 29164 7800 29170
rect 7748 29106 7800 29112
rect 7760 28762 7788 29106
rect 7656 28756 7708 28762
rect 7656 28698 7708 28704
rect 7748 28756 7800 28762
rect 7748 28698 7800 28704
rect 7668 28150 7696 28698
rect 7656 28144 7708 28150
rect 7656 28086 7708 28092
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7380 27940 7432 27946
rect 7380 27882 7432 27888
rect 7196 27532 7248 27538
rect 7196 27474 7248 27480
rect 7104 27328 7156 27334
rect 7104 27270 7156 27276
rect 7116 27130 7144 27270
rect 7104 27124 7156 27130
rect 7104 27066 7156 27072
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 7024 25294 7052 26182
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 7012 24880 7064 24886
rect 7116 24834 7144 26930
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7064 24828 7144 24834
rect 7012 24822 7144 24828
rect 7024 24806 7144 24822
rect 7116 24410 7144 24806
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 6918 24304 6974 24313
rect 6918 24239 6974 24248
rect 6828 24200 6880 24206
rect 6826 24168 6828 24177
rect 6880 24168 6882 24177
rect 6644 24132 6696 24138
rect 6826 24103 6882 24112
rect 6644 24074 6696 24080
rect 6656 23798 6684 24074
rect 7116 23798 7144 24346
rect 7208 24274 7236 25638
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7300 24410 7328 24686
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 6644 23792 6696 23798
rect 6644 23734 6696 23740
rect 7104 23792 7156 23798
rect 7156 23740 7236 23746
rect 7104 23734 7236 23740
rect 6656 22642 6684 23734
rect 7116 23718 7236 23734
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 7024 23186 7052 23598
rect 7208 23526 7236 23718
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6644 22160 6696 22166
rect 6644 22102 6696 22108
rect 6656 21418 6684 22102
rect 6748 22098 6776 22510
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6840 22030 6868 22646
rect 7300 22273 7328 22714
rect 7286 22264 7342 22273
rect 7286 22199 7342 22208
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6552 20528 6604 20534
rect 6552 20470 6604 20476
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 5920 15706 5948 15982
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6472 15502 6500 15846
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5736 14074 5764 14418
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 14074 6408 14350
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 5736 13326 5764 13874
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12306 5764 12854
rect 5920 12850 5948 13806
rect 6104 13530 6132 13874
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6380 13326 6408 14010
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5920 12220 5948 12786
rect 6104 12434 6132 13262
rect 6564 12434 6592 20470
rect 6656 20466 6684 21354
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7024 20942 7052 21082
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6656 19786 6684 20402
rect 6748 20330 6776 20470
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6840 19854 6868 20402
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6932 18970 6960 20402
rect 7024 20058 7052 20878
rect 7116 20534 7144 21490
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7208 20330 7236 20878
rect 7196 20324 7248 20330
rect 7196 20266 7248 20272
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7116 19922 7144 20198
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7024 18290 7052 19314
rect 7116 18766 7144 19654
rect 7300 18834 7328 22199
rect 7392 21010 7420 27882
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 7484 26994 7512 27474
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7576 27130 7604 27270
rect 7564 27124 7616 27130
rect 7760 27112 7788 28698
rect 7564 27066 7616 27072
rect 7668 27084 7788 27112
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7668 26926 7696 27084
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7656 26920 7708 26926
rect 7656 26862 7708 26868
rect 7668 26450 7696 26862
rect 7760 26586 7788 26930
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7656 26444 7708 26450
rect 7656 26386 7708 26392
rect 7668 25362 7696 26386
rect 7852 25945 7880 30602
rect 8036 30394 8064 31622
rect 8220 31346 8248 31758
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8220 30666 8248 31282
rect 8404 30870 8432 32524
rect 8484 32506 8536 32512
rect 8852 32564 8904 32570
rect 8852 32506 8904 32512
rect 8484 31884 8536 31890
rect 8484 31826 8536 31832
rect 8496 31210 8524 31826
rect 8760 31680 8812 31686
rect 8760 31622 8812 31628
rect 8484 31204 8536 31210
rect 8484 31146 8536 31152
rect 8392 30864 8444 30870
rect 8392 30806 8444 30812
rect 8208 30660 8260 30666
rect 8208 30602 8260 30608
rect 8024 30388 8076 30394
rect 8024 30330 8076 30336
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 8024 29776 8076 29782
rect 8024 29718 8076 29724
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 7944 27538 7972 29582
rect 8036 29306 8064 29718
rect 8128 29578 8156 29990
rect 8220 29714 8248 30602
rect 8496 30258 8524 31146
rect 8576 30864 8628 30870
rect 8576 30806 8628 30812
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 8312 29646 8340 30126
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8392 29640 8444 29646
rect 8392 29582 8444 29588
rect 8116 29572 8168 29578
rect 8116 29514 8168 29520
rect 8298 29336 8354 29345
rect 8024 29300 8076 29306
rect 8298 29271 8354 29280
rect 8024 29242 8076 29248
rect 8312 29170 8340 29271
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 8024 29028 8076 29034
rect 8024 28970 8076 28976
rect 8036 27674 8064 28970
rect 8404 28762 8432 29582
rect 8116 28756 8168 28762
rect 8116 28698 8168 28704
rect 8392 28756 8444 28762
rect 8392 28698 8444 28704
rect 8128 28558 8156 28698
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 8036 27130 8064 27610
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 8024 26784 8076 26790
rect 8128 26772 8156 27406
rect 8076 26744 8156 26772
rect 8024 26726 8076 26732
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7838 25936 7894 25945
rect 7838 25871 7894 25880
rect 7944 25702 7972 26318
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 8036 25226 8064 26386
rect 8220 26042 8248 27406
rect 8312 26450 8340 28494
rect 8496 28218 8524 30194
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8588 28098 8616 30806
rect 8772 30394 8800 31622
rect 8864 30598 8892 32506
rect 9140 31686 9168 32710
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9310 32328 9366 32337
rect 9310 32263 9312 32272
rect 9364 32263 9366 32272
rect 9312 32234 9364 32240
rect 9416 31686 9444 32370
rect 9508 32026 9536 33526
rect 9692 33114 9720 33798
rect 9784 33658 9812 33798
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 10152 33289 10180 33934
rect 10232 33856 10284 33862
rect 10232 33798 10284 33804
rect 10244 33454 10272 33798
rect 10232 33448 10284 33454
rect 10232 33390 10284 33396
rect 10138 33280 10194 33289
rect 10138 33215 10194 33224
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9588 32428 9640 32434
rect 9588 32370 9640 32376
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 9600 32026 9628 32370
rect 9680 32292 9732 32298
rect 9680 32234 9732 32240
rect 9496 32020 9548 32026
rect 9496 31962 9548 31968
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 9220 31680 9272 31686
rect 9220 31622 9272 31628
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9494 31648 9550 31657
rect 9232 31498 9260 31622
rect 9140 31470 9260 31498
rect 9310 31512 9366 31521
rect 9140 31385 9168 31470
rect 9310 31447 9366 31456
rect 9126 31376 9182 31385
rect 9324 31346 9352 31447
rect 9416 31362 9444 31622
rect 9494 31583 9550 31592
rect 9508 31482 9536 31583
rect 9496 31476 9548 31482
rect 9496 31418 9548 31424
rect 9126 31311 9182 31320
rect 9220 31340 9272 31346
rect 8944 31272 8996 31278
rect 8944 31214 8996 31220
rect 8956 30938 8984 31214
rect 9036 31136 9088 31142
rect 9036 31078 9088 31084
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 9048 30841 9076 31078
rect 9140 30870 9168 31311
rect 9220 31282 9272 31288
rect 9312 31340 9364 31346
rect 9416 31334 9536 31362
rect 9312 31282 9364 31288
rect 9232 31142 9260 31282
rect 9312 31204 9364 31210
rect 9312 31146 9364 31152
rect 9220 31136 9272 31142
rect 9220 31078 9272 31084
rect 9128 30864 9180 30870
rect 9034 30832 9090 30841
rect 9128 30806 9180 30812
rect 9034 30767 9090 30776
rect 9128 30728 9180 30734
rect 9128 30670 9180 30676
rect 8852 30592 8904 30598
rect 8852 30534 8904 30540
rect 8760 30388 8812 30394
rect 8760 30330 8812 30336
rect 8668 29640 8720 29646
rect 8668 29582 8720 29588
rect 8680 28966 8708 29582
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8392 28076 8444 28082
rect 8392 28018 8444 28024
rect 8496 28070 8616 28098
rect 8404 26586 8432 28018
rect 8496 27334 8524 28070
rect 8576 27464 8628 27470
rect 8576 27406 8628 27412
rect 8484 27328 8536 27334
rect 8484 27270 8536 27276
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8312 25906 8340 26386
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 8496 25786 8524 27270
rect 8588 26994 8616 27406
rect 8576 26988 8628 26994
rect 8680 26976 8708 28902
rect 8772 27538 8800 30330
rect 8852 30252 8904 30258
rect 8852 30194 8904 30200
rect 8864 28370 8892 30194
rect 9140 30054 9168 30670
rect 9232 30394 9260 31078
rect 9324 30938 9352 31146
rect 9312 30932 9364 30938
rect 9312 30874 9364 30880
rect 9220 30388 9272 30394
rect 9220 30330 9272 30336
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9128 30048 9180 30054
rect 9128 29990 9180 29996
rect 9416 29730 9444 30262
rect 9508 30258 9536 31334
rect 9600 30734 9628 31962
rect 9692 31958 9720 32234
rect 10048 32020 10100 32026
rect 10048 31962 10100 31968
rect 9680 31952 9732 31958
rect 9680 31894 9732 31900
rect 10060 31754 10088 31962
rect 10152 31754 10180 32370
rect 10048 31748 10100 31754
rect 10048 31690 10100 31696
rect 10140 31748 10192 31754
rect 10140 31690 10192 31696
rect 9770 31648 9826 31657
rect 10152 31634 10180 31690
rect 9826 31606 10180 31634
rect 9770 31583 9826 31592
rect 9784 30734 9812 31583
rect 10140 31408 10192 31414
rect 10140 31350 10192 31356
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 9968 31142 9996 31282
rect 9956 31136 10008 31142
rect 10008 31096 10088 31124
rect 9956 31078 10008 31084
rect 10060 30802 10088 31096
rect 10048 30796 10100 30802
rect 10048 30738 10100 30744
rect 9588 30728 9640 30734
rect 9588 30670 9640 30676
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9862 30696 9918 30705
rect 9680 30660 9732 30666
rect 9862 30631 9918 30640
rect 9956 30660 10008 30666
rect 9680 30602 9732 30608
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9496 30048 9548 30054
rect 9692 30036 9720 30602
rect 9548 30008 9720 30036
rect 9496 29990 9548 29996
rect 9048 29702 9444 29730
rect 9048 29306 9076 29702
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9126 29336 9182 29345
rect 9036 29300 9088 29306
rect 9182 29294 9260 29322
rect 9324 29306 9352 29582
rect 9126 29271 9182 29280
rect 9036 29242 9088 29248
rect 8944 29164 8996 29170
rect 9128 29164 9180 29170
rect 8944 29106 8996 29112
rect 9048 29124 9128 29152
rect 8956 28937 8984 29106
rect 8942 28928 8998 28937
rect 8942 28863 8998 28872
rect 9048 28490 9076 29124
rect 9128 29106 9180 29112
rect 9232 29034 9260 29294
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9404 29232 9456 29238
rect 9404 29174 9456 29180
rect 9220 29028 9272 29034
rect 9416 28994 9444 29174
rect 9220 28970 9272 28976
rect 9324 28966 9444 28994
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 8864 28342 9076 28370
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8956 27674 8984 28018
rect 8852 27668 8904 27674
rect 8852 27610 8904 27616
rect 8944 27668 8996 27674
rect 8944 27610 8996 27616
rect 8760 27532 8812 27538
rect 8760 27474 8812 27480
rect 8864 27334 8892 27610
rect 8852 27328 8904 27334
rect 8852 27270 8904 27276
rect 8760 26988 8812 26994
rect 8680 26948 8760 26976
rect 8576 26930 8628 26936
rect 8760 26930 8812 26936
rect 8850 26888 8906 26897
rect 8850 26823 8906 26832
rect 8864 26790 8892 26823
rect 8852 26784 8904 26790
rect 8852 26726 8904 26732
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8312 25758 8524 25786
rect 8208 25356 8260 25362
rect 8208 25298 8260 25304
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 8116 25220 8168 25226
rect 8116 25162 8168 25168
rect 7748 25152 7800 25158
rect 7746 25120 7748 25129
rect 7840 25152 7892 25158
rect 7800 25120 7802 25129
rect 7840 25094 7892 25100
rect 7746 25055 7802 25064
rect 7852 24614 7880 25094
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7564 23180 7616 23186
rect 7564 23122 7616 23128
rect 7576 22778 7604 23122
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7656 22704 7708 22710
rect 7654 22672 7656 22681
rect 7708 22672 7710 22681
rect 7654 22607 7710 22616
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7484 22166 7512 22442
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7668 22098 7696 22374
rect 7760 22098 7788 23530
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7484 21146 7512 21966
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7378 20904 7434 20913
rect 7378 20839 7434 20848
rect 7392 20806 7420 20839
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7470 20632 7526 20641
rect 7576 20602 7604 21966
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7470 20567 7526 20576
rect 7564 20596 7616 20602
rect 7484 20534 7512 20567
rect 7564 20538 7616 20544
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18426 7144 18566
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6656 17338 6684 18226
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17814 6868 18158
rect 6828 17808 6880 17814
rect 6828 17750 6880 17756
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 7024 16182 7052 18226
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7300 17882 7328 18158
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7116 16794 7144 17818
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6932 15570 6960 15982
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6748 13462 6776 14962
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6104 12406 6224 12434
rect 6564 12406 6776 12434
rect 6092 12232 6144 12238
rect 5920 12192 6092 12220
rect 6092 12174 6144 12180
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 11354 5856 11562
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5920 11014 5948 11494
rect 6104 11150 6132 12174
rect 6196 11558 6224 12406
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5920 10742 5948 10950
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5906 10160 5962 10169
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4620 10124 4672 10130
rect 5906 10095 5962 10104
rect 4620 10066 4672 10072
rect 4080 9518 4108 10066
rect 5920 10062 5948 10095
rect 5724 10056 5776 10062
rect 5908 10056 5960 10062
rect 5776 10016 5856 10044
rect 5724 9998 5776 10004
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 8974 4108 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 938 4176 994 4185
rect 4080 4146 4108 8910
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4816 8634 4844 8842
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5736 8430 5764 9862
rect 5828 9586 5856 10016
rect 5908 9998 5960 10004
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9042 5856 9522
rect 5920 9178 5948 9998
rect 6012 9926 6040 10746
rect 6288 10266 6316 11290
rect 6472 11150 6500 11630
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6564 10674 6592 12038
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6656 10674 6684 11222
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6564 10266 6592 10610
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6092 10192 6144 10198
rect 6090 10160 6092 10169
rect 6748 10169 6776 12406
rect 6840 10962 6868 14418
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12782 6960 13126
rect 7024 12850 7052 16118
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7116 14618 7144 16050
rect 7208 15162 7236 17546
rect 7300 17202 7328 17682
rect 7392 17610 7420 18158
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7484 16454 7512 20470
rect 7760 20058 7788 20946
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7852 18970 7880 24210
rect 8036 24206 8064 24550
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 23254 8064 23462
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 8024 22976 8076 22982
rect 8024 22918 8076 22924
rect 7932 22704 7984 22710
rect 7932 22646 7984 22652
rect 7944 22438 7972 22646
rect 8036 22642 8064 22918
rect 8128 22778 8156 25162
rect 8220 24750 8248 25298
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8220 23118 8248 23462
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8312 22778 8340 25758
rect 8482 25528 8538 25537
rect 8482 25463 8538 25472
rect 8496 25430 8524 25463
rect 8484 25424 8536 25430
rect 8484 25366 8536 25372
rect 8390 24848 8446 24857
rect 8390 24783 8446 24792
rect 8404 24342 8432 24783
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8392 24336 8444 24342
rect 8392 24278 8444 24284
rect 8496 24138 8524 24550
rect 8588 24177 8616 26318
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 8852 26240 8904 26246
rect 8852 26182 8904 26188
rect 8758 26072 8814 26081
rect 8758 26007 8814 26016
rect 8772 25906 8800 26007
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8668 25764 8720 25770
rect 8668 25706 8720 25712
rect 8574 24168 8630 24177
rect 8484 24132 8536 24138
rect 8574 24103 8630 24112
rect 8484 24074 8536 24080
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 23526 8432 24006
rect 8680 23866 8708 25706
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 22982 8432 23462
rect 8864 23186 8892 26182
rect 8956 25430 8984 26250
rect 8944 25424 8996 25430
rect 8944 25366 8996 25372
rect 9048 25242 9076 28342
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 9232 25809 9260 26454
rect 9324 26314 9352 28966
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9416 26518 9444 27270
rect 9404 26512 9456 26518
rect 9404 26454 9456 26460
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9324 25838 9352 26250
rect 9312 25832 9364 25838
rect 9218 25800 9274 25809
rect 9312 25774 9364 25780
rect 9218 25735 9274 25744
rect 8956 25214 9076 25242
rect 9128 25288 9180 25294
rect 9128 25230 9180 25236
rect 8852 23180 8904 23186
rect 8852 23122 8904 23128
rect 8956 23066 8984 25214
rect 9036 24948 9088 24954
rect 9036 24890 9088 24896
rect 8772 23038 8984 23066
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8484 22704 8536 22710
rect 8484 22646 8536 22652
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 8036 22234 8064 22578
rect 8024 22228 8076 22234
rect 8024 22170 8076 22176
rect 8300 22228 8352 22234
rect 8300 22170 8352 22176
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21690 7972 21830
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 8312 21554 8340 22170
rect 8496 22166 8524 22646
rect 8484 22160 8536 22166
rect 8484 22102 8536 22108
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8022 21176 8078 21185
rect 8022 21111 8024 21120
rect 8076 21111 8078 21120
rect 8024 21082 8076 21088
rect 8312 21010 8340 21490
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8024 20800 8076 20806
rect 8024 20742 8076 20748
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8036 20602 8064 20742
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 8036 19922 8064 20538
rect 8220 20398 8248 20742
rect 8312 20534 8340 20946
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8128 19922 8156 20266
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8312 18970 8340 19722
rect 8484 19508 8536 19514
rect 8484 19450 8536 19456
rect 8392 19236 8444 19242
rect 8392 19178 8444 19184
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8404 18834 8432 19178
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 7472 16448 7524 16454
rect 7472 16390 7524 16396
rect 7484 16250 7512 16390
rect 7576 16250 7604 18770
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8128 17746 8156 18702
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 16726 8064 17138
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 8036 16454 8064 16662
rect 8220 16538 8248 18362
rect 8128 16510 8248 16538
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7760 15570 7788 16390
rect 8036 16114 8064 16390
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7196 15156 7248 15162
rect 7472 15156 7524 15162
rect 7196 15098 7248 15104
rect 7392 15116 7472 15144
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7208 14482 7236 14962
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7208 12918 7236 14418
rect 7392 13938 7420 15116
rect 7472 15098 7524 15104
rect 7668 14482 7696 15302
rect 7760 15162 7788 15506
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7840 14952 7892 14958
rect 8024 14952 8076 14958
rect 7840 14894 7892 14900
rect 8022 14920 8024 14929
rect 8076 14920 8078 14929
rect 7852 14618 7880 14894
rect 7932 14884 7984 14890
rect 8022 14855 8078 14864
rect 7932 14826 7984 14832
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7484 13938 7512 14282
rect 7668 13938 7696 14418
rect 7944 13938 7972 14826
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14006 8064 14758
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7024 12306 7052 12786
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6932 11218 6960 12106
rect 7484 11762 7512 12718
rect 7576 12306 7604 12718
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 11898 7604 12106
rect 7668 11898 7696 12854
rect 8128 12850 8156 16510
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 15638 8248 16390
rect 8496 16114 8524 19450
rect 8588 18970 8616 20402
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8680 18630 8708 22918
rect 8772 22094 8800 23038
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 8772 22066 8892 22094
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8772 21894 8800 21966
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8772 21554 8800 21830
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8772 21010 8800 21490
rect 8760 21004 8812 21010
rect 8760 20946 8812 20952
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 8772 20466 8800 20810
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8772 18970 8800 19246
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 17542 8708 18566
rect 8772 18086 8800 18702
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8772 17746 8800 18022
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8864 17338 8892 22066
rect 8956 17338 8984 22714
rect 9048 21010 9076 24890
rect 9140 24682 9168 25230
rect 9232 24834 9260 25735
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9324 25498 9352 25638
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 9232 24806 9352 24834
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9128 24676 9180 24682
rect 9128 24618 9180 24624
rect 9232 23798 9260 24686
rect 9220 23792 9272 23798
rect 9220 23734 9272 23740
rect 9128 23724 9180 23730
rect 9128 23666 9180 23672
rect 9140 21622 9168 23666
rect 9220 23656 9272 23662
rect 9218 23624 9220 23633
rect 9272 23624 9274 23633
rect 9218 23559 9274 23568
rect 9232 22930 9260 23559
rect 9324 23050 9352 24806
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9232 22902 9352 22930
rect 9324 22166 9352 22902
rect 9416 22778 9444 23054
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9312 22160 9364 22166
rect 9312 22102 9364 22108
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9128 21616 9180 21622
rect 9232 21593 9260 21898
rect 9416 21894 9444 21966
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9128 21558 9180 21564
rect 9218 21584 9274 21593
rect 9508 21570 9536 29990
rect 9680 29844 9732 29850
rect 9680 29786 9732 29792
rect 9588 29164 9640 29170
rect 9588 29106 9640 29112
rect 9600 29073 9628 29106
rect 9586 29064 9642 29073
rect 9586 28999 9642 29008
rect 9692 28665 9720 29786
rect 9770 29608 9826 29617
rect 9770 29543 9826 29552
rect 9678 28656 9734 28665
rect 9678 28591 9734 28600
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9600 24954 9628 28494
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9692 28218 9720 28426
rect 9784 28422 9812 29543
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 9784 28098 9812 28358
rect 9692 28070 9812 28098
rect 9692 25922 9720 28070
rect 9770 27568 9826 27577
rect 9770 27503 9826 27512
rect 9784 26382 9812 27503
rect 9876 26586 9904 30631
rect 10152 30648 10180 31350
rect 10008 30620 10180 30648
rect 9956 30602 10008 30608
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 10060 29782 10088 30194
rect 10140 30116 10192 30122
rect 10140 30058 10192 30064
rect 10048 29776 10100 29782
rect 10048 29718 10100 29724
rect 10152 29510 10180 30058
rect 10140 29504 10192 29510
rect 10140 29446 10192 29452
rect 10244 29306 10272 33390
rect 10336 32502 10364 39039
rect 10980 37262 11008 39039
rect 11624 37262 11652 39039
rect 12268 37262 12296 39039
rect 12912 38978 12940 39039
rect 13004 38978 13032 39086
rect 12912 38950 13032 38978
rect 10968 37256 11020 37262
rect 10968 37198 11020 37204
rect 11612 37256 11664 37262
rect 11612 37198 11664 37204
rect 12256 37256 12308 37262
rect 12256 37198 12308 37204
rect 10784 37188 10836 37194
rect 10784 37130 10836 37136
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 10612 36242 10640 37062
rect 10692 36712 10744 36718
rect 10692 36654 10744 36660
rect 10600 36236 10652 36242
rect 10600 36178 10652 36184
rect 10600 36100 10652 36106
rect 10704 36088 10732 36654
rect 10652 36060 10732 36088
rect 10600 36042 10652 36048
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10324 32496 10376 32502
rect 10324 32438 10376 32444
rect 10324 32360 10376 32366
rect 10324 32302 10376 32308
rect 10336 31822 10364 32302
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10428 31822 10456 32166
rect 10324 31816 10376 31822
rect 10324 31758 10376 31764
rect 10416 31816 10468 31822
rect 10416 31758 10468 31764
rect 10336 30666 10364 31758
rect 10520 31668 10548 34478
rect 10612 31793 10640 36042
rect 10690 35048 10746 35057
rect 10796 35034 10824 37130
rect 10876 37120 10928 37126
rect 10876 37062 10928 37068
rect 10746 35006 10824 35034
rect 10690 34983 10746 34992
rect 10704 33114 10732 34983
rect 10888 34474 10916 37062
rect 10980 36854 11008 37198
rect 10968 36848 11020 36854
rect 11624 36836 11652 37198
rect 11888 37120 11940 37126
rect 11888 37062 11940 37068
rect 11900 36854 11928 37062
rect 11888 36848 11940 36854
rect 11624 36808 11744 36836
rect 10968 36790 11020 36796
rect 11716 36310 11744 36808
rect 11888 36790 11940 36796
rect 12164 36848 12216 36854
rect 12164 36790 12216 36796
rect 11704 36304 11756 36310
rect 11704 36246 11756 36252
rect 12176 36174 12204 36790
rect 12268 36718 12296 37198
rect 12348 37120 12400 37126
rect 12348 37062 12400 37068
rect 12256 36712 12308 36718
rect 12256 36654 12308 36660
rect 12360 36564 12388 37062
rect 12268 36536 12388 36564
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 12164 35692 12216 35698
rect 12164 35634 12216 35640
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 11612 35148 11664 35154
rect 11612 35090 11664 35096
rect 11532 34746 11560 35090
rect 11520 34740 11572 34746
rect 11520 34682 11572 34688
rect 11060 34536 11112 34542
rect 11060 34478 11112 34484
rect 10876 34468 10928 34474
rect 10876 34410 10928 34416
rect 10888 34134 10916 34410
rect 10876 34128 10928 34134
rect 10876 34070 10928 34076
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10692 33108 10744 33114
rect 10692 33050 10744 33056
rect 10796 33096 10824 33934
rect 10888 33590 10916 34070
rect 11072 33658 11100 34478
rect 11624 33998 11652 35090
rect 12176 35057 12204 35634
rect 12268 35630 12296 36536
rect 13268 36304 13320 36310
rect 13268 36246 13320 36252
rect 12624 36168 12676 36174
rect 12624 36110 12676 36116
rect 12532 35692 12584 35698
rect 12452 35652 12532 35680
rect 12256 35624 12308 35630
rect 12256 35566 12308 35572
rect 12268 35154 12296 35566
rect 12256 35148 12308 35154
rect 12256 35090 12308 35096
rect 12348 35080 12400 35086
rect 12162 35048 12218 35057
rect 12348 35022 12400 35028
rect 12162 34983 12218 34992
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11796 34944 11848 34950
rect 11796 34886 11848 34892
rect 11716 34678 11744 34886
rect 11704 34672 11756 34678
rect 11704 34614 11756 34620
rect 11808 34610 11836 34886
rect 12360 34610 12388 35022
rect 12452 35018 12480 35652
rect 12532 35634 12584 35640
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12440 35012 12492 35018
rect 12440 34954 12492 34960
rect 11796 34604 11848 34610
rect 11796 34546 11848 34552
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 12348 34604 12400 34610
rect 12348 34546 12400 34552
rect 11900 34406 11928 34546
rect 11888 34400 11940 34406
rect 11808 34360 11888 34388
rect 11612 33992 11664 33998
rect 11164 33930 11376 33946
rect 11612 33934 11664 33940
rect 11164 33924 11388 33930
rect 11164 33918 11336 33924
rect 11060 33652 11112 33658
rect 11060 33594 11112 33600
rect 10876 33584 10928 33590
rect 10876 33526 10928 33532
rect 11072 33522 11100 33594
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10968 33312 11020 33318
rect 10968 33254 11020 33260
rect 10876 33108 10928 33114
rect 10796 33068 10876 33096
rect 10598 31784 10654 31793
rect 10598 31719 10654 31728
rect 10428 31640 10548 31668
rect 10324 30660 10376 30666
rect 10324 30602 10376 30608
rect 10324 29640 10376 29646
rect 10322 29608 10324 29617
rect 10376 29608 10378 29617
rect 10322 29543 10378 29552
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10324 29300 10376 29306
rect 10324 29242 10376 29248
rect 10336 29186 10364 29242
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 10152 29158 10364 29186
rect 10060 29073 10088 29106
rect 10152 29102 10180 29158
rect 10140 29096 10192 29102
rect 10046 29064 10102 29073
rect 10140 29038 10192 29044
rect 10046 28999 10102 29008
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 10244 28937 10272 28970
rect 10324 28960 10376 28966
rect 10230 28928 10286 28937
rect 10324 28902 10376 28908
rect 10230 28863 10286 28872
rect 10232 28688 10284 28694
rect 10230 28656 10232 28665
rect 10284 28656 10286 28665
rect 10230 28591 10286 28600
rect 10232 28484 10284 28490
rect 10232 28426 10284 28432
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 10048 27532 10100 27538
rect 10048 27474 10100 27480
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9968 26994 9996 27406
rect 10060 27305 10088 27474
rect 10046 27296 10102 27305
rect 10046 27231 10102 27240
rect 10046 27160 10102 27169
rect 10046 27095 10102 27104
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9968 26586 9996 26930
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 9772 26376 9824 26382
rect 9772 26318 9824 26324
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9784 26042 9812 26182
rect 9772 26036 9824 26042
rect 9772 25978 9824 25984
rect 9692 25894 9812 25922
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9678 24848 9734 24857
rect 9784 24818 9812 25894
rect 9876 25498 9904 26318
rect 9956 26308 10008 26314
rect 9956 26250 10008 26256
rect 9968 26217 9996 26250
rect 9954 26208 10010 26217
rect 9954 26143 10010 26152
rect 9956 25900 10008 25906
rect 9956 25842 10008 25848
rect 9864 25492 9916 25498
rect 9864 25434 9916 25440
rect 9968 25294 9996 25842
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9678 24783 9680 24792
rect 9732 24783 9734 24792
rect 9772 24812 9824 24818
rect 9680 24754 9732 24760
rect 9772 24754 9824 24760
rect 9692 23866 9720 24754
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9678 23352 9734 23361
rect 9784 23322 9812 24142
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9876 23594 9904 24074
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9678 23287 9680 23296
rect 9732 23287 9734 23296
rect 9772 23316 9824 23322
rect 9680 23258 9732 23264
rect 9772 23258 9824 23264
rect 9876 22574 9904 23530
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9600 22030 9628 22170
rect 9876 22166 9904 22510
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9218 21519 9220 21528
rect 9272 21519 9274 21528
rect 9312 21548 9364 21554
rect 9220 21490 9272 21496
rect 9312 21490 9364 21496
rect 9416 21542 9536 21570
rect 9036 21004 9088 21010
rect 9036 20946 9088 20952
rect 9232 20942 9260 21490
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9324 20806 9352 21490
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 9048 18358 9076 19722
rect 9416 19666 9444 21542
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 9600 20806 9628 21354
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9508 20534 9536 20742
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 9600 20262 9628 20742
rect 9784 20466 9812 21626
rect 9876 21457 9904 21966
rect 9968 21622 9996 25230
rect 10060 25208 10088 27095
rect 10152 26897 10180 27950
rect 10244 26994 10272 28426
rect 10336 28422 10364 28902
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10322 27704 10378 27713
rect 10322 27639 10378 27648
rect 10336 27470 10364 27639
rect 10428 27606 10456 31640
rect 10506 31376 10562 31385
rect 10506 31311 10508 31320
rect 10560 31311 10562 31320
rect 10508 31282 10560 31288
rect 10704 29850 10732 33050
rect 10796 32026 10824 33068
rect 10876 33050 10928 33056
rect 10888 33017 10916 33050
rect 10874 33008 10930 33017
rect 10980 32994 11008 33254
rect 11072 33114 11100 33458
rect 11164 33386 11192 33918
rect 11336 33866 11388 33872
rect 11244 33856 11296 33862
rect 11244 33798 11296 33804
rect 11152 33380 11204 33386
rect 11152 33322 11204 33328
rect 11256 33114 11284 33798
rect 11520 33584 11572 33590
rect 11348 33532 11520 33538
rect 11348 33526 11572 33532
rect 11348 33522 11560 33526
rect 11336 33516 11560 33522
rect 11388 33510 11560 33516
rect 11336 33458 11388 33464
rect 11808 33318 11836 34360
rect 11888 34342 11940 34348
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 12072 33992 12124 33998
rect 12072 33934 12124 33940
rect 11900 33386 11928 33934
rect 11980 33924 12032 33930
rect 11980 33866 12032 33872
rect 11992 33538 12020 33866
rect 12084 33658 12112 33934
rect 12360 33930 12388 34546
rect 12452 34202 12480 34954
rect 12544 34474 12572 35226
rect 12636 35086 12664 36110
rect 12898 35864 12954 35873
rect 12898 35799 12900 35808
rect 12952 35799 12954 35808
rect 13176 35828 13228 35834
rect 12900 35770 12952 35776
rect 13176 35770 13228 35776
rect 12992 35692 13044 35698
rect 13188 35680 13216 35770
rect 13044 35652 13216 35680
rect 12992 35634 13044 35640
rect 12808 35488 12860 35494
rect 12714 35456 12770 35465
rect 12808 35430 12860 35436
rect 12714 35391 12770 35400
rect 12728 35290 12756 35391
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 12624 35080 12676 35086
rect 12622 35048 12624 35057
rect 12676 35048 12678 35057
rect 12622 34983 12678 34992
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12728 34678 12756 34886
rect 12716 34672 12768 34678
rect 12716 34614 12768 34620
rect 12820 34610 12848 35430
rect 13004 35290 13032 35634
rect 12992 35284 13044 35290
rect 12992 35226 13044 35232
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 12900 34944 12952 34950
rect 12900 34886 12952 34892
rect 12912 34746 12940 34886
rect 13004 34746 13032 35022
rect 12900 34740 12952 34746
rect 12900 34682 12952 34688
rect 12992 34740 13044 34746
rect 12992 34682 13044 34688
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12532 34468 12584 34474
rect 12532 34410 12584 34416
rect 12624 34400 12676 34406
rect 12624 34342 12676 34348
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12348 33924 12400 33930
rect 12348 33866 12400 33872
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 12636 33590 12664 34342
rect 12624 33584 12676 33590
rect 11992 33510 12112 33538
rect 12624 33526 12676 33532
rect 11888 33380 11940 33386
rect 11888 33322 11940 33328
rect 11796 33312 11848 33318
rect 11796 33254 11848 33260
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 11244 33108 11296 33114
rect 11244 33050 11296 33056
rect 10980 32966 11468 32994
rect 10874 32943 10930 32952
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10782 31512 10838 31521
rect 10782 31447 10838 31456
rect 10796 31414 10824 31447
rect 10784 31408 10836 31414
rect 10784 31350 10836 31356
rect 10796 30870 10824 31350
rect 10784 30864 10836 30870
rect 10784 30806 10836 30812
rect 10888 30258 10916 32846
rect 11060 32836 11112 32842
rect 11060 32778 11112 32784
rect 11072 32570 11100 32778
rect 11060 32564 11112 32570
rect 11060 32506 11112 32512
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 11244 32428 11296 32434
rect 11244 32370 11296 32376
rect 10966 31784 11022 31793
rect 11072 31754 11100 32370
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11164 31890 11192 32166
rect 11256 31906 11284 32370
rect 11336 32292 11388 32298
rect 11336 32234 11388 32240
rect 11348 32026 11376 32234
rect 11336 32020 11388 32026
rect 11336 31962 11388 31968
rect 11152 31884 11204 31890
rect 11256 31878 11376 31906
rect 11152 31826 11204 31832
rect 10966 31719 11022 31728
rect 11060 31748 11112 31754
rect 10980 30938 11008 31719
rect 11060 31690 11112 31696
rect 11072 31346 11100 31690
rect 11060 31340 11112 31346
rect 11060 31282 11112 31288
rect 10968 30932 11020 30938
rect 10968 30874 11020 30880
rect 11164 30734 11192 31826
rect 11348 31414 11376 31878
rect 11336 31408 11388 31414
rect 11336 31350 11388 31356
rect 11244 31340 11296 31346
rect 11244 31282 11296 31288
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 11164 30394 11192 30670
rect 11256 30598 11284 31282
rect 11244 30592 11296 30598
rect 11242 30560 11244 30569
rect 11296 30560 11298 30569
rect 11242 30495 11298 30504
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11440 30297 11468 32966
rect 11808 32570 11836 33254
rect 11796 32564 11848 32570
rect 11796 32506 11848 32512
rect 11520 32428 11572 32434
rect 11704 32428 11756 32434
rect 11572 32388 11652 32416
rect 11520 32370 11572 32376
rect 11520 31884 11572 31890
rect 11520 31826 11572 31832
rect 11532 31414 11560 31826
rect 11624 31822 11652 32388
rect 11704 32370 11756 32376
rect 11612 31816 11664 31822
rect 11612 31758 11664 31764
rect 11624 31414 11652 31758
rect 11716 31754 11744 32370
rect 11980 32360 12032 32366
rect 11980 32302 12032 32308
rect 11992 32026 12020 32302
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 12084 31906 12112 33510
rect 12348 33516 12400 33522
rect 12348 33458 12400 33464
rect 11992 31878 12112 31906
rect 11716 31726 11836 31754
rect 11520 31408 11572 31414
rect 11520 31350 11572 31356
rect 11612 31408 11664 31414
rect 11612 31350 11664 31356
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11716 30433 11744 30874
rect 11702 30424 11758 30433
rect 11702 30359 11758 30368
rect 11426 30288 11482 30297
rect 10876 30252 10928 30258
rect 11426 30223 11482 30232
rect 10876 30194 10928 30200
rect 11808 30054 11836 31726
rect 11888 31680 11940 31686
rect 11888 31622 11940 31628
rect 11900 31482 11928 31622
rect 11888 31476 11940 31482
rect 11888 31418 11940 31424
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11900 30938 11928 31282
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 11796 30048 11848 30054
rect 11796 29990 11848 29996
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10520 28082 10548 29582
rect 10600 29572 10652 29578
rect 10600 29514 10652 29520
rect 10612 29170 10640 29514
rect 10888 29170 10916 29582
rect 10968 29572 11020 29578
rect 10968 29514 11020 29520
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 10416 27464 10468 27470
rect 10416 27406 10468 27412
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10336 27062 10364 27270
rect 10324 27056 10376 27062
rect 10324 26998 10376 27004
rect 10232 26988 10284 26994
rect 10232 26930 10284 26936
rect 10138 26888 10194 26897
rect 10138 26823 10194 26832
rect 10244 25974 10272 26930
rect 10322 26888 10378 26897
rect 10322 26823 10378 26832
rect 10336 26234 10364 26823
rect 10428 26382 10456 27406
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10336 26206 10456 26234
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10232 25968 10284 25974
rect 10232 25910 10284 25916
rect 10140 25764 10192 25770
rect 10192 25724 10272 25752
rect 10140 25706 10192 25712
rect 10244 25294 10272 25724
rect 10336 25362 10364 25978
rect 10428 25838 10456 26206
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10232 25288 10284 25294
rect 10428 25242 10456 25774
rect 10232 25230 10284 25236
rect 10140 25220 10192 25226
rect 10060 25180 10140 25208
rect 10060 24954 10088 25180
rect 10140 25162 10192 25168
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 10060 24070 10088 24890
rect 10244 24750 10272 25230
rect 10336 25214 10456 25242
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 10140 24336 10192 24342
rect 10138 24304 10140 24313
rect 10192 24304 10194 24313
rect 10138 24239 10194 24248
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 10060 23225 10088 24006
rect 10152 23866 10180 24142
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 10152 23254 10180 23530
rect 10140 23248 10192 23254
rect 10046 23216 10102 23225
rect 10140 23190 10192 23196
rect 10046 23151 10048 23160
rect 10100 23151 10102 23160
rect 10048 23122 10100 23128
rect 10244 23118 10272 24686
rect 10336 24342 10364 25214
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10324 24336 10376 24342
rect 10324 24278 10376 24284
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10336 23866 10364 24142
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10322 23760 10378 23769
rect 10322 23695 10378 23704
rect 10140 23112 10192 23118
rect 10046 23080 10102 23089
rect 10140 23054 10192 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10046 23015 10048 23024
rect 10100 23015 10102 23024
rect 10048 22986 10100 22992
rect 10152 22794 10180 23054
rect 10244 22982 10272 23054
rect 10232 22976 10284 22982
rect 10232 22918 10284 22924
rect 10152 22766 10272 22794
rect 10244 22642 10272 22766
rect 10232 22636 10284 22642
rect 10232 22578 10284 22584
rect 10336 22438 10364 23695
rect 10428 23662 10456 24550
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 9862 21448 9918 21457
rect 9862 21383 9918 21392
rect 9876 20942 9904 21383
rect 10060 21049 10088 21966
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10152 21570 10180 21830
rect 10152 21542 10272 21570
rect 10244 21350 10272 21542
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10046 21040 10102 21049
rect 10244 21010 10272 21286
rect 10046 20975 10102 20984
rect 10232 21004 10284 21010
rect 10060 20942 10088 20975
rect 10232 20946 10284 20952
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9678 20088 9734 20097
rect 9678 20023 9734 20032
rect 9692 19990 9720 20023
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 10048 19712 10100 19718
rect 9416 19638 9536 19666
rect 10048 19654 10100 19660
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9416 18834 9444 19450
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9508 18358 9536 19638
rect 10060 19446 10088 19654
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 10336 19310 10364 22374
rect 10428 20913 10456 23598
rect 10520 21146 10548 28018
rect 10612 27470 10640 29106
rect 10784 29096 10836 29102
rect 10690 29064 10746 29073
rect 10784 29038 10836 29044
rect 10690 28999 10692 29008
rect 10744 28999 10746 29008
rect 10692 28970 10744 28976
rect 10796 28626 10824 29038
rect 10784 28620 10836 28626
rect 10784 28562 10836 28568
rect 10692 28144 10744 28150
rect 10692 28086 10744 28092
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10704 27130 10732 28086
rect 10784 27464 10836 27470
rect 10888 27452 10916 29106
rect 10980 29102 11008 29514
rect 10968 29096 11020 29102
rect 10968 29038 11020 29044
rect 10980 27538 11008 29038
rect 11072 28150 11100 29650
rect 11244 29572 11296 29578
rect 11244 29514 11296 29520
rect 11256 29238 11284 29514
rect 11336 29504 11388 29510
rect 11336 29446 11388 29452
rect 11348 29238 11376 29446
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11244 29232 11296 29238
rect 11244 29174 11296 29180
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 11520 29164 11572 29170
rect 11520 29106 11572 29112
rect 11244 28688 11296 28694
rect 11532 28665 11560 29106
rect 11244 28630 11296 28636
rect 11518 28656 11574 28665
rect 11152 28620 11204 28626
rect 11152 28562 11204 28568
rect 11060 28144 11112 28150
rect 11060 28086 11112 28092
rect 11164 28014 11192 28562
rect 11256 28082 11284 28630
rect 11518 28591 11520 28600
rect 11572 28591 11574 28600
rect 11520 28562 11572 28568
rect 11624 28490 11652 29242
rect 11808 29073 11836 29990
rect 11888 29096 11940 29102
rect 11794 29064 11850 29073
rect 11888 29038 11940 29044
rect 11794 28999 11850 29008
rect 11900 28558 11928 29038
rect 11888 28552 11940 28558
rect 11888 28494 11940 28500
rect 11520 28484 11572 28490
rect 11520 28426 11572 28432
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11428 28416 11480 28422
rect 11428 28358 11480 28364
rect 11244 28076 11296 28082
rect 11244 28018 11296 28024
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 10968 27532 11020 27538
rect 10968 27474 11020 27480
rect 10836 27424 10916 27452
rect 10784 27406 10836 27412
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10704 26897 10732 26930
rect 10690 26888 10746 26897
rect 10690 26823 10746 26832
rect 10796 26466 10824 27406
rect 10980 27169 11008 27474
rect 11152 27396 11204 27402
rect 11152 27338 11204 27344
rect 10966 27160 11022 27169
rect 10876 27124 10928 27130
rect 10966 27095 11022 27104
rect 10876 27066 10928 27072
rect 10704 26438 10824 26466
rect 10600 26240 10652 26246
rect 10600 26182 10652 26188
rect 10612 25650 10640 26182
rect 10704 25770 10732 26438
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 10796 25974 10824 26318
rect 10784 25968 10836 25974
rect 10784 25910 10836 25916
rect 10888 25906 10916 27066
rect 11164 26994 11192 27338
rect 11152 26988 11204 26994
rect 11152 26930 11204 26936
rect 11164 26897 11192 26930
rect 11150 26888 11206 26897
rect 11256 26874 11284 27814
rect 11336 27464 11388 27470
rect 11336 27406 11388 27412
rect 11348 27062 11376 27406
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11256 26858 11376 26874
rect 11256 26852 11388 26858
rect 11256 26846 11336 26852
rect 11150 26823 11206 26832
rect 11336 26794 11388 26800
rect 11060 26784 11112 26790
rect 10966 26752 11022 26761
rect 11244 26784 11296 26790
rect 11060 26726 11112 26732
rect 11150 26752 11206 26761
rect 10966 26687 11022 26696
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10692 25764 10744 25770
rect 10692 25706 10744 25712
rect 10612 25622 10732 25650
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 10612 25158 10640 25434
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10612 23730 10640 24006
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10612 22778 10640 23666
rect 10600 22772 10652 22778
rect 10600 22714 10652 22720
rect 10612 21962 10640 22714
rect 10704 22624 10732 25622
rect 10782 25528 10838 25537
rect 10782 25463 10838 25472
rect 10796 25158 10824 25463
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10888 24970 10916 25842
rect 10796 24942 10916 24970
rect 10796 24070 10824 24942
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10782 23216 10838 23225
rect 10782 23151 10838 23160
rect 10796 23118 10824 23151
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10704 22596 10824 22624
rect 10692 22500 10744 22506
rect 10692 22442 10744 22448
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10704 21690 10732 22442
rect 10796 22438 10824 22596
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10888 22386 10916 24210
rect 10980 22506 11008 26687
rect 11072 26489 11100 26726
rect 11244 26726 11296 26732
rect 11150 26687 11206 26696
rect 11058 26480 11114 26489
rect 11058 26415 11114 26424
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 11072 23594 11100 26250
rect 11164 26246 11192 26687
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11256 26042 11284 26726
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 11164 25226 11192 25774
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 11072 22574 11100 23530
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 11060 22432 11112 22438
rect 10888 22358 11008 22386
rect 11060 22374 11112 22380
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10888 21622 10916 21966
rect 10876 21616 10928 21622
rect 10598 21584 10654 21593
rect 10876 21558 10928 21564
rect 10598 21519 10600 21528
rect 10652 21519 10654 21528
rect 10600 21490 10652 21496
rect 10600 21412 10652 21418
rect 10600 21354 10652 21360
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10520 21010 10548 21082
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10414 20904 10470 20913
rect 10414 20839 10416 20848
rect 10468 20839 10470 20848
rect 10416 20810 10468 20816
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 19514 10456 19790
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10416 18896 10468 18902
rect 10414 18864 10416 18873
rect 10468 18864 10470 18873
rect 10414 18799 10470 18808
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9496 18352 9548 18358
rect 9496 18294 9548 18300
rect 9784 18057 9812 18634
rect 9968 18222 9996 18634
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9770 18048 9826 18057
rect 9770 17983 9826 17992
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16590 8616 16934
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8220 14414 8248 15574
rect 8312 15502 8340 15846
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 13802 8248 14214
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8312 12850 8340 15438
rect 8404 15366 8432 15574
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8404 14414 8432 15098
rect 8496 14482 8524 15302
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8484 14340 8536 14346
rect 8484 14282 8536 14288
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 14074 8432 14214
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8496 13938 8524 14282
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8128 12434 8156 12786
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 12442 8248 12718
rect 8036 12406 8156 12434
rect 8208 12436 8260 12442
rect 8036 12238 8064 12406
rect 8208 12378 8260 12384
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6840 10934 7144 10962
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7024 10674 7052 10746
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 10266 6960 10542
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6144 10160 6146 10169
rect 6090 10095 6146 10104
rect 6734 10160 6790 10169
rect 7024 10130 7052 10610
rect 7116 10130 7144 10934
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 6734 10095 6790 10104
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7208 10062 7236 10406
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9586 6040 9862
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6196 9489 6224 9590
rect 6182 9480 6238 9489
rect 6182 9415 6184 9424
rect 6236 9415 6238 9424
rect 6184 9386 6236 9392
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 6840 8974 6868 9998
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6932 9178 6960 9522
rect 7116 9178 7144 9522
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6828 8968 6880 8974
rect 6748 8928 6828 8956
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 6656 7954 6684 8774
rect 6748 8498 6776 8928
rect 6828 8910 6880 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6932 7818 6960 8366
rect 7116 8090 7144 8434
rect 7208 8430 7236 8910
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7300 8294 7328 11494
rect 7484 11082 7512 11698
rect 7668 11354 7696 11834
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7760 10674 7788 11494
rect 7852 11082 7880 11834
rect 8128 11150 8156 12038
rect 8220 11898 8248 12378
rect 8312 12306 8340 12786
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12374 8432 12582
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11898 8432 12174
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8496 11778 8524 12922
rect 8588 12646 8616 15642
rect 8680 12850 8708 17002
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8944 16584 8996 16590
rect 8942 16552 8944 16561
rect 8996 16552 8998 16561
rect 8942 16487 8998 16496
rect 8758 15600 8814 15609
rect 8758 15535 8760 15544
rect 8812 15535 8814 15544
rect 8760 15506 8812 15512
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8772 12850 8800 15098
rect 8864 14822 8892 15438
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8864 13938 8892 14418
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8956 13190 8984 15438
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12889 8984 13126
rect 9048 12986 9076 16934
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9416 16590 9444 16730
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9600 16522 9628 17478
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9692 16794 9720 17070
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9784 16590 9812 17983
rect 9968 17202 9996 18158
rect 10060 18154 10088 18702
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10244 18358 10272 18566
rect 10336 18426 10364 18566
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9956 16652 10008 16658
rect 9876 16612 9956 16640
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8942 12880 8998 12889
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8760 12844 8812 12850
rect 8942 12815 8998 12824
rect 9036 12844 9088 12850
rect 8760 12786 8812 12792
rect 9036 12786 9088 12792
rect 8680 12753 8708 12786
rect 8666 12744 8722 12753
rect 8772 12730 8800 12786
rect 8772 12702 8984 12730
rect 8666 12679 8668 12688
rect 8720 12679 8722 12688
rect 8668 12650 8720 12656
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8666 12472 8722 12481
rect 8666 12407 8722 12416
rect 8574 12336 8630 12345
rect 8574 12271 8630 12280
rect 8588 12238 8616 12271
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8220 11762 8524 11778
rect 8680 11762 8708 12407
rect 8208 11756 8524 11762
rect 8260 11750 8524 11756
rect 8668 11756 8720 11762
rect 8208 11698 8260 11704
rect 8668 11698 8720 11704
rect 8220 11626 8616 11642
rect 8208 11620 8616 11626
rect 8260 11614 8616 11620
rect 8208 11562 8260 11568
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7668 10470 7696 10610
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7392 8906 7420 10406
rect 7944 10266 7972 11018
rect 8220 10810 8248 11562
rect 8588 11558 8616 11614
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8496 11150 8524 11494
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10538 8064 10610
rect 8496 10606 8524 11086
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9586 7512 9862
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 8312 9110 8340 10406
rect 8772 10266 8800 12582
rect 8956 12374 8984 12702
rect 9048 12442 9076 12786
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 9140 12306 9168 16390
rect 9232 15026 9260 16390
rect 9600 16114 9628 16458
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9692 16046 9720 16526
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9402 15600 9458 15609
rect 9402 15535 9404 15544
rect 9456 15535 9458 15544
rect 9404 15506 9456 15512
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9324 14550 9352 15438
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9416 14346 9444 15302
rect 9692 15094 9720 15438
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9508 14929 9536 14962
rect 9588 14952 9640 14958
rect 9494 14920 9550 14929
rect 9588 14894 9640 14900
rect 9494 14855 9550 14864
rect 9600 14822 9628 14894
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9692 14414 9720 15030
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9416 13938 9444 14282
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9416 13410 9444 13874
rect 9508 13530 9536 13874
rect 9588 13864 9640 13870
rect 9692 13818 9720 14350
rect 9784 14074 9812 14350
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9770 13968 9826 13977
rect 9770 13903 9772 13912
rect 9824 13903 9826 13912
rect 9772 13874 9824 13880
rect 9640 13812 9720 13818
rect 9588 13806 9720 13812
rect 9600 13790 9720 13806
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9416 13382 9536 13410
rect 9508 13326 9536 13382
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9232 12714 9260 12786
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9218 12336 9274 12345
rect 9128 12300 9180 12306
rect 9324 12306 9352 12650
rect 9416 12442 9444 13262
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9692 12918 9720 13194
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9218 12271 9274 12280
rect 9312 12300 9364 12306
rect 9128 12242 9180 12248
rect 9232 11762 9260 12271
rect 9312 12242 9364 12248
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9324 11626 9352 12106
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11286 9168 11494
rect 9416 11286 9444 12242
rect 9508 12170 9536 12582
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9508 11694 9536 11834
rect 9600 11778 9628 12650
rect 9692 12238 9720 12854
rect 9876 12442 9904 16612
rect 9956 16594 10008 16600
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 15502 9996 16390
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9968 13938 9996 14350
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10060 13818 10088 16662
rect 10152 15638 10180 18022
rect 10244 17270 10272 18294
rect 10428 18290 10456 18702
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10520 16658 10548 16730
rect 10612 16726 10640 21354
rect 10888 20942 10916 21558
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10980 20466 11008 22358
rect 11072 22030 11100 22374
rect 11164 22030 11192 24754
rect 11244 23112 11296 23118
rect 11242 23080 11244 23089
rect 11296 23080 11298 23089
rect 11242 23015 11298 23024
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11072 21554 11100 21830
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10704 15994 10732 19314
rect 11072 18834 11100 21082
rect 11164 21010 11192 21830
rect 11348 21552 11376 26794
rect 11440 25378 11468 28358
rect 11532 28218 11560 28426
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11624 27946 11652 28426
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11532 25537 11560 25842
rect 11518 25528 11574 25537
rect 11518 25463 11574 25472
rect 11612 25424 11664 25430
rect 11610 25392 11612 25401
rect 11664 25392 11666 25401
rect 11440 25350 11560 25378
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11440 24410 11468 24686
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11532 24290 11560 25350
rect 11610 25327 11666 25336
rect 11612 25288 11664 25294
rect 11612 25230 11664 25236
rect 11624 24410 11652 25230
rect 11716 24614 11744 27950
rect 11900 26042 11928 28494
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11888 25832 11940 25838
rect 11808 25792 11888 25820
rect 11808 25158 11836 25792
rect 11888 25774 11940 25780
rect 11888 25288 11940 25294
rect 11888 25230 11940 25236
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11808 24834 11836 25094
rect 11900 24954 11928 25230
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 11808 24806 11928 24834
rect 11900 24750 11928 24806
rect 11992 24750 12020 31878
rect 12072 31816 12124 31822
rect 12070 31784 12072 31793
rect 12124 31784 12126 31793
rect 12360 31754 12388 33458
rect 12636 32978 12664 33526
rect 13082 33144 13138 33153
rect 13082 33079 13138 33088
rect 12624 32972 12676 32978
rect 12624 32914 12676 32920
rect 12900 32360 12952 32366
rect 12900 32302 12952 32308
rect 12532 32224 12584 32230
rect 12532 32166 12584 32172
rect 12544 32026 12572 32166
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12070 31719 12126 31728
rect 12176 31726 12388 31754
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 12084 30870 12112 31282
rect 12072 30864 12124 30870
rect 12072 30806 12124 30812
rect 12070 29472 12126 29481
rect 12070 29407 12126 29416
rect 12084 29170 12112 29407
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 12176 29050 12204 31726
rect 12912 31210 12940 32302
rect 12900 31204 12952 31210
rect 12900 31146 12952 31152
rect 12716 30048 12768 30054
rect 12716 29990 12768 29996
rect 12440 29708 12492 29714
rect 12440 29650 12492 29656
rect 12348 29164 12400 29170
rect 12348 29106 12400 29112
rect 12084 29022 12204 29050
rect 12084 26024 12112 29022
rect 12164 28960 12216 28966
rect 12164 28902 12216 28908
rect 12176 28626 12204 28902
rect 12360 28778 12388 29106
rect 12452 28937 12480 29650
rect 12728 29646 12756 29990
rect 13096 29646 13124 33079
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13188 32230 13216 32370
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13188 31346 13216 32166
rect 13176 31340 13228 31346
rect 13176 31282 13228 31288
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 12716 29640 12768 29646
rect 13084 29640 13136 29646
rect 12716 29582 12768 29588
rect 13004 29600 13084 29628
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12544 29073 12572 29446
rect 12636 29345 12664 29514
rect 12622 29336 12678 29345
rect 12622 29271 12678 29280
rect 12530 29064 12586 29073
rect 12530 28999 12586 29008
rect 12438 28928 12494 28937
rect 12438 28863 12494 28872
rect 12268 28750 12388 28778
rect 12268 28694 12296 28750
rect 12256 28688 12308 28694
rect 12532 28688 12584 28694
rect 12256 28630 12308 28636
rect 12530 28656 12532 28665
rect 12584 28656 12586 28665
rect 12164 28620 12216 28626
rect 12530 28591 12586 28600
rect 12164 28562 12216 28568
rect 12728 28558 12756 29582
rect 12898 29472 12954 29481
rect 12898 29407 12954 29416
rect 12912 29170 12940 29407
rect 13004 29238 13032 29600
rect 13084 29582 13136 29588
rect 13084 29300 13136 29306
rect 13084 29242 13136 29248
rect 12992 29232 13044 29238
rect 12992 29174 13044 29180
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 12912 29050 12940 29106
rect 12990 29064 13046 29073
rect 12912 29022 12990 29050
rect 12990 28999 13046 29008
rect 12808 28960 12860 28966
rect 12808 28902 12860 28908
rect 12256 28552 12308 28558
rect 12256 28494 12308 28500
rect 12348 28552 12400 28558
rect 12716 28552 12768 28558
rect 12348 28494 12400 28500
rect 12636 28512 12716 28540
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 12176 26994 12204 28358
rect 12268 28218 12296 28494
rect 12256 28212 12308 28218
rect 12256 28154 12308 28160
rect 12360 28082 12388 28494
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12530 27568 12586 27577
rect 12530 27503 12586 27512
rect 12544 27470 12572 27503
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12636 27316 12664 28512
rect 12716 28494 12768 28500
rect 12820 28014 12848 28902
rect 12808 28008 12860 28014
rect 12808 27950 12860 27956
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12912 27674 12940 27950
rect 12900 27668 12952 27674
rect 12900 27610 12952 27616
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 12544 27288 12664 27316
rect 12716 27328 12768 27334
rect 12544 26994 12572 27288
rect 12716 27270 12768 27276
rect 12728 27130 12756 27270
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12622 26888 12678 26897
rect 12622 26823 12678 26832
rect 12530 26616 12586 26625
rect 12530 26551 12586 26560
rect 12544 26382 12572 26551
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12544 26081 12572 26318
rect 12636 26314 12664 26823
rect 12728 26382 12756 27066
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12820 26790 12848 26930
rect 12912 26858 12940 27406
rect 13004 27169 13032 28999
rect 13096 28994 13124 29242
rect 13188 29170 13216 29990
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 13280 28994 13308 36246
rect 13372 34406 13400 39086
rect 21270 39039 21326 39839
rect 17224 37324 17276 37330
rect 17224 37266 17276 37272
rect 18144 37324 18196 37330
rect 18144 37266 18196 37272
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 13820 36916 13872 36922
rect 13820 36858 13872 36864
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13464 35562 13492 36314
rect 13636 35760 13688 35766
rect 13636 35702 13688 35708
rect 13452 35556 13504 35562
rect 13452 35498 13504 35504
rect 13648 35465 13676 35702
rect 13728 35624 13780 35630
rect 13728 35566 13780 35572
rect 13634 35456 13690 35465
rect 13634 35391 13690 35400
rect 13740 35154 13768 35566
rect 13728 35148 13780 35154
rect 13728 35090 13780 35096
rect 13360 34400 13412 34406
rect 13360 34342 13412 34348
rect 13360 33924 13412 33930
rect 13360 33866 13412 33872
rect 13372 29714 13400 33866
rect 13728 33584 13780 33590
rect 13728 33526 13780 33532
rect 13740 31793 13768 33526
rect 13832 32502 13860 36858
rect 14740 36848 14792 36854
rect 14740 36790 14792 36796
rect 16948 36848 17000 36854
rect 16948 36790 17000 36796
rect 14280 36712 14332 36718
rect 14280 36654 14332 36660
rect 14004 36576 14056 36582
rect 14004 36518 14056 36524
rect 14016 36310 14044 36518
rect 14004 36304 14056 36310
rect 14004 36246 14056 36252
rect 14186 35728 14242 35737
rect 14186 35663 14242 35672
rect 14200 35630 14228 35663
rect 14188 35624 14240 35630
rect 14016 35584 14188 35612
rect 14016 35086 14044 35584
rect 14188 35566 14240 35572
rect 14188 35488 14240 35494
rect 14188 35430 14240 35436
rect 14200 35290 14228 35430
rect 14292 35290 14320 36654
rect 14648 36576 14700 36582
rect 14648 36518 14700 36524
rect 14660 36174 14688 36518
rect 14752 36378 14780 36790
rect 15016 36712 15068 36718
rect 15016 36654 15068 36660
rect 14740 36372 14792 36378
rect 14740 36314 14792 36320
rect 14924 36236 14976 36242
rect 14924 36178 14976 36184
rect 14648 36168 14700 36174
rect 14648 36110 14700 36116
rect 14740 36168 14792 36174
rect 14740 36110 14792 36116
rect 14372 36032 14424 36038
rect 14372 35974 14424 35980
rect 14188 35284 14240 35290
rect 14188 35226 14240 35232
rect 14280 35284 14332 35290
rect 14280 35226 14332 35232
rect 14384 35086 14412 35974
rect 14556 35760 14608 35766
rect 14556 35702 14608 35708
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14004 33448 14056 33454
rect 14004 33390 14056 33396
rect 14016 33114 14044 33390
rect 14004 33108 14056 33114
rect 14004 33050 14056 33056
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13832 31822 13860 32438
rect 13820 31816 13872 31822
rect 13726 31784 13782 31793
rect 13820 31758 13872 31764
rect 14004 31816 14056 31822
rect 14004 31758 14056 31764
rect 13726 31719 13782 31728
rect 13740 31346 13768 31719
rect 14016 31414 14044 31758
rect 14476 31754 14504 34682
rect 14568 33930 14596 35702
rect 14752 35698 14780 36110
rect 14936 35766 14964 36178
rect 15028 36174 15056 36654
rect 16580 36576 16632 36582
rect 16580 36518 16632 36524
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 15292 36100 15344 36106
rect 15292 36042 15344 36048
rect 15384 36100 15436 36106
rect 15384 36042 15436 36048
rect 14924 35760 14976 35766
rect 14924 35702 14976 35708
rect 15304 35698 15332 36042
rect 15396 35834 15424 36042
rect 15384 35828 15436 35834
rect 15384 35770 15436 35776
rect 15658 35728 15714 35737
rect 14740 35692 14792 35698
rect 14740 35634 14792 35640
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 15292 35692 15344 35698
rect 15658 35663 15714 35672
rect 15936 35692 15988 35698
rect 15292 35634 15344 35640
rect 14738 35320 14794 35329
rect 14738 35255 14794 35264
rect 14752 35222 14780 35255
rect 14740 35216 14792 35222
rect 14740 35158 14792 35164
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 14832 34468 14884 34474
rect 14832 34410 14884 34416
rect 14740 33992 14792 33998
rect 14740 33934 14792 33940
rect 14556 33924 14608 33930
rect 14556 33866 14608 33872
rect 14556 33516 14608 33522
rect 14556 33458 14608 33464
rect 14568 32910 14596 33458
rect 14648 33380 14700 33386
rect 14648 33322 14700 33328
rect 14556 32904 14608 32910
rect 14556 32846 14608 32852
rect 14568 31890 14596 32846
rect 14660 32774 14688 33322
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14660 32502 14688 32710
rect 14752 32570 14780 33934
rect 14844 33658 14872 34410
rect 14924 33992 14976 33998
rect 14924 33934 14976 33940
rect 14832 33652 14884 33658
rect 14832 33594 14884 33600
rect 14844 32910 14872 33594
rect 14936 33318 14964 33934
rect 14924 33312 14976 33318
rect 14924 33254 14976 33260
rect 15028 33046 15056 34546
rect 15212 33998 15240 35634
rect 15672 35630 15700 35663
rect 15936 35634 15988 35640
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 15384 34400 15436 34406
rect 15384 34342 15436 34348
rect 15476 34400 15528 34406
rect 15476 34342 15528 34348
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15200 33992 15252 33998
rect 15200 33934 15252 33940
rect 15120 33658 15148 33934
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15212 33454 15240 33934
rect 15396 33590 15424 34342
rect 15384 33584 15436 33590
rect 15384 33526 15436 33532
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 15488 33386 15516 34342
rect 15476 33380 15528 33386
rect 15476 33322 15528 33328
rect 15568 33380 15620 33386
rect 15568 33322 15620 33328
rect 15580 33266 15608 33322
rect 15672 33318 15700 35566
rect 15948 35086 15976 35634
rect 15936 35080 15988 35086
rect 15936 35022 15988 35028
rect 15844 33924 15896 33930
rect 15844 33866 15896 33872
rect 15856 33454 15884 33866
rect 15844 33448 15896 33454
rect 15844 33390 15896 33396
rect 15488 33238 15608 33266
rect 15660 33312 15712 33318
rect 15660 33254 15712 33260
rect 15016 33040 15068 33046
rect 15016 32982 15068 32988
rect 15028 32910 15056 32982
rect 15488 32910 15516 33238
rect 15568 32972 15620 32978
rect 15620 32932 15792 32960
rect 15568 32914 15620 32920
rect 14832 32904 14884 32910
rect 14832 32846 14884 32852
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 14740 32564 14792 32570
rect 14740 32506 14792 32512
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14660 32026 14688 32438
rect 15120 32434 15148 32710
rect 15212 32434 15240 32778
rect 15396 32502 15424 32846
rect 15660 32768 15712 32774
rect 15660 32710 15712 32716
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 14740 32428 14792 32434
rect 14740 32370 14792 32376
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 15200 32428 15252 32434
rect 15200 32370 15252 32376
rect 14648 32020 14700 32026
rect 14648 31962 14700 31968
rect 14556 31884 14608 31890
rect 14556 31826 14608 31832
rect 14292 31726 14504 31754
rect 14004 31408 14056 31414
rect 14004 31350 14056 31356
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13912 30592 13964 30598
rect 13912 30534 13964 30540
rect 13452 30048 13504 30054
rect 13452 29990 13504 29996
rect 13464 29714 13492 29990
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 13452 29708 13504 29714
rect 13452 29650 13504 29656
rect 13096 28966 13308 28994
rect 13280 28626 13308 28966
rect 13268 28620 13320 28626
rect 13268 28562 13320 28568
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 12990 27160 13046 27169
rect 12990 27095 13046 27104
rect 12900 26852 12952 26858
rect 12900 26794 12952 26800
rect 12808 26784 12860 26790
rect 12808 26726 12860 26732
rect 12806 26480 12862 26489
rect 12806 26415 12862 26424
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12530 26072 12586 26081
rect 12084 25996 12204 26024
rect 12530 26007 12586 26016
rect 12176 25906 12204 25996
rect 12636 25974 12664 26250
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12084 25673 12112 25842
rect 12164 25764 12216 25770
rect 12216 25724 12296 25752
rect 12164 25706 12216 25712
rect 12070 25664 12126 25673
rect 12070 25599 12126 25608
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11888 24744 11940 24750
rect 11888 24686 11940 24692
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11612 24404 11664 24410
rect 11612 24346 11664 24352
rect 11532 24262 11652 24290
rect 11518 24168 11574 24177
rect 11518 24103 11574 24112
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11440 23118 11468 23666
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11336 21546 11388 21552
rect 11336 21488 11388 21494
rect 11532 21162 11560 24103
rect 11624 23186 11652 24262
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11716 23066 11744 24142
rect 11808 23526 11836 24686
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11992 24274 12020 24550
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11900 23730 11928 24006
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11992 23254 12020 24006
rect 12084 23662 12112 25230
rect 12164 24676 12216 24682
rect 12164 24618 12216 24624
rect 12176 24138 12204 24618
rect 12268 24614 12296 25724
rect 12544 25702 12572 25842
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12532 25696 12584 25702
rect 12346 25664 12402 25673
rect 12532 25638 12584 25644
rect 12346 25599 12402 25608
rect 12360 24818 12388 25599
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12440 25152 12492 25158
rect 12440 25094 12492 25100
rect 12452 24818 12480 25094
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12256 24608 12308 24614
rect 12544 24585 12572 25298
rect 12256 24550 12308 24556
rect 12530 24576 12586 24585
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23662 12204 24074
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12084 23322 12112 23598
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 11980 23248 12032 23254
rect 11978 23216 11980 23225
rect 12032 23216 12034 23225
rect 11796 23180 11848 23186
rect 11978 23151 12034 23160
rect 11796 23122 11848 23128
rect 11624 23038 11744 23066
rect 11624 22982 11652 23038
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11624 21894 11652 22918
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11612 21412 11664 21418
rect 11612 21354 11664 21360
rect 11348 21134 11560 21162
rect 11624 21146 11652 21354
rect 11612 21140 11664 21146
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11072 18737 11100 18770
rect 11058 18728 11114 18737
rect 11058 18663 11114 18672
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10888 18426 10916 18566
rect 10966 18456 11022 18465
rect 10876 18420 10928 18426
rect 10966 18391 10968 18400
rect 10876 18362 10928 18368
rect 11020 18391 11022 18400
rect 10968 18362 11020 18368
rect 11164 18034 11192 20742
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11256 18766 11284 19858
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11164 18006 11284 18034
rect 11150 17912 11206 17921
rect 11150 17847 11206 17856
rect 11164 17678 11192 17847
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 10980 17338 11008 17614
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 16590 10824 17138
rect 10888 16658 10916 17206
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 11072 16590 11100 17478
rect 11152 17128 11204 17134
rect 11256 17116 11284 18006
rect 11204 17088 11284 17116
rect 11152 17070 11204 17076
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10152 15502 10180 15574
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 9968 13790 10088 13818
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9772 12368 9824 12374
rect 9968 12322 9996 13790
rect 10152 13530 10180 13874
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 13258 10272 14758
rect 10336 13802 10364 15030
rect 10428 15026 10456 15438
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10520 14482 10548 15438
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10612 14362 10640 15982
rect 10704 15966 10916 15994
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15502 10732 15846
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10888 15450 10916 15966
rect 10980 15570 11008 16390
rect 11072 16114 11100 16526
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10704 15026 10732 15438
rect 10888 15422 11008 15450
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10520 14334 10640 14362
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10138 12880 10194 12889
rect 10336 12866 10364 13738
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10138 12815 10140 12824
rect 10192 12815 10194 12824
rect 10244 12838 10364 12866
rect 10140 12786 10192 12792
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9772 12310 9824 12316
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9784 12102 9812 12310
rect 9876 12294 9996 12322
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9600 11762 9720 11778
rect 9600 11756 9732 11762
rect 9600 11750 9680 11756
rect 9680 11698 9732 11704
rect 9784 11694 9812 12038
rect 9876 11778 9904 12294
rect 10060 12238 10088 12582
rect 10244 12434 10272 12838
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 12646 10364 12718
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10152 12406 10272 12434
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9968 11898 9996 12174
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9876 11750 10088 11778
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8666 10160 8722 10169
rect 8666 10095 8668 10104
rect 8720 10095 8722 10104
rect 8668 10066 8720 10072
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7300 7970 7328 8230
rect 7300 7942 7420 7970
rect 7392 7886 7420 7942
rect 8128 7886 8156 8842
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 8220 7750 8248 8910
rect 8312 8498 8340 9046
rect 8404 8906 8432 9998
rect 8956 9518 8984 9998
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8496 8090 8524 8978
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8498 8708 8774
rect 9048 8634 9076 8910
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9140 8566 9168 9930
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 9140 7886 9168 8502
rect 9324 8362 9352 11086
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10130 9444 11018
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10674 9720 10950
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9692 10169 9720 10406
rect 9784 10198 9812 10406
rect 9772 10192 9824 10198
rect 9678 10160 9734 10169
rect 9404 10124 9456 10130
rect 9772 10134 9824 10140
rect 9678 10095 9680 10104
rect 9404 10066 9456 10072
rect 9732 10095 9734 10104
rect 9680 10066 9732 10072
rect 9588 10056 9640 10062
rect 9876 10010 9904 11630
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10266 9996 10542
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9968 10062 9996 10202
rect 9640 10004 9904 10010
rect 9588 9998 9904 10004
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9600 9982 9904 9998
rect 9876 8974 9904 9982
rect 10060 9042 10088 11750
rect 10152 11218 10180 12406
rect 10232 12368 10284 12374
rect 10230 12336 10232 12345
rect 10284 12336 10286 12345
rect 10230 12271 10286 12280
rect 10336 12102 10364 12582
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10428 11762 10456 12922
rect 10520 12764 10548 14334
rect 10704 14006 10732 14962
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10796 13326 10824 14758
rect 10888 14414 10916 15302
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10888 13938 10916 14350
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10980 12986 11008 15422
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11072 14006 11100 14554
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13326 11100 13670
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10980 12850 11008 12922
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10600 12776 10652 12782
rect 10520 12736 10600 12764
rect 10600 12718 10652 12724
rect 10968 12640 11020 12646
rect 11164 12617 11192 17070
rect 11348 16289 11376 21134
rect 11612 21082 11664 21088
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 19854 11468 20198
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11440 19446 11468 19790
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11532 18834 11560 21014
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20466 11652 20878
rect 11716 20618 11744 22374
rect 11808 20806 11836 23122
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11900 22710 11928 22918
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 12084 22574 12112 23258
rect 12268 22778 12296 24550
rect 12530 24511 12586 24520
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 23769 12388 24142
rect 12346 23760 12402 23769
rect 12346 23695 12402 23704
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 12084 22030 12112 22510
rect 12176 22166 12204 22578
rect 12256 22500 12308 22506
rect 12256 22442 12308 22448
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12084 21486 12112 21626
rect 12176 21554 12204 22102
rect 12268 21690 12296 22442
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12072 21480 12124 21486
rect 12072 21422 12124 21428
rect 12268 21078 12296 21626
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11716 20590 11836 20618
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11702 20360 11758 20369
rect 11702 20295 11758 20304
rect 11716 19378 11744 20295
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11808 19258 11836 20590
rect 12360 19854 12388 23462
rect 12452 22982 12480 23666
rect 12544 23254 12572 24346
rect 12636 24313 12664 25774
rect 12728 25770 12756 25842
rect 12716 25764 12768 25770
rect 12716 25706 12768 25712
rect 12820 25242 12848 26415
rect 12912 26382 12940 26794
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 13004 25906 13032 27095
rect 13188 26976 13216 27406
rect 13280 27169 13308 27406
rect 13266 27160 13322 27169
rect 13266 27095 13322 27104
rect 13268 26988 13320 26994
rect 13096 26948 13268 26976
rect 13096 26382 13124 26948
rect 13268 26930 13320 26936
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 13280 26382 13308 26454
rect 13084 26376 13136 26382
rect 13268 26376 13320 26382
rect 13084 26318 13136 26324
rect 13266 26344 13268 26353
rect 13320 26344 13322 26353
rect 13266 26279 13322 26288
rect 13268 26240 13320 26246
rect 13266 26208 13268 26217
rect 13320 26208 13322 26217
rect 13266 26143 13322 26152
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 13372 25786 13400 29650
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 13648 29170 13676 29582
rect 13728 29572 13780 29578
rect 13728 29514 13780 29520
rect 13740 29238 13768 29514
rect 13820 29504 13872 29510
rect 13820 29446 13872 29452
rect 13832 29306 13860 29446
rect 13820 29300 13872 29306
rect 13820 29242 13872 29248
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 13452 29164 13504 29170
rect 13636 29164 13688 29170
rect 13504 29124 13584 29152
rect 13452 29106 13504 29112
rect 13556 29034 13584 29124
rect 13636 29106 13688 29112
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 13544 29028 13596 29034
rect 13544 28970 13596 28976
rect 13280 25758 13400 25786
rect 12728 25226 12848 25242
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 12716 25220 12848 25226
rect 12768 25214 12848 25220
rect 12716 25162 12768 25168
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12716 24812 12768 24818
rect 12716 24754 12768 24760
rect 12728 24342 12756 24754
rect 12716 24336 12768 24342
rect 12622 24304 12678 24313
rect 12716 24278 12768 24284
rect 12622 24239 12678 24248
rect 12636 24188 12664 24239
rect 12716 24200 12768 24206
rect 12636 24160 12716 24188
rect 12716 24142 12768 24148
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22642 12480 22918
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12544 22642 12572 22714
rect 12636 22642 12664 23054
rect 12728 22778 12756 24006
rect 12820 23186 12848 25094
rect 12900 24744 12952 24750
rect 13004 24732 13032 25230
rect 13096 24886 13124 25230
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 13280 24800 13308 25758
rect 13360 25696 13412 25702
rect 13360 25638 13412 25644
rect 13372 25294 13400 25638
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13372 24954 13400 25094
rect 13360 24948 13412 24954
rect 13360 24890 13412 24896
rect 13464 24818 13492 28970
rect 13556 27402 13584 28970
rect 13648 28558 13676 29106
rect 13636 28552 13688 28558
rect 13636 28494 13688 28500
rect 13740 28490 13768 29174
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13634 27432 13690 27441
rect 13544 27396 13596 27402
rect 13634 27367 13690 27376
rect 13544 27338 13596 27344
rect 13556 27146 13584 27338
rect 13648 27334 13676 27367
rect 13636 27328 13688 27334
rect 13636 27270 13688 27276
rect 13556 27118 13676 27146
rect 13542 27024 13598 27033
rect 13648 26994 13676 27118
rect 13542 26959 13544 26968
rect 13596 26959 13598 26968
rect 13636 26988 13688 26994
rect 13544 26930 13596 26936
rect 13636 26930 13688 26936
rect 13648 26234 13676 26930
rect 13726 26616 13782 26625
rect 13726 26551 13782 26560
rect 13556 26206 13676 26234
rect 13556 25770 13584 26206
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13544 25764 13596 25770
rect 13544 25706 13596 25712
rect 13556 24954 13584 25706
rect 13648 25498 13676 25842
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13360 24812 13412 24818
rect 13280 24772 13360 24800
rect 13004 24704 13124 24732
rect 12900 24686 12952 24692
rect 12912 24070 12940 24686
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 12808 23180 12860 23186
rect 12808 23122 12860 23128
rect 12912 22964 12940 23666
rect 13004 23118 13032 24550
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 12992 22976 13044 22982
rect 12912 22936 12992 22964
rect 12992 22918 13044 22924
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12452 21962 12480 22578
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12544 20058 12572 20334
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12544 19961 12572 19994
rect 12530 19952 12586 19961
rect 12530 19887 12586 19896
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11624 19230 11836 19258
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11532 18737 11560 18770
rect 11518 18728 11574 18737
rect 11518 18663 11574 18672
rect 11624 18578 11652 19230
rect 11704 18692 11756 18698
rect 11704 18634 11756 18640
rect 11440 18550 11652 18578
rect 11440 18290 11468 18550
rect 11716 18358 11744 18634
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11334 16280 11390 16289
rect 11334 16215 11390 16224
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13258 11284 14214
rect 11348 14074 11376 14418
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 10968 12582 11020 12588
rect 11150 12608 11206 12617
rect 10980 12434 11008 12582
rect 11150 12543 11206 12552
rect 10980 12406 11100 12434
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10508 12096 10560 12102
rect 10612 12084 10640 12242
rect 10692 12096 10744 12102
rect 10612 12056 10692 12084
rect 10508 12038 10560 12044
rect 10692 12038 10744 12044
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10152 10674 10180 11154
rect 10244 10674 10272 11494
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10232 10668 10284 10674
rect 10284 10628 10364 10656
rect 10232 10610 10284 10616
rect 10336 10198 10364 10628
rect 10324 10192 10376 10198
rect 10230 10160 10286 10169
rect 10324 10134 10376 10140
rect 10230 10095 10232 10104
rect 10284 10095 10286 10104
rect 10232 10066 10284 10072
rect 10244 9586 10272 10066
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9586 10456 9998
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9416 8022 9444 8434
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 8090 9536 8366
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10152 8090 10180 8298
rect 10244 8090 10272 8298
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9876 7886 9904 8026
rect 10336 7886 10364 9454
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 7886 10456 8774
rect 10520 8566 10548 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10796 11762 10824 11834
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10782 10704 10838 10713
rect 10692 10668 10744 10674
rect 10888 10674 10916 12310
rect 10980 12170 11008 12310
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 11072 12050 11100 12406
rect 11152 12368 11204 12374
rect 11150 12336 11152 12345
rect 11204 12336 11206 12345
rect 11348 12306 11376 12786
rect 11440 12714 11468 18226
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11532 16590 11560 16934
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 16114 11560 16526
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11624 15994 11652 18090
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11532 15966 11652 15994
rect 11428 12708 11480 12714
rect 11428 12650 11480 12656
rect 11426 12608 11482 12617
rect 11426 12543 11482 12552
rect 11150 12271 11206 12280
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10980 12022 11100 12050
rect 10980 11762 11008 12022
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11060 11688 11112 11694
rect 10980 11636 11060 11642
rect 10980 11630 11112 11636
rect 10980 11614 11100 11630
rect 10980 11014 11008 11614
rect 11164 11354 11192 12174
rect 11256 11898 11284 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10782 10639 10784 10648
rect 10692 10610 10744 10616
rect 10836 10639 10838 10648
rect 10876 10668 10928 10674
rect 10784 10610 10836 10616
rect 10876 10610 10928 10616
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10704 10266 10732 10610
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 11164 10062 11192 10610
rect 11256 10062 11284 11698
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11348 10266 11376 10678
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10968 10056 11020 10062
rect 11152 10056 11204 10062
rect 11020 10016 11100 10044
rect 10968 9998 11020 10004
rect 10612 9722 10640 9998
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 11072 9654 11100 10016
rect 11244 10056 11296 10062
rect 11152 9998 11204 10004
rect 11242 10024 11244 10033
rect 11296 10024 11298 10033
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11072 8974 11100 9590
rect 11164 9586 11192 9998
rect 11242 9959 11298 9968
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11348 9518 11376 10202
rect 11336 9512 11388 9518
rect 11336 9454 11388 9460
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10888 8430 10916 8774
rect 11348 8498 11376 9454
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 7886 10732 8230
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10980 7750 11008 8434
rect 11242 8120 11298 8129
rect 11242 8055 11244 8064
rect 11296 8055 11298 8064
rect 11244 8026 11296 8032
rect 11150 7984 11206 7993
rect 11150 7919 11206 7928
rect 11164 7886 11192 7919
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 938 4111 994 4120
rect 4068 4140 4120 4146
rect 952 4010 980 4111
rect 4068 4082 4120 4088
rect 940 4004 992 4010
rect 940 3946 992 3952
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 10980 3534 11008 3878
rect 11256 3534 11284 8026
rect 11440 7970 11468 12543
rect 11532 10810 11560 15966
rect 11716 15094 11744 16526
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14929 11652 14962
rect 11610 14920 11666 14929
rect 11610 14855 11666 14864
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11624 10282 11652 14214
rect 11808 12866 11836 18566
rect 11900 18426 11928 19314
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11992 17202 12020 19654
rect 12360 19446 12388 19790
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12084 18970 12112 19314
rect 12624 19304 12676 19310
rect 12254 19272 12310 19281
rect 12624 19246 12676 19252
rect 12254 19207 12310 19216
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18426 12112 18702
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12176 18306 12204 19110
rect 12268 18834 12296 19207
rect 12636 18834 12664 19246
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12360 18426 12388 18566
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12084 18278 12204 18306
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11980 17196 12032 17202
rect 11980 17138 12032 17144
rect 11900 17082 11928 17138
rect 12084 17082 12112 18278
rect 12636 18154 12664 18770
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17202 12204 17614
rect 12360 17270 12388 17682
rect 12636 17678 12664 18090
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 11900 17054 12112 17082
rect 11900 14278 11928 17054
rect 12176 16658 12204 17138
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 16250 12020 16390
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12452 16114 12480 17002
rect 12544 16590 12572 17478
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12636 16504 12664 17206
rect 12728 17134 12756 22374
rect 12820 22098 12848 22442
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 13004 20942 13032 22918
rect 13096 22506 13124 24704
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 13188 23730 13216 24006
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 13280 22094 13308 24772
rect 13360 24754 13412 24760
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13556 24274 13584 24890
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13648 24206 13676 25434
rect 13740 25226 13768 26551
rect 13728 25220 13780 25226
rect 13728 25162 13780 25168
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13832 24138 13860 29038
rect 13924 27130 13952 30534
rect 13912 27124 13964 27130
rect 13912 27066 13964 27072
rect 13910 27024 13966 27033
rect 13910 26959 13912 26968
rect 13964 26959 13966 26968
rect 13912 26930 13964 26936
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 13924 26382 13952 26726
rect 13912 26376 13964 26382
rect 13910 26344 13912 26353
rect 13964 26344 13966 26353
rect 14016 26314 14044 31350
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 14200 30734 14228 31078
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 14292 30546 14320 31726
rect 14556 31272 14608 31278
rect 14556 31214 14608 31220
rect 14568 30938 14596 31214
rect 14464 30932 14516 30938
rect 14464 30874 14516 30880
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14200 30518 14320 30546
rect 14094 29200 14150 29209
rect 14094 29135 14096 29144
rect 14148 29135 14150 29144
rect 14096 29106 14148 29112
rect 14200 29102 14228 30518
rect 14476 30394 14504 30874
rect 14554 30832 14610 30841
rect 14554 30767 14556 30776
rect 14608 30767 14610 30776
rect 14556 30738 14608 30744
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14464 29504 14516 29510
rect 14516 29464 14596 29492
rect 14464 29446 14516 29452
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14188 29096 14240 29102
rect 14476 29073 14504 29106
rect 14188 29038 14240 29044
rect 14462 29064 14518 29073
rect 14462 28999 14518 29008
rect 14568 28694 14596 29464
rect 14556 28688 14608 28694
rect 14556 28630 14608 28636
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 14094 27296 14150 27305
rect 14094 27231 14150 27240
rect 14108 27130 14136 27231
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14108 26382 14136 26726
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 13910 26279 13966 26288
rect 14004 26308 14056 26314
rect 14004 26250 14056 26256
rect 14200 25378 14228 28562
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 14372 26852 14424 26858
rect 14372 26794 14424 26800
rect 14384 26586 14412 26794
rect 14372 26580 14424 26586
rect 14372 26522 14424 26528
rect 14280 26512 14332 26518
rect 14280 26454 14332 26460
rect 14016 25350 14228 25378
rect 13910 24576 13966 24585
rect 13910 24511 13966 24520
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13818 23896 13874 23905
rect 13818 23831 13874 23840
rect 13832 23798 13860 23831
rect 13820 23792 13872 23798
rect 13820 23734 13872 23740
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13372 23186 13400 23666
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13372 22642 13400 23122
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13280 22066 13400 22094
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21486 13124 21966
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 13372 21146 13400 22066
rect 13556 22030 13584 23258
rect 13924 23118 13952 24511
rect 13912 23112 13964 23118
rect 13832 23072 13912 23100
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13832 21894 13860 23072
rect 13912 23054 13964 23060
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13924 22030 13952 22578
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13372 20942 13400 21082
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13084 20868 13136 20874
rect 13084 20810 13136 20816
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12912 17882 12940 18226
rect 13096 18222 13124 20810
rect 13280 20534 13308 20878
rect 13464 20754 13492 21014
rect 13372 20726 13492 20754
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13280 20058 13308 20470
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12716 16516 12768 16522
rect 12636 16476 12716 16504
rect 12716 16458 12768 16464
rect 12728 16114 12756 16458
rect 12820 16250 12848 17478
rect 12912 17338 12940 17818
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 13004 17066 13032 18158
rect 13084 17672 13136 17678
rect 13188 17660 13216 18158
rect 13136 17632 13216 17660
rect 13084 17614 13136 17620
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 11980 15020 12032 15026
rect 12032 14980 12204 15008
rect 11980 14962 12032 14968
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11716 12850 11836 12866
rect 11716 12844 11848 12850
rect 11716 12838 11796 12844
rect 11716 12238 11744 12838
rect 11796 12786 11848 12792
rect 11900 12238 11928 13738
rect 12084 13394 12112 14758
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12918 12112 13330
rect 12072 12912 12124 12918
rect 12176 12889 12204 14980
rect 12254 14920 12310 14929
rect 12254 14855 12256 14864
rect 12308 14855 12310 14864
rect 12256 14826 12308 14832
rect 12254 13968 12310 13977
rect 12254 13903 12310 13912
rect 12072 12854 12124 12860
rect 12162 12880 12218 12889
rect 12084 12764 12112 12854
rect 12162 12815 12218 12824
rect 12084 12736 12204 12764
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11978 12472 12034 12481
rect 11978 12407 12034 12416
rect 11992 12238 12020 12407
rect 12084 12306 12112 12582
rect 12176 12306 12204 12736
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 11704 12232 11756 12238
rect 11888 12232 11940 12238
rect 11704 12174 11756 12180
rect 11808 12192 11888 12220
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 10674 11744 12038
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11704 10532 11756 10538
rect 11808 10520 11836 12192
rect 11888 12174 11940 12180
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12084 11762 12112 12242
rect 12268 11762 12296 13903
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11756 10492 11836 10520
rect 11704 10474 11756 10480
rect 11624 10254 11836 10282
rect 11520 10056 11572 10062
rect 11612 10056 11664 10062
rect 11520 9998 11572 10004
rect 11610 10024 11612 10033
rect 11664 10024 11666 10033
rect 11532 9674 11560 9998
rect 11610 9959 11666 9968
rect 11808 9674 11836 10254
rect 11900 10062 11928 11630
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12268 11150 12296 11562
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12360 10554 12388 15914
rect 12728 15706 12756 16050
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12452 14618 12480 15438
rect 12544 15162 12572 15438
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12636 14550 12664 15574
rect 12820 15570 12848 15914
rect 12912 15706 12940 16526
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12452 14278 12480 14350
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12452 12238 12480 14214
rect 12544 13734 12572 14350
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12636 13938 12664 14282
rect 12728 14074 12756 15098
rect 12820 14278 12848 15506
rect 12912 14958 12940 15642
rect 13004 15502 13032 15846
rect 13096 15722 13124 17614
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13188 16590 13216 16934
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13188 16114 13216 16526
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13280 16046 13308 17478
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13372 15994 13400 20726
rect 13648 20466 13676 20742
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13648 19922 13676 20198
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13740 19786 13768 20470
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13832 19718 13860 20334
rect 13820 19712 13872 19718
rect 13924 19700 13952 21966
rect 14016 21010 14044 25350
rect 14292 25294 14320 26454
rect 14372 26376 14424 26382
rect 14370 26344 14372 26353
rect 14424 26344 14426 26353
rect 14370 26279 14426 26288
rect 14476 25294 14504 26862
rect 14660 26489 14688 31962
rect 14752 31686 14780 32370
rect 15396 32230 15424 32438
rect 15672 32230 15700 32710
rect 15764 32502 15792 32932
rect 15752 32496 15804 32502
rect 15752 32438 15804 32444
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15384 32224 15436 32230
rect 15384 32166 15436 32172
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15752 32224 15804 32230
rect 15752 32166 15804 32172
rect 15396 32026 15424 32166
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15764 31822 15792 32166
rect 15016 31816 15068 31822
rect 15016 31758 15068 31764
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15752 31816 15804 31822
rect 15752 31758 15804 31764
rect 14740 31680 14792 31686
rect 14740 31622 14792 31628
rect 14752 31482 14780 31622
rect 14740 31476 14792 31482
rect 14740 31418 14792 31424
rect 15028 31278 15056 31758
rect 15108 31748 15160 31754
rect 15108 31690 15160 31696
rect 15120 31346 15148 31690
rect 15304 31414 15332 31758
rect 15660 31680 15712 31686
rect 15660 31622 15712 31628
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15108 31340 15160 31346
rect 15108 31282 15160 31288
rect 15016 31272 15068 31278
rect 15016 31214 15068 31220
rect 15120 31210 15148 31282
rect 15108 31204 15160 31210
rect 15108 31146 15160 31152
rect 15672 30734 15700 31622
rect 15856 31482 15884 32370
rect 15844 31476 15896 31482
rect 15844 31418 15896 31424
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15304 29702 15792 29730
rect 15948 29714 15976 35022
rect 16500 33930 16528 36110
rect 16592 35562 16620 36518
rect 16764 36100 16816 36106
rect 16764 36042 16816 36048
rect 16776 35766 16804 36042
rect 16856 36032 16908 36038
rect 16856 35974 16908 35980
rect 16764 35760 16816 35766
rect 16764 35702 16816 35708
rect 16868 35698 16896 35974
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16580 35556 16632 35562
rect 16580 35498 16632 35504
rect 16856 35488 16908 35494
rect 16960 35476 16988 36790
rect 17052 36718 17080 37198
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 17052 36174 17080 36654
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 17052 35698 17080 36110
rect 17236 35698 17264 37266
rect 18156 36786 18184 37266
rect 19892 36848 19944 36854
rect 19892 36790 19944 36796
rect 20168 36848 20220 36854
rect 20168 36790 20220 36796
rect 20352 36848 20404 36854
rect 20352 36790 20404 36796
rect 17408 36780 17460 36786
rect 17408 36722 17460 36728
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 19524 36780 19576 36786
rect 19524 36722 19576 36728
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 16908 35448 16988 35476
rect 17224 35488 17276 35494
rect 16856 35430 16908 35436
rect 17224 35430 17276 35436
rect 16868 34746 16896 35430
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17236 34610 17264 35430
rect 17328 35086 17356 36110
rect 17420 35154 17448 36722
rect 17500 36712 17552 36718
rect 17500 36654 17552 36660
rect 17512 36378 17540 36654
rect 17500 36372 17552 36378
rect 17500 36314 17552 36320
rect 18156 36174 18184 36722
rect 18236 36712 18288 36718
rect 18236 36654 18288 36660
rect 19340 36712 19392 36718
rect 19340 36654 19392 36660
rect 18248 36310 18276 36654
rect 18236 36304 18288 36310
rect 18236 36246 18288 36252
rect 19352 36174 19380 36654
rect 19536 36258 19564 36722
rect 19536 36242 19656 36258
rect 19536 36236 19668 36242
rect 19536 36230 19616 36236
rect 19616 36178 19668 36184
rect 18144 36168 18196 36174
rect 18144 36110 18196 36116
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 18052 35828 18104 35834
rect 18156 35816 18184 36110
rect 18104 35788 18184 35816
rect 18234 35864 18290 35873
rect 19260 35834 19288 36110
rect 18234 35799 18290 35808
rect 19248 35828 19300 35834
rect 18052 35770 18104 35776
rect 18248 35766 18276 35799
rect 19248 35770 19300 35776
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 17776 35692 17828 35698
rect 17776 35634 17828 35640
rect 17868 35692 17920 35698
rect 17868 35634 17920 35640
rect 17408 35148 17460 35154
rect 17408 35090 17460 35096
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 16764 34604 16816 34610
rect 16764 34546 16816 34552
rect 17224 34604 17276 34610
rect 17224 34546 17276 34552
rect 16488 33924 16540 33930
rect 16488 33866 16540 33872
rect 16776 33658 16804 34546
rect 17236 34202 17264 34546
rect 17328 34542 17356 35022
rect 17316 34536 17368 34542
rect 17316 34478 17368 34484
rect 17224 34196 17276 34202
rect 17224 34138 17276 34144
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 16028 33516 16080 33522
rect 16028 33458 16080 33464
rect 16948 33516 17000 33522
rect 17052 33504 17080 33594
rect 17000 33476 17080 33504
rect 16948 33458 17000 33464
rect 16040 31482 16068 33458
rect 16120 33380 16172 33386
rect 16120 33322 16172 33328
rect 16132 32434 16160 33322
rect 16580 32836 16632 32842
rect 16580 32778 16632 32784
rect 16120 32428 16172 32434
rect 16120 32370 16172 32376
rect 16304 32360 16356 32366
rect 16304 32302 16356 32308
rect 16120 32224 16172 32230
rect 16120 32166 16172 32172
rect 16132 31822 16160 32166
rect 16316 31958 16344 32302
rect 16304 31952 16356 31958
rect 16304 31894 16356 31900
rect 16120 31816 16172 31822
rect 16120 31758 16172 31764
rect 16028 31476 16080 31482
rect 16028 31418 16080 31424
rect 14738 29608 14794 29617
rect 14738 29543 14794 29552
rect 14752 29170 14780 29543
rect 15014 29336 15070 29345
rect 15014 29271 15070 29280
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14832 29164 14884 29170
rect 14832 29106 14884 29112
rect 14844 28150 14872 29106
rect 15028 28994 15056 29271
rect 15212 29238 15240 29650
rect 15304 29578 15332 29702
rect 15764 29646 15792 29702
rect 15936 29708 15988 29714
rect 15936 29650 15988 29656
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15292 29572 15344 29578
rect 15292 29514 15344 29520
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 15396 29238 15424 29446
rect 15580 29306 15608 29582
rect 15660 29572 15712 29578
rect 15660 29514 15712 29520
rect 15568 29300 15620 29306
rect 15568 29242 15620 29248
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15384 29096 15436 29102
rect 15384 29038 15436 29044
rect 15028 28966 15148 28994
rect 14832 28144 14884 28150
rect 14832 28086 14884 28092
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14646 26480 14702 26489
rect 14646 26415 14702 26424
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14660 25702 14688 26318
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14108 24410 14136 24754
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14292 24206 14320 25230
rect 14476 24410 14504 25230
rect 14660 24993 14688 25230
rect 14646 24984 14702 24993
rect 14646 24919 14702 24928
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14476 24206 14504 24346
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14292 23866 14320 24142
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14476 23798 14504 24142
rect 14464 23792 14516 23798
rect 14464 23734 14516 23740
rect 14096 23724 14148 23730
rect 14096 23666 14148 23672
rect 14108 23633 14136 23666
rect 14094 23624 14150 23633
rect 14094 23559 14150 23568
rect 14660 23497 14688 24142
rect 14646 23488 14702 23497
rect 14646 23423 14702 23432
rect 14186 23216 14242 23225
rect 14186 23151 14242 23160
rect 14200 22642 14228 23151
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14188 22636 14240 22642
rect 14108 22596 14188 22624
rect 14108 21554 14136 22596
rect 14188 22578 14240 22584
rect 14292 22506 14320 22918
rect 14280 22500 14332 22506
rect 14280 22442 14332 22448
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14200 22234 14228 22374
rect 14292 22234 14320 22442
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14384 22166 14412 23054
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 14384 21690 14412 22102
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 14384 20806 14412 21422
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14004 20392 14056 20398
rect 14004 20334 14056 20340
rect 14016 19854 14044 20334
rect 14200 19854 14228 20742
rect 14004 19848 14056 19854
rect 14188 19848 14240 19854
rect 14056 19808 14136 19836
rect 14004 19790 14056 19796
rect 13924 19672 14044 19700
rect 13820 19654 13872 19660
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13556 17746 13584 19382
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16114 13492 16934
rect 13556 16590 13584 17478
rect 13634 17368 13690 17377
rect 13634 17303 13636 17312
rect 13688 17303 13690 17312
rect 13636 17274 13688 17280
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 17105 13676 17138
rect 13634 17096 13690 17105
rect 13634 17031 13690 17040
rect 13740 16697 13768 17750
rect 13832 17746 13860 18294
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13726 16688 13782 16697
rect 13726 16623 13782 16632
rect 13832 16590 13860 17682
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13924 16998 13952 17614
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16726 13952 16934
rect 14016 16794 14044 19672
rect 14108 18766 14136 19808
rect 14188 19790 14240 19796
rect 14186 19272 14242 19281
rect 14186 19207 14242 19216
rect 14096 18760 14148 18766
rect 14094 18728 14096 18737
rect 14148 18728 14150 18737
rect 14094 18663 14150 18672
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13556 16182 13584 16526
rect 13832 16250 13860 16526
rect 13910 16280 13966 16289
rect 13820 16244 13872 16250
rect 13910 16215 13966 16224
rect 13820 16186 13872 16192
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13726 16144 13782 16153
rect 13452 16108 13504 16114
rect 13924 16114 13952 16215
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13912 16108 13964 16114
rect 13726 16079 13782 16088
rect 13452 16050 13504 16056
rect 13372 15966 13584 15994
rect 13096 15694 13216 15722
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13004 15026 13032 15438
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 14618 12940 14894
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12912 14414 12940 14554
rect 13004 14414 13032 14962
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12808 14272 12860 14278
rect 13096 14226 13124 15574
rect 12808 14214 12860 14220
rect 12912 14198 13124 14226
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12268 10526 12388 10554
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11532 9646 11744 9674
rect 11808 9646 12020 9674
rect 11716 9586 11744 9646
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11532 8430 11560 8910
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11348 7942 11468 7970
rect 11348 7886 11376 7942
rect 11532 7886 11560 8366
rect 11992 7936 12020 9646
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12084 8634 12112 8842
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11992 7908 12112 7936
rect 11336 7880 11388 7886
rect 11520 7880 11572 7886
rect 11336 7822 11388 7828
rect 11440 7828 11520 7834
rect 11440 7822 11572 7828
rect 11440 7806 11560 7822
rect 11980 7812 12032 7818
rect 11440 6798 11468 7806
rect 11980 7754 12032 7760
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11532 7478 11560 7686
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11520 7472 11572 7478
rect 11624 7449 11652 7482
rect 11520 7414 11572 7420
rect 11610 7440 11666 7449
rect 11610 7375 11666 7384
rect 11808 7324 11836 7686
rect 11900 7478 11928 7686
rect 11992 7546 12020 7754
rect 12084 7546 12112 7908
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12072 7540 12124 7546
rect 12124 7500 12204 7528
rect 12072 7482 12124 7488
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11808 7296 12020 7324
rect 12084 7313 12112 7346
rect 11796 7200 11848 7206
rect 11794 7168 11796 7177
rect 11848 7168 11850 7177
rect 11794 7103 11850 7112
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11440 5778 11468 6734
rect 11704 6724 11756 6730
rect 11704 6666 11756 6672
rect 11716 6458 11744 6666
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11992 6322 12020 7296
rect 12070 7304 12126 7313
rect 12070 7239 12126 7248
rect 12084 6322 12112 7239
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11440 4554 11468 5714
rect 11900 5574 11928 6190
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4554 11560 4966
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 9876 3126 9904 3334
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 11348 2990 11376 4014
rect 11440 3534 11468 4490
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11440 3194 11468 3470
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11716 3194 11744 3402
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 11348 2514 11376 2926
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11900 2446 11928 5510
rect 11992 3058 12020 6258
rect 12176 5370 12204 7500
rect 12268 7177 12296 10526
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12360 10062 12388 10406
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12544 9586 12572 12650
rect 12912 12374 12940 14198
rect 13188 14090 13216 15694
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13096 14062 13216 14090
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 13004 12186 13032 13670
rect 13096 12646 13124 14062
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13188 13433 13216 13874
rect 13174 13424 13230 13433
rect 13174 13359 13230 13368
rect 13188 13326 13216 13359
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12636 12158 13032 12186
rect 12636 11014 12664 12158
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12728 10674 12756 12038
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12636 9450 12664 9998
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12530 7440 12586 7449
rect 12728 7410 12756 8978
rect 12820 8974 12848 11766
rect 12912 11150 12940 11834
rect 12992 11756 13044 11762
rect 13096 11744 13124 12582
rect 13188 11898 13216 12650
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13280 11762 13308 14826
rect 13372 13462 13400 15370
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13464 14618 13492 14894
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13938 13492 14214
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13372 12714 13400 13398
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13556 12434 13584 15966
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13648 13870 13676 14350
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13740 13394 13768 16079
rect 13832 16068 13912 16096
rect 13832 14958 13860 16068
rect 13912 16050 13964 16056
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13820 14952 13872 14958
rect 13818 14920 13820 14929
rect 13872 14920 13874 14929
rect 13818 14855 13874 14864
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13832 13938 13860 14350
rect 13924 14006 13952 15098
rect 14016 14822 14044 16118
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14108 14657 14136 18566
rect 14200 17338 14228 19207
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 14384 18426 14412 18634
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14094 14648 14150 14657
rect 14094 14583 14150 14592
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14108 13938 14136 14486
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13556 12406 13676 12434
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13044 11716 13124 11744
rect 13268 11756 13320 11762
rect 12992 11698 13044 11704
rect 13268 11698 13320 11704
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12990 11248 13046 11257
rect 13096 11218 13124 11562
rect 13464 11354 13492 12310
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13556 11286 13584 12038
rect 13648 11393 13676 12406
rect 13740 12294 14044 12322
rect 13740 12102 13768 12294
rect 14016 12238 14044 12294
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13740 11665 13768 11766
rect 13832 11694 13860 12174
rect 13820 11688 13872 11694
rect 13726 11656 13782 11665
rect 13820 11630 13872 11636
rect 13726 11591 13782 11600
rect 13634 11384 13690 11393
rect 13634 11319 13690 11328
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 12990 11183 13046 11192
rect 13084 11212 13136 11218
rect 13004 11150 13032 11183
rect 13084 11154 13136 11160
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12912 10713 12940 11086
rect 12898 10704 12954 10713
rect 12898 10639 12954 10648
rect 12912 9926 12940 10639
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12820 8566 12848 8910
rect 12808 8560 12860 8566
rect 12808 8502 12860 8508
rect 12716 7404 12768 7410
rect 12530 7375 12532 7384
rect 12584 7375 12586 7384
rect 12532 7346 12584 7352
rect 12636 7364 12716 7392
rect 12254 7168 12310 7177
rect 12254 7103 12310 7112
rect 12636 5846 12664 7364
rect 12716 7346 12768 7352
rect 13004 6866 13032 11086
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13280 10674 13308 10950
rect 13464 10674 13492 11154
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13280 10130 13308 10610
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13372 9926 13400 10474
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13464 9722 13492 9998
rect 13556 9994 13584 10406
rect 13924 10130 13952 10610
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 8566 13400 8774
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13450 8120 13506 8129
rect 13648 8090 13676 9522
rect 13450 8055 13452 8064
rect 13504 8055 13506 8064
rect 13636 8084 13688 8090
rect 13452 8026 13504 8032
rect 13636 8026 13688 8032
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13280 6390 13308 7278
rect 13464 7206 13492 8026
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13832 6866 13860 9862
rect 14016 9489 14044 12174
rect 14108 10674 14136 13330
rect 14200 12918 14228 16730
rect 14292 14804 14320 18090
rect 14476 17338 14504 22986
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14568 22166 14596 22442
rect 14556 22160 14608 22166
rect 14556 22102 14608 22108
rect 14568 22030 14596 22102
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14384 16153 14412 16186
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 14958 14412 15302
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14292 14776 14412 14804
rect 14278 14648 14334 14657
rect 14278 14583 14334 14592
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 9654 14228 10542
rect 14188 9648 14240 9654
rect 14094 9616 14150 9625
rect 14188 9590 14240 9596
rect 14094 9551 14150 9560
rect 14108 9518 14136 9551
rect 14096 9512 14148 9518
rect 14002 9480 14058 9489
rect 14096 9454 14148 9460
rect 14002 9415 14058 9424
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7410 13952 8230
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14016 7313 14044 7482
rect 14188 7336 14240 7342
rect 14002 7304 14058 7313
rect 14188 7278 14240 7284
rect 14002 7239 14058 7248
rect 14200 6934 14228 7278
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6390 13400 6598
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12176 4282 12204 5170
rect 12268 5166 12296 5646
rect 12820 5642 12848 6054
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12268 3738 12296 5102
rect 13096 4690 13124 6190
rect 13648 5778 13676 6734
rect 13740 5914 13768 6734
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 6254 14044 6598
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13832 5370 13860 5646
rect 14016 5574 14044 6190
rect 14292 5914 14320 14583
rect 14384 8820 14412 14776
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14476 13938 14504 14418
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14568 13818 14596 21490
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14660 20058 14688 20334
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14660 19310 14688 19790
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14660 17898 14688 19246
rect 14752 18057 14780 27406
rect 14844 26296 14872 28086
rect 15014 27568 15070 27577
rect 15014 27503 15070 27512
rect 14924 27464 14976 27470
rect 14924 27406 14976 27412
rect 14936 26586 14964 27406
rect 15028 27402 15056 27503
rect 15016 27396 15068 27402
rect 15016 27338 15068 27344
rect 15028 26926 15056 27338
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15014 26752 15070 26761
rect 15014 26687 15070 26696
rect 14924 26580 14976 26586
rect 14924 26522 14976 26528
rect 15028 26466 15056 26687
rect 14936 26450 15056 26466
rect 14924 26444 15056 26450
rect 14976 26438 15056 26444
rect 14924 26386 14976 26392
rect 14924 26308 14976 26314
rect 14844 26268 14924 26296
rect 14924 26250 14976 26256
rect 14936 22982 14964 26250
rect 15120 25786 15148 28966
rect 15292 28416 15344 28422
rect 15292 28358 15344 28364
rect 15028 25758 15148 25786
rect 15028 24138 15056 25758
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 15120 24886 15148 25638
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15108 24880 15160 24886
rect 15108 24822 15160 24828
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15212 23730 15240 25434
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15108 23248 15160 23254
rect 15108 23190 15160 23196
rect 14924 22976 14976 22982
rect 14924 22918 14976 22924
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 15028 22094 15056 22918
rect 14936 22066 15056 22094
rect 14936 21350 14964 22066
rect 15014 21720 15070 21729
rect 15014 21655 15070 21664
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14924 20868 14976 20874
rect 14924 20810 14976 20816
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14844 19854 14872 20742
rect 14936 19990 14964 20810
rect 14924 19984 14976 19990
rect 14924 19926 14976 19932
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14844 18222 14872 19654
rect 15028 18630 15056 21655
rect 15120 21554 15148 23190
rect 15212 23186 15240 23666
rect 15304 23662 15332 28358
rect 15396 27606 15424 29038
rect 15488 28994 15516 29106
rect 15672 29102 15700 29514
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15488 28966 15608 28994
rect 15384 27600 15436 27606
rect 15384 27542 15436 27548
rect 15580 27538 15608 28966
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 15580 26382 15608 27474
rect 15672 27402 15700 29038
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15948 28762 15976 28902
rect 15936 28756 15988 28762
rect 15936 28698 15988 28704
rect 15842 27704 15898 27713
rect 15842 27639 15898 27648
rect 15936 27668 15988 27674
rect 15856 27402 15884 27639
rect 15936 27610 15988 27616
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15844 27396 15896 27402
rect 15844 27338 15896 27344
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 15568 26376 15620 26382
rect 15568 26318 15620 26324
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15384 25424 15436 25430
rect 15384 25366 15436 25372
rect 15396 24954 15424 25366
rect 15488 25294 15516 25434
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15212 22778 15240 23122
rect 15396 23050 15424 24890
rect 15476 24608 15528 24614
rect 15580 24596 15608 26318
rect 15764 25906 15792 26930
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15672 24818 15700 25094
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15660 24608 15712 24614
rect 15580 24568 15660 24596
rect 15476 24550 15528 24556
rect 15660 24550 15712 24556
rect 15488 24342 15516 24550
rect 15476 24336 15528 24342
rect 15672 24313 15700 24550
rect 15476 24278 15528 24284
rect 15658 24304 15714 24313
rect 15658 24239 15714 24248
rect 15672 23866 15700 24239
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15660 23724 15712 23730
rect 15764 23712 15792 25842
rect 15856 24954 15884 26386
rect 15948 25906 15976 27610
rect 15936 25900 15988 25906
rect 15936 25842 15988 25848
rect 16040 25809 16068 31418
rect 16592 30433 16620 32778
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16684 31929 16712 32370
rect 16764 32224 16816 32230
rect 16764 32166 16816 32172
rect 16776 32026 16804 32166
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16868 31958 16896 32370
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 16856 31952 16908 31958
rect 16670 31920 16726 31929
rect 16856 31894 16908 31900
rect 16670 31855 16672 31864
rect 16724 31855 16726 31864
rect 16672 31826 16724 31832
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16868 31346 16896 31758
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16684 30734 16712 31078
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16578 30424 16634 30433
rect 16578 30359 16634 30368
rect 16684 29628 16712 30670
rect 16776 30666 16804 31078
rect 16960 30920 16988 32302
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17040 30932 17092 30938
rect 16960 30892 17040 30920
rect 17040 30874 17092 30880
rect 17144 30734 17172 31758
rect 17132 30728 17184 30734
rect 17132 30670 17184 30676
rect 16764 30660 16816 30666
rect 16764 30602 16816 30608
rect 17236 30580 17264 34138
rect 17328 33017 17356 34478
rect 17788 33998 17816 35634
rect 17880 35086 17908 35634
rect 18328 35488 18380 35494
rect 18328 35430 18380 35436
rect 18340 35086 18368 35430
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 18144 35080 18196 35086
rect 18144 35022 18196 35028
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18512 35080 18564 35086
rect 18512 35022 18564 35028
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17972 34202 18000 34614
rect 18156 34542 18184 35022
rect 18144 34536 18196 34542
rect 18144 34478 18196 34484
rect 18524 34490 18552 35022
rect 18616 34746 18644 35022
rect 19260 34746 19288 35770
rect 19352 35698 19380 36110
rect 19628 35698 19656 36178
rect 19904 36174 19932 36790
rect 19984 36712 20036 36718
rect 20180 36700 20208 36790
rect 20260 36712 20312 36718
rect 20180 36672 20260 36700
rect 19984 36654 20036 36660
rect 20260 36654 20312 36660
rect 19996 36378 20024 36654
rect 19984 36372 20036 36378
rect 19984 36314 20036 36320
rect 20364 36174 20392 36790
rect 20996 36236 21048 36242
rect 20996 36178 21048 36184
rect 19708 36168 19760 36174
rect 19708 36110 19760 36116
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 20352 36168 20404 36174
rect 20352 36110 20404 36116
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 19616 35692 19668 35698
rect 19616 35634 19668 35640
rect 19352 35086 19380 35634
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19628 34746 19656 35634
rect 19720 35630 19748 36110
rect 19904 36038 19932 36110
rect 19892 36032 19944 36038
rect 19892 35974 19944 35980
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 19708 35624 19760 35630
rect 19708 35566 19760 35572
rect 18604 34740 18656 34746
rect 18604 34682 18656 34688
rect 18972 34740 19024 34746
rect 18972 34682 19024 34688
rect 19248 34740 19300 34746
rect 19248 34682 19300 34688
rect 19616 34740 19668 34746
rect 19616 34682 19668 34688
rect 18984 34610 19012 34682
rect 18788 34604 18840 34610
rect 18788 34546 18840 34552
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 19064 34604 19116 34610
rect 19064 34546 19116 34552
rect 18524 34474 18644 34490
rect 18524 34468 18656 34474
rect 18524 34462 18604 34468
rect 18604 34410 18656 34416
rect 18420 34400 18472 34406
rect 18420 34342 18472 34348
rect 17960 34196 18012 34202
rect 17960 34138 18012 34144
rect 18328 34196 18380 34202
rect 18328 34138 18380 34144
rect 18340 34066 18368 34138
rect 18328 34060 18380 34066
rect 18328 34002 18380 34008
rect 18432 33998 18460 34342
rect 17592 33992 17644 33998
rect 17592 33934 17644 33940
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 18420 33992 18472 33998
rect 18420 33934 18472 33940
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 17500 33856 17552 33862
rect 17500 33798 17552 33804
rect 17314 33008 17370 33017
rect 17314 32943 17370 32952
rect 17328 32570 17356 32943
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17328 31822 17356 32506
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 17512 31686 17540 33798
rect 17604 33522 17632 33934
rect 17788 33658 17816 33934
rect 18524 33658 18552 33934
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 17592 33516 17644 33522
rect 17592 33458 17644 33464
rect 17788 32434 17816 33594
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 17868 32904 17920 32910
rect 17866 32872 17868 32881
rect 17920 32872 17922 32881
rect 17866 32807 17922 32816
rect 17776 32428 17828 32434
rect 17696 32388 17776 32416
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17604 31822 17632 32166
rect 17696 31958 17724 32388
rect 17776 32370 17828 32376
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17684 31952 17736 31958
rect 17684 31894 17736 31900
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17788 31754 17816 32234
rect 17868 31952 17920 31958
rect 17866 31920 17868 31929
rect 17920 31920 17922 31929
rect 17866 31855 17922 31864
rect 17972 31822 18000 32914
rect 18156 32910 18184 33254
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18144 32904 18196 32910
rect 18196 32864 18276 32892
rect 18144 32846 18196 32852
rect 18064 32337 18092 32846
rect 18144 32768 18196 32774
rect 18142 32736 18144 32745
rect 18196 32736 18198 32745
rect 18142 32671 18198 32680
rect 18050 32328 18106 32337
rect 18050 32263 18106 32272
rect 18144 32224 18196 32230
rect 18144 32166 18196 32172
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17776 31748 17828 31754
rect 17776 31690 17828 31696
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17328 30734 17356 31418
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 17512 30598 17540 31622
rect 18156 31414 18184 32166
rect 17684 31408 17736 31414
rect 17684 31350 17736 31356
rect 18144 31408 18196 31414
rect 18144 31350 18196 31356
rect 17696 31278 17724 31350
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17696 30938 17724 31214
rect 17684 30932 17736 30938
rect 17684 30874 17736 30880
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 17052 30552 17264 30580
rect 17500 30592 17552 30598
rect 16948 30116 17000 30122
rect 16948 30058 17000 30064
rect 16684 29600 16804 29628
rect 16212 29572 16264 29578
rect 16212 29514 16264 29520
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16132 28121 16160 29106
rect 16224 28490 16252 29514
rect 16304 29164 16356 29170
rect 16580 29164 16632 29170
rect 16356 29124 16580 29152
rect 16304 29106 16356 29112
rect 16580 29106 16632 29112
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 16118 28112 16174 28121
rect 16118 28047 16174 28056
rect 16224 27334 16252 28426
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16408 27538 16436 27814
rect 16592 27674 16620 28698
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 16396 27532 16448 27538
rect 16396 27474 16448 27480
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 16212 27328 16264 27334
rect 16396 27328 16448 27334
rect 16212 27270 16264 27276
rect 16394 27296 16396 27305
rect 16448 27296 16450 27305
rect 16224 26994 16252 27270
rect 16394 27231 16450 27240
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16488 26920 16540 26926
rect 16488 26862 16540 26868
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 16316 25906 16344 26182
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 16304 25900 16356 25906
rect 16304 25842 16356 25848
rect 16026 25800 16082 25809
rect 16026 25735 16082 25744
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 16040 24154 16068 25735
rect 15712 23684 15792 23712
rect 15856 24126 16068 24154
rect 16132 24138 16160 25842
rect 16396 25764 16448 25770
rect 16396 25706 16448 25712
rect 16408 25673 16436 25706
rect 16394 25664 16450 25673
rect 16394 25599 16450 25608
rect 16396 24404 16448 24410
rect 16396 24346 16448 24352
rect 16120 24132 16172 24138
rect 15660 23666 15712 23672
rect 15476 23656 15528 23662
rect 15476 23598 15528 23604
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15488 23322 15516 23598
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15384 23044 15436 23050
rect 15384 22986 15436 22992
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15488 22234 15516 23258
rect 15580 22964 15608 23598
rect 15672 23322 15700 23666
rect 15856 23662 15884 24126
rect 16120 24074 16172 24080
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 15844 23656 15896 23662
rect 15844 23598 15896 23604
rect 15936 23588 15988 23594
rect 15936 23530 15988 23536
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15672 23118 15700 23258
rect 15948 23254 15976 23530
rect 16040 23526 16068 24006
rect 16132 23798 16160 24074
rect 16408 23866 16436 24346
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16316 23594 16344 23666
rect 16304 23588 16356 23594
rect 16304 23530 16356 23536
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15580 22936 15700 22964
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 15474 21584 15530 21593
rect 15108 21548 15160 21554
rect 15474 21519 15530 21528
rect 15108 21490 15160 21496
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15016 18352 15068 18358
rect 15120 18340 15148 21490
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15200 20800 15252 20806
rect 15200 20742 15252 20748
rect 15212 20602 15240 20742
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 15304 20058 15332 21422
rect 15488 20942 15516 21519
rect 15580 21146 15608 22578
rect 15672 21434 15700 22936
rect 15764 22642 15792 23054
rect 15844 23044 15896 23050
rect 15844 22986 15896 22992
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15764 22166 15792 22578
rect 15856 22574 15884 22986
rect 15948 22642 15976 23190
rect 15936 22636 15988 22642
rect 15936 22578 15988 22584
rect 15844 22568 15896 22574
rect 15896 22516 15976 22522
rect 15844 22510 15976 22516
rect 15856 22494 15976 22510
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15948 22030 15976 22494
rect 16040 22098 16068 23462
rect 16408 23254 16436 23666
rect 16396 23248 16448 23254
rect 16396 23190 16448 23196
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16028 22092 16080 22098
rect 16028 22034 16080 22040
rect 16132 22030 16160 23054
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16316 22506 16344 22986
rect 16304 22500 16356 22506
rect 16304 22442 16356 22448
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15672 21406 15792 21434
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15580 20602 15608 20810
rect 15568 20596 15620 20602
rect 15488 20556 15568 20584
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15198 19952 15254 19961
rect 15198 19887 15254 19896
rect 15212 19854 15240 19887
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15068 18312 15148 18340
rect 15016 18294 15068 18300
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14738 18048 14794 18057
rect 14738 17983 14794 17992
rect 14660 17870 14780 17898
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14660 16726 14688 17546
rect 14752 17202 14780 17870
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14844 16946 14872 18158
rect 15304 18034 15332 19994
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15396 18057 15424 18634
rect 15212 18006 15332 18034
rect 15382 18048 15438 18057
rect 14924 17808 14976 17814
rect 15212 17762 15240 18006
rect 15382 17983 15438 17992
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 14924 17750 14976 17756
rect 14936 17678 14964 17750
rect 15120 17734 15240 17762
rect 15120 17678 15148 17734
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 14936 17066 14964 17478
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14660 16289 14688 16526
rect 14646 16280 14702 16289
rect 14646 16215 14702 16224
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14660 15026 14688 15642
rect 14752 15638 14780 16934
rect 14844 16918 14964 16946
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14844 15094 14872 15914
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14844 14822 14872 15030
rect 14648 14816 14700 14822
rect 14646 14784 14648 14793
rect 14740 14816 14792 14822
rect 14700 14784 14702 14793
rect 14740 14758 14792 14764
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14646 14719 14702 14728
rect 14660 14074 14688 14719
rect 14752 14550 14780 14758
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14752 13977 14780 14282
rect 14738 13968 14794 13977
rect 14844 13938 14872 14554
rect 14738 13903 14794 13912
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14568 13790 14780 13818
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12238 14596 12718
rect 14752 12442 14780 13790
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14660 12322 14688 12378
rect 14844 12322 14872 13874
rect 14936 12434 14964 16918
rect 15028 15706 15056 17478
rect 15120 17202 15148 17614
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15120 15042 15148 17002
rect 15212 16794 15240 17614
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15212 15094 15240 16390
rect 15028 15014 15148 15042
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15028 14414 15056 15014
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15120 14226 15148 14894
rect 15212 14414 15240 15030
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15028 13988 15056 14214
rect 15120 14198 15240 14226
rect 15108 14000 15160 14006
rect 15028 13960 15108 13988
rect 15108 13942 15160 13948
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15028 12850 15056 13194
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15212 12714 15240 14198
rect 15304 12986 15332 17818
rect 15384 17196 15436 17202
rect 15488 17184 15516 20556
rect 15568 20538 15620 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15580 19854 15608 20402
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15580 18034 15608 19790
rect 15672 18222 15700 21286
rect 15764 20806 15792 21406
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15764 20262 15792 20334
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 19786 15792 20198
rect 15752 19780 15804 19786
rect 15752 19722 15804 19728
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15580 18006 15792 18034
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15436 17156 15516 17184
rect 15384 17138 15436 17144
rect 15488 17066 15516 17156
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15396 16776 15424 17002
rect 15476 16788 15528 16794
rect 15396 16748 15476 16776
rect 15476 16730 15528 16736
rect 15580 16590 15608 17478
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15568 16108 15620 16114
rect 15672 16096 15700 17138
rect 15764 16726 15792 18006
rect 15856 17134 15884 21626
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16026 21312 16082 21321
rect 16026 21247 16082 21256
rect 16040 20806 16068 21247
rect 16224 21185 16252 21490
rect 16316 21418 16344 21898
rect 16304 21412 16356 21418
rect 16304 21354 16356 21360
rect 16210 21176 16266 21185
rect 16210 21111 16266 21120
rect 16224 21010 16252 21111
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16040 20466 16068 20742
rect 16132 20466 16160 20878
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16224 19334 16252 20946
rect 16408 20806 16436 23190
rect 16500 21690 16528 26862
rect 16592 26042 16620 27474
rect 16684 27470 16712 28018
rect 16776 27713 16804 29600
rect 16856 29572 16908 29578
rect 16856 29514 16908 29520
rect 16868 29238 16896 29514
rect 16856 29232 16908 29238
rect 16856 29174 16908 29180
rect 16854 28656 16910 28665
rect 16960 28626 16988 30058
rect 16854 28591 16856 28600
rect 16908 28591 16910 28600
rect 16948 28620 17000 28626
rect 16856 28562 16908 28568
rect 16948 28562 17000 28568
rect 16946 28520 17002 28529
rect 16946 28455 16948 28464
rect 17000 28455 17002 28464
rect 16948 28426 17000 28432
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16762 27704 16818 27713
rect 16762 27639 16818 27648
rect 16868 27577 16896 27814
rect 16854 27568 16910 27577
rect 16854 27503 16910 27512
rect 16868 27470 16896 27503
rect 16672 27464 16724 27470
rect 16764 27464 16816 27470
rect 16672 27406 16724 27412
rect 16762 27432 16764 27441
rect 16856 27464 16908 27470
rect 16816 27432 16818 27441
rect 16856 27406 16908 27412
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 16762 27367 16818 27376
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16684 26382 16712 26930
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 16578 25528 16634 25537
rect 16578 25463 16634 25472
rect 16592 25430 16620 25463
rect 16580 25424 16632 25430
rect 16580 25366 16632 25372
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16316 19854 16344 20470
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16592 19446 16620 25366
rect 16684 22574 16712 26318
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 25294 16804 26182
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16868 25129 16896 25162
rect 16854 25120 16910 25129
rect 16854 25055 16910 25064
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16776 23497 16804 24142
rect 16960 23866 16988 27406
rect 17052 25838 17080 30552
rect 17500 30534 17552 30540
rect 17880 30433 17908 30874
rect 17866 30424 17922 30433
rect 17866 30359 17922 30368
rect 17498 30288 17554 30297
rect 17498 30223 17554 30232
rect 17512 29850 17540 30223
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17224 29776 17276 29782
rect 17224 29718 17276 29724
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 17144 27334 17172 29038
rect 17236 28762 17264 29718
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17420 29034 17448 29650
rect 17696 29646 17724 30126
rect 17960 30116 18012 30122
rect 17960 30058 18012 30064
rect 17972 29782 18000 30058
rect 17960 29776 18012 29782
rect 17960 29718 18012 29724
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 17684 29640 17736 29646
rect 17684 29582 17736 29588
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 17512 29238 17540 29582
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17500 29232 17552 29238
rect 17500 29174 17552 29180
rect 17316 29028 17368 29034
rect 17316 28970 17368 28976
rect 17408 29028 17460 29034
rect 17408 28970 17460 28976
rect 17224 28756 17276 28762
rect 17224 28698 17276 28704
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17236 28393 17264 28494
rect 17222 28384 17278 28393
rect 17222 28319 17278 28328
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17236 27985 17264 28018
rect 17222 27976 17278 27985
rect 17222 27911 17278 27920
rect 17328 27656 17356 28970
rect 17408 28416 17460 28422
rect 17408 28358 17460 28364
rect 17420 28082 17448 28358
rect 17408 28076 17460 28082
rect 17408 28018 17460 28024
rect 17408 27668 17460 27674
rect 17328 27628 17408 27656
rect 17408 27610 17460 27616
rect 17420 27470 17448 27610
rect 17512 27606 17540 29174
rect 17604 28490 17632 29242
rect 17592 28484 17644 28490
rect 17592 28426 17644 28432
rect 17500 27600 17552 27606
rect 17500 27542 17552 27548
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17224 27328 17276 27334
rect 17328 27305 17356 27406
rect 17224 27270 17276 27276
rect 17314 27296 17370 27305
rect 17144 26382 17172 27270
rect 17236 26790 17264 27270
rect 17314 27231 17370 27240
rect 17420 26994 17448 27406
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 17052 25362 17080 25774
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 16948 23860 17000 23866
rect 16948 23802 17000 23808
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16762 23488 16818 23497
rect 16762 23423 16818 23432
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16776 22166 16804 22918
rect 16868 22642 16896 23054
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16684 19990 16712 21490
rect 16672 19984 16724 19990
rect 16672 19926 16724 19932
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16684 19378 16712 19926
rect 16132 19306 16252 19334
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 15948 18426 15976 18566
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15948 17338 15976 17818
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16040 16998 16068 18566
rect 16132 17610 16160 19306
rect 16500 18970 16528 19314
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16500 17746 16528 18906
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16592 18426 16620 18702
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16684 17814 16712 19314
rect 16868 18902 16896 22034
rect 16960 22030 16988 23666
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17052 21622 17080 24346
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 16960 21350 16988 21558
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 17052 20602 17080 21354
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17144 20058 17172 26318
rect 17236 24206 17264 26318
rect 17316 26240 17368 26246
rect 17420 26217 17448 26318
rect 17316 26182 17368 26188
rect 17406 26208 17462 26217
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17328 24154 17356 26182
rect 17406 26143 17462 26152
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17420 25378 17448 25842
rect 17512 25498 17540 26726
rect 17604 26450 17632 28426
rect 17696 28218 17724 29582
rect 17972 29306 18000 29582
rect 18064 29510 18092 31214
rect 18248 30870 18276 32864
rect 18236 30864 18288 30870
rect 18236 30806 18288 30812
rect 18144 30252 18196 30258
rect 18144 30194 18196 30200
rect 18156 29646 18184 30194
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 29646 18276 29990
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 18340 29510 18368 33050
rect 18524 33046 18552 33594
rect 18616 33590 18644 34410
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18800 33114 18828 34546
rect 19076 34377 19104 34546
rect 19156 34468 19208 34474
rect 19156 34410 19208 34416
rect 19062 34368 19118 34377
rect 19062 34303 19118 34312
rect 19064 34196 19116 34202
rect 19064 34138 19116 34144
rect 19076 34066 19104 34138
rect 19064 34060 19116 34066
rect 19064 34002 19116 34008
rect 19168 33153 19196 34410
rect 19720 34202 19748 35566
rect 19892 35488 19944 35494
rect 19892 35430 19944 35436
rect 19904 35154 19932 35430
rect 20088 35290 20116 35634
rect 20076 35284 20128 35290
rect 20076 35226 20128 35232
rect 19892 35148 19944 35154
rect 19892 35090 19944 35096
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 19708 34196 19760 34202
rect 19708 34138 19760 34144
rect 19432 33924 19484 33930
rect 19432 33866 19484 33872
rect 19800 33924 19852 33930
rect 19800 33866 19852 33872
rect 19340 33856 19392 33862
rect 19338 33824 19340 33833
rect 19392 33824 19394 33833
rect 19338 33759 19394 33768
rect 19444 33425 19472 33866
rect 19812 33833 19840 33866
rect 19798 33824 19854 33833
rect 19798 33759 19854 33768
rect 19430 33416 19486 33425
rect 19430 33351 19486 33360
rect 19154 33144 19210 33153
rect 18788 33108 18840 33114
rect 19154 33079 19210 33088
rect 18788 33050 18840 33056
rect 18512 33040 18564 33046
rect 18512 32982 18564 32988
rect 19432 33040 19484 33046
rect 19432 32982 19484 32988
rect 18788 32972 18840 32978
rect 18788 32914 18840 32920
rect 19156 32972 19208 32978
rect 19156 32914 19208 32920
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 18694 32872 18750 32881
rect 18432 32570 18460 32846
rect 18694 32807 18696 32816
rect 18748 32807 18750 32816
rect 18696 32778 18748 32784
rect 18604 32768 18656 32774
rect 18604 32710 18656 32716
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 18616 32230 18644 32710
rect 18696 32564 18748 32570
rect 18696 32506 18748 32512
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18604 31408 18656 31414
rect 18604 31350 18656 31356
rect 18616 30258 18644 31350
rect 18708 31210 18736 32506
rect 18800 32502 18828 32914
rect 18972 32904 19024 32910
rect 18972 32846 19024 32852
rect 18880 32768 18932 32774
rect 18878 32736 18880 32745
rect 18932 32736 18934 32745
rect 18878 32671 18934 32680
rect 18788 32496 18840 32502
rect 18788 32438 18840 32444
rect 18984 32026 19012 32846
rect 18972 32020 19024 32026
rect 18972 31962 19024 31968
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 19076 31906 19104 31962
rect 18892 31890 19104 31906
rect 18880 31884 19104 31890
rect 18932 31878 19104 31884
rect 18880 31826 18932 31832
rect 18892 31754 18920 31826
rect 18880 31748 18932 31754
rect 18880 31690 18932 31696
rect 18892 31482 18920 31690
rect 18880 31476 18932 31482
rect 18880 31418 18932 31424
rect 19168 31414 19196 32914
rect 19248 31952 19300 31958
rect 19248 31894 19300 31900
rect 19156 31408 19208 31414
rect 19156 31350 19208 31356
rect 19260 31278 19288 31894
rect 19340 31680 19392 31686
rect 19340 31622 19392 31628
rect 19352 31346 19380 31622
rect 19444 31482 19472 32982
rect 19524 32224 19576 32230
rect 19524 32166 19576 32172
rect 19536 31822 19564 32166
rect 19996 31822 20024 34682
rect 20260 33924 20312 33930
rect 20364 33912 20392 36110
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20456 35834 20484 35974
rect 20444 35828 20496 35834
rect 20444 35770 20496 35776
rect 20720 35760 20772 35766
rect 20720 35702 20772 35708
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20640 34950 20668 35566
rect 20732 34950 20760 35702
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20812 34196 20864 34202
rect 20812 34138 20864 34144
rect 20824 33998 20852 34138
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20312 33884 20392 33912
rect 20260 33866 20312 33872
rect 20076 32292 20128 32298
rect 20076 32234 20128 32240
rect 20088 31822 20116 32234
rect 19524 31816 19576 31822
rect 19524 31758 19576 31764
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 20076 31816 20128 31822
rect 20076 31758 20128 31764
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 19432 31340 19484 31346
rect 19536 31328 19564 31758
rect 19892 31748 19944 31754
rect 19892 31690 19944 31696
rect 19904 31482 19932 31690
rect 19996 31686 20024 31758
rect 19984 31680 20036 31686
rect 19984 31622 20036 31628
rect 19892 31476 19944 31482
rect 19892 31418 19944 31424
rect 19996 31414 20024 31622
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 19484 31300 19564 31328
rect 19892 31340 19944 31346
rect 19432 31282 19484 31288
rect 19892 31282 19944 31288
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 18696 31204 18748 31210
rect 18696 31146 18748 31152
rect 19904 30666 19932 31282
rect 20088 31210 20116 31758
rect 20076 31204 20128 31210
rect 20076 31146 20128 31152
rect 19892 30660 19944 30666
rect 19892 30602 19944 30608
rect 19904 30394 19932 30602
rect 19892 30388 19944 30394
rect 19892 30330 19944 30336
rect 18788 30320 18840 30326
rect 18788 30262 18840 30268
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 18432 29714 18460 30126
rect 18420 29708 18472 29714
rect 18420 29650 18472 29656
rect 18524 29578 18552 30194
rect 18800 29850 18828 30262
rect 19892 30184 19944 30190
rect 20088 30172 20116 31146
rect 20272 30326 20300 33866
rect 20904 33584 20956 33590
rect 20904 33526 20956 33532
rect 20916 33318 20944 33526
rect 20904 33312 20956 33318
rect 20904 33254 20956 33260
rect 21008 32858 21036 36178
rect 21180 34128 21232 34134
rect 21180 34070 21232 34076
rect 21192 33114 21220 34070
rect 21180 33108 21232 33114
rect 21180 33050 21232 33056
rect 20536 32836 20588 32842
rect 20536 32778 20588 32784
rect 20732 32830 21036 32858
rect 20548 32570 20576 32778
rect 20732 32774 20760 32830
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20812 32768 20864 32774
rect 20812 32710 20864 32716
rect 20824 32586 20852 32710
rect 20536 32564 20588 32570
rect 20536 32506 20588 32512
rect 20732 32558 20852 32586
rect 20444 32496 20496 32502
rect 20732 32450 20760 32558
rect 20496 32444 20760 32450
rect 20444 32438 20760 32444
rect 20456 32422 20760 32438
rect 20812 32428 20864 32434
rect 20812 32370 20864 32376
rect 20904 32428 20956 32434
rect 21008 32416 21036 32830
rect 20956 32388 21036 32416
rect 20904 32370 20956 32376
rect 20628 32224 20680 32230
rect 20628 32166 20680 32172
rect 20640 31958 20668 32166
rect 20824 32026 20852 32370
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 20720 31476 20772 31482
rect 20720 31418 20772 31424
rect 20352 30388 20404 30394
rect 20352 30330 20404 30336
rect 20260 30320 20312 30326
rect 20260 30262 20312 30268
rect 19944 30144 20116 30172
rect 19892 30126 19944 30132
rect 18604 29844 18656 29850
rect 18604 29786 18656 29792
rect 18788 29844 18840 29850
rect 18788 29786 18840 29792
rect 19892 29844 19944 29850
rect 19892 29786 19944 29792
rect 18512 29572 18564 29578
rect 18512 29514 18564 29520
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 18524 29238 18552 29514
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18236 29096 18288 29102
rect 18236 29038 18288 29044
rect 17868 29028 17920 29034
rect 17868 28970 17920 28976
rect 18144 29028 18196 29034
rect 18144 28970 18196 28976
rect 17776 28552 17828 28558
rect 17774 28520 17776 28529
rect 17828 28520 17830 28529
rect 17774 28455 17830 28464
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17684 28212 17736 28218
rect 17684 28154 17736 28160
rect 17682 28112 17738 28121
rect 17682 28047 17738 28056
rect 17696 26466 17724 28047
rect 17788 26926 17816 28358
rect 17880 27334 17908 28970
rect 18052 28552 18104 28558
rect 17972 28512 18052 28540
rect 17972 28121 18000 28512
rect 18052 28494 18104 28500
rect 18156 28257 18184 28970
rect 18142 28248 18198 28257
rect 18052 28212 18104 28218
rect 18142 28183 18198 28192
rect 18052 28154 18104 28160
rect 17958 28112 18014 28121
rect 18064 28082 18092 28154
rect 17958 28047 18014 28056
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17788 26586 17816 26726
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17592 26444 17644 26450
rect 17696 26438 17816 26466
rect 17592 26386 17644 26392
rect 17684 26308 17736 26314
rect 17604 26268 17684 26296
rect 17604 25906 17632 26268
rect 17684 26250 17736 26256
rect 17788 26217 17816 26438
rect 17774 26208 17830 26217
rect 17774 26143 17830 26152
rect 17788 25974 17816 26143
rect 17776 25968 17828 25974
rect 17776 25910 17828 25916
rect 17880 25906 17908 27270
rect 17592 25900 17644 25906
rect 17592 25842 17644 25848
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17420 25350 17540 25378
rect 17512 25158 17540 25350
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17420 24954 17448 25094
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17236 22642 17264 24142
rect 17328 24126 17448 24154
rect 17604 24138 17632 25842
rect 17776 25832 17828 25838
rect 17776 25774 17828 25780
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17696 24206 17724 24754
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 23730 17356 24006
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17224 22636 17276 22642
rect 17224 22578 17276 22584
rect 17420 22098 17448 24126
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17788 24018 17816 25774
rect 17880 25702 17908 25842
rect 17868 25696 17920 25702
rect 17868 25638 17920 25644
rect 17880 25498 17908 25638
rect 17868 25492 17920 25498
rect 17868 25434 17920 25440
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17604 23990 17816 24018
rect 17604 23100 17632 23990
rect 17684 23656 17736 23662
rect 17736 23616 17816 23644
rect 17684 23598 17736 23604
rect 17684 23112 17736 23118
rect 17604 23072 17684 23100
rect 17604 22642 17632 23072
rect 17684 23054 17736 23060
rect 17788 23050 17816 23616
rect 17880 23322 17908 24754
rect 17972 24614 18000 27814
rect 18064 27470 18092 28018
rect 18144 27940 18196 27946
rect 18144 27882 18196 27888
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18064 27130 18092 27406
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 18156 26858 18184 27882
rect 18248 27402 18276 29038
rect 18420 29028 18472 29034
rect 18420 28970 18472 28976
rect 18432 28762 18460 28970
rect 18420 28756 18472 28762
rect 18420 28698 18472 28704
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 18420 28076 18472 28082
rect 18420 28018 18472 28024
rect 18340 27606 18368 28018
rect 18432 27674 18460 28018
rect 18616 27690 18644 29786
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18708 28014 18736 29650
rect 19904 29170 19932 29786
rect 20364 29288 20392 30330
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20180 29260 20392 29288
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 18880 28484 18932 28490
rect 18880 28426 18932 28432
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18420 27668 18472 27674
rect 18420 27610 18472 27616
rect 18524 27662 18644 27690
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 18236 27396 18288 27402
rect 18236 27338 18288 27344
rect 18248 26858 18276 27338
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18144 26852 18196 26858
rect 18144 26794 18196 26800
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18052 26784 18104 26790
rect 18156 26761 18184 26794
rect 18052 26726 18104 26732
rect 18142 26752 18198 26761
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17972 23769 18000 23802
rect 17958 23760 18014 23769
rect 18064 23730 18092 26726
rect 18142 26687 18198 26696
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 18156 25838 18184 26250
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18248 25430 18276 25910
rect 18236 25424 18288 25430
rect 18142 25392 18198 25401
rect 18236 25366 18288 25372
rect 18142 25327 18198 25336
rect 18156 25226 18184 25327
rect 18144 25220 18196 25226
rect 18144 25162 18196 25168
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18156 24274 18184 24550
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18340 23730 18368 26930
rect 17958 23695 18014 23704
rect 18052 23724 18104 23730
rect 18328 23724 18380 23730
rect 18052 23666 18104 23672
rect 18248 23684 18328 23712
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 18144 23180 18196 23186
rect 18144 23122 18196 23128
rect 17776 23044 17828 23050
rect 17776 22986 17828 22992
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17408 21616 17460 21622
rect 17222 21584 17278 21593
rect 17408 21558 17460 21564
rect 17222 21519 17224 21528
rect 17276 21519 17278 21528
rect 17316 21548 17368 21554
rect 17224 21490 17276 21496
rect 17316 21490 17368 21496
rect 17328 21418 17356 21490
rect 17316 21412 17368 21418
rect 17316 21354 17368 21360
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 20330 17264 20878
rect 17224 20324 17276 20330
rect 17224 20266 17276 20272
rect 17420 20233 17448 21558
rect 17498 20904 17554 20913
rect 17498 20839 17500 20848
rect 17552 20839 17554 20848
rect 17592 20868 17644 20874
rect 17500 20810 17552 20816
rect 17592 20810 17644 20816
rect 17604 20754 17632 20810
rect 17512 20726 17632 20754
rect 17406 20224 17462 20233
rect 17406 20159 17462 20168
rect 17132 20052 17184 20058
rect 17132 19994 17184 20000
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17236 19514 17264 19790
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17420 19310 17448 20159
rect 17512 19854 17540 20726
rect 17592 20596 17644 20602
rect 17592 20538 17644 20544
rect 17500 19848 17552 19854
rect 17604 19825 17632 20538
rect 17500 19790 17552 19796
rect 17590 19816 17646 19825
rect 17590 19751 17646 19760
rect 17604 19446 17632 19751
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 16868 18766 16896 18838
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 16132 17270 16160 17546
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 16132 17134 16160 17206
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15752 16720 15804 16726
rect 15752 16662 15804 16668
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15620 16068 15700 16096
rect 15568 16050 15620 16056
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15502 15424 15846
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15488 15366 15516 15642
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15580 15201 15608 16050
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15764 15366 15792 15438
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15566 15192 15622 15201
rect 15672 15162 15700 15302
rect 15750 15192 15806 15201
rect 15566 15127 15622 15136
rect 15660 15156 15712 15162
rect 15750 15127 15806 15136
rect 15660 15098 15712 15104
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15396 13938 15424 14826
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15488 14074 15516 14554
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15488 12850 15516 13806
rect 15580 13802 15608 14894
rect 15672 14414 15700 14962
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15672 13530 15700 14350
rect 15764 14113 15792 15127
rect 15856 14890 15884 15438
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15750 14104 15806 14113
rect 15750 14039 15806 14048
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15672 12850 15700 13126
rect 15764 12986 15792 13466
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15476 12844 15528 12850
rect 15396 12804 15476 12832
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15212 12594 15240 12650
rect 15120 12566 15240 12594
rect 15120 12434 15148 12566
rect 15200 12436 15252 12442
rect 14936 12406 15056 12434
rect 15120 12406 15200 12434
rect 14660 12294 14872 12322
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14660 11898 14688 12106
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 14844 11694 14872 12294
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14752 10674 14780 11630
rect 14936 11014 14964 12174
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14556 8832 14608 8838
rect 14384 8792 14556 8820
rect 14556 8774 14608 8780
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14476 7818 14504 8434
rect 14464 7812 14516 7818
rect 14464 7754 14516 7760
rect 14476 6662 14504 7754
rect 14568 7750 14596 8774
rect 14660 8498 14688 10474
rect 14832 10056 14884 10062
rect 14884 10016 14964 10044
rect 14832 9998 14884 10004
rect 14936 9926 14964 10016
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14752 9586 14780 9862
rect 15028 9738 15056 12406
rect 15200 12378 15252 12384
rect 15396 11830 15424 12804
rect 15476 12786 15528 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15488 11286 15516 12174
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 14844 9710 15056 9738
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14844 9058 14872 9710
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 15014 9616 15070 9625
rect 14752 9030 14872 9058
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14752 8430 14780 9030
rect 14936 8974 14964 9590
rect 15014 9551 15070 9560
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14844 8537 14872 8842
rect 14830 8528 14886 8537
rect 14830 8463 14886 8472
rect 14844 8430 14872 8463
rect 14936 8430 14964 8910
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14832 8424 14884 8430
rect 14832 8366 14884 8372
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14752 8294 14780 8366
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 14016 5302 14044 5510
rect 14108 5302 14136 5510
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4078 13032 4422
rect 13188 4214 13216 4490
rect 13176 4208 13228 4214
rect 13176 4150 13228 4156
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12268 3602 12296 3674
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12268 2990 12296 3538
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 3194 12756 3334
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12820 2922 12848 3470
rect 12808 2916 12860 2922
rect 12808 2858 12860 2864
rect 13004 2446 13032 4014
rect 13084 3528 13136 3534
rect 13188 3516 13216 4150
rect 13832 3942 13860 4558
rect 14016 4554 14044 5238
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13136 3488 13216 3516
rect 13084 3470 13136 3476
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13464 3126 13492 3334
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13648 2446 13676 3538
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13740 3126 13768 3470
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13832 2446 13860 3878
rect 14568 3602 14596 7686
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14660 4554 14688 4966
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14752 4146 14780 8026
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 14844 7177 14872 7754
rect 14936 7546 14964 7754
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14830 7168 14886 7177
rect 14830 7103 14886 7112
rect 14844 6202 14872 7103
rect 14936 6322 14964 7482
rect 15028 6390 15056 9551
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 8838 15148 9454
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15198 9208 15254 9217
rect 15198 9143 15200 9152
rect 15252 9143 15254 9152
rect 15200 9114 15252 9120
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15108 8288 15160 8294
rect 15108 8230 15160 8236
rect 15120 7886 15148 8230
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15106 7712 15162 7721
rect 15106 7647 15162 7656
rect 15120 7478 15148 7647
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15120 7206 15148 7278
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15212 6866 15240 8570
rect 15304 7886 15332 9318
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7002 15332 7686
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14844 6174 14964 6202
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14660 2650 14688 3402
rect 14648 2644 14700 2650
rect 14648 2586 14700 2592
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 11624 800 11652 2246
rect 12268 800 12296 2246
rect 12912 800 12940 2246
rect 13556 800 13584 2246
rect 14200 800 14228 2246
rect 14844 800 14872 5510
rect 14936 5166 14964 6174
rect 15212 5794 15240 6802
rect 15212 5766 15332 5794
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15212 4690 15240 5646
rect 15304 5302 15332 5766
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15304 4690 15332 5238
rect 15396 5166 15424 11018
rect 15580 9586 15608 12786
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12442 15700 12582
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15764 11762 15792 12650
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15672 9518 15700 11494
rect 15856 11286 15884 14826
rect 15948 14550 15976 16526
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 14074 15976 14282
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16040 13326 16068 16934
rect 16224 16794 16252 17614
rect 16408 17134 16436 17682
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16224 16561 16252 16730
rect 16210 16552 16266 16561
rect 16120 16516 16172 16522
rect 16210 16487 16266 16496
rect 16120 16458 16172 16464
rect 16132 16250 16160 16458
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16224 16114 16252 16390
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16224 15502 16252 16050
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16132 15026 16160 15302
rect 16224 15162 16252 15302
rect 16316 15162 16344 15370
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16224 14770 16252 15098
rect 16408 15094 16436 15642
rect 16500 15638 16528 17682
rect 16684 17202 16712 17750
rect 16762 17368 16818 17377
rect 16762 17303 16818 17312
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16776 16182 16804 17303
rect 16960 16522 16988 19110
rect 17224 18896 17276 18902
rect 17130 18864 17186 18873
rect 17224 18838 17276 18844
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 17130 18799 17132 18808
rect 17184 18799 17186 18808
rect 17132 18770 17184 18776
rect 17236 18766 17264 18838
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 17052 17202 17080 17478
rect 17144 17202 17172 17546
rect 17328 17202 17356 18838
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17132 17196 17184 17202
rect 17316 17196 17368 17202
rect 17184 17156 17264 17184
rect 17132 17138 17184 17144
rect 17052 17066 17080 17138
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16684 15570 16712 15982
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16408 14793 16436 15030
rect 16580 14816 16632 14822
rect 16132 14742 16252 14770
rect 16394 14784 16450 14793
rect 16132 14278 16160 14742
rect 16580 14758 16632 14764
rect 16394 14719 16450 14728
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16132 12850 16160 14214
rect 16224 13326 16252 14554
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 16040 9722 16068 12786
rect 16132 12434 16160 12786
rect 16316 12646 16344 14350
rect 16408 13938 16436 14350
rect 16592 14346 16620 14758
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16592 14006 16620 14282
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16578 13832 16634 13841
rect 16578 13767 16634 13776
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16408 12434 16436 13631
rect 16132 12406 16252 12434
rect 16224 12238 16252 12406
rect 16316 12406 16528 12434
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16132 11898 16160 12174
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16224 10606 16252 11086
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16224 10266 16252 10542
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16210 10160 16266 10169
rect 16210 10095 16266 10104
rect 16224 10062 16252 10095
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15948 8974 15976 9522
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15842 7984 15898 7993
rect 16040 7954 16068 8230
rect 15842 7919 15898 7928
rect 16028 7948 16080 7954
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15764 7546 15792 7686
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15764 7342 15792 7482
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15856 6322 15884 7919
rect 16028 7890 16080 7896
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5778 15516 6054
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 4282 14964 4422
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 15212 3602 15240 4626
rect 15304 4214 15332 4626
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15304 3126 15332 4150
rect 15396 4078 15424 5102
rect 15856 4146 15884 6258
rect 16132 4826 16160 9114
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16224 8498 16252 8842
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16224 4486 16252 5102
rect 16316 5030 16344 12406
rect 16500 12238 16528 12406
rect 16592 12238 16620 13767
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16408 10962 16436 12106
rect 16684 11830 16712 15506
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16776 13802 16804 14962
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16672 11824 16724 11830
rect 16486 11792 16542 11801
rect 16672 11766 16724 11772
rect 16486 11727 16542 11736
rect 16500 11150 16528 11727
rect 16684 11558 16712 11766
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16762 11248 16818 11257
rect 16868 11218 16896 16390
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16960 13705 16988 16118
rect 17052 15638 17080 16526
rect 17144 15706 17172 16730
rect 17236 16572 17264 17156
rect 17316 17138 17368 17144
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16794 17356 16934
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17316 16584 17368 16590
rect 17236 16544 17316 16572
rect 17316 16526 17368 16532
rect 17224 16448 17276 16454
rect 17222 16416 17224 16425
rect 17276 16416 17278 16425
rect 17222 16351 17278 16360
rect 17420 16114 17448 18702
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17512 17610 17540 18362
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17604 17542 17632 18022
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17604 16833 17632 17478
rect 17590 16824 17646 16833
rect 17590 16759 17646 16768
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17512 16250 17540 16526
rect 17696 16454 17724 22714
rect 17788 22642 17816 22986
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17788 21146 17816 22578
rect 18064 22030 18092 22918
rect 18156 22574 18184 23122
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18156 22166 18184 22374
rect 18144 22160 18196 22166
rect 18144 22102 18196 22108
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17788 20602 17816 21082
rect 17880 20913 17908 21490
rect 17866 20904 17922 20913
rect 17866 20839 17922 20848
rect 17868 20800 17920 20806
rect 17972 20777 18000 21966
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18064 21010 18092 21490
rect 18156 21146 18184 21966
rect 18248 21729 18276 23684
rect 18328 23666 18380 23672
rect 18432 23526 18460 27270
rect 18524 27062 18552 27662
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18708 25702 18736 27542
rect 18892 27334 18920 28426
rect 19168 28218 19196 28902
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 18972 28008 19024 28014
rect 18970 27976 18972 27985
rect 19024 27976 19026 27985
rect 18970 27911 19026 27920
rect 19444 27470 19472 29106
rect 19996 28994 20024 29106
rect 19904 28966 20024 28994
rect 19708 28552 19760 28558
rect 19760 28512 19840 28540
rect 19708 28494 19760 28500
rect 19706 28248 19762 28257
rect 19706 28183 19762 28192
rect 19524 27872 19576 27878
rect 19524 27814 19576 27820
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 18880 27328 18932 27334
rect 18880 27270 18932 27276
rect 18892 26246 18920 27270
rect 19260 27062 19288 27338
rect 19444 27305 19472 27406
rect 19430 27296 19486 27305
rect 19430 27231 19486 27240
rect 19248 27056 19300 27062
rect 19248 26998 19300 27004
rect 19536 26994 19564 27814
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 18880 26240 18932 26246
rect 18880 26182 18932 26188
rect 19524 26036 19576 26042
rect 19524 25978 19576 25984
rect 18788 25900 18840 25906
rect 19064 25900 19116 25906
rect 18840 25860 18920 25888
rect 18788 25842 18840 25848
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18524 24818 18552 25230
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18708 24750 18736 25638
rect 18892 25294 18920 25860
rect 19064 25842 19116 25848
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18892 24954 18920 25230
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 18708 23730 18736 24550
rect 18696 23724 18748 23730
rect 18524 23684 18696 23712
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18234 21720 18290 21729
rect 18234 21655 18290 21664
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18248 21026 18276 21490
rect 18340 21350 18368 22578
rect 18524 22506 18552 23684
rect 18696 23666 18748 23672
rect 18788 23724 18840 23730
rect 18788 23666 18840 23672
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18616 23254 18644 23530
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18604 23248 18656 23254
rect 18604 23190 18656 23196
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18616 22012 18644 23190
rect 18524 21984 18644 22012
rect 18418 21856 18474 21865
rect 18418 21791 18474 21800
rect 18432 21486 18460 21791
rect 18420 21480 18472 21486
rect 18420 21422 18472 21428
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18340 21146 18368 21286
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18420 21072 18472 21078
rect 18248 21020 18420 21026
rect 18248 21014 18472 21020
rect 18052 21004 18104 21010
rect 18248 20998 18460 21014
rect 18052 20946 18104 20952
rect 17868 20742 17920 20748
rect 17958 20768 18014 20777
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17880 20448 17908 20742
rect 17958 20703 18014 20712
rect 18064 20466 18092 20946
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18328 20936 18380 20942
rect 18524 20924 18552 21984
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18380 20896 18552 20924
rect 18328 20878 18380 20884
rect 17788 20420 17908 20448
rect 18052 20460 18104 20466
rect 17788 18766 17816 20420
rect 18052 20402 18104 20408
rect 18064 20058 18092 20402
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18156 19990 18184 20878
rect 18248 20602 18276 20878
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 18144 19984 18196 19990
rect 18144 19926 18196 19932
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 19378 17908 19790
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17880 19145 17908 19314
rect 17972 19310 18000 19926
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 17866 19136 17922 19145
rect 17866 19071 17922 19080
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17880 17678 17908 19071
rect 17958 18456 18014 18465
rect 17958 18391 18014 18400
rect 17972 18290 18000 18391
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17880 16590 17908 17070
rect 17972 17066 18000 17614
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17958 16552 18014 16561
rect 17776 16516 17828 16522
rect 17958 16487 17960 16496
rect 17776 16458 17828 16464
rect 18012 16487 18014 16496
rect 17960 16458 18012 16464
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17408 16108 17460 16114
rect 17696 16096 17724 16186
rect 17460 16068 17724 16096
rect 17408 16050 17460 16056
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17040 15632 17092 15638
rect 17420 15586 17448 16050
rect 17040 15574 17092 15580
rect 17328 15558 17448 15586
rect 17590 15600 17646 15609
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 16946 13696 17002 13705
rect 16946 13631 17002 13640
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12306 16988 12582
rect 17052 12345 17080 14418
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17038 12336 17094 12345
rect 16948 12300 17000 12306
rect 17038 12271 17094 12280
rect 16948 12242 17000 12248
rect 17052 12238 17080 12271
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16960 11694 16988 12106
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17144 11626 17172 12174
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16762 11183 16818 11192
rect 16856 11212 16908 11218
rect 16776 11150 16804 11183
rect 16856 11154 16908 11160
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16764 11144 16816 11150
rect 16816 11092 16896 11098
rect 16764 11086 16896 11092
rect 16776 11070 16896 11086
rect 16408 10934 16528 10962
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16408 9586 16436 10134
rect 16500 10130 16528 10934
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16592 10266 16620 10678
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16684 9674 16712 10066
rect 16776 10033 16804 10406
rect 16762 10024 16818 10033
rect 16762 9959 16818 9968
rect 16684 9646 16804 9674
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16776 9489 16804 9646
rect 16762 9480 16818 9489
rect 16762 9415 16764 9424
rect 16816 9415 16818 9424
rect 16764 9386 16816 9392
rect 16868 9330 16896 11070
rect 16776 9302 16896 9330
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16592 7750 16620 7822
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6322 16712 7142
rect 16776 6798 16804 9302
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16868 8090 16896 8230
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16868 7392 16896 8026
rect 16960 7818 16988 11494
rect 17130 11248 17186 11257
rect 17130 11183 17186 11192
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17052 9518 17080 11086
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16948 7404 17000 7410
rect 16868 7364 16948 7392
rect 16868 7274 16896 7364
rect 16948 7346 17000 7352
rect 17052 7274 17080 8774
rect 17144 7886 17172 11183
rect 17236 10470 17264 14214
rect 17328 13841 17356 15558
rect 17590 15535 17646 15544
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17314 13832 17370 13841
rect 17314 13767 17370 13776
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 12986 17356 13670
rect 17420 13569 17448 15438
rect 17604 14958 17632 15535
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17406 13560 17462 13569
rect 17512 13530 17540 14826
rect 17788 14822 17816 16458
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17776 14816 17828 14822
rect 17590 14784 17646 14793
rect 17776 14758 17828 14764
rect 17590 14719 17646 14728
rect 17604 14550 17632 14719
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17592 14408 17644 14414
rect 17590 14376 17592 14385
rect 17644 14376 17646 14385
rect 17590 14311 17646 14320
rect 17696 14006 17724 14486
rect 17788 14074 17816 14758
rect 17880 14346 17908 16118
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15434 18000 16050
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15026 18000 15370
rect 18064 15065 18092 19722
rect 18144 19372 18196 19378
rect 18248 19360 18276 20538
rect 18340 19514 18368 20878
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18524 20369 18552 20470
rect 18510 20360 18566 20369
rect 18510 20295 18566 20304
rect 18512 20052 18564 20058
rect 18512 19994 18564 20000
rect 18524 19854 18552 19994
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18524 19378 18552 19790
rect 18196 19332 18276 19360
rect 18328 19372 18380 19378
rect 18144 19314 18196 19320
rect 18512 19372 18564 19378
rect 18380 19332 18460 19360
rect 18328 19314 18380 19320
rect 18142 19272 18198 19281
rect 18142 19207 18144 19216
rect 18196 19207 18198 19216
rect 18236 19236 18288 19242
rect 18144 19178 18196 19184
rect 18236 19178 18288 19184
rect 18248 18816 18276 19178
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18970 18368 19110
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18156 18788 18276 18816
rect 18156 18358 18184 18788
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18248 17814 18276 18090
rect 18236 17808 18288 17814
rect 18236 17750 18288 17756
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18156 17610 18184 17682
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 18156 16833 18184 17546
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18142 16824 18198 16833
rect 18142 16759 18198 16768
rect 18142 15600 18198 15609
rect 18142 15535 18144 15544
rect 18196 15535 18198 15544
rect 18144 15506 18196 15512
rect 18142 15328 18198 15337
rect 18142 15263 18198 15272
rect 18050 15056 18106 15065
rect 17960 15020 18012 15026
rect 18050 14991 18106 15000
rect 17960 14962 18012 14968
rect 18156 14890 18184 15263
rect 18248 15162 18276 17138
rect 18340 15162 18368 18906
rect 18432 18290 18460 19332
rect 18512 19314 18564 19320
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18432 17796 18460 18226
rect 18524 18154 18552 19314
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18512 17808 18564 17814
rect 18432 17768 18512 17796
rect 18512 17750 18564 17756
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18432 15065 18460 17478
rect 18524 17105 18552 17478
rect 18510 17096 18566 17105
rect 18510 17031 18566 17040
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 18524 16114 18552 16458
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18234 15056 18290 15065
rect 18234 14991 18236 15000
rect 18288 14991 18290 15000
rect 18418 15056 18474 15065
rect 18524 15026 18552 15506
rect 18418 14991 18474 15000
rect 18512 15020 18564 15026
rect 18236 14962 18288 14968
rect 18512 14962 18564 14968
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18156 14742 18552 14770
rect 18156 14414 18184 14742
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18340 14498 18368 14554
rect 18420 14544 18472 14550
rect 18340 14492 18420 14498
rect 18340 14486 18472 14492
rect 18340 14470 18460 14486
rect 18144 14408 18196 14414
rect 18328 14408 18380 14414
rect 18144 14350 18196 14356
rect 18326 14376 18328 14385
rect 18380 14376 18382 14385
rect 17868 14340 17920 14346
rect 17960 14340 18012 14346
rect 17920 14300 17960 14328
rect 17868 14282 17920 14288
rect 18012 14300 18092 14328
rect 18326 14311 18382 14320
rect 17960 14282 18012 14288
rect 18064 14260 18092 14300
rect 18524 14278 18552 14742
rect 18328 14272 18380 14278
rect 17958 14240 18014 14249
rect 18064 14232 18276 14260
rect 17958 14175 18014 14184
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17684 14000 17736 14006
rect 17868 14000 17920 14006
rect 17684 13942 17736 13948
rect 17788 13948 17868 13954
rect 17788 13942 17920 13948
rect 17788 13926 17908 13942
rect 17406 13495 17462 13504
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17604 13190 17632 13398
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17406 13016 17462 13025
rect 17316 12980 17368 12986
rect 17406 12951 17462 12960
rect 17316 12922 17368 12928
rect 17316 12844 17368 12850
rect 17420 12832 17448 12951
rect 17368 12804 17448 12832
rect 17316 12786 17368 12792
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17328 12442 17356 12650
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17314 12064 17370 12073
rect 17314 11999 17370 12008
rect 17328 11150 17356 11999
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17222 10160 17278 10169
rect 17328 10146 17356 10610
rect 17512 10266 17540 13126
rect 17788 12850 17816 13926
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17880 13326 17908 13738
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17774 12744 17830 12753
rect 17774 12679 17830 12688
rect 17788 12434 17816 12679
rect 17604 12406 17816 12434
rect 17500 10260 17552 10266
rect 17278 10118 17356 10146
rect 17420 10220 17500 10248
rect 17222 10095 17224 10104
rect 17276 10095 17278 10104
rect 17224 10066 17276 10072
rect 17316 10056 17368 10062
rect 17314 10024 17316 10033
rect 17368 10024 17370 10033
rect 17314 9959 17370 9968
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17328 8906 17356 9590
rect 17420 9178 17448 10220
rect 17500 10202 17552 10208
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17420 8974 17448 9114
rect 17512 9110 17540 9318
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17604 9058 17632 12406
rect 17880 12102 17908 12786
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11830 17908 12038
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17972 11354 18000 14175
rect 18050 13560 18106 13569
rect 18050 13495 18052 13504
rect 18104 13495 18106 13504
rect 18052 13466 18104 13472
rect 18050 13424 18106 13433
rect 18050 13359 18052 13368
rect 18104 13359 18106 13368
rect 18052 13330 18104 13336
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12442 18092 12786
rect 18156 12714 18184 13194
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18156 12238 18184 12650
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17972 10962 18000 11290
rect 18064 11150 18092 11630
rect 18156 11354 18184 11698
rect 18248 11354 18276 14232
rect 18328 14214 18380 14220
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18340 14074 18368 14214
rect 18418 14104 18474 14113
rect 18328 14068 18380 14074
rect 18418 14039 18474 14048
rect 18328 14010 18380 14016
rect 18326 13424 18382 13433
rect 18326 13359 18382 13368
rect 18340 13326 18368 13359
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18432 13190 18460 14039
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18432 12288 18460 13126
rect 18616 12986 18644 21830
rect 18708 17660 18736 23462
rect 18800 22778 18828 23666
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 18800 22030 18828 22442
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18800 21350 18828 21490
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18786 21176 18842 21185
rect 18892 21146 18920 24890
rect 18984 24818 19012 25366
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18970 24304 19026 24313
rect 19076 24274 19104 25842
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19156 25764 19208 25770
rect 19156 25706 19208 25712
rect 18970 24239 19026 24248
rect 19064 24268 19116 24274
rect 18984 23662 19012 24239
rect 19064 24210 19116 24216
rect 19062 24032 19118 24041
rect 19062 23967 19118 23976
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 18972 23316 19024 23322
rect 18972 23258 19024 23264
rect 18984 23118 19012 23258
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18984 22642 19012 23054
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 19076 22506 19104 23967
rect 19168 23798 19196 25706
rect 19444 25498 19472 25774
rect 19432 25492 19484 25498
rect 19432 25434 19484 25440
rect 19444 24886 19472 25434
rect 19536 25294 19564 25978
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 19522 24848 19578 24857
rect 19522 24783 19578 24792
rect 19536 24750 19564 24783
rect 19524 24744 19576 24750
rect 19524 24686 19576 24692
rect 19628 24698 19656 27814
rect 19720 27538 19748 28183
rect 19708 27532 19760 27538
rect 19708 27474 19760 27480
rect 19708 27396 19760 27402
rect 19708 27338 19760 27344
rect 19720 26994 19748 27338
rect 19708 26988 19760 26994
rect 19708 26930 19760 26936
rect 19708 25900 19760 25906
rect 19812 25888 19840 28512
rect 19904 28082 19932 28966
rect 19892 28076 19944 28082
rect 19892 28018 19944 28024
rect 19904 26994 19932 28018
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 19760 25860 19840 25888
rect 19708 25842 19760 25848
rect 19720 24857 19748 25842
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19812 25294 19840 25638
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19706 24848 19762 24857
rect 19904 24818 19932 26930
rect 19996 26489 20024 27270
rect 20076 26852 20128 26858
rect 20076 26794 20128 26800
rect 19982 26480 20038 26489
rect 20088 26450 20116 26794
rect 19982 26415 20038 26424
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 19984 25832 20036 25838
rect 19982 25800 19984 25809
rect 20036 25800 20038 25809
rect 19982 25735 20038 25744
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19706 24783 19762 24792
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19260 23662 19288 24618
rect 19432 24336 19484 24342
rect 19432 24278 19484 24284
rect 19536 24290 19564 24686
rect 19628 24670 19840 24698
rect 19628 24614 19656 24670
rect 19812 24614 19840 24670
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19708 24608 19760 24614
rect 19708 24550 19760 24556
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19720 24410 19748 24550
rect 19708 24404 19760 24410
rect 19708 24346 19760 24352
rect 19892 24336 19944 24342
rect 19444 24138 19472 24278
rect 19536 24262 19748 24290
rect 19892 24278 19944 24284
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19524 24064 19576 24070
rect 19524 24006 19576 24012
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19168 23225 19196 23462
rect 19260 23338 19288 23598
rect 19340 23520 19392 23526
rect 19338 23488 19340 23497
rect 19392 23488 19394 23497
rect 19338 23423 19394 23432
rect 19260 23310 19380 23338
rect 19154 23216 19210 23225
rect 19154 23151 19210 23160
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19260 23089 19288 23122
rect 19246 23080 19302 23089
rect 19156 23044 19208 23050
rect 19246 23015 19302 23024
rect 19156 22986 19208 22992
rect 19168 22778 19196 22986
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 19260 22710 19288 22918
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 18972 22160 19024 22166
rect 18972 22102 19024 22108
rect 18786 21111 18842 21120
rect 18880 21140 18932 21146
rect 18800 20874 18828 21111
rect 18880 21082 18932 21088
rect 18984 20942 19012 22102
rect 19168 21434 19196 22442
rect 19260 22273 19288 22510
rect 19246 22264 19302 22273
rect 19246 22199 19302 22208
rect 19352 22094 19380 23310
rect 19536 23118 19564 24006
rect 19628 23769 19656 24142
rect 19614 23760 19670 23769
rect 19614 23695 19670 23704
rect 19614 23624 19670 23633
rect 19614 23559 19670 23568
rect 19628 23526 19656 23559
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19432 23112 19484 23118
rect 19430 23080 19432 23089
rect 19524 23112 19576 23118
rect 19484 23080 19486 23089
rect 19720 23066 19748 24262
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19812 23662 19840 24006
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19904 23594 19932 24278
rect 19892 23588 19944 23594
rect 19892 23530 19944 23536
rect 19904 23186 19932 23530
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19524 23054 19576 23060
rect 19430 23015 19486 23024
rect 19628 23038 19748 23066
rect 19628 22438 19656 23038
rect 19708 22976 19760 22982
rect 19708 22918 19760 22924
rect 19800 22976 19852 22982
rect 19800 22918 19852 22924
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19352 22066 19564 22094
rect 19432 22024 19484 22030
rect 19430 21992 19432 22001
rect 19484 21992 19486 22001
rect 19430 21927 19486 21936
rect 19340 21888 19392 21894
rect 19260 21836 19340 21842
rect 19260 21830 19392 21836
rect 19260 21814 19380 21830
rect 19260 21622 19288 21814
rect 19430 21720 19486 21729
rect 19352 21664 19430 21672
rect 19352 21644 19432 21664
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19076 21406 19196 21434
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18788 20868 18840 20874
rect 18788 20810 18840 20816
rect 18788 20528 18840 20534
rect 18786 20496 18788 20505
rect 18840 20496 18842 20505
rect 18786 20431 18842 20440
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 18800 19378 18828 20266
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18800 18290 18828 19314
rect 18892 18426 18920 19314
rect 18984 18834 19012 20878
rect 19076 20466 19104 21406
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19168 20097 19196 21286
rect 19246 21040 19302 21049
rect 19246 20975 19248 20984
rect 19300 20975 19302 20984
rect 19248 20946 19300 20952
rect 19352 20942 19380 21644
rect 19484 21655 19486 21664
rect 19432 21626 19484 21632
rect 19536 21486 19564 22066
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 21185 19472 21286
rect 19430 21176 19486 21185
rect 19536 21146 19564 21422
rect 19430 21111 19486 21120
rect 19524 21140 19576 21146
rect 19340 20936 19392 20942
rect 19246 20904 19302 20913
rect 19340 20878 19392 20884
rect 19246 20839 19302 20848
rect 19154 20088 19210 20097
rect 19154 20023 19210 20032
rect 19260 19446 19288 20839
rect 19444 20262 19472 21111
rect 19524 21082 19576 21088
rect 19628 21049 19656 21626
rect 19720 21570 19748 22918
rect 19812 22642 19840 22918
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19720 21542 19840 21570
rect 19812 21400 19840 21542
rect 19720 21372 19840 21400
rect 19614 21040 19670 21049
rect 19614 20975 19670 20984
rect 19720 20942 19748 21372
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19338 19680 19394 19689
rect 19338 19615 19394 19624
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18800 18154 18828 18226
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 18878 17776 18934 17785
rect 18878 17711 18934 17720
rect 18892 17678 18920 17711
rect 18788 17672 18840 17678
rect 18708 17632 18788 17660
rect 18788 17614 18840 17620
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18878 17504 18934 17513
rect 18878 17439 18934 17448
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18708 16182 18736 16526
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18708 13530 18736 16118
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 15706 18828 15982
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14414 18828 14962
rect 18892 14521 18920 17439
rect 18984 16590 19012 18634
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 19076 16232 19104 19314
rect 19248 19304 19300 19310
rect 19246 19272 19248 19281
rect 19300 19272 19302 19281
rect 19246 19207 19302 19216
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19154 18456 19210 18465
rect 19154 18391 19210 18400
rect 19168 18358 19196 18391
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19168 17134 19196 18090
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19168 16522 19196 16934
rect 19260 16794 19288 18702
rect 19352 17610 19380 19615
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19444 18970 19472 19450
rect 19536 19378 19564 20878
rect 19628 20641 19656 20878
rect 19614 20632 19670 20641
rect 19614 20567 19670 20576
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19720 20233 19748 20334
rect 19706 20224 19762 20233
rect 19706 20159 19762 20168
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19628 18970 19656 19994
rect 19812 19825 19840 21082
rect 19798 19816 19854 19825
rect 19798 19751 19800 19760
rect 19852 19751 19854 19760
rect 19800 19722 19852 19728
rect 19708 19712 19760 19718
rect 19708 19654 19760 19660
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19720 18834 19748 19654
rect 19708 18828 19760 18834
rect 19760 18788 19840 18816
rect 19708 18770 19760 18776
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19536 18630 19564 18702
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19432 18624 19484 18630
rect 19430 18592 19432 18601
rect 19524 18624 19576 18630
rect 19484 18592 19486 18601
rect 19524 18566 19576 18572
rect 19430 18527 19486 18536
rect 19536 18358 19564 18566
rect 19524 18352 19576 18358
rect 19524 18294 19576 18300
rect 19720 18290 19748 18634
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19352 16998 19380 17138
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19156 16244 19208 16250
rect 19076 16204 19156 16232
rect 19156 16186 19208 16192
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19260 16153 19288 16186
rect 19246 16144 19302 16153
rect 18972 16108 19024 16114
rect 19246 16079 19302 16088
rect 18972 16050 19024 16056
rect 18984 15609 19012 16050
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 18970 15600 19026 15609
rect 18970 15535 19026 15544
rect 19062 15192 19118 15201
rect 19168 15162 19196 15982
rect 19352 15910 19380 16934
rect 19444 16590 19472 18090
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19444 15570 19472 16050
rect 19536 15638 19564 18022
rect 19812 17785 19840 18788
rect 19798 17776 19854 17785
rect 19798 17711 19854 17720
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19812 17202 19840 17478
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19062 15127 19064 15136
rect 19116 15127 19118 15136
rect 19156 15156 19208 15162
rect 19064 15098 19116 15104
rect 19156 15098 19208 15104
rect 19156 15020 19208 15026
rect 19156 14962 19208 14968
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18878 14512 18934 14521
rect 18878 14447 18934 14456
rect 18984 14414 19012 14758
rect 19062 14648 19118 14657
rect 19062 14583 19064 14592
rect 19116 14583 19118 14592
rect 19064 14554 19116 14560
rect 18788 14408 18840 14414
rect 18786 14376 18788 14385
rect 18880 14408 18932 14414
rect 18840 14376 18842 14385
rect 18880 14350 18932 14356
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18786 14311 18842 14320
rect 18788 14272 18840 14278
rect 18786 14240 18788 14249
rect 18840 14240 18842 14249
rect 18786 14175 18842 14184
rect 18892 14006 18920 14350
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18984 13870 19012 14350
rect 19168 14278 19196 14962
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19260 14550 19288 14826
rect 19352 14657 19380 14894
rect 19338 14648 19394 14657
rect 19338 14583 19394 14592
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 14074 19196 14214
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19444 14006 19472 15370
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19432 14000 19484 14006
rect 19338 13968 19394 13977
rect 19432 13942 19484 13948
rect 19338 13903 19394 13912
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 19352 13734 19380 13903
rect 19340 13728 19392 13734
rect 18878 13696 18934 13705
rect 19340 13670 19392 13676
rect 18878 13631 18934 13640
rect 18696 13524 18748 13530
rect 18696 13466 18748 13472
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18708 12442 18736 13466
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18604 12300 18656 12306
rect 18432 12260 18552 12288
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18432 11830 18460 12106
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18524 11694 18552 12260
rect 18604 12242 18656 12248
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18512 11552 18564 11558
rect 18326 11520 18382 11529
rect 18512 11494 18564 11500
rect 18326 11455 18382 11464
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18340 11150 18368 11455
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 17682 10296 17738 10305
rect 17788 10266 17816 10950
rect 17880 10742 17908 10950
rect 17972 10934 18092 10962
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17682 10231 17684 10240
rect 17736 10231 17738 10240
rect 17776 10260 17828 10266
rect 17684 10202 17736 10208
rect 17776 10202 17828 10208
rect 17972 9994 18000 10678
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17866 9208 17922 9217
rect 17866 9143 17922 9152
rect 17880 9110 17908 9143
rect 17868 9104 17920 9110
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17328 8090 17356 8842
rect 17420 8362 17448 8910
rect 17512 8498 17540 9046
rect 17604 9030 17816 9058
rect 17868 9046 17920 9052
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17604 8378 17632 8910
rect 17696 8634 17724 8910
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17512 8362 17632 8378
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17500 8356 17632 8362
rect 17552 8350 17632 8356
rect 17684 8356 17736 8362
rect 17500 8298 17552 8304
rect 17684 8298 17736 8304
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17696 7886 17724 8298
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 16856 7268 16908 7274
rect 16856 7210 16908 7216
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 17144 6866 17172 7822
rect 17314 7440 17370 7449
rect 17788 7410 17816 9030
rect 17972 8430 18000 9658
rect 18064 8498 18092 10934
rect 18524 10810 18552 11494
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18144 9988 18196 9994
rect 18144 9930 18196 9936
rect 18156 9722 18184 9930
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9217 18184 9318
rect 18142 9208 18198 9217
rect 18142 9143 18198 9152
rect 18052 8492 18104 8498
rect 18248 8480 18276 9658
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18340 8974 18368 9522
rect 18432 8974 18460 10066
rect 18524 9586 18552 10746
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18616 9382 18644 12242
rect 18892 12170 18920 13631
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18984 12306 19012 12378
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 19168 12170 19196 13194
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19260 12442 19288 12786
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19352 12306 19380 13466
rect 19432 13320 19484 13326
rect 19536 13308 19564 14962
rect 19484 13297 19564 13308
rect 19484 13288 19578 13297
rect 19484 13280 19522 13288
rect 19432 13262 19484 13268
rect 19522 13223 19578 13232
rect 19524 13184 19576 13190
rect 19430 13152 19486 13161
rect 19524 13126 19576 13132
rect 19430 13087 19486 13096
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 19062 11928 19118 11937
rect 19062 11863 19118 11872
rect 19076 11830 19104 11863
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18708 10198 18736 10542
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18708 9722 18736 10134
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18604 9376 18656 9382
rect 18524 9336 18604 9364
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18432 8566 18460 8910
rect 18524 8906 18552 9336
rect 18604 9318 18656 9324
rect 18602 9208 18658 9217
rect 18602 9143 18604 9152
rect 18656 9143 18658 9152
rect 18604 9114 18656 9120
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18616 8498 18644 8910
rect 18708 8634 18736 9522
rect 18800 8906 18828 11018
rect 18878 10704 18934 10713
rect 18878 10639 18934 10648
rect 18892 10198 18920 10639
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18892 9353 18920 9386
rect 18878 9344 18934 9353
rect 18878 9279 18934 9288
rect 18984 9042 19012 9522
rect 19076 9382 19104 11290
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18328 8492 18380 8498
rect 18248 8452 18328 8480
rect 18052 8434 18104 8440
rect 18328 8434 18380 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 18800 7478 18828 8842
rect 19076 8090 19104 8842
rect 19168 8566 19196 12106
rect 19352 11558 19380 12242
rect 19444 12102 19472 13087
rect 19536 12782 19564 13126
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11552 19392 11558
rect 19246 11520 19302 11529
rect 19340 11494 19392 11500
rect 19246 11455 19302 11464
rect 19260 11354 19288 11455
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19338 11248 19394 11257
rect 19338 11183 19340 11192
rect 19392 11183 19394 11192
rect 19340 11154 19392 11160
rect 19444 11150 19472 11698
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10810 19472 11086
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19338 10432 19394 10441
rect 19338 10367 19394 10376
rect 19352 9994 19380 10367
rect 19444 10062 19472 10610
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19444 9586 19472 9998
rect 19536 9761 19564 12718
rect 19628 11694 19656 17138
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19720 16522 19748 17002
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19706 16144 19762 16153
rect 19706 16079 19708 16088
rect 19760 16079 19762 16088
rect 19708 16050 19760 16056
rect 19812 15978 19840 16526
rect 19904 15978 19932 22578
rect 19996 18426 20024 25230
rect 20088 23118 20116 26386
rect 20180 26382 20208 29260
rect 20456 29238 20484 29582
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20260 29028 20312 29034
rect 20260 28970 20312 28976
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24313 20208 24754
rect 20166 24304 20222 24313
rect 20166 24239 20222 24248
rect 20180 24070 20208 24239
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20272 23746 20300 28970
rect 20364 28490 20392 29106
rect 20456 28762 20484 29174
rect 20640 29170 20668 29446
rect 20628 29164 20680 29170
rect 20628 29106 20680 29112
rect 20628 28960 20680 28966
rect 20628 28902 20680 28908
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 20640 28014 20668 28902
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20536 27328 20588 27334
rect 20536 27270 20588 27276
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20456 26790 20484 26930
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20456 26314 20484 26726
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 20364 24750 20392 25978
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20352 24744 20404 24750
rect 20352 24686 20404 24692
rect 20364 24206 20392 24686
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20272 23718 20392 23746
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 20272 23497 20300 23530
rect 20364 23526 20392 23718
rect 20352 23520 20404 23526
rect 20258 23488 20314 23497
rect 20352 23462 20404 23468
rect 20258 23423 20314 23432
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20088 21894 20116 22578
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20180 21729 20208 22578
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20272 22234 20300 22374
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20260 21888 20312 21894
rect 20364 21865 20392 23054
rect 20260 21830 20312 21836
rect 20350 21856 20406 21865
rect 20166 21720 20222 21729
rect 20166 21655 20222 21664
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20088 20466 20116 20878
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20534 20208 20810
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20076 20256 20128 20262
rect 20074 20224 20076 20233
rect 20128 20224 20130 20233
rect 20074 20159 20130 20168
rect 20180 20058 20208 20470
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20076 19168 20128 19174
rect 20272 19156 20300 21830
rect 20456 21842 20484 25230
rect 20548 24041 20576 27270
rect 20626 26208 20682 26217
rect 20732 26194 20760 31418
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20824 30870 20852 31282
rect 21008 30938 21036 31758
rect 21284 31754 21312 39039
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 22284 37392 22336 37398
rect 22284 37334 22336 37340
rect 22100 36032 22152 36038
rect 22100 35974 22152 35980
rect 21640 35760 21692 35766
rect 21640 35702 21692 35708
rect 21456 35692 21508 35698
rect 21456 35634 21508 35640
rect 21364 35624 21416 35630
rect 21364 35566 21416 35572
rect 21376 35018 21404 35566
rect 21468 35222 21496 35634
rect 21456 35216 21508 35222
rect 21456 35158 21508 35164
rect 21364 35012 21416 35018
rect 21364 34954 21416 34960
rect 21548 35012 21600 35018
rect 21548 34954 21600 34960
rect 21560 34610 21588 34954
rect 21548 34604 21600 34610
rect 21548 34546 21600 34552
rect 21652 34134 21680 35702
rect 22112 35680 22140 35974
rect 22192 35692 22244 35698
rect 22020 35652 22192 35680
rect 22020 35086 22048 35652
rect 22192 35634 22244 35640
rect 22100 35488 22152 35494
rect 22100 35430 22152 35436
rect 22192 35488 22244 35494
rect 22192 35430 22244 35436
rect 21916 35080 21968 35086
rect 21744 35040 21916 35068
rect 21744 34678 21772 35040
rect 21916 35022 21968 35028
rect 22008 35080 22060 35086
rect 22008 35022 22060 35028
rect 21732 34672 21784 34678
rect 21732 34614 21784 34620
rect 21916 34672 21968 34678
rect 21916 34614 21968 34620
rect 21640 34128 21692 34134
rect 21640 34070 21692 34076
rect 21928 33998 21956 34614
rect 22008 34536 22060 34542
rect 22008 34478 22060 34484
rect 21732 33992 21784 33998
rect 21732 33934 21784 33940
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 21548 33924 21600 33930
rect 21548 33866 21600 33872
rect 21560 33590 21588 33866
rect 21548 33584 21600 33590
rect 21548 33526 21600 33532
rect 21744 33454 21772 33934
rect 22020 33658 22048 34478
rect 22008 33652 22060 33658
rect 22008 33594 22060 33600
rect 21916 33584 21968 33590
rect 21916 33526 21968 33532
rect 21732 33448 21784 33454
rect 21362 33416 21418 33425
rect 21732 33390 21784 33396
rect 21822 33416 21878 33425
rect 21362 33351 21418 33360
rect 21822 33351 21824 33360
rect 21376 31822 21404 33351
rect 21876 33351 21878 33360
rect 21824 33322 21876 33328
rect 21732 33108 21784 33114
rect 21732 33050 21784 33056
rect 21744 32570 21772 33050
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21640 32564 21692 32570
rect 21640 32506 21692 32512
rect 21732 32564 21784 32570
rect 21732 32506 21784 32512
rect 21652 32434 21680 32506
rect 21640 32428 21692 32434
rect 21640 32370 21692 32376
rect 21456 32224 21508 32230
rect 21456 32166 21508 32172
rect 21468 31822 21496 32166
rect 21652 31822 21680 32370
rect 21732 32360 21784 32366
rect 21836 32348 21864 32710
rect 21784 32320 21864 32348
rect 21732 32302 21784 32308
rect 21928 32178 21956 33526
rect 22020 32434 22048 33594
rect 22112 32552 22140 35430
rect 22204 35018 22232 35430
rect 22192 35012 22244 35018
rect 22192 34954 22244 34960
rect 22204 34746 22232 34954
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 22204 34513 22232 34546
rect 22190 34504 22246 34513
rect 22190 34439 22246 34448
rect 22192 33856 22244 33862
rect 22192 33798 22244 33804
rect 22204 33318 22232 33798
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 22112 32524 22232 32552
rect 22204 32434 22232 32524
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 21744 32150 21956 32178
rect 21364 31816 21416 31822
rect 21364 31758 21416 31764
rect 21456 31816 21508 31822
rect 21456 31758 21508 31764
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21088 31748 21140 31754
rect 21088 31690 21140 31696
rect 21192 31726 21312 31754
rect 21548 31748 21600 31754
rect 21100 30938 21128 31690
rect 20996 30932 21048 30938
rect 20996 30874 21048 30880
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20812 30864 20864 30870
rect 20812 30806 20864 30812
rect 21192 30190 21220 31726
rect 21548 31690 21600 31696
rect 21364 31340 21416 31346
rect 21364 31282 21416 31288
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21272 31136 21324 31142
rect 21272 31078 21324 31084
rect 21284 30734 21312 31078
rect 21376 30802 21404 31282
rect 21468 31142 21496 31282
rect 21560 31278 21588 31690
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21456 31136 21508 31142
rect 21456 31078 21508 31084
rect 21468 30870 21496 31078
rect 21456 30864 21508 30870
rect 21456 30806 21508 30812
rect 21364 30796 21416 30802
rect 21364 30738 21416 30744
rect 21272 30728 21324 30734
rect 21272 30670 21324 30676
rect 21376 30297 21404 30738
rect 21362 30288 21418 30297
rect 21362 30223 21418 30232
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21640 29640 21692 29646
rect 21640 29582 21692 29588
rect 20916 29170 20944 29582
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21100 29073 21128 29106
rect 21086 29064 21142 29073
rect 21086 28999 21142 29008
rect 20902 28928 20958 28937
rect 20902 28863 20958 28872
rect 20916 28558 20944 28863
rect 21192 28626 21220 29106
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21284 28626 21312 28970
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 21272 28620 21324 28626
rect 21272 28562 21324 28568
rect 20904 28552 20956 28558
rect 20904 28494 20956 28500
rect 20916 27606 20944 28494
rect 21180 28484 21232 28490
rect 21180 28426 21232 28432
rect 21086 28248 21142 28257
rect 21086 28183 21142 28192
rect 21100 28082 21128 28183
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21192 27606 21220 28426
rect 20904 27600 20956 27606
rect 21180 27600 21232 27606
rect 20904 27542 20956 27548
rect 21008 27560 21180 27588
rect 20810 27296 20866 27305
rect 20810 27231 20866 27240
rect 20682 26166 20760 26194
rect 20626 26143 20682 26152
rect 20626 24984 20682 24993
rect 20626 24919 20682 24928
rect 20640 24818 20668 24919
rect 20824 24886 20852 27231
rect 20916 26994 20944 27542
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20916 24993 20944 26930
rect 21008 26586 21036 27560
rect 21180 27542 21232 27548
rect 21284 27470 21312 28562
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21364 28416 21416 28422
rect 21364 28358 21416 28364
rect 21376 27470 21404 28358
rect 21468 27470 21496 28494
rect 21548 28076 21600 28082
rect 21548 28018 21600 28024
rect 21560 27878 21588 28018
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21364 27464 21416 27470
rect 21364 27406 21416 27412
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21456 27328 21508 27334
rect 21456 27270 21508 27276
rect 21468 27130 21496 27270
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21548 27056 21600 27062
rect 21548 26998 21600 27004
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 21100 26314 21128 26930
rect 21560 26790 21588 26998
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 21088 26308 21140 26314
rect 21088 26250 21140 26256
rect 20902 24984 20958 24993
rect 20902 24919 20958 24928
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20628 24132 20680 24138
rect 20628 24074 20680 24080
rect 20534 24032 20590 24041
rect 20534 23967 20590 23976
rect 20536 23180 20588 23186
rect 20536 23122 20588 23128
rect 20548 22710 20576 23122
rect 20536 22704 20588 22710
rect 20536 22646 20588 22652
rect 20640 22438 20668 24074
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20640 22098 20668 22374
rect 20628 22092 20680 22098
rect 20628 22034 20680 22040
rect 20456 21814 20668 21842
rect 20350 21791 20406 21800
rect 20364 21554 20392 21791
rect 20442 21720 20498 21729
rect 20442 21655 20498 21664
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20456 21486 20484 21655
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20352 21344 20404 21350
rect 20444 21344 20496 21350
rect 20352 21286 20404 21292
rect 20442 21312 20444 21321
rect 20496 21312 20498 21321
rect 20364 20806 20392 21286
rect 20442 21247 20498 21256
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20128 19128 20300 19156
rect 20076 19110 20128 19116
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20088 18086 20116 19110
rect 20364 18834 20392 20402
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20456 18714 20484 21247
rect 20548 21146 20576 21490
rect 20640 21350 20668 21814
rect 20732 21690 20760 24754
rect 21192 23254 21220 26454
rect 21456 26308 21508 26314
rect 21456 26250 21508 26256
rect 21364 25424 21416 25430
rect 21364 25366 21416 25372
rect 21376 25294 21404 25366
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21376 24750 21404 25230
rect 21364 24744 21416 24750
rect 21364 24686 21416 24692
rect 21468 24614 21496 26250
rect 21546 25936 21602 25945
rect 21546 25871 21602 25880
rect 21560 25770 21588 25871
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21376 23633 21404 24550
rect 21560 23866 21588 24550
rect 21652 23866 21680 29582
rect 21744 28762 21772 32150
rect 22112 31414 22140 32370
rect 22204 31958 22232 32370
rect 22296 32065 22324 37334
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 26608 36916 26660 36922
rect 26608 36858 26660 36864
rect 23204 36712 23256 36718
rect 23204 36654 23256 36660
rect 24584 36712 24636 36718
rect 24584 36654 24636 36660
rect 24952 36712 25004 36718
rect 24952 36654 25004 36660
rect 25228 36712 25280 36718
rect 25228 36654 25280 36660
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 23124 36242 23152 36518
rect 23112 36236 23164 36242
rect 23112 36178 23164 36184
rect 23112 36100 23164 36106
rect 23112 36042 23164 36048
rect 23124 35834 23152 36042
rect 23216 35834 23244 36654
rect 24596 36174 24624 36654
rect 24964 36242 24992 36654
rect 25240 36378 25268 36654
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25228 36372 25280 36378
rect 25228 36314 25280 36320
rect 25976 36242 26004 36518
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 25688 36236 25740 36242
rect 25688 36178 25740 36184
rect 25964 36236 26016 36242
rect 25964 36178 26016 36184
rect 24216 36168 24268 36174
rect 24216 36110 24268 36116
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24124 36100 24176 36106
rect 24124 36042 24176 36048
rect 23112 35828 23164 35834
rect 23112 35770 23164 35776
rect 23204 35828 23256 35834
rect 23204 35770 23256 35776
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 22466 35728 22522 35737
rect 23018 35728 23074 35737
rect 22466 35663 22468 35672
rect 22520 35663 22522 35672
rect 22560 35692 22612 35698
rect 22468 35634 22520 35640
rect 22560 35634 22612 35640
rect 22928 35692 22980 35698
rect 23018 35663 23020 35672
rect 22928 35634 22980 35640
rect 23072 35663 23074 35672
rect 23020 35634 23072 35640
rect 22480 34610 22508 35634
rect 22572 35290 22600 35634
rect 22940 35578 22968 35634
rect 23676 35578 23704 35770
rect 24136 35698 24164 36042
rect 24228 35834 24256 36110
rect 24676 36032 24728 36038
rect 24676 35974 24728 35980
rect 24860 36032 24912 36038
rect 24860 35974 24912 35980
rect 24216 35828 24268 35834
rect 24216 35770 24268 35776
rect 24688 35698 24716 35974
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 23940 35692 23992 35698
rect 24124 35692 24176 35698
rect 23940 35634 23992 35640
rect 24044 35652 24124 35680
rect 22652 35556 22704 35562
rect 22652 35498 22704 35504
rect 22940 35550 23704 35578
rect 22664 35290 22692 35498
rect 22560 35284 22612 35290
rect 22560 35226 22612 35232
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 22468 34604 22520 34610
rect 22468 34546 22520 34552
rect 22836 34604 22888 34610
rect 22836 34546 22888 34552
rect 22468 34060 22520 34066
rect 22468 34002 22520 34008
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 22282 32056 22338 32065
rect 22282 31991 22338 32000
rect 22388 31958 22416 33458
rect 22480 33114 22508 34002
rect 22560 33992 22612 33998
rect 22560 33934 22612 33940
rect 22468 33108 22520 33114
rect 22468 33050 22520 33056
rect 22572 32858 22600 33934
rect 22848 33522 22876 34546
rect 22652 33516 22704 33522
rect 22652 33458 22704 33464
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22480 32830 22600 32858
rect 22480 32065 22508 32830
rect 22560 32768 22612 32774
rect 22560 32710 22612 32716
rect 22466 32056 22522 32065
rect 22466 31991 22522 32000
rect 22192 31952 22244 31958
rect 22376 31952 22428 31958
rect 22244 31900 22324 31906
rect 22192 31894 22324 31900
rect 22376 31894 22428 31900
rect 22204 31878 22324 31894
rect 22190 31784 22246 31793
rect 22190 31719 22246 31728
rect 22100 31408 22152 31414
rect 22100 31350 22152 31356
rect 22204 30682 22232 31719
rect 22296 30938 22324 31878
rect 22468 31816 22520 31822
rect 22468 31758 22520 31764
rect 22480 31346 22508 31758
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 22572 31278 22600 32710
rect 22664 32570 22692 33458
rect 22744 33448 22796 33454
rect 22848 33425 22876 33458
rect 22744 33390 22796 33396
rect 22834 33416 22890 33425
rect 22756 33318 22784 33390
rect 22834 33351 22890 33360
rect 22744 33312 22796 33318
rect 22744 33254 22796 33260
rect 22744 32972 22796 32978
rect 22744 32914 22796 32920
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22756 32450 22784 32914
rect 22664 32422 22784 32450
rect 22664 32366 22692 32422
rect 22652 32360 22704 32366
rect 22652 32302 22704 32308
rect 22940 32314 22968 35550
rect 23112 35488 23164 35494
rect 23112 35430 23164 35436
rect 23124 35086 23152 35430
rect 23952 35290 23980 35634
rect 23940 35284 23992 35290
rect 23940 35226 23992 35232
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 23480 34604 23532 34610
rect 23480 34546 23532 34552
rect 23216 34202 23244 34546
rect 23204 34196 23256 34202
rect 23204 34138 23256 34144
rect 23020 34128 23072 34134
rect 23020 34070 23072 34076
rect 23032 33522 23060 34070
rect 23492 33658 23520 34546
rect 23664 34400 23716 34406
rect 23664 34342 23716 34348
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23480 33652 23532 33658
rect 23480 33594 23532 33600
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 23584 33368 23612 33798
rect 23676 33590 23704 34342
rect 23860 33862 23888 34886
rect 24044 33862 24072 35652
rect 24124 35634 24176 35640
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24136 35562 24164 35634
rect 24124 35556 24176 35562
rect 24124 35498 24176 35504
rect 24780 35086 24808 35770
rect 24872 35766 24900 35974
rect 24860 35760 24912 35766
rect 24860 35702 24912 35708
rect 24872 35086 24900 35702
rect 24768 35080 24820 35086
rect 24768 35022 24820 35028
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24964 34134 24992 36178
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 25320 36032 25372 36038
rect 25320 35974 25372 35980
rect 25044 35692 25096 35698
rect 25044 35634 25096 35640
rect 25332 35680 25360 35974
rect 25412 35692 25464 35698
rect 25332 35652 25412 35680
rect 25056 35290 25084 35634
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25044 35284 25096 35290
rect 25044 35226 25096 35232
rect 25148 34542 25176 35566
rect 25136 34536 25188 34542
rect 25136 34478 25188 34484
rect 24952 34128 25004 34134
rect 24952 34070 25004 34076
rect 24124 33924 24176 33930
rect 24124 33866 24176 33872
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 24032 33856 24084 33862
rect 24032 33798 24084 33804
rect 23664 33584 23716 33590
rect 23664 33526 23716 33532
rect 23492 33340 23612 33368
rect 23018 32464 23074 32473
rect 23074 32408 23152 32416
rect 23018 32399 23020 32408
rect 23072 32388 23152 32408
rect 23020 32370 23072 32376
rect 22664 32026 22692 32302
rect 22940 32286 23060 32314
rect 22926 32056 22982 32065
rect 22756 32026 22876 32042
rect 22652 32020 22704 32026
rect 22652 31962 22704 31968
rect 22756 32020 22888 32026
rect 22756 32014 22836 32020
rect 22756 31822 22784 32014
rect 22926 31991 22982 32000
rect 22836 31962 22888 31968
rect 22836 31884 22888 31890
rect 22836 31826 22888 31832
rect 22744 31816 22796 31822
rect 22744 31758 22796 31764
rect 22848 31346 22876 31826
rect 22940 31754 22968 31991
rect 22928 31748 22980 31754
rect 22928 31690 22980 31696
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22284 30932 22336 30938
rect 22284 30874 22336 30880
rect 22940 30802 22968 31690
rect 22928 30796 22980 30802
rect 22928 30738 22980 30744
rect 22204 30654 22508 30682
rect 21822 30016 21878 30025
rect 21822 29951 21878 29960
rect 21836 29782 21864 29951
rect 21824 29776 21876 29782
rect 21824 29718 21876 29724
rect 21916 29776 21968 29782
rect 21916 29718 21968 29724
rect 21824 29504 21876 29510
rect 21824 29446 21876 29452
rect 21836 29238 21864 29446
rect 21824 29232 21876 29238
rect 21824 29174 21876 29180
rect 21928 29073 21956 29718
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 22204 29702 22416 29730
rect 22480 29714 22508 30654
rect 22928 30660 22980 30666
rect 22928 30602 22980 30608
rect 22940 30258 22968 30602
rect 23032 30598 23060 32286
rect 23124 31822 23152 32388
rect 23204 32224 23256 32230
rect 23204 32166 23256 32172
rect 23216 31822 23244 32166
rect 23112 31816 23164 31822
rect 23112 31758 23164 31764
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 23124 30818 23152 31758
rect 23124 30790 23336 30818
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22560 29776 22612 29782
rect 22560 29718 22612 29724
rect 22112 29510 22140 29650
rect 22204 29646 22232 29702
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22204 29322 22232 29446
rect 22112 29306 22232 29322
rect 22100 29300 22232 29306
rect 22152 29294 22232 29300
rect 22100 29242 22152 29248
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 21914 29064 21970 29073
rect 21914 28999 21970 29008
rect 21732 28756 21784 28762
rect 21732 28698 21784 28704
rect 21730 28656 21786 28665
rect 21730 28591 21732 28600
rect 21784 28591 21786 28600
rect 21732 28562 21784 28568
rect 21732 27600 21784 27606
rect 21732 27542 21784 27548
rect 21744 27402 21772 27542
rect 21732 27396 21784 27402
rect 21784 27356 21864 27384
rect 21732 27338 21784 27344
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21744 26450 21772 26726
rect 21836 26450 21864 27356
rect 21928 26761 21956 28999
rect 22020 28626 22048 29106
rect 22192 29096 22244 29102
rect 22190 29064 22192 29073
rect 22244 29064 22246 29073
rect 22296 29034 22324 29582
rect 22190 28999 22246 29008
rect 22284 29028 22336 29034
rect 22284 28970 22336 28976
rect 22388 28966 22416 29702
rect 22468 29708 22520 29714
rect 22468 29650 22520 29656
rect 22468 29572 22520 29578
rect 22468 29514 22520 29520
rect 22376 28960 22428 28966
rect 22376 28902 22428 28908
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 22192 28552 22244 28558
rect 22388 28540 22416 28902
rect 22244 28512 22416 28540
rect 22192 28494 22244 28500
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 21914 26752 21970 26761
rect 21970 26710 22048 26738
rect 21914 26687 21970 26696
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 21732 26444 21784 26450
rect 21732 26386 21784 26392
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 21836 24886 21864 26386
rect 21732 24880 21784 24886
rect 21730 24848 21732 24857
rect 21824 24880 21876 24886
rect 21784 24848 21786 24857
rect 21824 24822 21876 24828
rect 21730 24783 21786 24792
rect 21732 24744 21784 24750
rect 21730 24712 21732 24721
rect 21784 24712 21786 24721
rect 21730 24647 21786 24656
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 21640 23724 21692 23730
rect 21640 23666 21692 23672
rect 21362 23624 21418 23633
rect 21362 23559 21418 23568
rect 21180 23248 21232 23254
rect 21180 23190 21232 23196
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 20916 22778 20944 23054
rect 20996 22976 21048 22982
rect 20996 22918 21048 22924
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 21008 22642 21036 22918
rect 21284 22710 21312 23054
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21272 22704 21324 22710
rect 21272 22646 21324 22652
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20812 21072 20864 21078
rect 20812 21014 20864 21020
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20640 20466 20668 20946
rect 20824 20602 20852 21014
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20916 20466 20944 20878
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20640 20369 20668 20402
rect 20626 20360 20682 20369
rect 20626 20295 20682 20304
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20548 19378 20576 19926
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20640 19310 20668 19926
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20456 18686 20576 18714
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 20074 17232 20130 17241
rect 20074 17167 20130 17176
rect 20088 17134 20116 17167
rect 20180 17134 20208 18294
rect 20456 18290 20484 18566
rect 20548 18465 20576 18686
rect 20534 18456 20590 18465
rect 20534 18391 20590 18400
rect 20640 18340 20668 18770
rect 20732 18698 20760 20266
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20824 19514 20852 19722
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20916 19446 20944 20402
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20824 18766 20852 18838
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20548 18312 20668 18340
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19708 15904 19760 15910
rect 19708 15846 19760 15852
rect 19720 15366 19748 15846
rect 19812 15638 19840 15914
rect 19800 15632 19852 15638
rect 19800 15574 19852 15580
rect 19996 15502 20024 16730
rect 20088 16590 20116 17070
rect 20272 16658 20300 17682
rect 20548 17610 20576 18312
rect 20732 17814 20760 18634
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20548 17377 20576 17546
rect 20534 17368 20590 17377
rect 20534 17303 20590 17312
rect 20640 17202 20668 17614
rect 20732 17542 20760 17750
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20732 17270 20760 17478
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20916 17202 20944 18566
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16726 20392 16934
rect 20352 16720 20404 16726
rect 20352 16662 20404 16668
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20076 16584 20128 16590
rect 20168 16584 20220 16590
rect 20076 16526 20128 16532
rect 20166 16552 20168 16561
rect 20220 16552 20222 16561
rect 20166 16487 20222 16496
rect 20076 16176 20128 16182
rect 20180 16153 20208 16487
rect 20076 16118 20128 16124
rect 20166 16144 20222 16153
rect 20088 16028 20116 16118
rect 20166 16079 20222 16088
rect 20168 16040 20220 16046
rect 20088 16000 20168 16028
rect 20168 15982 20220 15988
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19800 15496 19852 15502
rect 19798 15464 19800 15473
rect 19984 15496 20036 15502
rect 19852 15464 19854 15473
rect 19984 15438 20036 15444
rect 19798 15399 19854 15408
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 14346 19840 15302
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19904 14498 19932 14962
rect 19996 14822 20024 15438
rect 20088 14890 20116 15846
rect 20180 15026 20208 15982
rect 20272 15609 20300 16594
rect 20456 15722 20484 17002
rect 20640 16590 20668 17138
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20640 16454 20668 16526
rect 20536 16448 20588 16454
rect 20534 16416 20536 16425
rect 20628 16448 20680 16454
rect 20588 16416 20590 16425
rect 20628 16390 20680 16396
rect 20534 16351 20590 16360
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20548 15881 20576 16186
rect 20534 15872 20590 15881
rect 20534 15807 20590 15816
rect 20456 15694 20576 15722
rect 20258 15600 20314 15609
rect 20258 15535 20314 15544
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20272 15042 20300 15438
rect 20168 15020 20220 15026
rect 20272 15014 20392 15042
rect 20168 14962 20220 14968
rect 20260 14952 20312 14958
rect 20260 14894 20312 14900
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19982 14648 20038 14657
rect 19982 14583 19984 14592
rect 20036 14583 20038 14592
rect 19984 14554 20036 14560
rect 19904 14470 20024 14498
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19798 14240 19854 14249
rect 19798 14175 19854 14184
rect 19708 14000 19760 14006
rect 19708 13942 19760 13948
rect 19720 13870 19748 13942
rect 19812 13938 19840 14175
rect 19892 14000 19944 14006
rect 19996 13988 20024 14470
rect 20088 14249 20116 14826
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20074 14240 20130 14249
rect 20074 14175 20130 14184
rect 19944 13960 20024 13988
rect 19892 13942 19944 13948
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19883 13728 19935 13734
rect 19935 13696 19946 13705
rect 19883 13670 19890 13676
rect 19890 13631 19946 13640
rect 19996 13410 20024 13960
rect 19904 13382 20024 13410
rect 20180 13394 20208 14758
rect 20272 14521 20300 14894
rect 20258 14512 20314 14521
rect 20258 14447 20314 14456
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20272 14249 20300 14350
rect 20258 14240 20314 14249
rect 20258 14175 20314 14184
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20168 13388 20220 13394
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19720 12986 19748 13262
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19904 12850 19932 13382
rect 20168 13330 20220 13336
rect 20272 13326 20300 14010
rect 20364 13530 20392 15014
rect 20548 14482 20576 15694
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20456 14074 20484 14350
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20364 13326 20392 13466
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19706 12744 19762 12753
rect 19706 12679 19762 12688
rect 19720 12374 19748 12679
rect 19812 12374 19840 12786
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19800 12368 19852 12374
rect 19800 12310 19852 12316
rect 19798 12200 19854 12209
rect 19904 12170 19932 12786
rect 19798 12135 19800 12144
rect 19852 12135 19854 12144
rect 19892 12164 19944 12170
rect 19800 12106 19852 12112
rect 19892 12106 19944 12112
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19628 11082 19656 11630
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19522 9752 19578 9761
rect 19522 9687 19578 9696
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19156 8560 19208 8566
rect 19156 8502 19208 8508
rect 19168 8265 19196 8502
rect 19154 8256 19210 8265
rect 19154 8191 19210 8200
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 17314 7375 17316 7384
rect 17368 7375 17370 7384
rect 17776 7404 17828 7410
rect 17316 7346 17368 7352
rect 17776 7346 17828 7352
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 17052 6322 17080 6666
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 6118 17264 6258
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 16776 5642 16804 6054
rect 17328 5914 17356 7346
rect 19168 7206 19196 7754
rect 19260 7410 19288 9007
rect 19352 8537 19380 9114
rect 19444 8974 19472 9522
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19338 8528 19394 8537
rect 19338 8463 19340 8472
rect 19392 8463 19394 8472
rect 19340 8434 19392 8440
rect 19444 8090 19472 8570
rect 19536 8566 19564 9687
rect 19628 9586 19656 10134
rect 19720 10130 19748 11222
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19720 9926 19748 10066
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19812 9518 19840 12106
rect 19996 11354 20024 12922
rect 20088 12424 20116 13194
rect 20180 13161 20208 13194
rect 20260 13184 20312 13190
rect 20166 13152 20222 13161
rect 20260 13126 20312 13132
rect 20166 13087 20222 13096
rect 20168 12436 20220 12442
rect 20088 12396 20168 12424
rect 20168 12378 20220 12384
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19904 11257 19932 11290
rect 19890 11248 19946 11257
rect 19890 11183 19946 11192
rect 20088 11150 20116 12106
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19904 9994 19932 11086
rect 20180 10996 20208 11222
rect 20088 10968 20208 10996
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19996 10062 20024 10610
rect 20088 10305 20116 10968
rect 20272 10674 20300 13126
rect 20364 11830 20392 13262
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20350 11520 20406 11529
rect 20350 11455 20406 11464
rect 20364 11286 20392 11455
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 20350 11112 20406 11121
rect 20350 11047 20406 11056
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20074 10296 20130 10305
rect 20180 10266 20208 10610
rect 20258 10432 20314 10441
rect 20258 10367 20314 10376
rect 20074 10231 20130 10240
rect 20168 10260 20220 10266
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19522 8392 19578 8401
rect 19522 8327 19524 8336
rect 19576 8327 19578 8336
rect 19524 8298 19576 8304
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19338 7984 19394 7993
rect 19338 7919 19340 7928
rect 19392 7919 19394 7928
rect 19340 7890 19392 7896
rect 19536 7886 19564 8298
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19628 7886 19656 8230
rect 19904 7993 19932 9930
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19996 8106 20024 8910
rect 20088 8294 20116 10231
rect 20168 10202 20220 10208
rect 20272 10062 20300 10367
rect 20260 10056 20312 10062
rect 20166 10024 20222 10033
rect 20260 9998 20312 10004
rect 20166 9959 20168 9968
rect 20220 9959 20222 9968
rect 20168 9930 20220 9936
rect 20258 9072 20314 9081
rect 20258 9007 20314 9016
rect 20272 8974 20300 9007
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8809 20300 8910
rect 20258 8800 20314 8809
rect 20258 8735 20314 8744
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19996 8078 20208 8106
rect 19890 7984 19946 7993
rect 19890 7919 19946 7928
rect 19524 7880 19576 7886
rect 19430 7848 19486 7857
rect 19524 7822 19576 7828
rect 19616 7880 19668 7886
rect 19708 7880 19760 7886
rect 19616 7822 19668 7828
rect 19706 7848 19708 7857
rect 19984 7880 20036 7886
rect 19760 7848 19762 7857
rect 19430 7783 19486 7792
rect 19706 7783 19762 7792
rect 19812 7840 19984 7868
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7449 19380 7686
rect 19338 7440 19394 7449
rect 19248 7404 19300 7410
rect 19444 7410 19472 7783
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19524 7472 19576 7478
rect 19628 7449 19656 7686
rect 19524 7414 19576 7420
rect 19614 7440 19670 7449
rect 19338 7375 19340 7384
rect 19248 7346 19300 7352
rect 19392 7375 19394 7384
rect 19432 7404 19484 7410
rect 19340 7346 19392 7352
rect 19432 7346 19484 7352
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 17774 6896 17830 6905
rect 17774 6831 17830 6840
rect 17788 6798 17816 6831
rect 19536 6798 19564 7414
rect 19812 7410 19840 7840
rect 20180 7857 20208 8078
rect 19984 7822 20036 7828
rect 20166 7848 20222 7857
rect 20166 7783 20222 7792
rect 19614 7375 19670 7384
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19628 6798 19656 7210
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 6390 17632 6598
rect 17696 6458 17724 6734
rect 20088 6730 20116 7278
rect 20180 6934 20208 7278
rect 20364 7274 20392 11047
rect 20456 8945 20484 13330
rect 20548 12900 20576 13806
rect 20640 13326 20668 16390
rect 20916 15706 20944 17138
rect 21008 16776 21036 21490
rect 21192 20874 21220 22578
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21192 20584 21220 20810
rect 21100 20556 21220 20584
rect 21100 20330 21128 20556
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21088 20324 21140 20330
rect 21088 20266 21140 20272
rect 21192 19990 21220 20402
rect 21284 20330 21312 21558
rect 21272 20324 21324 20330
rect 21272 20266 21324 20272
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21180 19780 21232 19786
rect 21180 19722 21232 19728
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 19281 21128 19654
rect 21086 19272 21142 19281
rect 21086 19207 21142 19216
rect 21088 18760 21140 18766
rect 21086 18728 21088 18737
rect 21140 18728 21142 18737
rect 21086 18663 21142 18672
rect 21100 17882 21128 18663
rect 21192 18601 21220 19722
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 18766 21312 19654
rect 21376 19360 21404 22918
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21468 22545 21496 22578
rect 21454 22536 21510 22545
rect 21454 22471 21510 22480
rect 21454 20496 21510 20505
rect 21560 20466 21588 23666
rect 21652 23186 21680 23666
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21744 22642 21772 24647
rect 21836 24070 21864 24822
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21836 21690 21864 23598
rect 21928 23254 21956 26522
rect 22020 23798 22048 26710
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22112 26042 22140 26318
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22204 25430 22232 28358
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22296 27334 22324 27814
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 26994 22324 27270
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 22388 26364 22416 28512
rect 22480 28404 22508 29514
rect 22572 29306 22600 29718
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22652 29232 22704 29238
rect 22652 29174 22704 29180
rect 22664 29073 22692 29174
rect 22650 29064 22706 29073
rect 22560 29028 22612 29034
rect 22650 28999 22706 29008
rect 22560 28970 22612 28976
rect 22572 28558 22600 28970
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22560 28416 22612 28422
rect 22480 28376 22560 28404
rect 22560 28358 22612 28364
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22480 27130 22508 27338
rect 22468 27124 22520 27130
rect 22468 27066 22520 27072
rect 22572 27033 22600 28358
rect 22756 28082 22784 29650
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 27062 22784 27270
rect 22744 27056 22796 27062
rect 22558 27024 22614 27033
rect 22744 26998 22796 27004
rect 22558 26959 22614 26968
rect 22572 26926 22600 26959
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22468 26376 22520 26382
rect 22388 26336 22468 26364
rect 22468 26318 22520 26324
rect 22572 26228 22600 26862
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22296 26200 22600 26228
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 22296 24206 22324 26200
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22376 24676 22428 24682
rect 22376 24618 22428 24624
rect 22388 24410 22416 24618
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22284 24200 22336 24206
rect 22388 24177 22416 24346
rect 22284 24142 22336 24148
rect 22374 24168 22430 24177
rect 22374 24103 22430 24112
rect 22480 24070 22508 25230
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 22192 23656 22244 23662
rect 22006 23624 22062 23633
rect 22192 23598 22244 23604
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22006 23559 22062 23568
rect 22020 23526 22048 23559
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 22020 23100 22048 23190
rect 21928 23072 22048 23100
rect 22204 23100 22232 23598
rect 22296 23526 22324 23598
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 22388 23186 22416 23666
rect 22572 23633 22600 23666
rect 22558 23624 22614 23633
rect 22558 23559 22614 23568
rect 22468 23248 22520 23254
rect 22520 23208 22600 23236
rect 22468 23190 22520 23196
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22284 23112 22336 23118
rect 22204 23072 22284 23100
rect 21928 22642 21956 23072
rect 22204 23066 22232 23072
rect 22112 23038 22232 23066
rect 22284 23054 22336 23060
rect 22376 23044 22428 23050
rect 22006 22944 22062 22953
rect 22006 22879 22062 22888
rect 22020 22710 22048 22879
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21652 20806 21680 20946
rect 21928 20942 21956 22578
rect 22112 22506 22140 23038
rect 22376 22986 22428 22992
rect 22388 22506 22416 22986
rect 22466 22944 22522 22953
rect 22466 22879 22522 22888
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22376 22500 22428 22506
rect 22376 22442 22428 22448
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22020 21010 22048 21898
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21454 20431 21510 20440
rect 21548 20460 21600 20466
rect 21468 20330 21496 20431
rect 21548 20402 21600 20408
rect 21652 20398 21680 20742
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21652 19786 21680 20334
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 21456 19372 21508 19378
rect 21376 19332 21456 19360
rect 21376 18902 21404 19332
rect 21456 19314 21508 19320
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21468 18766 21496 19178
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21178 18592 21234 18601
rect 21178 18527 21234 18536
rect 21192 18306 21220 18527
rect 21468 18426 21496 18702
rect 21560 18698 21588 19450
rect 21732 19440 21784 19446
rect 21732 19382 21784 19388
rect 21744 18902 21772 19382
rect 21836 19378 21864 19654
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 21836 19009 21864 19314
rect 21822 19000 21878 19009
rect 21822 18935 21878 18944
rect 21732 18896 21784 18902
rect 21732 18838 21784 18844
rect 21744 18766 21772 18838
rect 21732 18760 21784 18766
rect 21652 18720 21732 18748
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21560 18601 21588 18634
rect 21546 18592 21602 18601
rect 21546 18527 21602 18536
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21192 18278 21312 18306
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21192 17610 21220 18158
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21192 17202 21220 17274
rect 21284 17202 21312 18278
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21456 18284 21508 18290
rect 21652 18272 21680 18720
rect 21732 18702 21784 18708
rect 21822 18456 21878 18465
rect 21732 18420 21784 18426
rect 21822 18391 21878 18400
rect 21732 18362 21784 18368
rect 21508 18244 21680 18272
rect 21456 18226 21508 18232
rect 21376 17678 21404 18226
rect 21468 17814 21496 18226
rect 21638 18184 21694 18193
rect 21638 18119 21694 18128
rect 21652 18086 21680 18119
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21376 17338 21404 17614
rect 21652 17610 21680 18022
rect 21744 17610 21772 18362
rect 21836 18154 21864 18391
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21640 17604 21692 17610
rect 21640 17546 21692 17552
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21454 17504 21510 17513
rect 21454 17439 21510 17448
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21100 17066 21128 17138
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21180 16788 21232 16794
rect 21008 16748 21180 16776
rect 21008 16114 21036 16748
rect 21180 16730 21232 16736
rect 21284 16674 21312 17138
rect 21192 16646 21312 16674
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20732 13870 20760 15030
rect 20824 13977 20852 15438
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20916 15065 20944 15098
rect 20902 15056 20958 15065
rect 20902 14991 20958 15000
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20810 13968 20866 13977
rect 20810 13903 20866 13912
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20628 12912 20680 12918
rect 20548 12872 20628 12900
rect 20628 12854 20680 12860
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 11558 20576 12582
rect 20640 12170 20668 12854
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11937 20760 12038
rect 20718 11928 20774 11937
rect 20718 11863 20774 11872
rect 20824 11880 20852 12378
rect 20916 12050 20944 14350
rect 21008 12918 21036 14962
rect 21192 14822 21220 16646
rect 21468 16454 21496 17439
rect 21546 17368 21602 17377
rect 21546 17303 21602 17312
rect 21560 17202 21588 17303
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21652 16572 21680 17546
rect 21744 17134 21772 17546
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21732 16720 21784 16726
rect 21732 16662 21784 16668
rect 21560 16544 21680 16572
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 14074 21220 14214
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21284 13546 21312 16390
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21376 14618 21404 15438
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21468 15026 21496 15098
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14618 21496 14758
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21376 14278 21404 14418
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21192 13518 21312 13546
rect 21100 13433 21128 13466
rect 21086 13424 21142 13433
rect 21086 13359 21142 13368
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 21100 12374 21128 13194
rect 21192 12986 21220 13518
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21284 12832 21312 13262
rect 21376 13025 21404 14214
rect 21454 13968 21510 13977
rect 21454 13903 21510 13912
rect 21362 13016 21418 13025
rect 21362 12951 21418 12960
rect 21192 12804 21312 12832
rect 21364 12844 21416 12850
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21192 12322 21220 12804
rect 21364 12786 21416 12792
rect 21376 12442 21404 12786
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21100 12170 21128 12310
rect 21192 12294 21312 12322
rect 21284 12238 21312 12294
rect 21468 12288 21496 13903
rect 21560 13462 21588 16544
rect 21744 16454 21772 16662
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21824 16040 21876 16046
rect 21730 16008 21786 16017
rect 21824 15982 21876 15988
rect 21730 15943 21786 15952
rect 21638 15736 21694 15745
rect 21638 15671 21694 15680
rect 21652 14958 21680 15671
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21652 13326 21680 13670
rect 21640 13320 21692 13326
rect 21560 13280 21640 13308
rect 21560 12345 21588 13280
rect 21640 13262 21692 13268
rect 21744 13002 21772 15943
rect 21836 15502 21864 15982
rect 21928 15706 21956 20878
rect 22204 20602 22232 21558
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22020 19417 22048 20402
rect 22006 19408 22062 19417
rect 22006 19343 22062 19352
rect 22020 18426 22048 19343
rect 22098 19272 22154 19281
rect 22098 19207 22154 19216
rect 22112 19174 22140 19207
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22112 18850 22140 19110
rect 22192 18964 22244 18970
rect 22296 18952 22324 21626
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22244 18924 22324 18952
rect 22192 18906 22244 18912
rect 22112 18834 22232 18850
rect 22112 18828 22244 18834
rect 22112 18822 22192 18828
rect 22192 18770 22244 18776
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22112 18601 22140 18702
rect 22098 18592 22154 18601
rect 22098 18527 22154 18536
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22112 18306 22140 18527
rect 22020 18278 22140 18306
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21914 15192 21970 15201
rect 21914 15127 21970 15136
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14618 21864 14758
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21928 13410 21956 15127
rect 22020 14890 22048 18278
rect 22204 17066 22232 18770
rect 22282 18456 22338 18465
rect 22282 18391 22338 18400
rect 22296 18290 22324 18391
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22388 17882 22416 20878
rect 22480 19334 22508 22879
rect 22572 21672 22600 23208
rect 22664 22778 22692 26726
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22756 24750 22784 25366
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22756 23066 22784 24142
rect 22848 23322 22876 29582
rect 22940 27713 22968 30194
rect 23124 30122 23152 30670
rect 23216 30258 23244 30670
rect 23308 30394 23336 30790
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23112 30116 23164 30122
rect 23112 30058 23164 30064
rect 23018 29472 23074 29481
rect 23018 29407 23074 29416
rect 23032 29034 23060 29407
rect 23124 29306 23152 30058
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23112 29096 23164 29102
rect 23110 29064 23112 29073
rect 23164 29064 23166 29073
rect 23020 29028 23072 29034
rect 23110 28999 23166 29008
rect 23020 28970 23072 28976
rect 23124 28529 23152 28999
rect 23110 28520 23166 28529
rect 23110 28455 23166 28464
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 22926 27704 22982 27713
rect 22926 27639 22982 27648
rect 22940 26382 22968 27639
rect 23124 27606 23152 28358
rect 23112 27600 23164 27606
rect 23112 27542 23164 27548
rect 23020 27464 23072 27470
rect 23018 27432 23020 27441
rect 23216 27452 23244 30194
rect 23492 30190 23520 33340
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23584 31822 23612 32846
rect 23860 32026 23888 32846
rect 24044 32366 24072 33798
rect 24032 32360 24084 32366
rect 24032 32302 24084 32308
rect 24136 32298 24164 33866
rect 24676 33584 24728 33590
rect 24676 33526 24728 33532
rect 24400 33448 24452 33454
rect 24400 33390 24452 33396
rect 24216 32836 24268 32842
rect 24216 32778 24268 32784
rect 24308 32836 24360 32842
rect 24308 32778 24360 32784
rect 24228 32434 24256 32778
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24124 32292 24176 32298
rect 24124 32234 24176 32240
rect 23848 32020 23900 32026
rect 23848 31962 23900 31968
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23572 31816 23624 31822
rect 23572 31758 23624 31764
rect 23860 31414 23888 31962
rect 23952 31890 23980 31962
rect 23940 31884 23992 31890
rect 23940 31826 23992 31832
rect 24136 31414 24164 32234
rect 24228 31793 24256 32370
rect 24320 32314 24348 32778
rect 24412 32434 24440 33390
rect 24688 32978 24716 33526
rect 24676 32972 24728 32978
rect 24676 32914 24728 32920
rect 24400 32428 24452 32434
rect 24400 32370 24452 32376
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24320 32298 24440 32314
rect 24320 32292 24452 32298
rect 24320 32286 24400 32292
rect 24320 31822 24348 32286
rect 24400 32234 24452 32240
rect 24308 31816 24360 31822
rect 24214 31784 24270 31793
rect 24308 31758 24360 31764
rect 24214 31719 24270 31728
rect 24228 31482 24256 31719
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 23848 31408 23900 31414
rect 23848 31350 23900 31356
rect 24124 31408 24176 31414
rect 24124 31350 24176 31356
rect 24412 31346 24440 31622
rect 24596 31414 24624 32370
rect 24688 31498 24716 32914
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24872 32366 24900 32710
rect 24964 32570 24992 34070
rect 25148 33590 25176 34478
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 25056 33318 25084 33458
rect 25044 33312 25096 33318
rect 25044 33254 25096 33260
rect 24952 32564 25004 32570
rect 24952 32506 25004 32512
rect 25056 32434 25084 33254
rect 25148 32978 25176 33526
rect 25136 32972 25188 32978
rect 25136 32914 25188 32920
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 24860 32360 24912 32366
rect 24860 32302 24912 32308
rect 24768 32020 24820 32026
rect 24768 31962 24820 31968
rect 24780 31686 24808 31962
rect 24860 31816 24912 31822
rect 24860 31758 24912 31764
rect 24872 31686 24900 31758
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24860 31680 24912 31686
rect 24860 31622 24912 31628
rect 24688 31482 24808 31498
rect 24688 31476 24820 31482
rect 24688 31470 24768 31476
rect 24768 31418 24820 31424
rect 24584 31408 24636 31414
rect 24584 31350 24636 31356
rect 24872 31346 24900 31622
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 24228 31249 24256 31282
rect 24214 31240 24270 31249
rect 24214 31175 24270 31184
rect 23572 30864 23624 30870
rect 23572 30806 23624 30812
rect 23480 30184 23532 30190
rect 23480 30126 23532 30132
rect 23584 30054 23612 30806
rect 23756 30660 23808 30666
rect 23756 30602 23808 30608
rect 23664 30592 23716 30598
rect 23664 30534 23716 30540
rect 23676 30394 23704 30534
rect 23664 30388 23716 30394
rect 23664 30330 23716 30336
rect 23676 30258 23704 30330
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 23572 30048 23624 30054
rect 23572 29990 23624 29996
rect 23296 29164 23348 29170
rect 23348 29124 23520 29152
rect 23296 29106 23348 29112
rect 23492 28966 23520 29124
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23388 28552 23440 28558
rect 23072 27432 23074 27441
rect 23018 27367 23074 27376
rect 23124 27424 23244 27452
rect 23308 28512 23388 28540
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 23032 25514 23060 27367
rect 22940 25486 23060 25514
rect 22940 25226 22968 25486
rect 23020 25356 23072 25362
rect 23020 25298 23072 25304
rect 22928 25220 22980 25226
rect 22928 25162 22980 25168
rect 22940 25129 22968 25162
rect 22926 25120 22982 25129
rect 22926 25055 22982 25064
rect 23032 24750 23060 25298
rect 23020 24744 23072 24750
rect 23020 24686 23072 24692
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 22940 24138 22968 24346
rect 23032 24206 23060 24686
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22928 24132 22980 24138
rect 22928 24074 22980 24080
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 22756 23050 22876 23066
rect 22756 23044 22888 23050
rect 22756 23038 22836 23044
rect 22836 22986 22888 22992
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22650 22672 22706 22681
rect 22650 22607 22652 22616
rect 22704 22607 22706 22616
rect 22652 22578 22704 22584
rect 22756 22574 22784 22918
rect 22744 22568 22796 22574
rect 22742 22536 22744 22545
rect 22796 22536 22798 22545
rect 22742 22471 22798 22480
rect 22940 22094 22968 24074
rect 22848 22066 22968 22094
rect 22744 21684 22796 21690
rect 22572 21644 22744 21672
rect 22744 21626 22796 21632
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22572 20942 22600 21490
rect 22848 21146 22876 22066
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22652 21140 22704 21146
rect 22836 21140 22888 21146
rect 22704 21100 22784 21128
rect 22652 21082 22704 21088
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22480 19306 22600 19334
rect 22468 18692 22520 18698
rect 22468 18634 22520 18640
rect 22480 18358 22508 18634
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22480 17882 22508 18294
rect 22572 18290 22600 19306
rect 22664 18698 22692 20402
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22284 17808 22336 17814
rect 22572 17762 22600 18226
rect 22664 18086 22692 18634
rect 22756 18358 22784 21100
rect 22836 21082 22888 21088
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22848 19446 22876 20470
rect 22836 19440 22888 19446
rect 22836 19382 22888 19388
rect 22940 18816 22968 21966
rect 23124 21418 23152 27424
rect 23308 26042 23336 28512
rect 23388 28494 23440 28500
rect 23388 28416 23440 28422
rect 23386 28384 23388 28393
rect 23440 28384 23442 28393
rect 23386 28319 23442 28328
rect 23388 28008 23440 28014
rect 23388 27950 23440 27956
rect 23400 27470 23428 27950
rect 23492 27538 23520 28902
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23296 26036 23348 26042
rect 23296 25978 23348 25984
rect 23204 25934 23256 25940
rect 23400 25922 23428 27270
rect 23492 27130 23520 27270
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23584 26042 23612 29990
rect 23664 29572 23716 29578
rect 23664 29514 23716 29520
rect 23676 27946 23704 29514
rect 23768 29209 23796 30602
rect 24216 30048 24268 30054
rect 24214 30016 24216 30025
rect 24268 30016 24270 30025
rect 24214 29951 24270 29960
rect 24228 29714 24256 29951
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 24308 29640 24360 29646
rect 24308 29582 24360 29588
rect 23940 29504 23992 29510
rect 23940 29446 23992 29452
rect 23754 29200 23810 29209
rect 23952 29170 23980 29446
rect 24320 29306 24348 29582
rect 24308 29300 24360 29306
rect 24308 29242 24360 29248
rect 24124 29232 24176 29238
rect 24124 29174 24176 29180
rect 23754 29135 23810 29144
rect 23940 29164 23992 29170
rect 23664 27940 23716 27946
rect 23664 27882 23716 27888
rect 23768 27520 23796 29135
rect 23940 29106 23992 29112
rect 23952 28994 23980 29106
rect 24136 29050 24164 29174
rect 24044 29034 24164 29050
rect 23860 28966 23980 28994
rect 24032 29028 24164 29034
rect 24084 29022 24164 29028
rect 24032 28970 24084 28976
rect 23860 28422 23888 28966
rect 23848 28416 23900 28422
rect 23848 28358 23900 28364
rect 23676 27492 23796 27520
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23676 25945 23704 27492
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23204 25876 23256 25882
rect 23308 25894 23428 25922
rect 23662 25936 23718 25945
rect 23216 25158 23244 25876
rect 23308 25702 23336 25894
rect 23662 25871 23718 25880
rect 23768 25770 23796 27338
rect 23860 26858 23888 28358
rect 24306 28112 24362 28121
rect 23940 28076 23992 28082
rect 24306 28047 24308 28056
rect 23940 28018 23992 28024
rect 24360 28047 24362 28056
rect 24308 28018 24360 28024
rect 23848 26852 23900 26858
rect 23848 26794 23900 26800
rect 23846 26752 23902 26761
rect 23846 26687 23902 26696
rect 23860 26042 23888 26687
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23848 25900 23900 25906
rect 23848 25842 23900 25848
rect 23756 25764 23808 25770
rect 23756 25706 23808 25712
rect 23296 25696 23348 25702
rect 23296 25638 23348 25644
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23664 25696 23716 25702
rect 23664 25638 23716 25644
rect 23400 25158 23428 25638
rect 23676 25362 23704 25638
rect 23860 25498 23888 25842
rect 23848 25492 23900 25498
rect 23848 25434 23900 25440
rect 23664 25356 23716 25362
rect 23664 25298 23716 25304
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23388 25152 23440 25158
rect 23388 25094 23440 25100
rect 23216 23361 23244 25094
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23308 24274 23336 24754
rect 23400 24410 23428 24754
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23308 23798 23336 24210
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 23202 23352 23258 23361
rect 23202 23287 23258 23296
rect 23216 22760 23244 23287
rect 23308 22964 23336 23734
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23400 23322 23428 23666
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23492 23254 23520 25230
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23584 23050 23612 24754
rect 23756 24132 23808 24138
rect 23756 24074 23808 24080
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23388 22976 23440 22982
rect 23308 22936 23388 22964
rect 23388 22918 23440 22924
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23400 22778 23428 22918
rect 23388 22772 23440 22778
rect 23216 22732 23336 22760
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23216 22137 23244 22578
rect 23202 22128 23258 22137
rect 23202 22063 23258 22072
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23032 20398 23060 20742
rect 23124 20602 23152 20742
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23020 20392 23072 20398
rect 23020 20334 23072 20340
rect 22848 18788 22968 18816
rect 22848 18426 22876 18788
rect 22928 18692 22980 18698
rect 22928 18634 22980 18640
rect 22940 18426 22968 18634
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 22744 18352 22796 18358
rect 22744 18294 22796 18300
rect 22756 18222 22784 18294
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22284 17750 22336 17756
rect 22296 17542 22324 17750
rect 22480 17734 22600 17762
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 17202 22324 17478
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22282 16144 22338 16153
rect 22282 16079 22284 16088
rect 22336 16079 22338 16088
rect 22284 16050 22336 16056
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22296 15638 22324 15914
rect 22376 15700 22428 15706
rect 22376 15642 22428 15648
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22112 15026 22140 15438
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22204 14618 22232 15438
rect 22296 15026 22324 15574
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22388 14906 22416 15642
rect 22296 14878 22416 14906
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22190 14512 22246 14521
rect 22190 14447 22246 14456
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21652 12974 21772 13002
rect 21836 13382 21956 13410
rect 21376 12260 21496 12288
rect 21546 12336 21602 12345
rect 21546 12271 21548 12280
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21088 12164 21140 12170
rect 21088 12106 21140 12112
rect 21180 12096 21232 12102
rect 20916 12022 21036 12050
rect 21180 12038 21232 12044
rect 20732 11830 20760 11863
rect 20824 11852 20944 11880
rect 20628 11824 20680 11830
rect 20626 11792 20628 11801
rect 20720 11824 20772 11830
rect 20680 11792 20682 11801
rect 20772 11784 20852 11812
rect 20720 11766 20772 11772
rect 20626 11727 20682 11736
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 11354 20760 11494
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20824 11286 20852 11784
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20916 11218 20944 11852
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20548 9110 20576 11154
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20720 11144 20772 11150
rect 20772 11104 20852 11132
rect 20720 11086 20772 11092
rect 20640 10248 20668 11086
rect 20720 10260 20772 10266
rect 20640 10220 20720 10248
rect 20720 10202 20772 10208
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20640 9586 20668 9998
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20442 8936 20498 8945
rect 20442 8871 20498 8880
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20352 7268 20404 7274
rect 20352 7210 20404 7216
rect 20456 7206 20484 8434
rect 20548 8362 20576 9046
rect 20640 9042 20668 9522
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20640 8498 20668 8978
rect 20732 8566 20760 10202
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 20626 8256 20682 8265
rect 20626 8191 20682 8200
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20168 6928 20220 6934
rect 20168 6870 20220 6876
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17328 5642 17356 5850
rect 16764 5636 16816 5642
rect 16764 5578 16816 5584
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 16868 5166 16896 5510
rect 17512 5234 17540 5510
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4690 16528 4966
rect 16868 4690 16896 5102
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15396 3466 15424 4014
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 2514 15240 2790
rect 15488 2514 15516 3538
rect 15580 3466 15608 3878
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16132 3058 16160 3402
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 16224 2446 16252 4422
rect 17604 4214 17632 5306
rect 17696 5234 17724 6394
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17696 4282 17724 5170
rect 17788 5166 17816 6054
rect 18892 5914 18920 6326
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18984 5710 19012 6258
rect 19352 6254 19380 6666
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17866 5400 17922 5409
rect 17866 5335 17868 5344
rect 17920 5335 17922 5344
rect 17868 5306 17920 5312
rect 17972 5302 18000 5510
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17604 4049 17632 4150
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17590 4040 17646 4049
rect 16948 4004 17000 4010
rect 17590 3975 17646 3984
rect 16948 3946 17000 3952
rect 16960 3738 16988 3946
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17604 3670 17632 3975
rect 17696 3738 17724 4082
rect 17788 4078 17816 5102
rect 18432 4758 18460 5646
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18156 4214 18184 4422
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 2990 16804 3470
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 17052 2514 17080 3334
rect 17144 3126 17172 3334
rect 17788 3194 17816 4014
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 18156 2854 18184 3334
rect 18248 3058 18276 4490
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 15488 800 15516 2246
rect 16132 800 16160 2246
rect 16762 1864 16818 1873
rect 16762 1799 16818 1808
rect 16776 800 16804 1799
rect 17512 1170 17540 2586
rect 18248 2378 18276 2994
rect 18432 2582 18460 3470
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 18524 2446 18552 4014
rect 18708 3942 18736 4558
rect 19076 4554 19104 5850
rect 19168 5710 19196 6190
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 19076 4214 19104 4490
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 18616 1873 18644 3538
rect 19168 3534 19196 5646
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19248 5160 19300 5166
rect 19248 5102 19300 5108
rect 19260 4622 19288 5102
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18602 1864 18658 1873
rect 18800 1850 18828 3470
rect 19352 3108 19380 5238
rect 19444 4146 19472 6054
rect 19536 5710 19564 6190
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5846 19656 6054
rect 19616 5840 19668 5846
rect 19616 5782 19668 5788
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 5370 19564 5646
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19628 5234 19656 5306
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19524 4072 19576 4078
rect 19522 4040 19524 4049
rect 19576 4040 19578 4049
rect 19522 3975 19578 3984
rect 19628 3618 19656 4762
rect 19720 4010 19748 6598
rect 20534 6488 20590 6497
rect 20534 6423 20590 6432
rect 20548 6390 20576 6423
rect 20444 6384 20496 6390
rect 20444 6326 20496 6332
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 19800 6180 19852 6186
rect 19800 6122 19852 6128
rect 19812 4078 19840 6122
rect 20352 5296 20404 5302
rect 20350 5264 20352 5273
rect 20404 5264 20406 5273
rect 20350 5199 20406 5208
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20364 4826 20392 5102
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 19892 4616 19944 4622
rect 19892 4558 19944 4564
rect 19904 4282 19932 4558
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 20272 4146 20300 4694
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20364 3670 20392 3878
rect 19536 3590 19656 3618
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 19536 3534 19564 3590
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19432 3120 19484 3126
rect 19352 3080 19432 3108
rect 19432 3062 19484 3068
rect 20456 2990 20484 6326
rect 20640 5846 20668 8191
rect 20732 6730 20760 8366
rect 20824 7206 20852 11104
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20916 10985 20944 11018
rect 20902 10976 20958 10985
rect 20902 10911 20958 10920
rect 21008 10033 21036 12022
rect 21192 11762 21220 12038
rect 21376 11762 21404 12260
rect 21600 12271 21602 12280
rect 21548 12242 21600 12248
rect 21456 12164 21508 12170
rect 21456 12106 21508 12112
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21272 11552 21324 11558
rect 21270 11520 21272 11529
rect 21324 11520 21326 11529
rect 21270 11455 21326 11464
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21180 11280 21232 11286
rect 21178 11248 21180 11257
rect 21232 11248 21234 11257
rect 21178 11183 21234 11192
rect 21178 10976 21234 10985
rect 21178 10911 21234 10920
rect 20994 10024 21050 10033
rect 20916 9982 20994 10010
rect 20916 8362 20944 9982
rect 20994 9959 21050 9968
rect 20994 9344 21050 9353
rect 20994 9279 21050 9288
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 21008 8090 21036 9279
rect 21086 9208 21142 9217
rect 21086 9143 21142 9152
rect 21100 8498 21128 9143
rect 21192 8634 21220 10911
rect 21284 10470 21312 11290
rect 21376 11257 21404 11698
rect 21468 11354 21496 12106
rect 21546 11792 21602 11801
rect 21546 11727 21602 11736
rect 21560 11354 21588 11727
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21362 11248 21418 11257
rect 21362 11183 21418 11192
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21376 10742 21404 11086
rect 21560 11014 21588 11086
rect 21652 11014 21680 12974
rect 21732 12912 21784 12918
rect 21732 12854 21784 12860
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21560 10742 21588 10950
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 21548 10736 21600 10742
rect 21548 10678 21600 10684
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21468 10062 21496 10474
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21284 9654 21312 9930
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21376 9178 21404 9862
rect 21454 9208 21510 9217
rect 21364 9172 21416 9178
rect 21454 9143 21456 9152
rect 21364 9114 21416 9120
rect 21508 9143 21510 9152
rect 21456 9114 21508 9120
rect 21560 9058 21588 10678
rect 21652 10169 21680 10950
rect 21638 10160 21694 10169
rect 21638 10095 21694 10104
rect 21560 9030 21680 9058
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21086 8392 21142 8401
rect 21086 8327 21142 8336
rect 21192 8344 21220 8570
rect 21284 8537 21312 8774
rect 21468 8566 21496 8910
rect 21456 8560 21508 8566
rect 21270 8528 21326 8537
rect 21456 8502 21508 8508
rect 21270 8463 21326 8472
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21100 7886 21128 8327
rect 21192 8316 21312 8344
rect 21178 8256 21234 8265
rect 21178 8191 21234 8200
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 20916 7274 20944 7414
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20916 5692 20944 7210
rect 21192 7002 21220 8191
rect 21284 7410 21312 8316
rect 21468 7886 21496 8502
rect 21560 8430 21588 8910
rect 21652 8634 21680 9030
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21560 8090 21588 8366
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21652 7478 21680 8570
rect 21744 8106 21772 12854
rect 21836 9926 21864 13382
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21928 12458 21956 13262
rect 22020 12628 22048 14350
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22112 12850 22140 13466
rect 22204 13172 22232 14447
rect 22296 14414 22324 14878
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22284 13184 22336 13190
rect 22204 13144 22284 13172
rect 22284 13126 22336 13132
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22020 12600 22232 12628
rect 21928 12430 22140 12458
rect 21914 12200 21970 12209
rect 21914 12135 21916 12144
rect 21968 12135 21970 12144
rect 21916 12106 21968 12112
rect 21928 10266 21956 12106
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11286 22048 11698
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 22020 10146 22048 10610
rect 21928 10118 22048 10146
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 21836 8242 21864 9862
rect 21928 8838 21956 10118
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 22020 9178 22048 9998
rect 22112 9674 22140 12430
rect 22204 11150 22232 12600
rect 22296 12481 22324 13126
rect 22282 12472 22338 12481
rect 22282 12407 22338 12416
rect 22388 12356 22416 14758
rect 22480 14521 22508 17734
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 17338 22600 17478
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22560 17128 22612 17134
rect 22558 17096 22560 17105
rect 22612 17096 22614 17105
rect 22558 17031 22614 17040
rect 22572 15745 22600 17031
rect 22664 16998 22692 17614
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22756 17338 22784 17546
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22558 15736 22614 15745
rect 22558 15671 22614 15680
rect 22664 15620 22692 16934
rect 22756 16522 22784 17138
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22848 16182 22876 18362
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22572 15592 22692 15620
rect 22572 15162 22600 15592
rect 22848 15502 22876 16118
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22466 14512 22522 14521
rect 22466 14447 22522 14456
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22480 12442 22508 14350
rect 22572 14278 22600 14962
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22558 12880 22614 12889
rect 22558 12815 22560 12824
rect 22612 12815 22614 12824
rect 22560 12786 22612 12792
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22296 12328 22416 12356
rect 22296 11694 22324 12328
rect 22572 12322 22600 12786
rect 22480 12306 22600 12322
rect 22480 12300 22612 12306
rect 22480 12294 22560 12300
rect 22480 12220 22508 12294
rect 22560 12242 22612 12248
rect 22388 12192 22508 12220
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22192 11144 22244 11150
rect 22296 11121 22324 11290
rect 22192 11086 22244 11092
rect 22282 11112 22338 11121
rect 22282 11047 22284 11056
rect 22336 11047 22338 11056
rect 22284 11018 22336 11024
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22204 10266 22232 10406
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22112 9646 22232 9674
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 22008 8424 22060 8430
rect 22060 8384 22140 8412
rect 22008 8366 22060 8372
rect 22008 8288 22060 8294
rect 22006 8256 22008 8265
rect 22060 8256 22062 8265
rect 21836 8214 21956 8242
rect 21744 8078 21864 8106
rect 21732 8016 21784 8022
rect 21730 7984 21732 7993
rect 21784 7984 21786 7993
rect 21730 7919 21786 7928
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21560 6730 21588 7346
rect 21836 7274 21864 8078
rect 21928 7750 21956 8214
rect 22006 8191 22062 8200
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21916 7540 21968 7546
rect 21916 7482 21968 7488
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21638 7032 21694 7041
rect 21638 6967 21694 6976
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21652 6322 21680 6967
rect 21928 6633 21956 7482
rect 22020 7478 22048 8191
rect 22112 8022 22140 8384
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22112 7857 22140 7958
rect 22098 7848 22154 7857
rect 22098 7783 22154 7792
rect 22204 7546 22232 9646
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22008 7472 22060 7478
rect 22008 7414 22060 7420
rect 22100 7472 22152 7478
rect 22100 7414 22152 7420
rect 22020 7002 22048 7414
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 21914 6624 21970 6633
rect 21914 6559 21970 6568
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21824 5840 21876 5846
rect 21824 5782 21876 5788
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20996 5704 21048 5710
rect 20916 5664 20996 5692
rect 20996 5646 21048 5652
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 4078 20760 5510
rect 20824 4622 20852 5578
rect 21008 5030 21036 5646
rect 21100 5098 21128 5714
rect 21744 5710 21772 5782
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 21100 4554 21128 5034
rect 21284 4690 21312 5646
rect 21836 5642 21864 5782
rect 21928 5692 21956 6258
rect 22020 6118 22048 6938
rect 22112 6798 22140 7414
rect 22296 7002 22324 8434
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 22008 6112 22060 6118
rect 22008 6054 22060 6060
rect 22098 5808 22154 5817
rect 22098 5743 22154 5752
rect 22112 5710 22140 5743
rect 22008 5704 22060 5710
rect 21928 5664 22008 5692
rect 21824 5636 21876 5642
rect 21824 5578 21876 5584
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21928 4622 21956 5664
rect 22008 5646 22060 5652
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22112 5166 22140 5510
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 22112 3194 22140 4626
rect 22296 4554 22324 5510
rect 22388 5302 22416 12192
rect 22560 12164 22612 12170
rect 22560 12106 22612 12112
rect 22572 12073 22600 12106
rect 22558 12064 22614 12073
rect 22558 11999 22614 12008
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22480 11150 22508 11494
rect 22664 11336 22692 15438
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22756 12646 22784 15370
rect 22940 15366 22968 18158
rect 23032 16561 23060 20334
rect 23110 18728 23166 18737
rect 23110 18663 23166 18672
rect 23018 16552 23074 16561
rect 23018 16487 23074 16496
rect 23124 15706 23152 18663
rect 23216 18086 23244 22063
rect 23308 21185 23336 22732
rect 23388 22714 23440 22720
rect 23294 21176 23350 21185
rect 23492 21146 23520 22918
rect 23570 21992 23626 22001
rect 23570 21927 23626 21936
rect 23584 21894 23612 21927
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23294 21111 23350 21120
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23386 20768 23442 20777
rect 23386 20703 23442 20712
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 23308 20398 23336 20470
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23308 18222 23336 20198
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 23018 15192 23074 15201
rect 23018 15127 23020 15136
rect 23072 15127 23074 15136
rect 23020 15098 23072 15104
rect 23216 15094 23244 18022
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23308 17377 23336 17546
rect 23294 17368 23350 17377
rect 23294 17303 23296 17312
rect 23348 17303 23350 17312
rect 23296 17274 23348 17280
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23308 16590 23336 17002
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23400 16250 23428 20703
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23492 20262 23520 20402
rect 23480 20256 23532 20262
rect 23480 20198 23532 20204
rect 23480 19236 23532 19242
rect 23480 19178 23532 19184
rect 23492 17082 23520 19178
rect 23584 17678 23612 21558
rect 23676 20262 23704 24006
rect 23768 23798 23796 24074
rect 23756 23792 23808 23798
rect 23756 23734 23808 23740
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23664 19984 23716 19990
rect 23664 19926 23716 19932
rect 23676 19854 23704 19926
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23676 17814 23704 19790
rect 23768 19514 23796 23054
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23860 21622 23888 21898
rect 23848 21616 23900 21622
rect 23848 21558 23900 21564
rect 23848 21480 23900 21486
rect 23846 21448 23848 21457
rect 23900 21448 23902 21457
rect 23846 21383 23902 21392
rect 23952 21332 23980 28018
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24214 27704 24270 27713
rect 24214 27639 24270 27648
rect 24228 27538 24256 27639
rect 24320 27606 24348 27814
rect 24308 27600 24360 27606
rect 24308 27542 24360 27548
rect 24216 27532 24268 27538
rect 24216 27474 24268 27480
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24044 27130 24072 27406
rect 24124 27396 24176 27402
rect 24124 27338 24176 27344
rect 24032 27124 24084 27130
rect 24032 27066 24084 27072
rect 24032 26920 24084 26926
rect 24032 26862 24084 26868
rect 24044 22030 24072 26862
rect 24136 24750 24164 27338
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24228 26994 24256 27066
rect 24306 27024 24362 27033
rect 24216 26988 24268 26994
rect 24306 26959 24308 26968
rect 24216 26930 24268 26936
rect 24360 26959 24362 26968
rect 24308 26930 24360 26936
rect 24216 26852 24268 26858
rect 24216 26794 24268 26800
rect 24228 25888 24256 26794
rect 24308 26512 24360 26518
rect 24308 26454 24360 26460
rect 24320 26353 24348 26454
rect 24306 26344 24362 26353
rect 24306 26279 24362 26288
rect 24308 25900 24360 25906
rect 24228 25860 24308 25888
rect 24308 25842 24360 25848
rect 24412 25498 24440 31282
rect 24872 30938 24900 31282
rect 25332 30977 25360 35652
rect 25412 35634 25464 35640
rect 25516 35290 25544 36110
rect 25596 35488 25648 35494
rect 25596 35430 25648 35436
rect 25504 35284 25556 35290
rect 25504 35226 25556 35232
rect 25608 35154 25636 35430
rect 25596 35148 25648 35154
rect 25596 35090 25648 35096
rect 25700 34474 25728 36178
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26148 36032 26200 36038
rect 26148 35974 26200 35980
rect 26160 35494 26188 35974
rect 26252 35834 26280 36110
rect 26240 35828 26292 35834
rect 26240 35770 26292 35776
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 26160 35222 26188 35430
rect 26148 35216 26200 35222
rect 26148 35158 26200 35164
rect 26252 35086 26280 35770
rect 26344 35698 26372 36110
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 25872 35012 25924 35018
rect 25872 34954 25924 34960
rect 25884 34746 25912 34954
rect 26240 34944 26292 34950
rect 26240 34886 26292 34892
rect 25872 34740 25924 34746
rect 25872 34682 25924 34688
rect 26252 34610 26280 34886
rect 26344 34678 26372 35634
rect 26516 35556 26568 35562
rect 26516 35498 26568 35504
rect 26528 35290 26556 35498
rect 26516 35284 26568 35290
rect 26516 35226 26568 35232
rect 26332 34672 26384 34678
rect 26332 34614 26384 34620
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 25688 34468 25740 34474
rect 25688 34410 25740 34416
rect 25700 33590 25728 34410
rect 26056 34400 26108 34406
rect 26056 34342 26108 34348
rect 26068 34066 26096 34342
rect 26056 34060 26108 34066
rect 26056 34002 26108 34008
rect 26620 33930 26648 36858
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 26792 35148 26844 35154
rect 26792 35090 26844 35096
rect 26804 34542 26832 35090
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 26792 34536 26844 34542
rect 26792 34478 26844 34484
rect 27528 34468 27580 34474
rect 27528 34410 27580 34416
rect 27540 34202 27568 34410
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 27528 34196 27580 34202
rect 27528 34138 27580 34144
rect 26608 33924 26660 33930
rect 26608 33866 26660 33872
rect 25688 33584 25740 33590
rect 25688 33526 25740 33532
rect 25688 33448 25740 33454
rect 25688 33390 25740 33396
rect 25504 32768 25556 32774
rect 25556 32728 25636 32756
rect 25504 32710 25556 32716
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25424 31958 25452 32370
rect 25504 32224 25556 32230
rect 25504 32166 25556 32172
rect 25412 31952 25464 31958
rect 25412 31894 25464 31900
rect 25516 31754 25544 32166
rect 25504 31748 25556 31754
rect 25504 31690 25556 31696
rect 25608 31278 25636 32728
rect 25700 32434 25728 33390
rect 26620 32842 26648 33866
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 30196 32972 30248 32978
rect 30196 32914 30248 32920
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 25964 32836 26016 32842
rect 25964 32778 26016 32784
rect 26608 32836 26660 32842
rect 26608 32778 26660 32784
rect 27344 32836 27396 32842
rect 27344 32778 27396 32784
rect 25976 32473 26004 32778
rect 25962 32464 26018 32473
rect 25688 32428 25740 32434
rect 25962 32399 25964 32408
rect 25688 32370 25740 32376
rect 26016 32399 26018 32408
rect 25964 32370 26016 32376
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25792 31890 25820 32302
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 25780 31884 25832 31890
rect 25780 31826 25832 31832
rect 25596 31272 25648 31278
rect 25596 31214 25648 31220
rect 25688 31272 25740 31278
rect 25688 31214 25740 31220
rect 25318 30968 25374 30977
rect 24860 30932 24912 30938
rect 25318 30903 25374 30912
rect 24860 30874 24912 30880
rect 25700 30734 25728 31214
rect 25792 30802 25820 31826
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25976 30802 26004 31078
rect 26160 30802 26188 31282
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25964 30796 26016 30802
rect 25964 30738 26016 30744
rect 26148 30796 26200 30802
rect 26148 30738 26200 30744
rect 24676 30728 24728 30734
rect 24674 30696 24676 30705
rect 24860 30728 24912 30734
rect 24728 30696 24730 30705
rect 24860 30670 24912 30676
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 25688 30728 25740 30734
rect 25688 30670 25740 30676
rect 24674 30631 24730 30640
rect 24768 30388 24820 30394
rect 24768 30330 24820 30336
rect 24780 29646 24808 30330
rect 24872 29714 24900 30670
rect 25240 30297 25268 30670
rect 26252 30326 26280 32166
rect 26620 31142 26648 32778
rect 27356 32570 27384 32778
rect 28172 32768 28224 32774
rect 28172 32710 28224 32716
rect 27344 32564 27396 32570
rect 27344 32506 27396 32512
rect 27252 32360 27304 32366
rect 27252 32302 27304 32308
rect 27264 32026 27292 32302
rect 27252 32020 27304 32026
rect 27528 32020 27580 32026
rect 27252 31962 27304 31968
rect 27448 31980 27528 32008
rect 26608 31136 26660 31142
rect 26608 31078 26660 31084
rect 26976 31136 27028 31142
rect 26976 31078 27028 31084
rect 26988 30666 27016 31078
rect 26976 30660 27028 30666
rect 26976 30602 27028 30608
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 26240 30320 26292 30326
rect 25226 30288 25282 30297
rect 26240 30262 26292 30268
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 25226 30223 25282 30232
rect 24952 30184 25004 30190
rect 24952 30126 25004 30132
rect 24964 29850 24992 30126
rect 25320 30048 25372 30054
rect 25320 29990 25372 29996
rect 25502 30016 25558 30025
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 25136 29300 25188 29306
rect 25136 29242 25188 29248
rect 24492 29164 24544 29170
rect 24492 29106 24544 29112
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24504 28626 24532 29106
rect 24596 28966 24624 29106
rect 24780 29073 24808 29106
rect 25044 29096 25096 29102
rect 24766 29064 24822 29073
rect 25044 29038 25096 29044
rect 24766 28999 24822 29008
rect 24584 28960 24636 28966
rect 24584 28902 24636 28908
rect 24952 28960 25004 28966
rect 24952 28902 25004 28908
rect 24492 28620 24544 28626
rect 24492 28562 24544 28568
rect 24504 27130 24532 28562
rect 24584 28008 24636 28014
rect 24584 27950 24636 27956
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24596 27062 24624 27950
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24872 27674 24900 27814
rect 24860 27668 24912 27674
rect 24860 27610 24912 27616
rect 24676 27464 24728 27470
rect 24860 27464 24912 27470
rect 24728 27424 24808 27452
rect 24676 27406 24728 27412
rect 24780 27334 24808 27424
rect 24860 27406 24912 27412
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 24584 27056 24636 27062
rect 24584 26998 24636 27004
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24688 26353 24716 26930
rect 24674 26344 24730 26353
rect 24780 26314 24808 27270
rect 24674 26279 24730 26288
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24676 26240 24728 26246
rect 24676 26182 24728 26188
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24504 25770 24532 25842
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24492 25764 24544 25770
rect 24492 25706 24544 25712
rect 24400 25492 24452 25498
rect 24400 25434 24452 25440
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24124 24608 24176 24614
rect 24124 24550 24176 24556
rect 24136 22642 24164 24550
rect 24504 23798 24532 25230
rect 24596 24041 24624 25774
rect 24688 25498 24716 26182
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24780 25430 24808 25706
rect 24768 25424 24820 25430
rect 24768 25366 24820 25372
rect 24872 25294 24900 27406
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 24766 24984 24822 24993
rect 24766 24919 24822 24928
rect 24780 24886 24808 24919
rect 24768 24880 24820 24886
rect 24768 24822 24820 24828
rect 24964 24206 24992 28902
rect 25056 28762 25084 29038
rect 25044 28756 25096 28762
rect 25044 28698 25096 28704
rect 25148 28626 25176 29242
rect 25332 29170 25360 29990
rect 25502 29951 25558 29960
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 25136 28620 25188 28626
rect 25056 28580 25136 28608
rect 25056 24614 25084 28580
rect 25136 28562 25188 28568
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25148 27062 25176 27406
rect 25136 27056 25188 27062
rect 25240 27033 25268 29106
rect 25332 29073 25360 29106
rect 25318 29064 25374 29073
rect 25318 28999 25374 29008
rect 25320 28008 25372 28014
rect 25320 27950 25372 27956
rect 25136 26998 25188 27004
rect 25226 27024 25282 27033
rect 25148 26042 25176 26998
rect 25226 26959 25282 26968
rect 25136 26036 25188 26042
rect 25136 25978 25188 25984
rect 25332 25906 25360 27950
rect 25412 27940 25464 27946
rect 25412 27882 25464 27888
rect 25424 26840 25452 27882
rect 25516 27470 25544 29951
rect 26056 29572 26108 29578
rect 26056 29514 26108 29520
rect 26068 29238 26096 29514
rect 26056 29232 26108 29238
rect 26056 29174 26108 29180
rect 26068 28558 26096 29174
rect 26252 29170 26280 30262
rect 26332 30048 26384 30054
rect 26332 29990 26384 29996
rect 26344 29782 26372 29990
rect 26332 29776 26384 29782
rect 26384 29736 26464 29764
rect 26332 29718 26384 29724
rect 26240 29164 26292 29170
rect 26240 29106 26292 29112
rect 26332 29164 26384 29170
rect 26332 29106 26384 29112
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 26252 28762 26280 28902
rect 26344 28762 26372 29106
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 25872 28552 25924 28558
rect 25872 28494 25924 28500
rect 26056 28552 26108 28558
rect 26240 28552 26292 28558
rect 26056 28494 26108 28500
rect 26160 28500 26240 28506
rect 26160 28494 26292 28500
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25780 28416 25832 28422
rect 25780 28358 25832 28364
rect 25608 28082 25636 28358
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25792 27674 25820 28358
rect 25884 28014 25912 28494
rect 26160 28478 26280 28494
rect 25964 28076 26016 28082
rect 25964 28018 26016 28024
rect 25872 28008 25924 28014
rect 25872 27950 25924 27956
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 25780 27668 25832 27674
rect 25780 27610 25832 27616
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25778 27432 25834 27441
rect 25778 27367 25780 27376
rect 25832 27367 25834 27376
rect 25780 27338 25832 27344
rect 25688 27328 25740 27334
rect 25594 27296 25650 27305
rect 25688 27270 25740 27276
rect 25594 27231 25650 27240
rect 25608 26926 25636 27231
rect 25596 26920 25648 26926
rect 25596 26862 25648 26868
rect 25504 26852 25556 26858
rect 25424 26812 25504 26840
rect 25504 26794 25556 26800
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25412 25832 25464 25838
rect 25134 25800 25190 25809
rect 25412 25774 25464 25780
rect 25134 25735 25136 25744
rect 25188 25735 25190 25744
rect 25136 25706 25188 25712
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25240 24721 25268 24754
rect 25226 24712 25282 24721
rect 25148 24670 25226 24698
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 25148 24206 25176 24670
rect 25226 24647 25282 24656
rect 25332 24596 25360 25230
rect 25424 25226 25452 25774
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25240 24568 25360 24596
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 25136 24200 25188 24206
rect 25136 24142 25188 24148
rect 24582 24032 24638 24041
rect 24582 23967 24638 23976
rect 24492 23792 24544 23798
rect 24490 23760 24492 23769
rect 24544 23760 24546 23769
rect 24688 23730 24716 24142
rect 24872 23730 24900 24142
rect 24950 23760 25006 23769
rect 24490 23695 24546 23704
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24860 23724 24912 23730
rect 25056 23746 25084 24142
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25006 23718 25084 23746
rect 24950 23695 24952 23704
rect 24860 23666 24912 23672
rect 25004 23695 25006 23704
rect 24952 23666 25004 23672
rect 25056 23118 25084 23718
rect 25148 23254 25176 24006
rect 25240 23730 25268 24568
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24400 22636 24452 22642
rect 24400 22578 24452 22584
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24136 22438 24164 22578
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 24044 21350 24072 21830
rect 23860 21304 23980 21332
rect 24032 21344 24084 21350
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23768 18426 23796 18566
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23768 18086 23796 18226
rect 23860 18222 23888 21304
rect 24032 21286 24084 21292
rect 24136 21146 24164 21966
rect 24228 21554 24256 22578
rect 24412 21894 24440 22578
rect 24492 22432 24544 22438
rect 24492 22374 24544 22380
rect 24308 21888 24360 21894
rect 24306 21856 24308 21865
rect 24400 21888 24452 21894
rect 24360 21856 24362 21865
rect 24400 21830 24452 21836
rect 24306 21791 24362 21800
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23952 20058 23980 20402
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23940 19372 23992 19378
rect 24044 19360 24072 20266
rect 23992 19332 24072 19360
rect 23940 19314 23992 19320
rect 23938 19272 23994 19281
rect 23938 19207 23994 19216
rect 23952 18290 23980 19207
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23664 17808 23716 17814
rect 23664 17750 23716 17756
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23584 17338 23612 17614
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23676 17202 23704 17750
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23492 17054 23612 17082
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23492 16046 23520 16934
rect 23584 16590 23612 17054
rect 23572 16584 23624 16590
rect 23664 16584 23716 16590
rect 23572 16526 23624 16532
rect 23662 16552 23664 16561
rect 23716 16552 23718 16561
rect 23296 16040 23348 16046
rect 23480 16040 23532 16046
rect 23348 16000 23428 16028
rect 23296 15982 23348 15988
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23204 15088 23256 15094
rect 22926 15056 22982 15065
rect 23204 15030 23256 15036
rect 22926 14991 22928 15000
rect 22980 14991 22982 15000
rect 22928 14962 22980 14968
rect 22940 13977 22968 14962
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22926 13968 22982 13977
rect 22926 13903 22982 13912
rect 23032 12782 23060 14758
rect 23112 14476 23164 14482
rect 23112 14418 23164 14424
rect 23124 13462 23152 14418
rect 23216 14414 23244 15030
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23204 13796 23256 13802
rect 23204 13738 23256 13744
rect 23112 13456 23164 13462
rect 23112 13398 23164 13404
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 23216 12442 23244 13738
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 23032 12186 23060 12378
rect 22940 12158 23060 12186
rect 22834 11384 22890 11393
rect 22664 11308 22784 11336
rect 22834 11319 22836 11328
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22756 11082 22784 11308
rect 22888 11319 22890 11328
rect 22836 11290 22888 11296
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22744 11076 22796 11082
rect 22744 11018 22796 11024
rect 22652 11008 22704 11014
rect 22704 10956 22784 10962
rect 22652 10950 22784 10956
rect 22664 10934 22784 10950
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22480 10418 22508 10542
rect 22480 10390 22600 10418
rect 22572 9586 22600 10390
rect 22650 9616 22706 9625
rect 22560 9580 22612 9586
rect 22650 9551 22706 9560
rect 22560 9522 22612 9528
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22480 8498 22508 9318
rect 22572 9217 22600 9386
rect 22558 9208 22614 9217
rect 22664 9178 22692 9551
rect 22756 9178 22784 10934
rect 22848 10266 22876 11154
rect 22940 11082 22968 12158
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11354 23060 12038
rect 23308 11880 23336 15302
rect 23400 15026 23428 16000
rect 23480 15982 23532 15988
rect 23584 15162 23612 16526
rect 23662 16487 23718 16496
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23400 14074 23428 14962
rect 23480 14952 23532 14958
rect 23480 14894 23532 14900
rect 23492 14822 23520 14894
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23676 14618 23704 16050
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23400 12442 23428 14010
rect 23492 12730 23520 14350
rect 23768 14113 23796 18022
rect 23860 15570 23888 18158
rect 24044 17882 24072 19332
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24136 17762 24164 21082
rect 24214 20632 24270 20641
rect 24214 20567 24270 20576
rect 24228 20398 24256 20567
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24228 18086 24256 19790
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24044 17734 24164 17762
rect 24044 17066 24072 17734
rect 24228 17678 24256 18022
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 24044 16794 24072 17002
rect 24136 16833 24164 17002
rect 24122 16824 24178 16833
rect 24032 16788 24084 16794
rect 24122 16759 24178 16768
rect 24032 16730 24084 16736
rect 24032 16516 24084 16522
rect 24032 16458 24084 16464
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 24044 15162 24072 16458
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24136 15881 24164 16050
rect 24320 15978 24348 21490
rect 24412 21332 24440 21830
rect 24504 21690 24532 22374
rect 24584 22092 24636 22098
rect 24584 22034 24636 22040
rect 24596 22001 24624 22034
rect 24582 21992 24638 22001
rect 24582 21927 24638 21936
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24688 21554 24716 22578
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24674 21448 24730 21457
rect 24674 21383 24730 21392
rect 24492 21344 24544 21350
rect 24412 21312 24492 21332
rect 24544 21312 24546 21321
rect 24412 21304 24490 21312
rect 24490 21247 24546 21256
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24584 19848 24636 19854
rect 24584 19790 24636 19796
rect 24412 19514 24440 19790
rect 24490 19680 24546 19689
rect 24490 19615 24546 19624
rect 24400 19508 24452 19514
rect 24400 19450 24452 19456
rect 24398 19408 24454 19417
rect 24504 19378 24532 19615
rect 24398 19343 24400 19352
rect 24452 19343 24454 19352
rect 24492 19372 24544 19378
rect 24400 19314 24452 19320
rect 24492 19314 24544 19320
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18766 24440 19110
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24504 18426 24532 18566
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24596 18057 24624 19790
rect 24688 19292 24716 21383
rect 24780 20466 24808 22374
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24872 22030 24900 22170
rect 25042 22128 25098 22137
rect 25042 22063 25098 22072
rect 25056 22030 25084 22063
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 24952 21956 25004 21962
rect 24952 21898 25004 21904
rect 24964 21729 24992 21898
rect 24950 21720 25006 21729
rect 24950 21655 25006 21664
rect 24950 21584 25006 21593
rect 24950 21519 25006 21528
rect 24964 21350 24992 21519
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24860 20256 24912 20262
rect 24912 20216 24992 20244
rect 24860 20198 24912 20204
rect 24860 20052 24912 20058
rect 24860 19994 24912 20000
rect 24766 19680 24822 19689
rect 24766 19615 24822 19624
rect 24780 19514 24808 19615
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24872 19378 24900 19994
rect 24964 19854 24992 20216
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24688 19264 24808 19292
rect 24674 19136 24730 19145
rect 24674 19071 24730 19080
rect 24688 18766 24716 19071
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24582 18048 24638 18057
rect 24582 17983 24638 17992
rect 24400 17196 24452 17202
rect 24400 17138 24452 17144
rect 24412 17105 24440 17138
rect 24398 17096 24454 17105
rect 24688 17066 24716 18702
rect 24780 18222 24808 19264
rect 24964 19258 24992 19790
rect 25056 19378 25084 20402
rect 25148 20330 25176 22986
rect 25240 22964 25268 23666
rect 25332 23118 25360 23666
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25320 22976 25372 22982
rect 25240 22936 25320 22964
rect 25240 21418 25268 22936
rect 25320 22918 25372 22924
rect 25424 21593 25452 25162
rect 25516 24138 25544 26794
rect 25700 26353 25728 27270
rect 25884 26382 25912 27814
rect 25976 27130 26004 28018
rect 26160 27826 26188 28478
rect 26344 28257 26372 28698
rect 26436 28490 26464 29736
rect 26620 29646 26648 30262
rect 27356 30258 27384 30534
rect 27344 30252 27396 30258
rect 27344 30194 27396 30200
rect 27448 29753 27476 31980
rect 27528 31962 27580 31968
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27632 31278 27660 31758
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27620 31272 27672 31278
rect 27620 31214 27672 31220
rect 27620 31136 27672 31142
rect 27620 31078 27672 31084
rect 27712 31136 27764 31142
rect 27712 31078 27764 31084
rect 27526 30288 27582 30297
rect 27526 30223 27528 30232
rect 27580 30223 27582 30232
rect 27528 30194 27580 30200
rect 27632 30122 27660 31078
rect 27724 30734 27752 31078
rect 27816 30870 27844 31690
rect 28080 31680 28132 31686
rect 28000 31628 28080 31634
rect 28000 31622 28132 31628
rect 28000 31606 28120 31622
rect 28000 31414 28028 31606
rect 28184 31498 28212 32710
rect 28828 32298 28856 32846
rect 28908 32496 28960 32502
rect 28908 32438 28960 32444
rect 28816 32292 28868 32298
rect 28816 32234 28868 32240
rect 28724 32224 28776 32230
rect 28724 32166 28776 32172
rect 28264 31952 28316 31958
rect 28264 31894 28316 31900
rect 28538 31920 28594 31929
rect 28092 31470 28212 31498
rect 28092 31414 28120 31470
rect 27988 31408 28040 31414
rect 27988 31350 28040 31356
rect 28080 31408 28132 31414
rect 28080 31350 28132 31356
rect 28276 31278 28304 31894
rect 28448 31884 28500 31890
rect 28538 31855 28594 31864
rect 28448 31826 28500 31832
rect 28460 31754 28488 31826
rect 28552 31788 28580 31855
rect 28368 31726 28488 31754
rect 28540 31782 28592 31788
rect 28368 31346 28396 31726
rect 28540 31724 28592 31730
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28356 31340 28408 31346
rect 28356 31282 28408 31288
rect 28264 31272 28316 31278
rect 28460 31226 28488 31622
rect 28736 31346 28764 32166
rect 28724 31340 28776 31346
rect 28724 31282 28776 31288
rect 28264 31214 28316 31220
rect 28368 31198 28488 31226
rect 27804 30864 27856 30870
rect 27804 30806 27856 30812
rect 28172 30796 28224 30802
rect 28172 30738 28224 30744
rect 27712 30728 27764 30734
rect 27712 30670 27764 30676
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 27620 30116 27672 30122
rect 27620 30058 27672 30064
rect 27896 30116 27948 30122
rect 27896 30058 27948 30064
rect 27988 30116 28040 30122
rect 27988 30058 28040 30064
rect 27802 30016 27858 30025
rect 27802 29951 27858 29960
rect 27620 29844 27672 29850
rect 27620 29786 27672 29792
rect 27434 29744 27490 29753
rect 26896 29714 27108 29730
rect 26884 29708 27108 29714
rect 26936 29702 27108 29708
rect 26884 29650 26936 29656
rect 26608 29640 26660 29646
rect 26660 29600 26740 29628
rect 26608 29582 26660 29588
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26528 28529 26556 29242
rect 26608 28620 26660 28626
rect 26608 28562 26660 28568
rect 26514 28520 26570 28529
rect 26424 28484 26476 28490
rect 26514 28455 26570 28464
rect 26424 28426 26476 28432
rect 26330 28248 26386 28257
rect 26330 28183 26386 28192
rect 26436 27878 26464 28426
rect 26516 28416 26568 28422
rect 26516 28358 26568 28364
rect 26424 27872 26476 27878
rect 26160 27798 26280 27826
rect 26424 27814 26476 27820
rect 26056 27396 26108 27402
rect 26056 27338 26108 27344
rect 25964 27124 26016 27130
rect 25964 27066 26016 27072
rect 26068 27033 26096 27338
rect 26252 27334 26280 27798
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26054 27024 26110 27033
rect 26054 26959 26110 26968
rect 26252 26790 26280 27270
rect 26332 27056 26384 27062
rect 26332 26998 26384 27004
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26148 26580 26200 26586
rect 26148 26522 26200 26528
rect 25872 26376 25924 26382
rect 25686 26344 25742 26353
rect 25872 26318 25924 26324
rect 25686 26279 25742 26288
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25504 23792 25556 23798
rect 25504 23734 25556 23740
rect 25516 23050 25544 23734
rect 25608 23730 25636 24006
rect 25700 23866 25728 25842
rect 25792 25430 25820 25978
rect 25780 25424 25832 25430
rect 25780 25366 25832 25372
rect 25884 24750 25912 26318
rect 25962 25936 26018 25945
rect 25962 25871 25964 25880
rect 26016 25871 26018 25880
rect 25964 25842 26016 25848
rect 25976 25294 26004 25842
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 25872 24744 25924 24750
rect 25872 24686 25924 24692
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25884 24206 25912 24550
rect 25976 24410 26004 24550
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 26068 24290 26096 25094
rect 25976 24262 26096 24290
rect 25780 24200 25832 24206
rect 25780 24142 25832 24148
rect 25872 24200 25924 24206
rect 25872 24142 25924 24148
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25686 23760 25742 23769
rect 25596 23724 25648 23730
rect 25686 23695 25688 23704
rect 25596 23666 25648 23672
rect 25740 23695 25742 23704
rect 25688 23666 25740 23672
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25504 23044 25556 23050
rect 25504 22986 25556 22992
rect 25516 22778 25544 22986
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25608 21842 25636 23190
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25700 22030 25728 23054
rect 25792 22094 25820 24142
rect 25792 22066 25912 22094
rect 25688 22024 25740 22030
rect 25686 21992 25688 22001
rect 25740 21992 25742 22001
rect 25686 21927 25742 21936
rect 25608 21814 25728 21842
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25608 21593 25636 21626
rect 25410 21584 25466 21593
rect 25410 21519 25466 21528
rect 25594 21584 25650 21593
rect 25594 21519 25650 21528
rect 25228 21412 25280 21418
rect 25228 21354 25280 21360
rect 25320 20392 25372 20398
rect 25320 20334 25372 20340
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25240 19378 25268 19722
rect 25332 19446 25360 20334
rect 25410 19952 25466 19961
rect 25410 19887 25412 19896
rect 25464 19887 25466 19896
rect 25412 19858 25464 19864
rect 25320 19440 25372 19446
rect 25320 19382 25372 19388
rect 25596 19440 25648 19446
rect 25596 19382 25648 19388
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 24872 19230 24992 19258
rect 24768 18216 24820 18222
rect 24766 18184 24768 18193
rect 24820 18184 24822 18193
rect 24766 18119 24822 18128
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24398 17031 24454 17040
rect 24676 17060 24728 17066
rect 24676 17002 24728 17008
rect 24398 16688 24454 16697
rect 24398 16623 24454 16632
rect 24412 16522 24440 16623
rect 24400 16516 24452 16522
rect 24400 16458 24452 16464
rect 24780 16250 24808 17274
rect 24872 16590 24900 19230
rect 25056 18970 25084 19314
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 25148 18850 25176 19246
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 25056 18822 25176 18850
rect 24964 18290 24992 18770
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24964 17678 24992 18226
rect 24952 17672 25004 17678
rect 25056 17649 25084 18822
rect 25228 18692 25280 18698
rect 25148 18652 25228 18680
rect 25148 18290 25176 18652
rect 25228 18634 25280 18640
rect 25332 18442 25360 19382
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25424 18970 25452 19314
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25516 18630 25544 19314
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25332 18414 25544 18442
rect 25320 18352 25372 18358
rect 25318 18320 25320 18329
rect 25372 18320 25374 18329
rect 25136 18284 25188 18290
rect 25318 18255 25374 18264
rect 25136 18226 25188 18232
rect 25320 18148 25372 18154
rect 25320 18090 25372 18096
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17882 25268 18022
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25240 17785 25268 17818
rect 25226 17776 25282 17785
rect 25226 17711 25282 17720
rect 24952 17614 25004 17620
rect 25042 17640 25098 17649
rect 25042 17575 25044 17584
rect 25096 17575 25098 17584
rect 25044 17546 25096 17552
rect 25240 17338 25268 17711
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 24950 17232 25006 17241
rect 24950 17167 25006 17176
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24492 16108 24544 16114
rect 24492 16050 24544 16056
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24504 16017 24532 16050
rect 24490 16008 24546 16017
rect 24308 15972 24360 15978
rect 24490 15943 24546 15952
rect 24308 15914 24360 15920
rect 24122 15872 24178 15881
rect 24122 15807 24178 15816
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 24044 14822 24072 15098
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23754 14104 23810 14113
rect 23754 14039 23810 14048
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23584 12850 23612 13126
rect 23676 12850 23704 13194
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23492 12702 23612 12730
rect 23388 12436 23440 12442
rect 23584 12434 23612 12702
rect 23768 12442 23796 14039
rect 23388 12378 23440 12384
rect 23492 12406 23612 12434
rect 23664 12436 23716 12442
rect 23386 12200 23442 12209
rect 23386 12135 23388 12144
rect 23440 12135 23442 12144
rect 23388 12106 23440 12112
rect 23216 11852 23336 11880
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 22928 10600 22980 10606
rect 22928 10542 22980 10548
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22940 10130 22968 10542
rect 23018 10432 23074 10441
rect 23018 10367 23074 10376
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 22940 9586 22968 9930
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 23032 9450 23060 10367
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 22836 9376 22888 9382
rect 22834 9344 22836 9353
rect 22888 9344 22890 9353
rect 22834 9279 22890 9288
rect 22558 9143 22614 9152
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22572 8634 22600 9046
rect 22756 8786 22784 9114
rect 23124 8974 23152 10950
rect 23216 9586 23244 11852
rect 23400 11830 23428 12106
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23296 11756 23348 11762
rect 23296 11698 23348 11704
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23112 8968 23164 8974
rect 22848 8906 23060 8922
rect 23112 8910 23164 8916
rect 22836 8900 23060 8906
rect 22888 8894 23060 8900
rect 22836 8842 22888 8848
rect 22664 8758 22784 8786
rect 22928 8832 22980 8838
rect 22928 8774 22980 8780
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22664 7478 22692 8758
rect 22742 8664 22798 8673
rect 22742 8599 22744 8608
rect 22796 8599 22798 8608
rect 22744 8570 22796 8576
rect 22940 7750 22968 8774
rect 23032 8673 23060 8894
rect 23018 8664 23074 8673
rect 23018 8599 23074 8608
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22940 7410 22968 7686
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 22664 7002 22692 7142
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23124 6458 23152 6734
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23020 6180 23072 6186
rect 23020 6122 23072 6128
rect 23032 5710 23060 6122
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22376 5296 22428 5302
rect 22560 5296 22612 5302
rect 22376 5238 22428 5244
rect 22558 5264 22560 5273
rect 22612 5264 22614 5273
rect 22558 5199 22614 5208
rect 22284 4548 22336 4554
rect 22572 4536 22600 5199
rect 22940 4826 22968 5646
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 23308 4706 23336 11698
rect 23400 11665 23428 11766
rect 23386 11656 23442 11665
rect 23386 11591 23442 11600
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 23400 9382 23428 11222
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23400 7002 23428 7414
rect 23388 6996 23440 7002
rect 23388 6938 23440 6944
rect 23492 6798 23520 12406
rect 23664 12378 23716 12384
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 23584 11218 23612 12106
rect 23676 11830 23704 12378
rect 23754 11928 23810 11937
rect 23754 11863 23810 11872
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23662 11520 23718 11529
rect 23662 11455 23718 11464
rect 23676 11354 23704 11455
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23584 10674 23612 11018
rect 23676 10674 23704 11290
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23664 10668 23716 10674
rect 23664 10610 23716 10616
rect 23768 10146 23796 11863
rect 23860 11694 23888 14554
rect 23938 14512 23994 14521
rect 23938 14447 23994 14456
rect 23952 14346 23980 14447
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 23952 13734 23980 14282
rect 23940 13728 23992 13734
rect 23940 13670 23992 13676
rect 24044 12481 24072 14758
rect 24030 12472 24086 12481
rect 24030 12407 24086 12416
rect 24044 12238 24072 12407
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 23940 12164 23992 12170
rect 23940 12106 23992 12112
rect 23952 11937 23980 12106
rect 23938 11928 23994 11937
rect 23938 11863 23994 11872
rect 23848 11688 23900 11694
rect 23848 11630 23900 11636
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23860 11121 23888 11494
rect 23938 11384 23994 11393
rect 23938 11319 23994 11328
rect 23846 11112 23902 11121
rect 23846 11047 23902 11056
rect 23860 11014 23888 11047
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23846 10840 23902 10849
rect 23846 10775 23902 10784
rect 23860 10742 23888 10775
rect 23848 10736 23900 10742
rect 23848 10678 23900 10684
rect 23952 10554 23980 11319
rect 23676 10118 23796 10146
rect 23860 10526 23980 10554
rect 23570 9480 23626 9489
rect 23570 9415 23572 9424
rect 23624 9415 23626 9424
rect 23572 9386 23624 9392
rect 23676 7546 23704 10118
rect 23860 10010 23888 10526
rect 23940 10464 23992 10470
rect 23938 10432 23940 10441
rect 23992 10432 23994 10441
rect 23938 10367 23994 10376
rect 23768 9982 23888 10010
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23768 7886 23796 9982
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23860 8566 23888 9590
rect 23952 8906 23980 9998
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23676 6882 23704 7482
rect 23768 7449 23796 7822
rect 23754 7440 23810 7449
rect 23754 7375 23810 7384
rect 23860 7342 23888 8502
rect 23952 8498 23980 8842
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23952 7478 23980 8434
rect 24044 8090 24072 12174
rect 24136 8430 24164 15807
rect 24596 15609 24624 16050
rect 24582 15600 24638 15609
rect 24582 15535 24638 15544
rect 24768 15496 24820 15502
rect 24768 15438 24820 15444
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24216 15088 24268 15094
rect 24214 15056 24216 15065
rect 24268 15056 24270 15065
rect 24214 14991 24270 15000
rect 24400 14952 24452 14958
rect 24400 14894 24452 14900
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24228 12850 24256 14758
rect 24412 14618 24440 14894
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24228 11529 24256 12650
rect 24412 12442 24440 12718
rect 24308 12436 24360 12442
rect 24308 12378 24360 12384
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24320 12238 24348 12378
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24400 12164 24452 12170
rect 24400 12106 24452 12112
rect 24214 11520 24270 11529
rect 24412 11506 24440 12106
rect 24504 11558 24532 15370
rect 24780 15026 24808 15438
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24858 14920 24914 14929
rect 24858 14855 24914 14864
rect 24768 14816 24820 14822
rect 24766 14784 24768 14793
rect 24820 14784 24822 14793
rect 24766 14719 24822 14728
rect 24872 14414 24900 14855
rect 24964 14498 24992 17167
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 25056 16182 25084 16934
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 25056 15570 25084 16118
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 25042 15192 25098 15201
rect 25042 15127 25098 15136
rect 25056 14958 25084 15127
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24964 14470 25084 14498
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24674 13696 24730 13705
rect 24674 13631 24730 13640
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24596 12594 24624 12854
rect 24688 12714 24716 13631
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 12782 24808 13262
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24676 12708 24728 12714
rect 24676 12650 24728 12656
rect 24596 12566 24716 12594
rect 24214 11455 24270 11464
rect 24320 11478 24440 11506
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24228 10674 24256 11290
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24320 9994 24348 11478
rect 24490 11248 24546 11257
rect 24490 11183 24546 11192
rect 24504 11150 24532 11183
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24596 11082 24624 11494
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24490 10840 24546 10849
rect 24490 10775 24546 10784
rect 24504 10742 24532 10775
rect 24492 10736 24544 10742
rect 24492 10678 24544 10684
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24308 9988 24360 9994
rect 24308 9930 24360 9936
rect 24412 9586 24440 10406
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24504 9466 24532 10678
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24596 9722 24624 10406
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24320 9438 24532 9466
rect 24124 8424 24176 8430
rect 24124 8366 24176 8372
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 23940 7472 23992 7478
rect 23940 7414 23992 7420
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 23584 6854 23704 6882
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23480 6656 23532 6662
rect 23584 6644 23612 6854
rect 23860 6730 23888 7142
rect 23664 6724 23716 6730
rect 23664 6666 23716 6672
rect 23848 6724 23900 6730
rect 23848 6666 23900 6672
rect 23532 6616 23612 6644
rect 23480 6598 23532 6604
rect 23676 6322 23704 6666
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23860 5914 23888 6666
rect 23952 6662 23980 7414
rect 24136 7410 24164 7890
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23952 6186 23980 6598
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23952 5846 23980 6122
rect 23940 5840 23992 5846
rect 23386 5808 23442 5817
rect 23940 5782 23992 5788
rect 23386 5743 23442 5752
rect 23400 5710 23428 5743
rect 23388 5704 23440 5710
rect 23388 5646 23440 5652
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23124 4690 23336 4706
rect 23112 4684 23336 4690
rect 23164 4678 23336 4684
rect 23112 4626 23164 4632
rect 22652 4548 22704 4554
rect 22572 4508 22652 4536
rect 22284 4490 22336 4496
rect 22652 4490 22704 4496
rect 22664 4214 22692 4490
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 23308 4146 23336 4678
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23308 3602 23336 4082
rect 23584 4078 23612 5510
rect 23952 4078 23980 5646
rect 24320 5250 24348 9438
rect 24596 9330 24624 9522
rect 24412 9302 24624 9330
rect 24412 9178 24440 9302
rect 24400 9172 24452 9178
rect 24688 9160 24716 12566
rect 24872 12102 24900 14350
rect 24964 13870 24992 14350
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24964 13705 24992 13806
rect 24950 13696 25006 13705
rect 24950 13631 25006 13640
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11756 24820 11762
rect 24768 11698 24820 11704
rect 24780 10674 24808 11698
rect 24872 11354 24900 11766
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24768 10668 24820 10674
rect 24820 10628 24900 10656
rect 24768 10610 24820 10616
rect 24400 9114 24452 9120
rect 24504 9132 24716 9160
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 24412 8498 24440 8570
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 24412 7721 24440 8298
rect 24398 7712 24454 7721
rect 24398 7647 24454 7656
rect 24504 7546 24532 9132
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24596 8498 24624 8774
rect 24688 8634 24716 8910
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24688 8004 24716 8434
rect 24596 7976 24716 8004
rect 24596 7886 24624 7976
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24412 6390 24440 7346
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 24596 6254 24624 7822
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24688 6798 24716 7754
rect 24780 7732 24808 8434
rect 24872 7886 24900 10628
rect 24860 7880 24912 7886
rect 24860 7822 24912 7828
rect 24780 7704 24900 7732
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24780 6934 24808 7278
rect 24768 6928 24820 6934
rect 24768 6870 24820 6876
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24768 6792 24820 6798
rect 24872 6780 24900 7704
rect 24820 6752 24900 6780
rect 24768 6734 24820 6740
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24674 5808 24730 5817
rect 24492 5772 24544 5778
rect 24674 5743 24730 5752
rect 24492 5714 24544 5720
rect 24504 5574 24532 5714
rect 24688 5710 24716 5743
rect 24780 5710 24808 6122
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 24320 5234 24440 5250
rect 24504 5234 24532 5510
rect 24780 5302 24808 5646
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24320 5228 24452 5234
rect 24320 5222 24400 5228
rect 24400 5170 24452 5176
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24412 5030 24440 5170
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24872 4690 24900 5170
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23940 3664 23992 3670
rect 23940 3606 23992 3612
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 23308 3126 23336 3538
rect 23296 3120 23348 3126
rect 23296 3062 23348 3068
rect 23952 3058 23980 3606
rect 24044 3466 24072 4150
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24032 3460 24084 3466
rect 24032 3402 24084 3408
rect 24044 3194 24072 3402
rect 24872 3194 24900 4082
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 18984 2650 19012 2926
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19720 2514 19748 2790
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 18602 1799 18658 1808
rect 18708 1822 18828 1850
rect 17420 1142 17540 1170
rect 17420 800 17448 1142
rect 18708 800 18736 1822
rect 23860 800 23888 2790
rect 24964 2446 24992 12650
rect 25056 12186 25084 14470
rect 25148 12345 25176 16186
rect 25240 14890 25268 17274
rect 25332 17270 25360 18090
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25332 15910 25360 17206
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25424 15706 25452 16526
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25516 15042 25544 18414
rect 25608 17066 25636 19382
rect 25700 18698 25728 21814
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25792 19718 25820 20266
rect 25884 19990 25912 22066
rect 25872 19984 25924 19990
rect 25872 19926 25924 19932
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25688 18352 25740 18358
rect 25686 18320 25688 18329
rect 25740 18320 25742 18329
rect 25686 18255 25742 18264
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25700 17678 25728 18022
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25596 17060 25648 17066
rect 25596 17002 25648 17008
rect 25608 16969 25636 17002
rect 25594 16960 25650 16969
rect 25594 16895 25650 16904
rect 25700 16590 25728 17138
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25700 16454 25728 16526
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25792 16402 25820 19314
rect 25870 19000 25926 19009
rect 25870 18935 25926 18944
rect 25884 18834 25912 18935
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25884 17338 25912 17614
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25976 16726 26004 24262
rect 26054 23760 26110 23769
rect 26054 23695 26056 23704
rect 26108 23695 26110 23704
rect 26056 23666 26108 23672
rect 26160 23322 26188 26522
rect 26344 26450 26372 26998
rect 26332 26444 26384 26450
rect 26332 26386 26384 26392
rect 26424 26376 26476 26382
rect 26424 26318 26476 26324
rect 26436 25974 26464 26318
rect 26424 25968 26476 25974
rect 26424 25910 26476 25916
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26252 24886 26280 25842
rect 26424 25288 26476 25294
rect 26424 25230 26476 25236
rect 26240 24880 26292 24886
rect 26240 24822 26292 24828
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26148 23316 26200 23322
rect 26148 23258 26200 23264
rect 26148 23112 26200 23118
rect 26146 23080 26148 23089
rect 26200 23080 26202 23089
rect 26146 23015 26202 23024
rect 26148 22772 26200 22778
rect 26148 22714 26200 22720
rect 26160 22098 26188 22714
rect 26252 22166 26280 24618
rect 26436 24449 26464 25230
rect 26422 24440 26478 24449
rect 26528 24410 26556 28358
rect 26620 26586 26648 28562
rect 26712 28558 26740 29600
rect 26884 29572 26936 29578
rect 26884 29514 26936 29520
rect 26790 29064 26846 29073
rect 26896 29034 26924 29514
rect 26976 29096 27028 29102
rect 26976 29038 27028 29044
rect 27080 29050 27108 29702
rect 27434 29679 27490 29688
rect 27252 29572 27304 29578
rect 27252 29514 27304 29520
rect 27160 29504 27212 29510
rect 27160 29446 27212 29452
rect 27172 29170 27200 29446
rect 27264 29306 27292 29514
rect 27252 29300 27304 29306
rect 27252 29242 27304 29248
rect 27160 29164 27212 29170
rect 27344 29164 27396 29170
rect 27160 29106 27212 29112
rect 27264 29124 27344 29152
rect 27264 29073 27292 29124
rect 27344 29106 27396 29112
rect 27250 29064 27306 29073
rect 26790 28999 26792 29008
rect 26844 28999 26846 29008
rect 26884 29028 26936 29034
rect 26792 28970 26844 28976
rect 26884 28970 26936 28976
rect 26896 28694 26924 28970
rect 26884 28688 26936 28694
rect 26884 28630 26936 28636
rect 26988 28558 27016 29038
rect 27080 29022 27200 29050
rect 26700 28552 26752 28558
rect 26700 28494 26752 28500
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 26804 28422 26832 28494
rect 26792 28416 26844 28422
rect 26792 28358 26844 28364
rect 26804 27470 26832 28358
rect 26884 28008 26936 28014
rect 26884 27950 26936 27956
rect 26896 27674 26924 27950
rect 26884 27668 26936 27674
rect 26884 27610 26936 27616
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26698 27024 26754 27033
rect 26698 26959 26754 26968
rect 26792 26988 26844 26994
rect 26608 26580 26660 26586
rect 26608 26522 26660 26528
rect 26620 26314 26648 26522
rect 26712 26314 26740 26959
rect 26792 26930 26844 26936
rect 26608 26308 26660 26314
rect 26608 26250 26660 26256
rect 26700 26308 26752 26314
rect 26700 26250 26752 26256
rect 26620 24818 26648 26250
rect 26804 25158 26832 26930
rect 26896 26450 26924 27610
rect 26988 27062 27016 28494
rect 27068 27396 27120 27402
rect 27068 27338 27120 27344
rect 26976 27056 27028 27062
rect 26976 26998 27028 27004
rect 26988 26586 27016 26998
rect 26976 26580 27028 26586
rect 26976 26522 27028 26528
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26884 25968 26936 25974
rect 26884 25910 26936 25916
rect 26792 25152 26844 25158
rect 26792 25094 26844 25100
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26700 24812 26752 24818
rect 26700 24754 26752 24760
rect 26422 24375 26478 24384
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26332 24200 26384 24206
rect 26332 24142 26384 24148
rect 26344 23322 26372 24142
rect 26516 23860 26568 23866
rect 26516 23802 26568 23808
rect 26332 23316 26384 23322
rect 26332 23258 26384 23264
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26240 22160 26292 22166
rect 26240 22102 26292 22108
rect 26148 22092 26200 22098
rect 26148 22034 26200 22040
rect 26056 21888 26108 21894
rect 26056 21830 26108 21836
rect 26068 19174 26096 21830
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26252 19854 26280 20198
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26252 19242 26280 19790
rect 26436 19258 26464 23054
rect 26528 22953 26556 23802
rect 26606 23352 26662 23361
rect 26606 23287 26662 23296
rect 26514 22944 26570 22953
rect 26514 22879 26570 22888
rect 26620 22760 26648 23287
rect 26712 23118 26740 24754
rect 26896 24018 26924 25910
rect 26988 25906 27016 26522
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 26988 24954 27016 25842
rect 27080 25401 27108 27338
rect 27066 25392 27122 25401
rect 27066 25327 27122 25336
rect 27080 25158 27108 25327
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 27172 24750 27200 29022
rect 27250 28999 27306 29008
rect 27160 24744 27212 24750
rect 27160 24686 27212 24692
rect 27172 24614 27200 24686
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26804 23990 26924 24018
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 26620 22732 26740 22760
rect 26608 22568 26660 22574
rect 26608 22510 26660 22516
rect 26620 22030 26648 22510
rect 26516 22024 26568 22030
rect 26516 21966 26568 21972
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26528 21078 26556 21966
rect 26620 21894 26648 21966
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26516 21072 26568 21078
rect 26516 21014 26568 21020
rect 26606 21040 26662 21049
rect 26606 20975 26662 20984
rect 26620 20924 26648 20975
rect 26528 20896 26648 20924
rect 26528 19718 26556 20896
rect 26606 20632 26662 20641
rect 26606 20567 26608 20576
rect 26660 20567 26662 20576
rect 26608 20538 26660 20544
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26516 19712 26568 19718
rect 26514 19680 26516 19689
rect 26568 19680 26570 19689
rect 26514 19615 26570 19624
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 26332 19236 26384 19242
rect 26436 19230 26556 19258
rect 26332 19178 26384 19184
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26056 18284 26108 18290
rect 26056 18226 26108 18232
rect 25964 16720 26016 16726
rect 25962 16688 25964 16697
rect 26016 16688 26018 16697
rect 25962 16623 26018 16632
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 25700 16114 25728 16390
rect 25792 16374 25912 16402
rect 25778 16280 25834 16289
rect 25778 16215 25780 16224
rect 25832 16215 25834 16224
rect 25780 16186 25832 16192
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 25700 15502 25728 16050
rect 25688 15496 25740 15502
rect 25688 15438 25740 15444
rect 25320 15020 25372 15026
rect 25516 15014 25820 15042
rect 25320 14962 25372 14968
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25240 12986 25268 14826
rect 25332 14793 25360 14962
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25318 14784 25374 14793
rect 25374 14742 25452 14770
rect 25318 14719 25374 14728
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25134 12336 25190 12345
rect 25134 12271 25190 12280
rect 25056 12158 25360 12186
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25056 11762 25084 12038
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25056 11218 25084 11698
rect 25148 11354 25176 11834
rect 25240 11762 25268 12038
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25240 11014 25268 11698
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25240 10674 25268 10950
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25240 10062 25268 10610
rect 25332 10606 25360 12158
rect 25424 11830 25452 14742
rect 25700 14414 25728 14894
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25608 13870 25636 14350
rect 25700 13938 25728 14350
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25700 13394 25728 13874
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25608 12850 25636 13262
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25516 11694 25544 12718
rect 25412 11688 25464 11694
rect 25412 11630 25464 11636
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25424 11354 25452 11630
rect 25412 11348 25464 11354
rect 25412 11290 25464 11296
rect 25424 10674 25452 11290
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25228 10056 25280 10062
rect 25228 9998 25280 10004
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 25136 9512 25188 9518
rect 25136 9454 25188 9460
rect 25056 9178 25084 9454
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25148 9058 25176 9454
rect 25056 9030 25176 9058
rect 25056 6458 25084 9030
rect 25240 6730 25268 9998
rect 25332 7410 25360 10542
rect 25412 10532 25464 10538
rect 25412 10474 25464 10480
rect 25424 10266 25452 10474
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25516 9586 25544 11630
rect 25608 11218 25636 12786
rect 25700 12782 25728 13330
rect 25688 12776 25740 12782
rect 25792 12753 25820 15014
rect 25884 14890 25912 16374
rect 25976 15978 26004 16526
rect 25964 15972 26016 15978
rect 25964 15914 26016 15920
rect 25976 15366 26004 15914
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25872 14884 25924 14890
rect 25872 14826 25924 14832
rect 25884 12918 25912 14826
rect 26068 14482 26096 18226
rect 26160 18086 26188 19110
rect 26344 18766 26372 19178
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26252 18426 26280 18702
rect 26436 18698 26464 19110
rect 26424 18692 26476 18698
rect 26424 18634 26476 18640
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 26160 17202 26188 18022
rect 26238 17912 26294 17921
rect 26344 17898 26372 18566
rect 26422 18456 26478 18465
rect 26422 18391 26424 18400
rect 26476 18391 26478 18400
rect 26424 18362 26476 18368
rect 26294 17870 26372 17898
rect 26238 17847 26294 17856
rect 26252 17746 26280 17847
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26332 16176 26384 16182
rect 26332 16118 26384 16124
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 15706 26188 15982
rect 26148 15700 26200 15706
rect 26148 15642 26200 15648
rect 26148 15360 26200 15366
rect 26344 15314 26372 16118
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26148 15302 26200 15308
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 26068 14385 26096 14418
rect 26054 14376 26110 14385
rect 26054 14311 26110 14320
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 25962 13424 26018 13433
rect 25962 13359 26018 13368
rect 25872 12912 25924 12918
rect 25872 12854 25924 12860
rect 25688 12718 25740 12724
rect 25778 12744 25834 12753
rect 25778 12679 25834 12688
rect 25872 12708 25924 12714
rect 25686 12336 25742 12345
rect 25686 12271 25742 12280
rect 25700 11370 25728 12271
rect 25792 11626 25820 12679
rect 25872 12650 25924 12656
rect 25884 12238 25912 12650
rect 25872 12232 25924 12238
rect 25872 12174 25924 12180
rect 25780 11620 25832 11626
rect 25780 11562 25832 11568
rect 25700 11342 25820 11370
rect 25596 11212 25648 11218
rect 25648 11172 25728 11200
rect 25596 11154 25648 11160
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 25608 10810 25636 11018
rect 25596 10804 25648 10810
rect 25596 10746 25648 10752
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25608 9994 25636 10610
rect 25700 10130 25728 11172
rect 25688 10124 25740 10130
rect 25688 10066 25740 10072
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25424 7546 25452 9318
rect 25516 8566 25544 9522
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 25504 8560 25556 8566
rect 25504 8502 25556 8508
rect 25504 8356 25556 8362
rect 25608 8344 25636 9046
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 25700 8673 25728 8978
rect 25686 8664 25742 8673
rect 25686 8599 25742 8608
rect 25556 8316 25636 8344
rect 25504 8298 25556 8304
rect 25516 8265 25544 8298
rect 25502 8256 25558 8265
rect 25502 8191 25558 8200
rect 25504 8016 25556 8022
rect 25504 7958 25556 7964
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25516 7410 25544 7958
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25608 7546 25636 7754
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 25148 6118 25176 6598
rect 25700 6118 25728 7822
rect 25792 7342 25820 11342
rect 25872 11280 25924 11286
rect 25872 11222 25924 11228
rect 25884 9450 25912 11222
rect 25976 9518 26004 13359
rect 26068 13326 26096 14214
rect 26056 13320 26108 13326
rect 26056 13262 26108 13268
rect 26160 12442 26188 15302
rect 26252 15286 26372 15314
rect 26252 13734 26280 15286
rect 26330 15192 26386 15201
rect 26330 15127 26332 15136
rect 26384 15127 26386 15136
rect 26332 15098 26384 15104
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26436 13530 26464 15438
rect 26528 14385 26556 19230
rect 26620 18601 26648 20402
rect 26606 18592 26662 18601
rect 26606 18527 26662 18536
rect 26712 16232 26740 22732
rect 26804 21894 26832 23990
rect 27172 23905 27200 24142
rect 27158 23896 27214 23905
rect 27158 23831 27214 23840
rect 27264 23798 27292 28999
rect 27448 27334 27476 29679
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27540 28762 27568 29106
rect 27528 28756 27580 28762
rect 27528 28698 27580 28704
rect 27632 28558 27660 29786
rect 27710 29608 27766 29617
rect 27710 29543 27766 29552
rect 27724 29170 27752 29543
rect 27816 29238 27844 29951
rect 27804 29232 27856 29238
rect 27804 29174 27856 29180
rect 27712 29164 27764 29170
rect 27712 29106 27764 29112
rect 27816 28966 27844 29174
rect 27804 28960 27856 28966
rect 27804 28902 27856 28908
rect 27712 28688 27764 28694
rect 27712 28630 27764 28636
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27436 27328 27488 27334
rect 27436 27270 27488 27276
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 26382 27476 26862
rect 27436 26376 27488 26382
rect 27436 26318 27488 26324
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27356 25362 27384 25638
rect 27344 25356 27396 25362
rect 27344 25298 27396 25304
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27252 23792 27304 23798
rect 27252 23734 27304 23740
rect 26976 23112 27028 23118
rect 27264 23089 27292 23734
rect 27356 23361 27384 24210
rect 27448 24154 27476 26318
rect 27620 25968 27672 25974
rect 27620 25910 27672 25916
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27540 24682 27568 25842
rect 27528 24676 27580 24682
rect 27528 24618 27580 24624
rect 27448 24126 27568 24154
rect 27342 23352 27398 23361
rect 27342 23287 27344 23296
rect 27396 23287 27398 23296
rect 27344 23258 27396 23264
rect 26976 23054 27028 23060
rect 27250 23080 27306 23089
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26896 22778 26924 22918
rect 26988 22778 27016 23054
rect 27160 23044 27212 23050
rect 27540 23050 27568 24126
rect 27250 23015 27306 23024
rect 27528 23044 27580 23050
rect 27160 22986 27212 22992
rect 27528 22986 27580 22992
rect 26884 22772 26936 22778
rect 26884 22714 26936 22720
rect 26976 22772 27028 22778
rect 26976 22714 27028 22720
rect 27068 22704 27120 22710
rect 27068 22646 27120 22652
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26882 22536 26938 22545
rect 26882 22471 26938 22480
rect 26896 22438 26924 22471
rect 26884 22432 26936 22438
rect 26884 22374 26936 22380
rect 26896 22098 26924 22374
rect 26884 22092 26936 22098
rect 26884 22034 26936 22040
rect 26884 21956 26936 21962
rect 26884 21898 26936 21904
rect 26792 21888 26844 21894
rect 26896 21865 26924 21898
rect 26792 21830 26844 21836
rect 26882 21856 26938 21865
rect 26804 17134 26832 21830
rect 26882 21791 26938 21800
rect 26882 21720 26938 21729
rect 26988 21706 27016 22578
rect 26938 21678 27016 21706
rect 26882 21655 26938 21664
rect 26896 20777 26924 21655
rect 26976 21344 27028 21350
rect 27080 21332 27108 22646
rect 27172 22574 27200 22986
rect 27540 22642 27568 22986
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27160 22568 27212 22574
rect 27160 22510 27212 22516
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 27172 22030 27200 22170
rect 27356 22166 27384 22578
rect 27528 22500 27580 22506
rect 27528 22442 27580 22448
rect 27344 22160 27396 22166
rect 27344 22102 27396 22108
rect 27160 22024 27212 22030
rect 27212 21984 27292 22012
rect 27160 21966 27212 21972
rect 27264 21486 27292 21984
rect 27356 21622 27384 22102
rect 27540 22012 27568 22442
rect 27632 22094 27660 25910
rect 27724 24138 27752 28630
rect 27804 28416 27856 28422
rect 27804 28358 27856 28364
rect 27816 28082 27844 28358
rect 27804 28076 27856 28082
rect 27804 28018 27856 28024
rect 27908 26586 27936 30058
rect 28000 29714 28028 30058
rect 27988 29708 28040 29714
rect 27988 29650 28040 29656
rect 27896 26580 27948 26586
rect 27896 26522 27948 26528
rect 27908 26382 27936 26522
rect 28092 26432 28120 30670
rect 28184 30569 28212 30738
rect 28170 30560 28226 30569
rect 28170 30495 28226 30504
rect 28184 30054 28212 30495
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28172 30048 28224 30054
rect 28172 29990 28224 29996
rect 28276 29850 28304 30126
rect 28264 29844 28316 29850
rect 28264 29786 28316 29792
rect 28172 29300 28224 29306
rect 28172 29242 28224 29248
rect 28184 28370 28212 29242
rect 28276 28490 28304 29786
rect 28368 29306 28396 31198
rect 28736 30410 28764 31282
rect 28816 31272 28868 31278
rect 28816 31214 28868 31220
rect 28828 30938 28856 31214
rect 28816 30932 28868 30938
rect 28816 30874 28868 30880
rect 28644 30394 28764 30410
rect 28632 30388 28764 30394
rect 28684 30382 28764 30388
rect 28632 30330 28684 30336
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28552 29578 28580 30194
rect 28632 30116 28684 30122
rect 28632 30058 28684 30064
rect 28540 29572 28592 29578
rect 28540 29514 28592 29520
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28448 29300 28500 29306
rect 28448 29242 28500 29248
rect 28368 29170 28396 29242
rect 28460 29170 28488 29242
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 28356 28484 28408 28490
rect 28356 28426 28408 28432
rect 28184 28342 28304 28370
rect 28172 27872 28224 27878
rect 28172 27814 28224 27820
rect 28184 27674 28212 27814
rect 28172 27668 28224 27674
rect 28172 27610 28224 27616
rect 28276 27577 28304 28342
rect 28368 28150 28396 28426
rect 28356 28144 28408 28150
rect 28356 28086 28408 28092
rect 28356 28008 28408 28014
rect 28460 27962 28488 29106
rect 28540 29028 28592 29034
rect 28540 28970 28592 28976
rect 28408 27956 28488 27962
rect 28356 27950 28488 27956
rect 28368 27934 28488 27950
rect 28262 27568 28318 27577
rect 28262 27503 28264 27512
rect 28316 27503 28318 27512
rect 28264 27474 28316 27480
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 28276 26489 28304 26930
rect 28262 26480 28318 26489
rect 28092 26404 28212 26432
rect 28262 26415 28318 26424
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 28080 26308 28132 26314
rect 28080 26250 28132 26256
rect 27988 26240 28040 26246
rect 27988 26182 28040 26188
rect 28000 25974 28028 26182
rect 27988 25968 28040 25974
rect 27988 25910 28040 25916
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27712 24132 27764 24138
rect 27712 24074 27764 24080
rect 27816 23662 27844 25230
rect 28092 24818 28120 26250
rect 28184 25770 28212 26404
rect 28368 26382 28396 27066
rect 28356 26376 28408 26382
rect 28356 26318 28408 26324
rect 28264 26308 28316 26314
rect 28264 26250 28316 26256
rect 28172 25764 28224 25770
rect 28172 25706 28224 25712
rect 28184 25498 28212 25706
rect 28172 25492 28224 25498
rect 28172 25434 28224 25440
rect 28276 24818 28304 26250
rect 28356 25152 28408 25158
rect 28356 25094 28408 25100
rect 28080 24812 28132 24818
rect 28000 24772 28080 24800
rect 27894 24712 27950 24721
rect 27894 24647 27950 24656
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 27908 22982 27936 24647
rect 28000 23526 28028 24772
rect 28080 24754 28132 24760
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 28184 24206 28212 24686
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28080 24064 28132 24070
rect 28080 24006 28132 24012
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 28092 23730 28120 24006
rect 28184 23866 28212 24006
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28080 23724 28132 23730
rect 28080 23666 28132 23672
rect 28172 23724 28224 23730
rect 28172 23666 28224 23672
rect 28092 23633 28120 23666
rect 28078 23624 28134 23633
rect 28078 23559 28134 23568
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 27896 22976 27948 22982
rect 27896 22918 27948 22924
rect 28184 22817 28212 23666
rect 28170 22808 28226 22817
rect 28170 22743 28226 22752
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 27632 22066 27752 22094
rect 27620 22024 27672 22030
rect 27540 21984 27620 22012
rect 27620 21966 27672 21972
rect 27344 21616 27396 21622
rect 27344 21558 27396 21564
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 27436 21480 27488 21486
rect 27436 21422 27488 21428
rect 27028 21304 27108 21332
rect 26976 21286 27028 21292
rect 26988 21146 27016 21286
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 26882 20768 26938 20777
rect 26882 20703 26938 20712
rect 26884 20528 26936 20534
rect 26884 20470 26936 20476
rect 26896 19854 26924 20470
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 26884 19848 26936 19854
rect 26882 19816 26884 19825
rect 26936 19816 26938 19825
rect 26882 19751 26938 19760
rect 26884 19372 26936 19378
rect 26884 19314 26936 19320
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 26620 16204 26740 16232
rect 26620 16114 26648 16204
rect 26804 16114 26832 17070
rect 26608 16108 26660 16114
rect 26608 16050 26660 16056
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 26792 16108 26844 16114
rect 26792 16050 26844 16056
rect 26608 15360 26660 15366
rect 26606 15328 26608 15337
rect 26660 15328 26662 15337
rect 26606 15263 26662 15272
rect 26606 14920 26662 14929
rect 26606 14855 26662 14864
rect 26514 14376 26570 14385
rect 26514 14311 26570 14320
rect 26620 14249 26648 14855
rect 26606 14240 26662 14249
rect 26606 14175 26662 14184
rect 26620 14074 26648 14175
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26620 13326 26648 13806
rect 26712 13530 26740 16050
rect 26792 15496 26844 15502
rect 26792 15438 26844 15444
rect 26804 14822 26832 15438
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26896 14532 26924 19314
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 26976 18760 27028 18766
rect 26974 18728 26976 18737
rect 27028 18728 27030 18737
rect 26974 18663 27030 18672
rect 27066 17912 27122 17921
rect 27066 17847 27122 17856
rect 27080 17746 27108 17847
rect 27068 17740 27120 17746
rect 27068 17682 27120 17688
rect 27080 17338 27108 17682
rect 27068 17332 27120 17338
rect 27068 17274 27120 17280
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26988 15337 27016 17138
rect 27172 15502 27200 19110
rect 27264 18698 27292 19246
rect 27252 18692 27304 18698
rect 27252 18634 27304 18640
rect 27160 15496 27212 15502
rect 27080 15456 27160 15484
rect 26974 15328 27030 15337
rect 26974 15263 27030 15272
rect 26976 15156 27028 15162
rect 26976 15098 27028 15104
rect 26804 14504 26924 14532
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 26252 12102 26280 12922
rect 26620 12918 26648 13262
rect 26712 12986 26740 13466
rect 26804 13190 26832 14504
rect 26988 14464 27016 15098
rect 26896 14436 27016 14464
rect 26896 13326 26924 14436
rect 26974 14376 27030 14385
rect 26974 14311 26976 14320
rect 27028 14311 27030 14320
rect 26976 14282 27028 14288
rect 26974 14104 27030 14113
rect 26974 14039 26976 14048
rect 27028 14039 27030 14048
rect 26976 14010 27028 14016
rect 26976 13796 27028 13802
rect 26976 13738 27028 13744
rect 26988 13326 27016 13738
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26608 12912 26660 12918
rect 26608 12854 26660 12860
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26332 12164 26384 12170
rect 26332 12106 26384 12112
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 26148 11756 26200 11762
rect 26148 11698 26200 11704
rect 26160 10674 26188 11698
rect 26252 10985 26280 12038
rect 26238 10976 26294 10985
rect 26238 10911 26294 10920
rect 26252 10674 26280 10911
rect 26148 10668 26200 10674
rect 26148 10610 26200 10616
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26344 10554 26372 12106
rect 26528 11830 26556 12242
rect 26620 12238 26648 12854
rect 26700 12844 26752 12850
rect 26700 12786 26752 12792
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26712 12084 26740 12786
rect 26804 12782 26832 13126
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26896 12714 26924 13262
rect 26884 12708 26936 12714
rect 26884 12650 26936 12656
rect 26790 12336 26846 12345
rect 26790 12271 26846 12280
rect 26884 12300 26936 12306
rect 26804 12238 26832 12271
rect 26884 12242 26936 12248
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26620 12056 26740 12084
rect 26516 11824 26568 11830
rect 26516 11766 26568 11772
rect 26422 10704 26478 10713
rect 26422 10639 26424 10648
rect 26476 10639 26478 10648
rect 26424 10610 26476 10616
rect 26252 10538 26372 10554
rect 26240 10532 26372 10538
rect 26292 10526 26372 10532
rect 26240 10474 26292 10480
rect 26252 10130 26280 10474
rect 26436 10305 26464 10610
rect 26422 10296 26478 10305
rect 26422 10231 26478 10240
rect 26422 10160 26478 10169
rect 26240 10124 26292 10130
rect 26422 10095 26424 10104
rect 26240 10066 26292 10072
rect 26476 10095 26478 10104
rect 26424 10066 26476 10072
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 26068 9586 26096 9930
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25872 9444 25924 9450
rect 25872 9386 25924 9392
rect 26332 9444 26384 9450
rect 26332 9386 26384 9392
rect 25884 8498 25912 9386
rect 26344 9353 26372 9386
rect 26330 9344 26386 9353
rect 26330 9279 26386 9288
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25976 8537 26004 9114
rect 26240 9104 26292 9110
rect 26240 9046 26292 9052
rect 26252 8974 26280 9046
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 25962 8528 26018 8537
rect 25872 8492 25924 8498
rect 25962 8463 26018 8472
rect 25872 8434 25924 8440
rect 26252 8430 26280 8910
rect 26240 8424 26292 8430
rect 26240 8366 26292 8372
rect 26252 8022 26280 8366
rect 26240 8016 26292 8022
rect 26240 7958 26292 7964
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 26068 7342 26096 7686
rect 26252 7342 26280 7958
rect 26436 7546 26464 10066
rect 26516 9988 26568 9994
rect 26620 9976 26648 12056
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26712 10577 26740 10610
rect 26698 10568 26754 10577
rect 26698 10503 26754 10512
rect 26700 10124 26752 10130
rect 26700 10066 26752 10072
rect 26568 9948 26648 9976
rect 26516 9930 26568 9936
rect 26712 9586 26740 10066
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26804 9110 26832 11834
rect 26896 11234 26924 12242
rect 26988 11898 27016 13262
rect 27080 12850 27108 15456
rect 27160 15438 27212 15444
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 27172 13841 27200 15302
rect 27158 13832 27214 13841
rect 27158 13767 27214 13776
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 27172 13258 27200 13670
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 27264 12918 27292 18634
rect 27356 17513 27384 20402
rect 27448 20398 27476 21422
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27448 19514 27476 20334
rect 27620 20256 27672 20262
rect 27620 20198 27672 20204
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27436 19508 27488 19514
rect 27436 19450 27488 19456
rect 27540 19174 27568 19790
rect 27632 19174 27660 20198
rect 27724 19922 27752 22066
rect 28092 21622 28120 22374
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 28080 21616 28132 21622
rect 28080 21558 28132 21564
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 27908 20602 27936 20878
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 27896 20596 27948 20602
rect 27896 20538 27948 20544
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27908 20369 27936 20402
rect 27894 20360 27950 20369
rect 27894 20295 27950 20304
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27528 19168 27580 19174
rect 27528 19110 27580 19116
rect 27620 19168 27672 19174
rect 27620 19110 27672 19116
rect 27632 18970 27660 19110
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27342 17504 27398 17513
rect 27342 17439 27398 17448
rect 27724 17270 27752 19450
rect 27816 18290 27844 20198
rect 28000 19378 28028 20742
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27804 18284 27856 18290
rect 27804 18226 27856 18232
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 27712 17264 27764 17270
rect 27434 17232 27490 17241
rect 27712 17206 27764 17212
rect 27434 17167 27490 17176
rect 27528 17196 27580 17202
rect 27448 16522 27476 17167
rect 27528 17138 27580 17144
rect 27436 16516 27488 16522
rect 27436 16458 27488 16464
rect 27436 15496 27488 15502
rect 27436 15438 27488 15444
rect 27448 15162 27476 15438
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 27344 15020 27396 15026
rect 27344 14962 27396 14968
rect 27356 14414 27384 14962
rect 27448 14550 27476 15098
rect 27540 15026 27568 17138
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27632 16250 27660 16526
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27620 16040 27672 16046
rect 27724 16028 27752 16934
rect 27816 16590 27844 18090
rect 27908 16590 27936 19246
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27804 16584 27856 16590
rect 27804 16526 27856 16532
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27672 16000 27752 16028
rect 27620 15982 27672 15988
rect 27618 15736 27674 15745
rect 27618 15671 27674 15680
rect 27632 15162 27660 15671
rect 27724 15366 27752 16000
rect 27712 15360 27764 15366
rect 27712 15302 27764 15308
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27816 15094 27844 16526
rect 27908 16250 27936 16526
rect 27896 16244 27948 16250
rect 27896 16186 27948 16192
rect 27896 16108 27948 16114
rect 27896 16050 27948 16056
rect 27908 15706 27936 16050
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 28000 15450 28028 18226
rect 28092 16674 28120 21558
rect 28184 21554 28212 21830
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 28170 21448 28226 21457
rect 28170 21383 28226 21392
rect 28184 19310 28212 21383
rect 28276 20534 28304 24754
rect 28368 24614 28396 25094
rect 28446 24848 28502 24857
rect 28552 24818 28580 28970
rect 28644 27538 28672 30058
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28736 29646 28764 29990
rect 28724 29640 28776 29646
rect 28828 29628 28856 30874
rect 28920 30258 28948 32438
rect 29092 32360 29144 32366
rect 29092 32302 29144 32308
rect 29000 32224 29052 32230
rect 29000 32166 29052 32172
rect 29012 32026 29040 32166
rect 29000 32020 29052 32026
rect 29000 31962 29052 31968
rect 29104 31482 29132 32302
rect 29736 31884 29788 31890
rect 29736 31826 29788 31832
rect 29552 31816 29604 31822
rect 29550 31784 29552 31793
rect 29604 31784 29606 31793
rect 29606 31728 29684 31754
rect 29550 31726 29684 31728
rect 29550 31719 29606 31726
rect 29092 31476 29144 31482
rect 29092 31418 29144 31424
rect 29184 31340 29236 31346
rect 29184 31282 29236 31288
rect 29092 31204 29144 31210
rect 29092 31146 29144 31152
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 29000 30184 29052 30190
rect 28906 30152 28962 30161
rect 29000 30126 29052 30132
rect 28906 30087 28908 30096
rect 28960 30087 28962 30096
rect 28908 30058 28960 30064
rect 29012 29714 29040 30126
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 28908 29640 28960 29646
rect 28828 29600 28908 29628
rect 28724 29582 28776 29588
rect 28908 29582 28960 29588
rect 28632 27532 28684 27538
rect 28632 27474 28684 27480
rect 28644 25362 28672 27474
rect 28736 26024 28764 29582
rect 28816 29504 28868 29510
rect 28816 29446 28868 29452
rect 28828 29170 28856 29446
rect 28920 29306 28948 29582
rect 29000 29572 29052 29578
rect 29000 29514 29052 29520
rect 28908 29300 28960 29306
rect 28908 29242 28960 29248
rect 28906 29200 28962 29209
rect 28816 29164 28868 29170
rect 28906 29135 28908 29144
rect 28816 29106 28868 29112
rect 28960 29135 28962 29144
rect 28908 29106 28960 29112
rect 28816 28960 28868 28966
rect 28816 28902 28868 28908
rect 28828 28762 28856 28902
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28908 28756 28960 28762
rect 28908 28698 28960 28704
rect 28920 28642 28948 28698
rect 28828 28614 28948 28642
rect 28828 28422 28856 28614
rect 28816 28416 28868 28422
rect 28816 28358 28868 28364
rect 28828 28218 28856 28358
rect 28816 28212 28868 28218
rect 28816 28154 28868 28160
rect 29012 28150 29040 29514
rect 29104 28218 29132 31146
rect 29196 30394 29224 31282
rect 29460 31272 29512 31278
rect 29460 31214 29512 31220
rect 29276 30864 29328 30870
rect 29276 30806 29328 30812
rect 29288 30394 29316 30806
rect 29472 30666 29500 31214
rect 29656 30666 29684 31726
rect 29748 31414 29776 31826
rect 29736 31408 29788 31414
rect 29736 31350 29788 31356
rect 29828 31272 29880 31278
rect 29828 31214 29880 31220
rect 29460 30660 29512 30666
rect 29460 30602 29512 30608
rect 29644 30660 29696 30666
rect 29644 30602 29696 30608
rect 29184 30388 29236 30394
rect 29184 30330 29236 30336
rect 29276 30388 29328 30394
rect 29276 30330 29328 30336
rect 29736 30320 29788 30326
rect 29458 30288 29514 30297
rect 29736 30262 29788 30268
rect 29458 30223 29514 30232
rect 29368 30184 29420 30190
rect 29368 30126 29420 30132
rect 29380 29850 29408 30126
rect 29276 29844 29328 29850
rect 29276 29786 29328 29792
rect 29368 29844 29420 29850
rect 29368 29786 29420 29792
rect 29288 29578 29316 29786
rect 29276 29572 29328 29578
rect 29276 29514 29328 29520
rect 29184 29096 29236 29102
rect 29184 29038 29236 29044
rect 29368 29096 29420 29102
rect 29368 29038 29420 29044
rect 29196 28558 29224 29038
rect 29276 28960 29328 28966
rect 29276 28902 29328 28908
rect 29184 28552 29236 28558
rect 29184 28494 29236 28500
rect 29196 28422 29224 28494
rect 29184 28416 29236 28422
rect 29184 28358 29236 28364
rect 29182 28248 29238 28257
rect 29092 28212 29144 28218
rect 29182 28183 29238 28192
rect 29092 28154 29144 28160
rect 29000 28144 29052 28150
rect 29000 28086 29052 28092
rect 29196 28082 29224 28183
rect 29288 28082 29316 28902
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 28920 27130 28948 28018
rect 29092 27872 29144 27878
rect 29092 27814 29144 27820
rect 28998 27432 29054 27441
rect 28998 27367 29000 27376
rect 29052 27367 29054 27376
rect 29000 27338 29052 27344
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 29000 27124 29052 27130
rect 29000 27066 29052 27072
rect 29012 26994 29040 27066
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 29000 26852 29052 26858
rect 29000 26794 29052 26800
rect 28908 26240 28960 26246
rect 28908 26182 28960 26188
rect 28736 25996 28856 26024
rect 28724 25900 28776 25906
rect 28724 25842 28776 25848
rect 28632 25356 28684 25362
rect 28632 25298 28684 25304
rect 28632 25152 28684 25158
rect 28632 25094 28684 25100
rect 28446 24783 28502 24792
rect 28540 24812 28592 24818
rect 28356 24608 28408 24614
rect 28356 24550 28408 24556
rect 28356 24404 28408 24410
rect 28356 24346 28408 24352
rect 28368 24313 28396 24346
rect 28354 24304 28410 24313
rect 28354 24239 28410 24248
rect 28356 24200 28408 24206
rect 28354 24168 28356 24177
rect 28408 24168 28410 24177
rect 28354 24103 28410 24112
rect 28460 23526 28488 24783
rect 28540 24754 28592 24760
rect 28552 23866 28580 24754
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 28540 23724 28592 23730
rect 28540 23666 28592 23672
rect 28552 23526 28580 23666
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28540 23520 28592 23526
rect 28540 23462 28592 23468
rect 28356 23248 28408 23254
rect 28356 23190 28408 23196
rect 28368 22710 28396 23190
rect 28460 23118 28488 23462
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 28552 23050 28580 23258
rect 28540 23044 28592 23050
rect 28540 22986 28592 22992
rect 28446 22808 28502 22817
rect 28446 22743 28502 22752
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28368 21894 28396 22646
rect 28460 22488 28488 22743
rect 28540 22500 28592 22506
rect 28460 22460 28540 22488
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28368 21332 28396 21830
rect 28460 21457 28488 22460
rect 28540 22442 28592 22448
rect 28644 22094 28672 25094
rect 28736 24886 28764 25842
rect 28828 24954 28856 25996
rect 28920 25673 28948 26182
rect 29012 25838 29040 26794
rect 29000 25832 29052 25838
rect 29000 25774 29052 25780
rect 28906 25664 28962 25673
rect 28906 25599 28962 25608
rect 28908 25424 28960 25430
rect 28908 25366 28960 25372
rect 28816 24948 28868 24954
rect 28816 24890 28868 24896
rect 28724 24880 28776 24886
rect 28724 24822 28776 24828
rect 28736 24206 28764 24822
rect 28724 24200 28776 24206
rect 28828 24177 28856 24890
rect 28724 24142 28776 24148
rect 28814 24168 28870 24177
rect 28814 24103 28870 24112
rect 28724 24064 28776 24070
rect 28722 24032 28724 24041
rect 28776 24032 28778 24041
rect 28722 23967 28778 23976
rect 28828 23712 28856 24103
rect 28828 23684 28865 23712
rect 28837 23594 28865 23684
rect 28816 23588 28868 23594
rect 28816 23530 28868 23536
rect 28816 23180 28868 23186
rect 28816 23122 28868 23128
rect 28552 22066 28672 22094
rect 28446 21448 28502 21457
rect 28446 21383 28502 21392
rect 28368 21304 28514 21332
rect 28354 21176 28410 21185
rect 28486 21162 28514 21304
rect 28354 21111 28410 21120
rect 28460 21134 28514 21162
rect 28368 20942 28396 21111
rect 28460 21010 28488 21134
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28264 20528 28316 20534
rect 28264 20470 28316 20476
rect 28276 19990 28304 20470
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28368 19836 28396 20878
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28460 20262 28488 20810
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28276 19808 28396 19836
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 28276 18358 28304 19808
rect 28354 19408 28410 19417
rect 28552 19394 28580 22066
rect 28724 22024 28776 22030
rect 28724 21966 28776 21972
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 28644 21457 28672 21626
rect 28630 21448 28686 21457
rect 28630 21383 28686 21392
rect 28736 21185 28764 21966
rect 28722 21176 28778 21185
rect 28722 21111 28724 21120
rect 28776 21111 28778 21120
rect 28724 21082 28776 21088
rect 28724 20936 28776 20942
rect 28724 20878 28776 20884
rect 28736 20602 28764 20878
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28724 20460 28776 20466
rect 28828 20448 28856 23122
rect 28920 22438 28948 25366
rect 29012 25362 29040 25774
rect 29000 25356 29052 25362
rect 29000 25298 29052 25304
rect 29000 25220 29052 25226
rect 29000 25162 29052 25168
rect 29012 24562 29040 25162
rect 29104 24818 29132 27814
rect 29196 26217 29224 28018
rect 29276 27328 29328 27334
rect 29276 27270 29328 27276
rect 29288 27169 29316 27270
rect 29274 27160 29330 27169
rect 29380 27130 29408 29038
rect 29472 29034 29500 30223
rect 29748 29170 29776 30262
rect 29840 29850 29868 31214
rect 29932 30938 29960 32846
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 30024 31686 30052 32710
rect 30208 32502 30236 32914
rect 30840 32836 30892 32842
rect 30840 32778 30892 32784
rect 30656 32768 30708 32774
rect 30656 32710 30708 32716
rect 30196 32496 30248 32502
rect 30196 32438 30248 32444
rect 30208 31890 30236 32438
rect 30668 32434 30696 32710
rect 30656 32428 30708 32434
rect 30656 32370 30708 32376
rect 30564 32292 30616 32298
rect 30564 32234 30616 32240
rect 30196 31884 30248 31890
rect 30196 31826 30248 31832
rect 30208 31754 30236 31826
rect 30208 31726 30328 31754
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 30104 31680 30156 31686
rect 30104 31622 30156 31628
rect 29920 30932 29972 30938
rect 29920 30874 29972 30880
rect 30024 30734 30052 31622
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 29920 30388 29972 30394
rect 29920 30330 29972 30336
rect 29828 29844 29880 29850
rect 29828 29786 29880 29792
rect 29552 29164 29604 29170
rect 29736 29164 29788 29170
rect 29552 29106 29604 29112
rect 29656 29124 29736 29152
rect 29460 29028 29512 29034
rect 29460 28970 29512 28976
rect 29564 28966 29592 29106
rect 29552 28960 29604 28966
rect 29552 28902 29604 28908
rect 29460 27940 29512 27946
rect 29460 27882 29512 27888
rect 29472 27577 29500 27882
rect 29552 27668 29604 27674
rect 29552 27610 29604 27616
rect 29458 27568 29514 27577
rect 29458 27503 29514 27512
rect 29460 27328 29512 27334
rect 29460 27270 29512 27276
rect 29274 27095 29330 27104
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 29472 27010 29500 27270
rect 29288 26994 29500 27010
rect 29288 26988 29512 26994
rect 29288 26982 29460 26988
rect 29182 26208 29238 26217
rect 29182 26143 29238 26152
rect 29288 25974 29316 26982
rect 29460 26930 29512 26936
rect 29564 26926 29592 27610
rect 29656 27169 29684 29124
rect 29736 29106 29788 29112
rect 29826 29064 29882 29073
rect 29932 29050 29960 30330
rect 30012 29708 30064 29714
rect 30012 29650 30064 29656
rect 29882 29022 29960 29050
rect 29826 28999 29882 29008
rect 29736 28416 29788 28422
rect 29736 28358 29788 28364
rect 29748 27402 29776 28358
rect 29840 27674 29868 28999
rect 30024 28994 30052 29650
rect 29932 28966 30052 28994
rect 29932 28150 29960 28966
rect 30010 28248 30066 28257
rect 30010 28183 30066 28192
rect 30024 28150 30052 28183
rect 29920 28144 29972 28150
rect 29920 28086 29972 28092
rect 30012 28144 30064 28150
rect 30116 28121 30144 31622
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30208 29866 30236 31078
rect 30300 30258 30328 31726
rect 30576 31686 30604 32234
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30656 31952 30708 31958
rect 30656 31894 30708 31900
rect 30564 31680 30616 31686
rect 30564 31622 30616 31628
rect 30668 30734 30696 31894
rect 30656 30728 30708 30734
rect 30656 30670 30708 30676
rect 30760 30326 30788 31962
rect 30852 31482 30880 32778
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 30932 32564 30984 32570
rect 30932 32506 30984 32512
rect 33324 32564 33376 32570
rect 33324 32506 33376 32512
rect 30944 31822 30972 32506
rect 31116 32428 31168 32434
rect 31116 32370 31168 32376
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 31484 32428 31536 32434
rect 31484 32370 31536 32376
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 31128 31686 31156 32370
rect 31312 32230 31340 32370
rect 31300 32224 31352 32230
rect 31300 32166 31352 32172
rect 31206 31920 31262 31929
rect 31206 31855 31262 31864
rect 31116 31680 31168 31686
rect 31116 31622 31168 31628
rect 30840 31476 30892 31482
rect 30840 31418 30892 31424
rect 30852 31362 30880 31418
rect 30852 31334 30972 31362
rect 30840 31272 30892 31278
rect 30840 31214 30892 31220
rect 30852 30802 30880 31214
rect 30944 30938 30972 31334
rect 31128 31210 31156 31622
rect 31116 31204 31168 31210
rect 31116 31146 31168 31152
rect 30932 30932 30984 30938
rect 30932 30874 30984 30880
rect 31024 30864 31076 30870
rect 31024 30806 31076 30812
rect 30840 30796 30892 30802
rect 30840 30738 30892 30744
rect 30748 30320 30800 30326
rect 30748 30262 30800 30268
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 30286 29880 30342 29889
rect 30208 29838 30286 29866
rect 30286 29815 30342 29824
rect 30196 29640 30248 29646
rect 30196 29582 30248 29588
rect 30208 29345 30236 29582
rect 30300 29510 30328 29815
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30378 29608 30434 29617
rect 30378 29543 30434 29552
rect 30288 29504 30340 29510
rect 30288 29446 30340 29452
rect 30194 29336 30250 29345
rect 30194 29271 30196 29280
rect 30248 29271 30250 29280
rect 30196 29242 30248 29248
rect 30392 29170 30420 29543
rect 30196 29164 30248 29170
rect 30196 29106 30248 29112
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30012 28086 30064 28092
rect 30102 28112 30158 28121
rect 29932 27849 29960 28086
rect 30102 28047 30158 28056
rect 30104 28008 30156 28014
rect 30010 27976 30066 27985
rect 30104 27950 30156 27956
rect 30010 27911 30066 27920
rect 29918 27840 29974 27849
rect 29918 27775 29974 27784
rect 29828 27668 29880 27674
rect 29828 27610 29880 27616
rect 29918 27432 29974 27441
rect 29736 27396 29788 27402
rect 29788 27356 29868 27384
rect 29918 27367 29920 27376
rect 29736 27338 29788 27344
rect 29642 27160 29698 27169
rect 29840 27146 29868 27356
rect 29972 27367 29974 27376
rect 29920 27338 29972 27344
rect 29840 27118 29960 27146
rect 29642 27095 29698 27104
rect 29552 26920 29604 26926
rect 29552 26862 29604 26868
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29472 25974 29500 26522
rect 29276 25968 29328 25974
rect 29276 25910 29328 25916
rect 29460 25968 29512 25974
rect 29460 25910 29512 25916
rect 29460 25764 29512 25770
rect 29460 25706 29512 25712
rect 29552 25764 29604 25770
rect 29552 25706 29604 25712
rect 29276 25696 29328 25702
rect 29276 25638 29328 25644
rect 29288 24993 29316 25638
rect 29274 24984 29330 24993
rect 29274 24919 29330 24928
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29184 24812 29236 24818
rect 29184 24754 29236 24760
rect 29012 24534 29132 24562
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 29012 21978 29040 24346
rect 29104 23798 29132 24534
rect 29196 24410 29224 24754
rect 29276 24608 29328 24614
rect 29276 24550 29328 24556
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 29288 24206 29316 24550
rect 29276 24200 29328 24206
rect 29276 24142 29328 24148
rect 29092 23792 29144 23798
rect 29092 23734 29144 23740
rect 29104 23322 29132 23734
rect 29092 23316 29144 23322
rect 29092 23258 29144 23264
rect 29184 23044 29236 23050
rect 29184 22986 29236 22992
rect 29092 22976 29144 22982
rect 29092 22918 29144 22924
rect 28920 21950 29040 21978
rect 28920 20788 28948 21950
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 29012 21554 29040 21830
rect 29000 21548 29052 21554
rect 29000 21490 29052 21496
rect 29012 20942 29040 21490
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28920 20760 29040 20788
rect 28828 20420 28948 20448
rect 28724 20402 28776 20408
rect 28632 20392 28684 20398
rect 28632 20334 28684 20340
rect 28410 19366 28580 19394
rect 28354 19343 28356 19352
rect 28408 19343 28410 19352
rect 28356 19314 28408 19320
rect 28540 19236 28592 19242
rect 28540 19178 28592 19184
rect 28264 18352 28316 18358
rect 28264 18294 28316 18300
rect 28276 18086 28304 18294
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28092 16646 28212 16674
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 28092 16182 28120 16526
rect 28080 16176 28132 16182
rect 28080 16118 28132 16124
rect 28000 15422 28120 15450
rect 27986 15328 28042 15337
rect 27986 15263 28042 15272
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27436 14544 27488 14550
rect 27436 14486 27488 14492
rect 27344 14408 27396 14414
rect 27396 14368 27476 14396
rect 27344 14350 27396 14356
rect 27448 14006 27476 14368
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27344 13456 27396 13462
rect 27344 13398 27396 13404
rect 27356 12918 27384 13398
rect 27252 12912 27304 12918
rect 27252 12854 27304 12860
rect 27344 12912 27396 12918
rect 27344 12854 27396 12860
rect 27448 12850 27476 13942
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 27080 11778 27108 12786
rect 27160 12776 27212 12782
rect 27160 12718 27212 12724
rect 27172 12238 27200 12718
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27344 12232 27396 12238
rect 27344 12174 27396 12180
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27172 11937 27200 12038
rect 27158 11928 27214 11937
rect 27158 11863 27214 11872
rect 27080 11750 27292 11778
rect 27356 11762 27384 12174
rect 27264 11694 27292 11750
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27068 11688 27120 11694
rect 27160 11688 27212 11694
rect 27068 11630 27120 11636
rect 27158 11656 27160 11665
rect 27252 11688 27304 11694
rect 27212 11656 27214 11665
rect 26896 11206 27016 11234
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26792 9104 26844 9110
rect 26792 9046 26844 9052
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26528 8294 26556 8842
rect 26712 8430 26740 8978
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26700 8424 26752 8430
rect 26700 8366 26752 8372
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 26528 8022 26556 8230
rect 26516 8016 26568 8022
rect 26568 7964 26648 7970
rect 26516 7958 26648 7964
rect 26528 7942 26648 7958
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 25780 7336 25832 7342
rect 25780 7278 25832 7284
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 25872 6996 25924 7002
rect 25872 6938 25924 6944
rect 25778 6352 25834 6361
rect 25884 6322 25912 6938
rect 26068 6866 26096 7278
rect 26252 6984 26280 7278
rect 26424 7200 26476 7206
rect 26424 7142 26476 7148
rect 26332 6996 26384 7002
rect 26252 6956 26332 6984
rect 26332 6938 26384 6944
rect 26344 6866 26372 6938
rect 26056 6860 26108 6866
rect 26056 6802 26108 6808
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 26436 6798 26464 7142
rect 26528 6798 26556 7346
rect 26620 7206 26648 7942
rect 26712 7750 26740 8366
rect 26804 8090 26832 8434
rect 26792 8084 26844 8090
rect 26792 8026 26844 8032
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26712 7256 26740 7686
rect 26804 7410 26832 8026
rect 26792 7404 26844 7410
rect 26792 7346 26844 7352
rect 26792 7268 26844 7274
rect 26712 7228 26792 7256
rect 26792 7210 26844 7216
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 26804 6798 26832 7210
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 26516 6792 26568 6798
rect 26516 6734 26568 6740
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 25778 6287 25780 6296
rect 25832 6287 25834 6296
rect 25872 6316 25924 6322
rect 25780 6258 25832 6264
rect 25872 6258 25924 6264
rect 26528 6118 26556 6734
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 26620 6458 26648 6598
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26700 6384 26752 6390
rect 26700 6326 26752 6332
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 25700 5710 25728 6054
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25320 5568 25372 5574
rect 25320 5510 25372 5516
rect 25136 5296 25188 5302
rect 25136 5238 25188 5244
rect 25148 4536 25176 5238
rect 25332 4690 25360 5510
rect 26424 5364 26476 5370
rect 26424 5306 26476 5312
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25228 4548 25280 4554
rect 25148 4508 25228 4536
rect 25148 3466 25176 4508
rect 25228 4490 25280 4496
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26344 3738 26372 4014
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 25136 3460 25188 3466
rect 25136 3402 25188 3408
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26252 3126 26280 3334
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 26436 3058 26464 5306
rect 26712 4826 26740 6326
rect 26804 6254 26832 6734
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26896 5370 26924 11086
rect 26988 10441 27016 11206
rect 27080 10674 27108 11630
rect 27252 11630 27304 11636
rect 27158 11591 27214 11600
rect 27172 11354 27200 11591
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27264 10742 27292 11630
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27252 10736 27304 10742
rect 27252 10678 27304 10684
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 26974 10432 27030 10441
rect 26974 10367 27030 10376
rect 26988 9654 27016 10367
rect 27080 9926 27108 10610
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 27068 9920 27120 9926
rect 27172 9897 27200 10406
rect 27068 9862 27120 9868
rect 27158 9888 27214 9897
rect 26976 9648 27028 9654
rect 26976 9590 27028 9596
rect 26976 9104 27028 9110
rect 26976 9046 27028 9052
rect 26988 8498 27016 9046
rect 26976 8492 27028 8498
rect 26976 8434 27028 8440
rect 27080 8090 27108 9862
rect 27158 9823 27214 9832
rect 27158 9616 27214 9625
rect 27158 9551 27160 9560
rect 27212 9551 27214 9560
rect 27160 9522 27212 9528
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 27066 6624 27122 6633
rect 27172 6610 27200 9522
rect 27264 8634 27292 10678
rect 27356 10606 27384 10746
rect 27448 10674 27476 12786
rect 27540 11694 27568 14962
rect 27618 14648 27674 14657
rect 27618 14583 27620 14592
rect 27672 14583 27674 14592
rect 27620 14554 27672 14560
rect 27816 14414 27844 15030
rect 28000 14414 28028 15263
rect 27804 14408 27856 14414
rect 27804 14350 27856 14356
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27618 13968 27674 13977
rect 27618 13903 27620 13912
rect 27672 13903 27674 13912
rect 27620 13874 27672 13880
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27632 12889 27660 13126
rect 27618 12880 27674 12889
rect 27618 12815 27674 12824
rect 27620 12776 27672 12782
rect 27620 12718 27672 12724
rect 27632 12306 27660 12718
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27618 12200 27674 12209
rect 27618 12135 27620 12144
rect 27672 12135 27674 12144
rect 27620 12106 27672 12112
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27356 10470 27384 10542
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27252 8628 27304 8634
rect 27252 8570 27304 8576
rect 27252 6928 27304 6934
rect 27356 6916 27384 9998
rect 27448 9518 27476 10610
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27448 7410 27476 7686
rect 27436 7404 27488 7410
rect 27436 7346 27488 7352
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 27304 6888 27384 6916
rect 27252 6870 27304 6876
rect 27448 6882 27476 7142
rect 27540 7002 27568 11630
rect 27620 11620 27672 11626
rect 27620 11562 27672 11568
rect 27632 8265 27660 11562
rect 27724 9450 27752 14214
rect 27816 11694 27844 14350
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27908 12850 27936 14282
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 28000 13977 28028 14010
rect 27986 13968 28042 13977
rect 27986 13903 28042 13912
rect 27988 13864 28040 13870
rect 27986 13832 27988 13841
rect 28040 13832 28042 13841
rect 27986 13767 28042 13776
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 27896 12844 27948 12850
rect 27896 12786 27948 12792
rect 27908 12753 27936 12786
rect 27894 12744 27950 12753
rect 27894 12679 27950 12688
rect 28000 12102 28028 13670
rect 28092 13394 28120 15422
rect 28184 14550 28212 16646
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28368 15910 28396 16594
rect 28448 16108 28500 16114
rect 28448 16050 28500 16056
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28264 15360 28316 15366
rect 28264 15302 28316 15308
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 28184 13938 28212 14350
rect 28276 13938 28304 15302
rect 28368 15026 28396 15302
rect 28356 15020 28408 15026
rect 28356 14962 28408 14968
rect 28172 13932 28224 13938
rect 28172 13874 28224 13880
rect 28264 13932 28316 13938
rect 28264 13874 28316 13880
rect 28356 13932 28408 13938
rect 28356 13874 28408 13880
rect 28184 13530 28212 13874
rect 28276 13734 28304 13874
rect 28264 13728 28316 13734
rect 28264 13670 28316 13676
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 28092 13002 28120 13330
rect 28092 12974 28212 13002
rect 28184 12918 28212 12974
rect 28172 12912 28224 12918
rect 28172 12854 28224 12860
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 28092 12714 28120 12786
rect 28184 12730 28212 12854
rect 28368 12832 28396 13874
rect 28460 13326 28488 16050
rect 28552 14822 28580 19178
rect 28644 16114 28672 20334
rect 28736 19718 28764 20402
rect 28816 20324 28868 20330
rect 28816 20266 28868 20272
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28736 19378 28764 19654
rect 28724 19372 28776 19378
rect 28724 19314 28776 19320
rect 28724 18896 28776 18902
rect 28722 18864 28724 18873
rect 28776 18864 28778 18873
rect 28722 18799 28778 18808
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28828 15858 28856 20266
rect 28920 16658 28948 20420
rect 29012 16998 29040 20760
rect 29104 20466 29132 22918
rect 29196 21554 29224 22986
rect 29366 22672 29422 22681
rect 29366 22607 29368 22616
rect 29420 22607 29422 22616
rect 29368 22578 29420 22584
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 29000 16992 29052 16998
rect 29000 16934 29052 16940
rect 28908 16652 28960 16658
rect 28908 16594 28960 16600
rect 28644 15830 28856 15858
rect 28644 15502 28672 15830
rect 29104 15688 29132 20266
rect 29196 20262 29224 21014
rect 29184 20256 29236 20262
rect 29184 20198 29236 20204
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 29196 18766 29224 19246
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 29196 17542 29224 18158
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29196 16998 29224 17478
rect 29288 17218 29316 22510
rect 29380 22234 29408 22578
rect 29368 22228 29420 22234
rect 29368 22170 29420 22176
rect 29368 21956 29420 21962
rect 29368 21898 29420 21904
rect 29380 21865 29408 21898
rect 29366 21856 29422 21865
rect 29366 21791 29422 21800
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29380 18902 29408 20742
rect 29368 18896 29420 18902
rect 29368 18838 29420 18844
rect 29368 18420 29420 18426
rect 29368 18362 29420 18368
rect 29380 17338 29408 18362
rect 29472 18154 29500 25706
rect 29564 22982 29592 25706
rect 29552 22976 29604 22982
rect 29552 22918 29604 22924
rect 29552 22704 29604 22710
rect 29552 22646 29604 22652
rect 29564 22438 29592 22646
rect 29552 22432 29604 22438
rect 29552 22374 29604 22380
rect 29552 21412 29604 21418
rect 29552 21354 29604 21360
rect 29564 20942 29592 21354
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29564 19553 29592 20878
rect 29656 20534 29684 27095
rect 29736 26580 29788 26586
rect 29736 26522 29788 26528
rect 29748 25702 29776 26522
rect 29828 26512 29880 26518
rect 29828 26454 29880 26460
rect 29736 25696 29788 25702
rect 29736 25638 29788 25644
rect 29748 25498 29776 25638
rect 29736 25492 29788 25498
rect 29736 25434 29788 25440
rect 29736 24880 29788 24886
rect 29736 24822 29788 24828
rect 29748 24138 29776 24822
rect 29736 24132 29788 24138
rect 29736 24074 29788 24080
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29748 22137 29776 23530
rect 29840 22982 29868 26454
rect 29932 26450 29960 27118
rect 29920 26444 29972 26450
rect 29920 26386 29972 26392
rect 29918 26072 29974 26081
rect 29918 26007 29974 26016
rect 29932 25906 29960 26007
rect 30024 25906 30052 27911
rect 30116 27674 30144 27950
rect 30104 27668 30156 27674
rect 30104 27610 30156 27616
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 30116 26897 30144 26998
rect 30102 26888 30158 26897
rect 30102 26823 30158 26832
rect 30104 26784 30156 26790
rect 30208 26772 30236 29106
rect 30484 28966 30512 29650
rect 30472 28960 30524 28966
rect 30472 28902 30524 28908
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 30484 28218 30512 28494
rect 30472 28212 30524 28218
rect 30472 28154 30524 28160
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30300 27402 30328 27814
rect 30378 27704 30434 27713
rect 30378 27639 30434 27648
rect 30392 27606 30420 27639
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30288 27396 30340 27402
rect 30288 27338 30340 27344
rect 30300 26790 30328 27338
rect 30392 26858 30420 27406
rect 30380 26852 30432 26858
rect 30380 26794 30432 26800
rect 30156 26744 30236 26772
rect 30288 26784 30340 26790
rect 30104 26726 30156 26732
rect 30288 26726 30340 26732
rect 29920 25900 29972 25906
rect 29920 25842 29972 25848
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 29932 25430 29960 25638
rect 29920 25424 29972 25430
rect 29920 25366 29972 25372
rect 29918 24168 29974 24177
rect 29918 24103 29974 24112
rect 29932 24070 29960 24103
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 30024 23322 30052 25842
rect 30012 23316 30064 23322
rect 30012 23258 30064 23264
rect 29828 22976 29880 22982
rect 29828 22918 29880 22924
rect 30012 22976 30064 22982
rect 30012 22918 30064 22924
rect 29734 22128 29790 22137
rect 29734 22063 29790 22072
rect 29736 20936 29788 20942
rect 29840 20924 29868 22918
rect 30024 22642 30052 22918
rect 29920 22636 29972 22642
rect 29920 22578 29972 22584
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 29932 21894 29960 22578
rect 30024 22234 30052 22578
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 30010 22128 30066 22137
rect 30010 22063 30066 22072
rect 29920 21888 29972 21894
rect 29920 21830 29972 21836
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29932 21078 29960 21490
rect 29920 21072 29972 21078
rect 29920 21014 29972 21020
rect 29788 20896 29868 20924
rect 29736 20878 29788 20884
rect 29644 20528 29696 20534
rect 29644 20470 29696 20476
rect 29828 20460 29880 20466
rect 29828 20402 29880 20408
rect 29840 20330 29868 20402
rect 29828 20324 29880 20330
rect 29828 20266 29880 20272
rect 30024 20210 30052 22063
rect 30116 20856 30144 26726
rect 30392 26450 30420 26794
rect 30484 26586 30512 27950
rect 30576 27878 30604 30126
rect 30668 29306 30696 30194
rect 30852 30161 30880 30738
rect 31036 30682 31064 30806
rect 30944 30654 31064 30682
rect 30944 30258 30972 30654
rect 31024 30592 31076 30598
rect 31116 30592 31168 30598
rect 31024 30534 31076 30540
rect 31114 30560 31116 30569
rect 31168 30560 31170 30569
rect 30932 30252 30984 30258
rect 30932 30194 30984 30200
rect 30838 30152 30894 30161
rect 30838 30087 30894 30096
rect 30748 29640 30800 29646
rect 30746 29608 30748 29617
rect 30840 29640 30892 29646
rect 30800 29608 30802 29617
rect 30840 29582 30892 29588
rect 30930 29608 30986 29617
rect 30746 29543 30802 29552
rect 30748 29504 30800 29510
rect 30748 29446 30800 29452
rect 30656 29300 30708 29306
rect 30656 29242 30708 29248
rect 30564 27872 30616 27878
rect 30564 27814 30616 27820
rect 30654 27840 30710 27849
rect 30654 27775 30710 27784
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 30472 26580 30524 26586
rect 30472 26522 30524 26528
rect 30196 26444 30248 26450
rect 30196 26386 30248 26392
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30208 25974 30236 26386
rect 30196 25968 30248 25974
rect 30248 25928 30328 25956
rect 30196 25910 30248 25916
rect 30196 24948 30248 24954
rect 30196 24890 30248 24896
rect 30208 23866 30236 24890
rect 30300 24290 30328 25928
rect 30576 25650 30604 27270
rect 30668 27062 30696 27775
rect 30760 27674 30788 29446
rect 30852 28422 30880 29582
rect 30930 29543 30986 29552
rect 30944 29306 30972 29543
rect 31036 29322 31064 30534
rect 31114 30495 31170 30504
rect 31220 29730 31248 31855
rect 31312 31142 31340 32166
rect 31496 32026 31524 32370
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 32496 32360 32548 32366
rect 32496 32302 32548 32308
rect 31484 32020 31536 32026
rect 31484 31962 31536 31968
rect 32324 31890 32352 32302
rect 31392 31884 31444 31890
rect 31392 31826 31444 31832
rect 32312 31884 32364 31890
rect 32312 31826 32364 31832
rect 31300 31136 31352 31142
rect 31300 31078 31352 31084
rect 31404 30326 31432 31826
rect 31668 31136 31720 31142
rect 31668 31078 31720 31084
rect 31392 30320 31444 30326
rect 31392 30262 31444 30268
rect 31484 30252 31536 30258
rect 31484 30194 31536 30200
rect 31496 29850 31524 30194
rect 31484 29844 31536 29850
rect 31484 29786 31536 29792
rect 31390 29744 31446 29753
rect 31220 29702 31340 29730
rect 31208 29640 31260 29646
rect 31208 29582 31260 29588
rect 30932 29300 30984 29306
rect 31036 29294 31156 29322
rect 30932 29242 30984 29248
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 31036 28626 31064 29106
rect 31128 29073 31156 29294
rect 31220 29238 31248 29582
rect 31208 29232 31260 29238
rect 31208 29174 31260 29180
rect 31114 29064 31170 29073
rect 31114 28999 31170 29008
rect 31024 28620 31076 28626
rect 31024 28562 31076 28568
rect 30840 28416 30892 28422
rect 30840 28358 30892 28364
rect 30932 28008 30984 28014
rect 30930 27976 30932 27985
rect 30984 27976 30986 27985
rect 30930 27911 30986 27920
rect 30840 27872 30892 27878
rect 30840 27814 30892 27820
rect 30748 27668 30800 27674
rect 30748 27610 30800 27616
rect 30656 27056 30708 27062
rect 30656 26998 30708 27004
rect 30760 26994 30788 27610
rect 30756 26988 30808 26994
rect 30756 26930 30808 26936
rect 30656 26852 30708 26858
rect 30656 26794 30708 26800
rect 30484 25622 30604 25650
rect 30380 24812 30432 24818
rect 30380 24754 30432 24760
rect 30392 24410 30420 24754
rect 30380 24404 30432 24410
rect 30380 24346 30432 24352
rect 30300 24262 30420 24290
rect 30196 23860 30248 23866
rect 30196 23802 30248 23808
rect 30208 23118 30236 23802
rect 30288 23520 30340 23526
rect 30288 23462 30340 23468
rect 30300 23118 30328 23462
rect 30392 23254 30420 24262
rect 30380 23248 30432 23254
rect 30380 23190 30432 23196
rect 30196 23112 30248 23118
rect 30196 23054 30248 23060
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30208 22642 30236 22918
rect 30300 22642 30328 23054
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30196 22500 30248 22506
rect 30196 22442 30248 22448
rect 30208 22166 30236 22442
rect 30392 22234 30420 23054
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30196 22160 30248 22166
rect 30196 22102 30248 22108
rect 30208 22030 30236 22102
rect 30196 22024 30248 22030
rect 30196 21966 30248 21972
rect 30288 21888 30340 21894
rect 30340 21836 30420 21842
rect 30288 21830 30420 21836
rect 30300 21814 30420 21830
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 30196 20868 30248 20874
rect 30116 20828 30196 20856
rect 30196 20810 30248 20816
rect 30300 20534 30328 21626
rect 30392 21010 30420 21814
rect 30380 21004 30432 21010
rect 30380 20946 30432 20952
rect 30288 20528 30340 20534
rect 30288 20470 30340 20476
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 29656 20182 30052 20210
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29550 19544 29606 19553
rect 29550 19479 29606 19488
rect 29564 19378 29592 19479
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29552 18692 29604 18698
rect 29552 18634 29604 18640
rect 29460 18148 29512 18154
rect 29460 18090 29512 18096
rect 29368 17332 29420 17338
rect 29564 17320 29592 18634
rect 29656 17610 29684 20182
rect 29828 20052 29880 20058
rect 29828 19994 29880 20000
rect 29920 20052 29972 20058
rect 29920 19994 29972 20000
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29748 19446 29776 19790
rect 29736 19440 29788 19446
rect 29840 19417 29868 19994
rect 29736 19382 29788 19388
rect 29826 19408 29882 19417
rect 29644 17604 29696 17610
rect 29644 17546 29696 17552
rect 29564 17292 29684 17320
rect 29368 17274 29420 17280
rect 29288 17190 29592 17218
rect 29276 17128 29328 17134
rect 29276 17070 29328 17076
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29182 16144 29238 16153
rect 29182 16079 29184 16088
rect 29236 16079 29238 16088
rect 29184 16050 29236 16056
rect 28920 15660 29132 15688
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28724 15428 28776 15434
rect 28724 15370 28776 15376
rect 28540 14816 28592 14822
rect 28540 14758 28592 14764
rect 28736 14550 28764 15370
rect 28828 15094 28856 15438
rect 28920 15162 28948 15660
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 28908 15156 28960 15162
rect 28908 15098 28960 15104
rect 28816 15088 28868 15094
rect 28816 15030 28868 15036
rect 29012 15026 29040 15506
rect 29288 15314 29316 17070
rect 29380 16590 29408 17070
rect 29368 16584 29420 16590
rect 29368 16526 29420 16532
rect 29380 16153 29408 16526
rect 29366 16144 29422 16153
rect 29366 16079 29368 16088
rect 29420 16079 29422 16088
rect 29368 16050 29420 16056
rect 29380 15570 29408 16050
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29196 15286 29316 15314
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 28816 14952 28868 14958
rect 28816 14894 28868 14900
rect 28828 14822 28856 14894
rect 28816 14816 28868 14822
rect 28920 14793 28948 14962
rect 28816 14758 28868 14764
rect 28906 14784 28962 14793
rect 28906 14719 28962 14728
rect 28632 14544 28684 14550
rect 28632 14486 28684 14492
rect 28724 14544 28776 14550
rect 28724 14486 28776 14492
rect 28644 13870 28672 14486
rect 28736 13938 28764 14486
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28920 13938 28948 14214
rect 28724 13932 28776 13938
rect 28724 13874 28776 13880
rect 28908 13932 28960 13938
rect 28908 13874 28960 13880
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 28632 13864 28684 13870
rect 28552 13824 28632 13852
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28368 12804 28488 12832
rect 28080 12708 28132 12714
rect 28184 12702 28396 12730
rect 28080 12650 28132 12656
rect 28264 12640 28316 12646
rect 28264 12582 28316 12588
rect 28170 12336 28226 12345
rect 28276 12306 28304 12582
rect 28170 12271 28226 12280
rect 28264 12300 28316 12306
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 27988 12096 28040 12102
rect 27988 12038 28040 12044
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 27802 10976 27858 10985
rect 27802 10911 27858 10920
rect 27816 10810 27844 10911
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27908 10606 27936 11290
rect 28000 10674 28028 11834
rect 28092 11150 28120 12106
rect 28184 11898 28212 12271
rect 28264 12242 28316 12248
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28276 11762 28304 12106
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28170 11384 28226 11393
rect 28170 11319 28226 11328
rect 28184 11150 28212 11319
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28184 10742 28212 11086
rect 28172 10736 28224 10742
rect 28172 10678 28224 10684
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 27896 10600 27948 10606
rect 27896 10542 27948 10548
rect 27804 10532 27856 10538
rect 27804 10474 27856 10480
rect 27816 9625 27844 10474
rect 27908 10198 27936 10542
rect 27896 10192 27948 10198
rect 27896 10134 27948 10140
rect 27896 10056 27948 10062
rect 27894 10024 27896 10033
rect 27948 10024 27950 10033
rect 27894 9959 27950 9968
rect 27802 9616 27858 9625
rect 27802 9551 27858 9560
rect 27804 9512 27856 9518
rect 27804 9454 27856 9460
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27816 8906 27844 9454
rect 28000 9042 28028 10610
rect 28080 10532 28132 10538
rect 28080 10474 28132 10480
rect 28092 10282 28120 10474
rect 28172 10464 28224 10470
rect 28170 10432 28172 10441
rect 28224 10432 28226 10441
rect 28170 10367 28226 10376
rect 28092 10254 28212 10282
rect 28078 10160 28134 10169
rect 28078 10095 28134 10104
rect 28092 9994 28120 10095
rect 28184 10062 28212 10254
rect 28172 10056 28224 10062
rect 28172 9998 28224 10004
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 27988 9036 28040 9042
rect 27988 8978 28040 8984
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27618 8256 27674 8265
rect 27618 8191 27674 8200
rect 27632 7274 27660 8191
rect 27724 7886 27752 8298
rect 27816 8022 27844 8842
rect 27908 8401 27936 8910
rect 27894 8392 27950 8401
rect 27894 8327 27950 8336
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 28000 7886 28028 8230
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 27908 7478 27936 7822
rect 27896 7472 27948 7478
rect 27896 7414 27948 7420
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 27528 6996 27580 7002
rect 27528 6938 27580 6944
rect 27122 6582 27200 6610
rect 27066 6559 27122 6568
rect 27080 6254 27108 6559
rect 27264 6322 27292 6870
rect 27448 6854 27568 6882
rect 27540 6798 27568 6854
rect 27344 6792 27396 6798
rect 27344 6734 27396 6740
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27356 6390 27384 6734
rect 27540 6458 27568 6734
rect 28092 6662 28120 7346
rect 28184 7342 28212 8910
rect 28172 7336 28224 7342
rect 28172 7278 28224 7284
rect 28080 6656 28132 6662
rect 28080 6598 28132 6604
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 27068 6248 27120 6254
rect 27068 6190 27120 6196
rect 27356 6118 27384 6326
rect 27540 6322 27568 6394
rect 28276 6322 28304 11698
rect 28368 11150 28396 12702
rect 28460 12442 28488 12804
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 28448 12300 28500 12306
rect 28448 12242 28500 12248
rect 28460 11558 28488 12242
rect 28552 11830 28580 13824
rect 28632 13806 28684 13812
rect 28906 13832 28962 13841
rect 28816 13796 28868 13802
rect 28906 13767 28908 13776
rect 28816 13738 28868 13744
rect 28960 13767 28962 13776
rect 28908 13738 28960 13744
rect 28828 13546 28856 13738
rect 29104 13546 29132 13874
rect 29196 13818 29224 15286
rect 29274 15192 29330 15201
rect 29274 15127 29330 15136
rect 29288 15094 29316 15127
rect 29276 15088 29328 15094
rect 29328 15048 29408 15076
rect 29276 15030 29328 15036
rect 29276 14952 29328 14958
rect 29276 14894 29328 14900
rect 29288 14482 29316 14894
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29380 13928 29408 15048
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 29472 14618 29500 14894
rect 29460 14612 29512 14618
rect 29460 14554 29512 14560
rect 29472 14482 29500 14554
rect 29460 14476 29512 14482
rect 29460 14418 29512 14424
rect 29460 14340 29512 14346
rect 29460 14282 29512 14288
rect 29368 13922 29420 13928
rect 29368 13864 29420 13870
rect 29196 13790 29408 13818
rect 29472 13802 29500 14282
rect 29564 13841 29592 17190
rect 29656 15094 29684 17292
rect 29748 15502 29776 19382
rect 29932 19378 29960 19994
rect 29826 19343 29882 19352
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29932 18426 29960 19314
rect 30116 18630 30144 20198
rect 30208 19378 30236 20402
rect 30288 20392 30340 20398
rect 30340 20340 30420 20346
rect 30288 20334 30420 20340
rect 30300 20318 30420 20334
rect 30286 19544 30342 19553
rect 30286 19479 30342 19488
rect 30300 19378 30328 19479
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30392 19334 30420 20318
rect 30484 19854 30512 25622
rect 30668 25537 30696 26794
rect 30748 26240 30800 26246
rect 30748 26182 30800 26188
rect 30760 25702 30788 26182
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30654 25528 30710 25537
rect 30654 25463 30710 25472
rect 30748 25152 30800 25158
rect 30748 25094 30800 25100
rect 30564 23520 30616 23526
rect 30564 23462 30616 23468
rect 30576 23118 30604 23462
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30576 22137 30604 22714
rect 30562 22128 30618 22137
rect 30562 22063 30618 22072
rect 30564 21956 30616 21962
rect 30564 21898 30616 21904
rect 30576 21622 30604 21898
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 30668 21486 30696 22918
rect 30656 21480 30708 21486
rect 30656 21422 30708 21428
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30576 20777 30604 20810
rect 30562 20768 30618 20777
rect 30562 20703 30618 20712
rect 30668 20262 30696 21422
rect 30760 20398 30788 25094
rect 30852 23118 30880 27814
rect 30932 27464 30984 27470
rect 31036 27452 31064 28562
rect 31116 28552 31168 28558
rect 31116 28494 31168 28500
rect 30984 27424 31064 27452
rect 30932 27406 30984 27412
rect 31036 27112 31064 27424
rect 30944 27084 31064 27112
rect 30944 26081 30972 27084
rect 31024 26988 31076 26994
rect 31024 26930 31076 26936
rect 31036 26353 31064 26930
rect 31022 26344 31078 26353
rect 31022 26279 31024 26288
rect 31076 26279 31078 26288
rect 31024 26250 31076 26256
rect 30930 26072 30986 26081
rect 30930 26007 30986 26016
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 30930 25528 30986 25537
rect 30930 25463 30986 25472
rect 30944 24954 30972 25463
rect 31036 25294 31064 25774
rect 31024 25288 31076 25294
rect 31024 25230 31076 25236
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 30944 24818 30972 24890
rect 30932 24812 30984 24818
rect 30932 24754 30984 24760
rect 30932 24608 30984 24614
rect 30932 24550 30984 24556
rect 31024 24608 31076 24614
rect 31024 24550 31076 24556
rect 30840 23112 30892 23118
rect 30944 23089 30972 24550
rect 30840 23054 30892 23060
rect 30930 23080 30986 23089
rect 30930 23015 30986 23024
rect 30932 22976 30984 22982
rect 30838 22944 30894 22953
rect 30932 22918 30984 22924
rect 30838 22879 30894 22888
rect 30852 22778 30880 22879
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30852 22098 30880 22578
rect 30840 22092 30892 22098
rect 30840 22034 30892 22040
rect 30852 21418 30880 22034
rect 30944 22030 30972 22918
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 31036 21570 31064 24550
rect 31128 24206 31156 28494
rect 31220 25294 31248 29174
rect 31312 28257 31340 29702
rect 31390 29679 31446 29688
rect 31404 29646 31432 29679
rect 31392 29640 31444 29646
rect 31392 29582 31444 29588
rect 31392 29096 31444 29102
rect 31392 29038 31444 29044
rect 31404 28937 31432 29038
rect 31390 28928 31446 28937
rect 31390 28863 31446 28872
rect 31392 28484 31444 28490
rect 31392 28426 31444 28432
rect 31404 28393 31432 28426
rect 31390 28384 31446 28393
rect 31390 28319 31446 28328
rect 31298 28248 31354 28257
rect 31496 28200 31524 29786
rect 31576 29776 31628 29782
rect 31576 29718 31628 29724
rect 31588 29238 31616 29718
rect 31680 29714 31708 31078
rect 32324 30802 32352 31826
rect 32404 31680 32456 31686
rect 32404 31622 32456 31628
rect 32416 31346 32444 31622
rect 32508 31482 32536 32302
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32496 31476 32548 31482
rect 32496 31418 32548 31424
rect 32404 31340 32456 31346
rect 32456 31300 32536 31328
rect 32404 31282 32456 31288
rect 32508 30870 32536 31300
rect 32496 30864 32548 30870
rect 32496 30806 32548 30812
rect 32312 30796 32364 30802
rect 32312 30738 32364 30744
rect 32404 30388 32456 30394
rect 32404 30330 32456 30336
rect 32220 30320 32272 30326
rect 32220 30262 32272 30268
rect 31760 30252 31812 30258
rect 31760 30194 31812 30200
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 31772 30161 31800 30194
rect 32140 30161 32168 30194
rect 31758 30152 31814 30161
rect 32126 30152 32182 30161
rect 31814 30122 31984 30138
rect 31814 30116 31996 30122
rect 31814 30110 31944 30116
rect 31758 30087 31814 30096
rect 32126 30087 32182 30096
rect 31944 30058 31996 30064
rect 31668 29708 31720 29714
rect 31668 29650 31720 29656
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 32140 29510 32168 29582
rect 32232 29510 32260 30262
rect 32416 30258 32444 30330
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32404 30252 32456 30258
rect 32404 30194 32456 30200
rect 32324 29782 32352 30194
rect 32312 29776 32364 29782
rect 32416 29753 32444 30194
rect 32312 29718 32364 29724
rect 32402 29744 32458 29753
rect 32402 29679 32458 29688
rect 32404 29640 32456 29646
rect 32310 29608 32366 29617
rect 32366 29588 32404 29594
rect 32366 29582 32456 29588
rect 32366 29566 32444 29582
rect 32310 29543 32366 29552
rect 32508 29560 32536 30806
rect 32600 30054 32628 31758
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 33048 31340 33100 31346
rect 33048 31282 33100 31288
rect 32692 30394 32720 31282
rect 32864 30660 32916 30666
rect 32864 30602 32916 30608
rect 32680 30388 32732 30394
rect 32680 30330 32732 30336
rect 32876 30326 32904 30602
rect 32864 30320 32916 30326
rect 32864 30262 32916 30268
rect 32772 30252 32824 30258
rect 32772 30194 32824 30200
rect 32956 30252 33008 30258
rect 32956 30194 33008 30200
rect 32588 30048 32640 30054
rect 32588 29990 32640 29996
rect 32680 29640 32732 29646
rect 32680 29582 32732 29588
rect 32588 29572 32640 29578
rect 31668 29504 31720 29510
rect 31668 29446 31720 29452
rect 32128 29504 32180 29510
rect 32128 29446 32180 29452
rect 32220 29504 32272 29510
rect 32220 29446 32272 29452
rect 31680 29306 31708 29446
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 32036 29300 32088 29306
rect 32036 29242 32088 29248
rect 31576 29232 31628 29238
rect 31576 29174 31628 29180
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 31576 29096 31628 29102
rect 31574 29064 31576 29073
rect 31628 29064 31630 29073
rect 31956 29034 31984 29106
rect 31574 28999 31630 29008
rect 31944 29028 31996 29034
rect 31944 28970 31996 28976
rect 31850 28792 31906 28801
rect 31850 28727 31906 28736
rect 31574 28520 31630 28529
rect 31574 28455 31630 28464
rect 31588 28422 31616 28455
rect 31576 28416 31628 28422
rect 31576 28358 31628 28364
rect 31588 28218 31616 28358
rect 31298 28183 31354 28192
rect 31312 28150 31340 28183
rect 31404 28172 31524 28200
rect 31576 28212 31628 28218
rect 31300 28144 31352 28150
rect 31300 28086 31352 28092
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31312 25294 31340 27814
rect 31208 25288 31260 25294
rect 31208 25230 31260 25236
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 31116 24200 31168 24206
rect 31116 24142 31168 24148
rect 31116 23520 31168 23526
rect 31220 23508 31248 25230
rect 31300 24880 31352 24886
rect 31298 24848 31300 24857
rect 31352 24848 31354 24857
rect 31298 24783 31354 24792
rect 31300 24608 31352 24614
rect 31300 24550 31352 24556
rect 31312 24449 31340 24550
rect 31298 24440 31354 24449
rect 31298 24375 31354 24384
rect 31404 23746 31432 28172
rect 31864 28200 31892 28727
rect 31944 28688 31996 28694
rect 31942 28656 31944 28665
rect 31996 28656 31998 28665
rect 31942 28591 31998 28600
rect 32048 28558 32076 29242
rect 32140 29238 32168 29446
rect 32128 29232 32180 29238
rect 32128 29174 32180 29180
rect 32140 28558 32168 29174
rect 32036 28552 32088 28558
rect 31576 28154 31628 28160
rect 31772 28172 31892 28200
rect 31956 28512 32036 28540
rect 31666 28112 31722 28121
rect 31484 28076 31536 28082
rect 31484 28018 31536 28024
rect 31576 28076 31628 28082
rect 31666 28047 31722 28056
rect 31576 28018 31628 28024
rect 31496 27538 31524 28018
rect 31588 27849 31616 28018
rect 31680 27946 31708 28047
rect 31772 27946 31800 28172
rect 31668 27940 31720 27946
rect 31668 27882 31720 27888
rect 31760 27940 31812 27946
rect 31760 27882 31812 27888
rect 31574 27840 31630 27849
rect 31956 27826 31984 28512
rect 32036 28494 32088 28500
rect 32128 28552 32180 28558
rect 32128 28494 32180 28500
rect 32036 28416 32088 28422
rect 32036 28358 32088 28364
rect 31574 27775 31630 27784
rect 31772 27798 31984 27826
rect 32048 28200 32076 28358
rect 32128 28212 32180 28218
rect 32048 28172 32128 28200
rect 31484 27532 31536 27538
rect 31484 27474 31536 27480
rect 31484 27328 31536 27334
rect 31484 27270 31536 27276
rect 31496 27130 31524 27270
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31496 24750 31524 27066
rect 31588 27062 31616 27775
rect 31772 27470 31800 27798
rect 31852 27668 31904 27674
rect 31852 27610 31904 27616
rect 31864 27470 31892 27610
rect 31760 27464 31812 27470
rect 31760 27406 31812 27412
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31668 27396 31720 27402
rect 31668 27338 31720 27344
rect 31576 27056 31628 27062
rect 31576 26998 31628 27004
rect 31484 24744 31536 24750
rect 31484 24686 31536 24692
rect 31588 23798 31616 26998
rect 31680 24410 31708 27338
rect 31772 26382 31800 27406
rect 32048 27334 32076 28172
rect 32128 28154 32180 28160
rect 32128 28008 32180 28014
rect 32128 27950 32180 27956
rect 32140 27674 32168 27950
rect 32128 27668 32180 27674
rect 32128 27610 32180 27616
rect 32232 27384 32260 29446
rect 32324 29306 32352 29543
rect 32508 29532 32588 29560
rect 32588 29514 32640 29520
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32416 29209 32444 29446
rect 32494 29336 32550 29345
rect 32494 29271 32550 29280
rect 32402 29200 32458 29209
rect 32402 29135 32404 29144
rect 32456 29135 32458 29144
rect 32404 29106 32456 29112
rect 32402 29064 32458 29073
rect 32402 28999 32458 29008
rect 32312 28960 32364 28966
rect 32312 28902 32364 28908
rect 32324 28393 32352 28902
rect 32310 28384 32366 28393
rect 32310 28319 32366 28328
rect 32324 27606 32352 28319
rect 32416 28064 32444 28999
rect 32508 28218 32536 29271
rect 32588 29164 32640 29170
rect 32588 29106 32640 29112
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32496 28076 32548 28082
rect 32416 28036 32496 28064
rect 32312 27600 32364 27606
rect 32312 27542 32364 27548
rect 32140 27356 32260 27384
rect 32036 27328 32088 27334
rect 32036 27270 32088 27276
rect 31852 27056 31904 27062
rect 31852 26998 31904 27004
rect 31760 26376 31812 26382
rect 31760 26318 31812 26324
rect 31760 25900 31812 25906
rect 31864 25888 31892 26998
rect 32140 26518 32168 27356
rect 32220 27124 32272 27130
rect 32220 27066 32272 27072
rect 32128 26512 32180 26518
rect 32128 26454 32180 26460
rect 32128 26308 32180 26314
rect 32128 26250 32180 26256
rect 31944 26240 31996 26246
rect 31944 26182 31996 26188
rect 31956 25906 31984 26182
rect 32034 26072 32090 26081
rect 32140 26042 32168 26250
rect 32034 26007 32036 26016
rect 32088 26007 32090 26016
rect 32128 26036 32180 26042
rect 32036 25978 32088 25984
rect 32128 25978 32180 25984
rect 31812 25860 31892 25888
rect 31760 25842 31812 25848
rect 31864 25786 31892 25860
rect 31944 25900 31996 25906
rect 31944 25842 31996 25848
rect 32128 25900 32180 25906
rect 32232 25888 32260 27066
rect 32416 27062 32444 28036
rect 32496 28018 32548 28024
rect 32600 27878 32628 29106
rect 32692 28694 32720 29582
rect 32784 29306 32812 30194
rect 32864 30048 32916 30054
rect 32864 29990 32916 29996
rect 32772 29300 32824 29306
rect 32772 29242 32824 29248
rect 32876 29186 32904 29990
rect 32784 29158 32904 29186
rect 32784 29102 32812 29158
rect 32772 29096 32824 29102
rect 32772 29038 32824 29044
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 32680 28688 32732 28694
rect 32680 28630 32732 28636
rect 32680 28552 32732 28558
rect 32678 28520 32680 28529
rect 32732 28520 32734 28529
rect 32678 28455 32734 28464
rect 32678 28112 32734 28121
rect 32678 28047 32734 28056
rect 32692 27878 32720 28047
rect 32588 27872 32640 27878
rect 32588 27814 32640 27820
rect 32680 27872 32732 27878
rect 32680 27814 32732 27820
rect 32494 27432 32550 27441
rect 32784 27402 32812 29038
rect 32876 28937 32904 29038
rect 32862 28928 32918 28937
rect 32862 28863 32918 28872
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32494 27367 32550 27376
rect 32772 27396 32824 27402
rect 32404 27056 32456 27062
rect 32404 26998 32456 27004
rect 32404 26784 32456 26790
rect 32404 26726 32456 26732
rect 32416 26246 32444 26726
rect 32508 26246 32536 27367
rect 32772 27338 32824 27344
rect 32784 27130 32812 27338
rect 32772 27124 32824 27130
rect 32772 27066 32824 27072
rect 32588 27056 32640 27062
rect 32588 26998 32640 27004
rect 32404 26240 32456 26246
rect 32404 26182 32456 26188
rect 32496 26240 32548 26246
rect 32496 26182 32548 26188
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32180 25860 32260 25888
rect 32128 25842 32180 25848
rect 31864 25758 31984 25786
rect 31852 25696 31904 25702
rect 31852 25638 31904 25644
rect 31864 25294 31892 25638
rect 31760 25288 31812 25294
rect 31758 25256 31760 25265
rect 31852 25288 31904 25294
rect 31812 25256 31814 25265
rect 31852 25230 31904 25236
rect 31758 25191 31814 25200
rect 31864 24954 31892 25230
rect 31852 24948 31904 24954
rect 31852 24890 31904 24896
rect 31760 24608 31812 24614
rect 31760 24550 31812 24556
rect 31668 24404 31720 24410
rect 31668 24346 31720 24352
rect 31680 24070 31708 24346
rect 31772 24138 31800 24550
rect 31760 24132 31812 24138
rect 31760 24074 31812 24080
rect 31668 24064 31720 24070
rect 31668 24006 31720 24012
rect 31576 23792 31628 23798
rect 31300 23724 31352 23730
rect 31404 23718 31524 23746
rect 31576 23734 31628 23740
rect 31300 23666 31352 23672
rect 31168 23480 31248 23508
rect 31116 23462 31168 23468
rect 31116 23248 31168 23254
rect 31116 23190 31168 23196
rect 31128 22710 31156 23190
rect 31208 23112 31260 23118
rect 31208 23054 31260 23060
rect 31220 22982 31248 23054
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 31116 22568 31168 22574
rect 31116 22510 31168 22516
rect 31128 22234 31156 22510
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 31220 22114 31248 22918
rect 31128 22086 31248 22114
rect 31128 21894 31156 22086
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31116 21888 31168 21894
rect 31116 21830 31168 21836
rect 30944 21542 31064 21570
rect 30840 21412 30892 21418
rect 30840 21354 30892 21360
rect 30840 20868 30892 20874
rect 30840 20810 30892 20816
rect 30852 20466 30880 20810
rect 30840 20460 30892 20466
rect 30840 20402 30892 20408
rect 30748 20392 30800 20398
rect 30748 20334 30800 20340
rect 30840 20324 30892 20330
rect 30840 20266 30892 20272
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30472 19848 30524 19854
rect 30472 19790 30524 19796
rect 30484 19446 30512 19790
rect 30852 19689 30880 20266
rect 30838 19680 30894 19689
rect 30838 19615 30894 19624
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 30472 19440 30524 19446
rect 30472 19382 30524 19388
rect 30392 19306 30604 19334
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 29920 18420 29972 18426
rect 29920 18362 29972 18368
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 29828 16652 29880 16658
rect 29828 16594 29880 16600
rect 29840 16250 29868 16594
rect 29828 16244 29880 16250
rect 29828 16186 29880 16192
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29644 15088 29696 15094
rect 29644 15030 29696 15036
rect 29840 15026 29868 16186
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 29644 14952 29696 14958
rect 29644 14894 29696 14900
rect 29656 14346 29684 14894
rect 29736 14612 29788 14618
rect 29736 14554 29788 14560
rect 29644 14340 29696 14346
rect 29644 14282 29696 14288
rect 29550 13832 29606 13841
rect 28828 13530 28948 13546
rect 28724 13524 28776 13530
rect 28828 13524 28960 13530
rect 28828 13518 28908 13524
rect 28724 13466 28776 13472
rect 28908 13466 28960 13472
rect 29012 13518 29132 13546
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28644 12628 28672 13262
rect 28736 12850 28764 13466
rect 29012 13394 29040 13518
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29000 13252 29052 13258
rect 29000 13194 29052 13200
rect 29012 12850 29040 13194
rect 28724 12844 28776 12850
rect 28724 12786 28776 12792
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 28724 12640 28776 12646
rect 28644 12600 28724 12628
rect 28540 11824 28592 11830
rect 28540 11766 28592 11772
rect 28448 11552 28500 11558
rect 28448 11494 28500 11500
rect 28460 11150 28488 11494
rect 28552 11354 28580 11766
rect 28540 11348 28592 11354
rect 28540 11290 28592 11296
rect 28356 11144 28408 11150
rect 28354 11112 28356 11121
rect 28448 11144 28500 11150
rect 28408 11112 28410 11121
rect 28448 11086 28500 11092
rect 28354 11047 28410 11056
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28368 10130 28396 10474
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28460 9518 28488 10950
rect 28552 10810 28580 11290
rect 28644 11150 28672 12600
rect 28724 12582 28776 12588
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 29092 12640 29144 12646
rect 29092 12582 29144 12588
rect 28828 12481 28856 12582
rect 28814 12472 28870 12481
rect 28724 12436 28776 12442
rect 28814 12407 28870 12416
rect 28724 12378 28776 12384
rect 28736 12186 28764 12378
rect 28828 12306 28856 12407
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28908 12232 28960 12238
rect 28736 12158 28856 12186
rect 28908 12174 28960 12180
rect 28724 12096 28776 12102
rect 28722 12064 28724 12073
rect 28776 12064 28778 12073
rect 28722 11999 28778 12008
rect 28828 11880 28856 12158
rect 28736 11852 28856 11880
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28632 11008 28684 11014
rect 28736 10996 28764 11852
rect 28920 11830 28948 12174
rect 28908 11824 28960 11830
rect 28908 11766 28960 11772
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 28828 11286 28856 11698
rect 28816 11280 28868 11286
rect 28816 11222 28868 11228
rect 28684 10968 28764 10996
rect 28632 10950 28684 10956
rect 28540 10804 28592 10810
rect 28540 10746 28592 10752
rect 28724 10736 28776 10742
rect 28644 10684 28724 10690
rect 28920 10724 28948 11766
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29012 11150 29040 11290
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 28644 10678 28776 10684
rect 28895 10696 28948 10724
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 28644 10662 28764 10678
rect 28552 10305 28580 10610
rect 28538 10296 28594 10305
rect 28538 10231 28594 10240
rect 28552 9722 28580 10231
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28356 8968 28408 8974
rect 28354 8936 28356 8945
rect 28408 8936 28410 8945
rect 28354 8871 28410 8880
rect 28368 6662 28396 8871
rect 28552 8634 28580 9658
rect 28644 8838 28672 10662
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28736 10198 28764 10542
rect 28895 10452 28923 10696
rect 28828 10424 28923 10452
rect 29104 10441 29132 12582
rect 29182 11656 29238 11665
rect 29288 11626 29316 13262
rect 29182 11591 29238 11600
rect 29276 11620 29328 11626
rect 29196 11558 29224 11591
rect 29276 11562 29328 11568
rect 29184 11552 29236 11558
rect 29184 11494 29236 11500
rect 29196 11354 29224 11494
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 29184 11144 29236 11150
rect 29184 11086 29236 11092
rect 29196 11014 29224 11086
rect 29184 11008 29236 11014
rect 29184 10950 29236 10956
rect 29274 10976 29330 10985
rect 29196 10810 29224 10950
rect 29274 10911 29330 10920
rect 29288 10810 29316 10911
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29276 10804 29328 10810
rect 29276 10746 29328 10752
rect 29090 10432 29146 10441
rect 28724 10192 28776 10198
rect 28724 10134 28776 10140
rect 28736 9761 28764 10134
rect 28722 9752 28778 9761
rect 28722 9687 28778 9696
rect 28736 9654 28764 9687
rect 28724 9648 28776 9654
rect 28724 9590 28776 9596
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28736 9217 28764 9318
rect 28722 9208 28778 9217
rect 28722 9143 28778 9152
rect 28828 8906 28856 10424
rect 29090 10367 29146 10376
rect 29288 10169 29316 10746
rect 29274 10160 29330 10169
rect 29274 10095 29330 10104
rect 29184 10056 29236 10062
rect 28908 10034 28960 10040
rect 28906 10024 28908 10033
rect 28960 10024 28962 10033
rect 29184 9998 29236 10004
rect 28906 9959 28962 9968
rect 28908 9512 28960 9518
rect 28960 9460 29040 9466
rect 28908 9454 29040 9460
rect 28920 9438 29040 9454
rect 28908 9376 28960 9382
rect 28908 9318 28960 9324
rect 28816 8900 28868 8906
rect 28816 8842 28868 8848
rect 28632 8832 28684 8838
rect 28632 8774 28684 8780
rect 28644 8634 28672 8774
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28828 8498 28856 8842
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28552 8294 28580 8366
rect 28644 8294 28672 8434
rect 28540 8288 28592 8294
rect 28540 8230 28592 8236
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28644 7954 28672 8230
rect 28828 8090 28856 8434
rect 28920 8430 28948 9318
rect 29012 8838 29040 9438
rect 29196 9042 29224 9998
rect 29274 9888 29330 9897
rect 29274 9823 29330 9832
rect 29288 9586 29316 9823
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29380 9110 29408 13790
rect 29460 13796 29512 13802
rect 29550 13767 29606 13776
rect 29460 13738 29512 13744
rect 29550 13560 29606 13569
rect 29550 13495 29606 13504
rect 29460 12844 29512 12850
rect 29460 12786 29512 12792
rect 29472 10266 29500 12786
rect 29564 12458 29592 13495
rect 29564 12430 29684 12458
rect 29552 11688 29604 11694
rect 29550 11656 29552 11665
rect 29604 11656 29606 11665
rect 29550 11591 29606 11600
rect 29550 11112 29606 11121
rect 29550 11047 29606 11056
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 29472 9654 29500 10202
rect 29564 10062 29592 11047
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29460 9648 29512 9654
rect 29460 9590 29512 9596
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29368 9104 29420 9110
rect 29368 9046 29420 9052
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 29012 8514 29040 8774
rect 29012 8486 29132 8514
rect 29104 8430 29132 8486
rect 28908 8424 28960 8430
rect 28908 8366 28960 8372
rect 29092 8424 29144 8430
rect 29092 8366 29144 8372
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28540 7268 28592 7274
rect 28540 7210 28592 7216
rect 28552 6746 28580 7210
rect 28644 6798 28672 7890
rect 28920 7886 28948 8366
rect 29196 8090 29224 8978
rect 29564 8974 29592 9590
rect 29656 8974 29684 12430
rect 29748 12374 29776 14554
rect 29828 14544 29880 14550
rect 29828 14486 29880 14492
rect 29736 12368 29788 12374
rect 29736 12310 29788 12316
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29748 9926 29776 10610
rect 29840 10062 29868 14486
rect 29932 14074 29960 15982
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 29920 13796 29972 13802
rect 29920 13738 29972 13744
rect 29932 13326 29960 13738
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29918 10704 29974 10713
rect 29918 10639 29920 10648
rect 29972 10639 29974 10648
rect 29920 10610 29972 10616
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 29736 9920 29788 9926
rect 29828 9920 29880 9926
rect 29736 9862 29788 9868
rect 29826 9888 29828 9897
rect 29880 9888 29882 9897
rect 29748 9110 29776 9862
rect 29826 9823 29882 9832
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29644 8968 29696 8974
rect 29644 8910 29696 8916
rect 29458 8256 29514 8265
rect 29458 8191 29514 8200
rect 29184 8084 29236 8090
rect 29184 8026 29236 8032
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28816 7812 28868 7818
rect 28816 7754 28868 7760
rect 28828 7478 28856 7754
rect 28816 7472 28868 7478
rect 28816 7414 28868 7420
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28460 6730 28580 6746
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28448 6724 28580 6730
rect 28500 6718 28580 6724
rect 28448 6666 28500 6672
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28460 6458 28488 6666
rect 28448 6452 28500 6458
rect 28448 6394 28500 6400
rect 28644 6390 28672 6734
rect 28736 6730 28764 7346
rect 28828 6934 28856 7414
rect 28920 7342 28948 7822
rect 29184 7812 29236 7818
rect 29184 7754 29236 7760
rect 28998 7576 29054 7585
rect 28998 7511 29000 7520
rect 29052 7511 29054 7520
rect 29000 7482 29052 7488
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 29196 7002 29224 7754
rect 29288 7750 29316 8026
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 29276 7744 29328 7750
rect 29276 7686 29328 7692
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 29380 6866 29408 7958
rect 29472 7818 29500 8191
rect 29460 7812 29512 7818
rect 29460 7754 29512 7760
rect 29368 6860 29420 6866
rect 29368 6802 29420 6808
rect 28724 6724 28776 6730
rect 28724 6666 28776 6672
rect 28722 6624 28778 6633
rect 28722 6559 28778 6568
rect 28736 6390 28764 6559
rect 28632 6384 28684 6390
rect 28632 6326 28684 6332
rect 28724 6384 28776 6390
rect 28724 6326 28776 6332
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 28264 6316 28316 6322
rect 28264 6258 28316 6264
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 28276 5778 28304 6258
rect 29380 6254 29408 6802
rect 29564 6730 29592 8910
rect 29552 6724 29604 6730
rect 29552 6666 29604 6672
rect 29368 6248 29420 6254
rect 29368 6190 29420 6196
rect 29656 5914 29684 8910
rect 29748 8022 29776 9046
rect 29840 8566 29868 9522
rect 29932 9382 29960 9930
rect 30024 9586 30052 18226
rect 30116 16590 30144 18566
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30300 17338 30328 18226
rect 30472 18080 30524 18086
rect 30472 18022 30524 18028
rect 30288 17332 30340 17338
rect 30288 17274 30340 17280
rect 30104 16584 30156 16590
rect 30104 16526 30156 16532
rect 30300 16522 30328 17274
rect 30288 16516 30340 16522
rect 30288 16458 30340 16464
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30196 16040 30248 16046
rect 30194 16008 30196 16017
rect 30248 16008 30250 16017
rect 30104 15972 30156 15978
rect 30194 15943 30250 15952
rect 30104 15914 30156 15920
rect 30116 15706 30144 15914
rect 30104 15700 30156 15706
rect 30104 15642 30156 15648
rect 30194 15464 30250 15473
rect 30194 15399 30250 15408
rect 30104 14272 30156 14278
rect 30104 14214 30156 14220
rect 30116 13938 30144 14214
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30208 13870 30236 15399
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30300 14414 30328 14894
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30196 13864 30248 13870
rect 30196 13806 30248 13812
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30104 11008 30156 11014
rect 30104 10950 30156 10956
rect 30116 10062 30144 10950
rect 30300 10538 30328 11698
rect 30392 11354 30420 16050
rect 30484 12850 30512 18022
rect 30576 16182 30604 19306
rect 30760 18358 30788 19450
rect 30748 18352 30800 18358
rect 30748 18294 30800 18300
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30564 16176 30616 16182
rect 30564 16118 30616 16124
rect 30564 16040 30616 16046
rect 30564 15982 30616 15988
rect 30576 14414 30604 15982
rect 30668 15910 30696 16390
rect 30748 16176 30800 16182
rect 30748 16118 30800 16124
rect 30656 15904 30708 15910
rect 30656 15846 30708 15852
rect 30760 15502 30788 16118
rect 30748 15496 30800 15502
rect 30748 15438 30800 15444
rect 30748 15156 30800 15162
rect 30748 15098 30800 15104
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30576 13433 30604 14214
rect 30668 13938 30696 14758
rect 30656 13932 30708 13938
rect 30656 13874 30708 13880
rect 30562 13424 30618 13433
rect 30562 13359 30618 13368
rect 30760 12850 30788 15098
rect 30472 12844 30524 12850
rect 30472 12786 30524 12792
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30746 12744 30802 12753
rect 30746 12679 30748 12688
rect 30800 12679 30802 12688
rect 30748 12650 30800 12656
rect 30746 12472 30802 12481
rect 30746 12407 30802 12416
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 30288 10532 30340 10538
rect 30288 10474 30340 10480
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30208 9926 30236 9998
rect 30392 9926 30420 11154
rect 30576 11150 30604 11698
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 30668 10606 30696 11018
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30760 10062 30788 12407
rect 30852 11014 30880 18158
rect 30944 18086 30972 21542
rect 31024 21412 31076 21418
rect 31024 21354 31076 21360
rect 31036 21146 31064 21354
rect 31116 21344 31168 21350
rect 31116 21286 31168 21292
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 31128 20942 31156 21286
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31024 20800 31076 20806
rect 31024 20742 31076 20748
rect 31036 18698 31064 20742
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 31024 18692 31076 18698
rect 31024 18634 31076 18640
rect 30932 18080 30984 18086
rect 30932 18022 30984 18028
rect 30930 17912 30986 17921
rect 30930 17847 30986 17856
rect 30944 16114 30972 17847
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 31036 15570 31064 17546
rect 31024 15564 31076 15570
rect 30944 15524 31024 15552
rect 30944 12714 30972 15524
rect 31024 15506 31076 15512
rect 31128 14482 31156 20334
rect 31220 18970 31248 21966
rect 31312 21418 31340 23666
rect 31392 23588 31444 23594
rect 31392 23530 31444 23536
rect 31404 22574 31432 23530
rect 31496 23118 31524 23718
rect 31668 23588 31720 23594
rect 31668 23530 31720 23536
rect 31576 23316 31628 23322
rect 31576 23258 31628 23264
rect 31484 23112 31536 23118
rect 31484 23054 31536 23060
rect 31484 22772 31536 22778
rect 31484 22714 31536 22720
rect 31392 22568 31444 22574
rect 31496 22545 31524 22714
rect 31588 22642 31616 23258
rect 31680 23186 31708 23530
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31760 23112 31812 23118
rect 31666 23080 31722 23089
rect 31864 23100 31892 24890
rect 31956 24886 31984 25758
rect 32220 25696 32272 25702
rect 32220 25638 32272 25644
rect 32232 25430 32260 25638
rect 32220 25424 32272 25430
rect 32220 25366 32272 25372
rect 32036 25356 32088 25362
rect 32088 25316 32168 25344
rect 32036 25298 32088 25304
rect 32034 25256 32090 25265
rect 32034 25191 32090 25200
rect 31944 24880 31996 24886
rect 31944 24822 31996 24828
rect 31956 24614 31984 24822
rect 31944 24608 31996 24614
rect 31944 24550 31996 24556
rect 31944 24132 31996 24138
rect 31944 24074 31996 24080
rect 31812 23072 31892 23100
rect 31760 23054 31812 23060
rect 31666 23015 31722 23024
rect 31576 22636 31628 22642
rect 31576 22578 31628 22584
rect 31392 22510 31444 22516
rect 31482 22536 31538 22545
rect 31482 22471 31538 22480
rect 31680 22438 31708 23015
rect 31576 22432 31628 22438
rect 31576 22374 31628 22380
rect 31668 22432 31720 22438
rect 31668 22374 31720 22380
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31404 21146 31432 21422
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31484 21004 31536 21010
rect 31484 20946 31536 20952
rect 31496 20641 31524 20946
rect 31588 20942 31616 22374
rect 31772 21690 31800 23054
rect 31850 22944 31906 22953
rect 31850 22879 31906 22888
rect 31864 22710 31892 22879
rect 31852 22704 31904 22710
rect 31852 22646 31904 22652
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31758 21040 31814 21049
rect 31758 20975 31814 20984
rect 31772 20942 31800 20975
rect 31576 20936 31628 20942
rect 31576 20878 31628 20884
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31576 20800 31628 20806
rect 31576 20742 31628 20748
rect 31668 20800 31720 20806
rect 31668 20742 31720 20748
rect 31482 20632 31538 20641
rect 31482 20567 31538 20576
rect 31298 20496 31354 20505
rect 31298 20431 31354 20440
rect 31312 19854 31340 20431
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 31300 19848 31352 19854
rect 31404 19825 31432 20334
rect 31484 20256 31536 20262
rect 31484 20198 31536 20204
rect 31300 19790 31352 19796
rect 31390 19816 31446 19825
rect 31312 19718 31340 19790
rect 31390 19751 31446 19760
rect 31300 19712 31352 19718
rect 31300 19654 31352 19660
rect 31390 19680 31446 19689
rect 31312 19446 31340 19654
rect 31390 19615 31446 19624
rect 31300 19440 31352 19446
rect 31300 19382 31352 19388
rect 31404 19292 31432 19615
rect 31312 19264 31432 19292
rect 31208 18964 31260 18970
rect 31208 18906 31260 18912
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 31220 18426 31248 18634
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31220 16289 31248 17138
rect 31206 16280 31262 16289
rect 31206 16215 31262 16224
rect 31220 16114 31248 16215
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 31312 15994 31340 19264
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31220 15966 31340 15994
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 31036 12850 31064 14350
rect 31024 12844 31076 12850
rect 31024 12786 31076 12792
rect 30932 12708 30984 12714
rect 30932 12650 30984 12656
rect 30944 11830 30972 12650
rect 31220 12434 31248 15966
rect 31404 15706 31432 16050
rect 31496 15706 31524 20198
rect 31588 18902 31616 20742
rect 31680 20505 31708 20742
rect 31666 20496 31722 20505
rect 31666 20431 31722 20440
rect 31668 20392 31720 20398
rect 31666 20360 31668 20369
rect 31720 20360 31722 20369
rect 31666 20295 31722 20304
rect 31668 20256 31720 20262
rect 31668 20198 31720 20204
rect 31680 20058 31708 20198
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31576 18896 31628 18902
rect 31576 18838 31628 18844
rect 31574 16144 31630 16153
rect 31574 16079 31576 16088
rect 31628 16079 31630 16088
rect 31576 16050 31628 16056
rect 31576 15904 31628 15910
rect 31576 15846 31628 15852
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31484 15700 31536 15706
rect 31484 15642 31536 15648
rect 31588 15502 31616 15846
rect 31668 15632 31720 15638
rect 31668 15574 31720 15580
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31576 15496 31628 15502
rect 31576 15438 31628 15444
rect 31300 15360 31352 15366
rect 31298 15328 31300 15337
rect 31352 15328 31354 15337
rect 31298 15263 31354 15272
rect 31220 12406 31340 12434
rect 30932 11824 30984 11830
rect 30932 11766 30984 11772
rect 30840 11008 30892 11014
rect 30840 10950 30892 10956
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30196 9920 30248 9926
rect 30196 9862 30248 9868
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30392 9654 30420 9862
rect 30380 9648 30432 9654
rect 30380 9590 30432 9596
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 29920 9376 29972 9382
rect 29920 9318 29972 9324
rect 29920 8832 29972 8838
rect 29920 8774 29972 8780
rect 29828 8560 29880 8566
rect 29828 8502 29880 8508
rect 29828 8424 29880 8430
rect 29826 8392 29828 8401
rect 29880 8392 29882 8401
rect 29826 8327 29882 8336
rect 29736 8016 29788 8022
rect 29736 7958 29788 7964
rect 29932 7954 29960 8774
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29932 7410 29960 7890
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 30024 6882 30052 9522
rect 30104 9376 30156 9382
rect 30104 9318 30156 9324
rect 30116 8498 30144 9318
rect 30196 8900 30248 8906
rect 30196 8842 30248 8848
rect 30208 8498 30236 8842
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30288 8560 30340 8566
rect 30288 8502 30340 8508
rect 30104 8492 30156 8498
rect 30104 8434 30156 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30196 7812 30248 7818
rect 30196 7754 30248 7760
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 7410 30144 7686
rect 30104 7404 30156 7410
rect 30104 7346 30156 7352
rect 30208 7041 30236 7754
rect 30300 7410 30328 8502
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 30392 7546 30420 7958
rect 30484 7954 30512 8570
rect 30562 7984 30618 7993
rect 30472 7948 30524 7954
rect 30562 7919 30618 7928
rect 30472 7890 30524 7896
rect 30380 7540 30432 7546
rect 30380 7482 30432 7488
rect 30288 7404 30340 7410
rect 30288 7346 30340 7352
rect 30576 7313 30604 7919
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30562 7304 30618 7313
rect 30562 7239 30618 7248
rect 30194 7032 30250 7041
rect 30194 6967 30250 6976
rect 29932 6866 30052 6882
rect 29920 6860 30052 6866
rect 29972 6854 30052 6860
rect 29920 6802 29972 6808
rect 30208 6458 30236 6967
rect 30576 6662 30604 7239
rect 30668 7002 30696 7686
rect 30760 7546 30788 9998
rect 30944 9994 30972 11766
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31114 11520 31170 11529
rect 31114 11455 31170 11464
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 31036 10266 31064 10610
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 30932 9988 30984 9994
rect 30932 9930 30984 9936
rect 31128 9926 31156 11455
rect 31220 10198 31248 11698
rect 31312 10742 31340 12406
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 31208 10192 31260 10198
rect 31208 10134 31260 10140
rect 31208 10056 31260 10062
rect 31206 10024 31208 10033
rect 31260 10024 31262 10033
rect 31206 9959 31262 9968
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 31220 8974 31248 9959
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 30944 8022 30972 8434
rect 31220 8362 31248 8570
rect 31208 8356 31260 8362
rect 31208 8298 31260 8304
rect 31024 8288 31076 8294
rect 31024 8230 31076 8236
rect 30932 8016 30984 8022
rect 30932 7958 30984 7964
rect 30840 7812 30892 7818
rect 30840 7754 30892 7760
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 30656 6996 30708 7002
rect 30656 6938 30708 6944
rect 30852 6866 30880 7754
rect 30944 7478 30972 7958
rect 31036 7886 31064 8230
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 30932 7472 30984 7478
rect 30932 7414 30984 7420
rect 30944 6866 30972 7414
rect 31036 7342 31064 7822
rect 31312 7478 31340 10678
rect 31404 10130 31432 15438
rect 31496 15314 31524 15438
rect 31680 15314 31708 15574
rect 31496 15286 31708 15314
rect 31484 14816 31536 14822
rect 31484 14758 31536 14764
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31496 14414 31524 14758
rect 31588 14550 31616 14758
rect 31576 14544 31628 14550
rect 31576 14486 31628 14492
rect 31484 14408 31536 14414
rect 31484 14350 31536 14356
rect 31680 14226 31708 15286
rect 31772 15094 31800 20878
rect 31852 20256 31904 20262
rect 31850 20224 31852 20233
rect 31904 20224 31906 20233
rect 31850 20159 31906 20168
rect 31852 16516 31904 16522
rect 31852 16458 31904 16464
rect 31864 15910 31892 16458
rect 31956 16250 31984 24074
rect 32048 23526 32076 25191
rect 32140 24818 32168 25316
rect 32218 25120 32274 25129
rect 32218 25055 32274 25064
rect 32128 24812 32180 24818
rect 32128 24754 32180 24760
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 32036 23520 32088 23526
rect 32036 23462 32088 23468
rect 32034 23352 32090 23361
rect 32034 23287 32090 23296
rect 32048 23254 32076 23287
rect 32036 23248 32088 23254
rect 32036 23190 32088 23196
rect 32048 22030 32076 23190
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32036 21344 32088 21350
rect 32036 21286 32088 21292
rect 32048 17202 32076 21286
rect 32140 20874 32168 24550
rect 32232 22574 32260 25055
rect 32324 24818 32352 25910
rect 32416 25362 32444 26182
rect 32496 26036 32548 26042
rect 32496 25978 32548 25984
rect 32508 25770 32536 25978
rect 32496 25764 32548 25770
rect 32496 25706 32548 25712
rect 32404 25356 32456 25362
rect 32404 25298 32456 25304
rect 32496 25288 32548 25294
rect 32600 25265 32628 26998
rect 32876 26874 32904 28358
rect 32968 27878 32996 30194
rect 33060 29510 33088 31282
rect 33336 31142 33364 32506
rect 34428 32360 34480 32366
rect 34428 32302 34480 32308
rect 34060 32224 34112 32230
rect 34060 32166 34112 32172
rect 33416 31884 33468 31890
rect 33416 31826 33468 31832
rect 33428 31482 33456 31826
rect 33968 31680 34020 31686
rect 33968 31622 34020 31628
rect 33416 31476 33468 31482
rect 33416 31418 33468 31424
rect 33980 31346 34008 31622
rect 34072 31414 34100 32166
rect 34336 31748 34388 31754
rect 34336 31690 34388 31696
rect 34060 31408 34112 31414
rect 34060 31350 34112 31356
rect 33876 31340 33928 31346
rect 33876 31282 33928 31288
rect 33968 31340 34020 31346
rect 33968 31282 34020 31288
rect 33324 31136 33376 31142
rect 33324 31078 33376 31084
rect 33232 30592 33284 30598
rect 33232 30534 33284 30540
rect 33244 30297 33272 30534
rect 33600 30320 33652 30326
rect 33230 30288 33286 30297
rect 33600 30262 33652 30268
rect 33230 30223 33286 30232
rect 33416 30252 33468 30258
rect 33048 29504 33100 29510
rect 33048 29446 33100 29452
rect 33060 29306 33180 29322
rect 33048 29300 33180 29306
rect 33100 29294 33180 29300
rect 33048 29242 33100 29248
rect 33048 28960 33100 28966
rect 33048 28902 33100 28908
rect 33060 28121 33088 28902
rect 33152 28801 33180 29294
rect 33244 29034 33272 30223
rect 33468 30212 33548 30240
rect 33416 30194 33468 30200
rect 33520 29889 33548 30212
rect 33506 29880 33562 29889
rect 33506 29815 33562 29824
rect 33414 29336 33470 29345
rect 33414 29271 33470 29280
rect 33428 29238 33456 29271
rect 33416 29232 33468 29238
rect 33416 29174 33468 29180
rect 33324 29096 33376 29102
rect 33324 29038 33376 29044
rect 33232 29028 33284 29034
rect 33232 28970 33284 28976
rect 33138 28792 33194 28801
rect 33138 28727 33194 28736
rect 33232 28756 33284 28762
rect 33336 28744 33364 29038
rect 33284 28716 33364 28744
rect 33232 28698 33284 28704
rect 33140 28688 33192 28694
rect 33140 28630 33192 28636
rect 33152 28393 33180 28630
rect 33244 28558 33272 28698
rect 33520 28642 33548 29815
rect 33612 29481 33640 30262
rect 33692 30252 33744 30258
rect 33692 30194 33744 30200
rect 33704 29850 33732 30194
rect 33692 29844 33744 29850
rect 33692 29786 33744 29792
rect 33784 29572 33836 29578
rect 33784 29514 33836 29520
rect 33598 29472 33654 29481
rect 33598 29407 33654 29416
rect 33796 29170 33824 29514
rect 33784 29164 33836 29170
rect 33784 29106 33836 29112
rect 33336 28614 33548 28642
rect 33600 28688 33652 28694
rect 33600 28630 33652 28636
rect 33690 28656 33746 28665
rect 33232 28552 33284 28558
rect 33232 28494 33284 28500
rect 33138 28384 33194 28393
rect 33138 28319 33194 28328
rect 33046 28112 33102 28121
rect 33046 28047 33102 28056
rect 33244 28014 33272 28494
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 32956 27872 33008 27878
rect 32956 27814 33008 27820
rect 33140 27872 33192 27878
rect 33140 27814 33192 27820
rect 32692 26846 32904 26874
rect 32692 25770 32720 26846
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32772 26580 32824 26586
rect 32772 26522 32824 26528
rect 32680 25764 32732 25770
rect 32680 25706 32732 25712
rect 32496 25230 32548 25236
rect 32586 25256 32642 25265
rect 32404 25220 32456 25226
rect 32404 25162 32456 25168
rect 32416 24993 32444 25162
rect 32402 24984 32458 24993
rect 32508 24954 32536 25230
rect 32784 25242 32812 26522
rect 32876 26382 32904 26726
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 32864 25764 32916 25770
rect 32864 25706 32916 25712
rect 32586 25191 32642 25200
rect 32692 25214 32812 25242
rect 32402 24919 32458 24928
rect 32496 24948 32548 24954
rect 32496 24890 32548 24896
rect 32494 24848 32550 24857
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32404 24812 32456 24818
rect 32494 24783 32550 24792
rect 32588 24812 32640 24818
rect 32404 24754 32456 24760
rect 32324 23730 32352 24754
rect 32416 24614 32444 24754
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32508 24206 32536 24783
rect 32588 24754 32640 24760
rect 32600 24614 32628 24754
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 32600 24138 32628 24550
rect 32588 24132 32640 24138
rect 32588 24074 32640 24080
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32588 23520 32640 23526
rect 32588 23462 32640 23468
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32324 22681 32352 23054
rect 32496 23044 32548 23050
rect 32496 22986 32548 22992
rect 32310 22672 32366 22681
rect 32310 22607 32366 22616
rect 32220 22568 32272 22574
rect 32220 22510 32272 22516
rect 32232 22234 32260 22510
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32310 22128 32366 22137
rect 32310 22063 32366 22072
rect 32128 20868 32180 20874
rect 32128 20810 32180 20816
rect 32324 20466 32352 22063
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 32416 20346 32444 22374
rect 32324 20318 32444 20346
rect 32128 19508 32180 19514
rect 32128 19450 32180 19456
rect 32036 17196 32088 17202
rect 32036 17138 32088 17144
rect 32036 17060 32088 17066
rect 32036 17002 32088 17008
rect 31944 16244 31996 16250
rect 31944 16186 31996 16192
rect 31852 15904 31904 15910
rect 31852 15846 31904 15852
rect 31760 15088 31812 15094
rect 31760 15030 31812 15036
rect 31680 14198 31800 14226
rect 31772 13734 31800 14198
rect 31760 13728 31812 13734
rect 31760 13670 31812 13676
rect 31588 13530 31800 13546
rect 31576 13524 31812 13530
rect 31628 13518 31760 13524
rect 31576 13466 31628 13472
rect 31760 13466 31812 13472
rect 31864 13394 31892 15846
rect 31944 14816 31996 14822
rect 31944 14758 31996 14764
rect 31956 14550 31984 14758
rect 31944 14544 31996 14550
rect 31944 14486 31996 14492
rect 31944 13864 31996 13870
rect 31944 13806 31996 13812
rect 31852 13388 31904 13394
rect 31852 13330 31904 13336
rect 31956 13326 31984 13806
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31668 13252 31720 13258
rect 31668 13194 31720 13200
rect 31680 12434 31708 13194
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31588 12406 31708 12434
rect 31484 12096 31536 12102
rect 31484 12038 31536 12044
rect 31496 11898 31524 12038
rect 31484 11892 31536 11898
rect 31484 11834 31536 11840
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31404 9042 31432 10066
rect 31484 9920 31536 9926
rect 31484 9862 31536 9868
rect 31392 9036 31444 9042
rect 31392 8978 31444 8984
rect 31392 8492 31444 8498
rect 31392 8434 31444 8440
rect 31404 7954 31432 8434
rect 31496 8430 31524 9862
rect 31588 9178 31616 12406
rect 31666 12336 31722 12345
rect 31666 12271 31722 12280
rect 31680 10062 31708 12271
rect 31772 11762 31800 12786
rect 32048 12102 32076 17002
rect 32140 14804 32168 19450
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32232 14958 32260 18702
rect 32324 17921 32352 20318
rect 32404 20256 32456 20262
rect 32404 20198 32456 20204
rect 32416 19417 32444 20198
rect 32402 19408 32458 19417
rect 32402 19343 32458 19352
rect 32508 19242 32536 22986
rect 32600 20262 32628 23462
rect 32692 21010 32720 25214
rect 32876 24970 32904 25706
rect 32968 25158 32996 27814
rect 33152 27538 33180 27814
rect 33140 27532 33192 27538
rect 33140 27474 33192 27480
rect 33140 27056 33192 27062
rect 33140 26998 33192 27004
rect 33336 27010 33364 28614
rect 33416 28552 33468 28558
rect 33468 28512 33548 28540
rect 33416 28494 33468 28500
rect 33416 28416 33468 28422
rect 33416 28358 33468 28364
rect 33428 28257 33456 28358
rect 33414 28248 33470 28257
rect 33414 28183 33470 28192
rect 33416 28144 33468 28150
rect 33520 28132 33548 28512
rect 33468 28104 33548 28132
rect 33416 28086 33468 28092
rect 33520 27946 33548 28104
rect 33508 27940 33560 27946
rect 33508 27882 33560 27888
rect 33612 27334 33640 28630
rect 33690 28591 33746 28600
rect 33704 28404 33732 28591
rect 33796 28558 33824 29106
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33704 28376 33824 28404
rect 33888 28393 33916 31282
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 34348 31226 34376 31690
rect 34440 31414 34468 32302
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34520 31884 34572 31890
rect 34520 31826 34572 31832
rect 34428 31408 34480 31414
rect 34428 31350 34480 31356
rect 34532 31346 34560 31826
rect 34704 31680 34756 31686
rect 34704 31622 34756 31628
rect 34716 31482 34744 31622
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34704 31476 34756 31482
rect 34704 31418 34756 31424
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34164 30190 34192 31214
rect 34348 31198 34468 31226
rect 34440 31142 34468 31198
rect 34428 31136 34480 31142
rect 34428 31078 34480 31084
rect 34336 30932 34388 30938
rect 34336 30874 34388 30880
rect 34152 30184 34204 30190
rect 34152 30126 34204 30132
rect 34060 29504 34112 29510
rect 34060 29446 34112 29452
rect 33968 28756 34020 28762
rect 33968 28698 34020 28704
rect 33692 28076 33744 28082
rect 33692 28018 33744 28024
rect 33704 27713 33732 28018
rect 33690 27704 33746 27713
rect 33690 27639 33746 27648
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33048 26784 33100 26790
rect 33048 26726 33100 26732
rect 33060 26450 33088 26726
rect 33152 26450 33180 26998
rect 33232 26988 33284 26994
rect 33336 26982 33548 27010
rect 33612 26994 33640 27270
rect 33690 27024 33746 27033
rect 33232 26930 33284 26936
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33140 26444 33192 26450
rect 33140 26386 33192 26392
rect 33244 26042 33272 26930
rect 33324 26376 33376 26382
rect 33324 26318 33376 26324
rect 33232 26036 33284 26042
rect 33232 25978 33284 25984
rect 33046 25936 33102 25945
rect 33046 25871 33102 25880
rect 33140 25900 33192 25906
rect 33060 25838 33088 25871
rect 33140 25842 33192 25848
rect 33048 25832 33100 25838
rect 33152 25809 33180 25842
rect 33048 25774 33100 25780
rect 33138 25800 33194 25809
rect 33138 25735 33194 25744
rect 33048 25492 33100 25498
rect 33048 25434 33100 25440
rect 32956 25152 33008 25158
rect 32956 25094 33008 25100
rect 32876 24942 32996 24970
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32770 24304 32826 24313
rect 32876 24274 32904 24754
rect 32770 24239 32826 24248
rect 32864 24268 32916 24274
rect 32784 24206 32812 24239
rect 32864 24210 32916 24216
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 32772 24064 32824 24070
rect 32824 24024 32904 24052
rect 32772 24006 32824 24012
rect 32876 22642 32904 24024
rect 32968 22982 32996 24942
rect 33060 24426 33088 25434
rect 33152 24954 33180 25735
rect 33244 25498 33272 25978
rect 33336 25906 33364 26318
rect 33324 25900 33376 25906
rect 33324 25842 33376 25848
rect 33416 25764 33468 25770
rect 33416 25706 33468 25712
rect 33322 25664 33378 25673
rect 33322 25599 33378 25608
rect 33232 25492 33284 25498
rect 33232 25434 33284 25440
rect 33232 25152 33284 25158
rect 33232 25094 33284 25100
rect 33140 24948 33192 24954
rect 33140 24890 33192 24896
rect 33244 24614 33272 25094
rect 33336 24818 33364 25599
rect 33428 25537 33456 25706
rect 33414 25528 33470 25537
rect 33414 25463 33470 25472
rect 33416 25424 33468 25430
rect 33416 25366 33468 25372
rect 33428 25129 33456 25366
rect 33414 25120 33470 25129
rect 33414 25055 33470 25064
rect 33324 24812 33376 24818
rect 33324 24754 33376 24760
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 33060 24398 33180 24426
rect 33048 24336 33100 24342
rect 33048 24278 33100 24284
rect 33060 23050 33088 24278
rect 33048 23044 33100 23050
rect 33048 22986 33100 22992
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32968 22817 32996 22918
rect 32954 22808 33010 22817
rect 32954 22743 33010 22752
rect 32956 22704 33008 22710
rect 32956 22646 33008 22652
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 32772 22228 32824 22234
rect 32772 22170 32824 22176
rect 32680 21004 32732 21010
rect 32680 20946 32732 20952
rect 32588 20256 32640 20262
rect 32588 20198 32640 20204
rect 32680 19780 32732 19786
rect 32680 19722 32732 19728
rect 32496 19236 32548 19242
rect 32496 19178 32548 19184
rect 32404 18828 32456 18834
rect 32404 18770 32456 18776
rect 32416 18193 32444 18770
rect 32692 18766 32720 19722
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32402 18184 32458 18193
rect 32402 18119 32458 18128
rect 32310 17912 32366 17921
rect 32310 17847 32366 17856
rect 32312 17604 32364 17610
rect 32312 17546 32364 17552
rect 32324 17202 32352 17546
rect 32312 17196 32364 17202
rect 32312 17138 32364 17144
rect 32404 16652 32456 16658
rect 32404 16594 32456 16600
rect 32220 14952 32272 14958
rect 32220 14894 32272 14900
rect 32416 14822 32444 16594
rect 32508 16454 32536 18702
rect 32784 16998 32812 22170
rect 32876 21350 32904 22578
rect 32864 21344 32916 21350
rect 32864 21286 32916 21292
rect 32864 20800 32916 20806
rect 32862 20768 32864 20777
rect 32916 20768 32918 20777
rect 32862 20703 32918 20712
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32876 18970 32904 20402
rect 32968 20097 32996 22646
rect 33060 22642 33088 22986
rect 33048 22636 33100 22642
rect 33048 22578 33100 22584
rect 33152 22234 33180 24398
rect 33324 24404 33376 24410
rect 33324 24346 33376 24352
rect 33336 23866 33364 24346
rect 33416 24132 33468 24138
rect 33416 24074 33468 24080
rect 33324 23860 33376 23866
rect 33324 23802 33376 23808
rect 33428 23594 33456 24074
rect 33520 24052 33548 26982
rect 33600 26988 33652 26994
rect 33690 26959 33746 26968
rect 33600 26930 33652 26936
rect 33612 26586 33640 26930
rect 33600 26580 33652 26586
rect 33600 26522 33652 26528
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33612 26042 33640 26318
rect 33600 26036 33652 26042
rect 33600 25978 33652 25984
rect 33600 25832 33652 25838
rect 33600 25774 33652 25780
rect 33612 24970 33640 25774
rect 33704 25673 33732 26959
rect 33796 26568 33824 28376
rect 33874 28384 33930 28393
rect 33874 28319 33930 28328
rect 33876 28212 33928 28218
rect 33876 28154 33928 28160
rect 33888 27849 33916 28154
rect 33980 27878 34008 28698
rect 34072 28626 34100 29446
rect 34164 29102 34192 30126
rect 34348 29510 34376 30874
rect 34440 30666 34468 31078
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34428 30660 34480 30666
rect 34428 30602 34480 30608
rect 34440 30054 34468 30602
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 36084 30252 36136 30258
rect 36084 30194 36136 30200
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34704 29776 34756 29782
rect 34704 29718 34756 29724
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34336 29504 34388 29510
rect 34336 29446 34388 29452
rect 34532 29306 34560 29582
rect 34520 29300 34572 29306
rect 34520 29242 34572 29248
rect 34152 29096 34204 29102
rect 34152 29038 34204 29044
rect 34428 29096 34480 29102
rect 34428 29038 34480 29044
rect 34060 28620 34112 28626
rect 34060 28562 34112 28568
rect 33968 27872 34020 27878
rect 33874 27840 33930 27849
rect 33968 27814 34020 27820
rect 33874 27775 33930 27784
rect 33980 27674 34008 27814
rect 33968 27668 34020 27674
rect 33968 27610 34020 27616
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 34072 26858 34100 27406
rect 33968 26852 34020 26858
rect 33968 26794 34020 26800
rect 34060 26852 34112 26858
rect 34060 26794 34112 26800
rect 33876 26580 33928 26586
rect 33796 26540 33876 26568
rect 33876 26522 33928 26528
rect 33876 26376 33928 26382
rect 33782 26344 33838 26353
rect 33876 26318 33928 26324
rect 33782 26279 33838 26288
rect 33690 25664 33746 25673
rect 33690 25599 33746 25608
rect 33692 25424 33744 25430
rect 33692 25366 33744 25372
rect 33704 25294 33732 25366
rect 33796 25294 33824 26279
rect 33692 25288 33744 25294
rect 33690 25256 33692 25265
rect 33784 25288 33836 25294
rect 33744 25256 33746 25265
rect 33784 25230 33836 25236
rect 33690 25191 33746 25200
rect 33796 25106 33824 25230
rect 33888 25226 33916 26318
rect 33980 25974 34008 26794
rect 34072 26518 34100 26794
rect 34060 26512 34112 26518
rect 34060 26454 34112 26460
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 33968 25968 34020 25974
rect 33968 25910 34020 25916
rect 34072 25906 34100 26318
rect 34060 25900 34112 25906
rect 34060 25842 34112 25848
rect 33968 25832 34020 25838
rect 33968 25774 34020 25780
rect 33876 25220 33928 25226
rect 33876 25162 33928 25168
rect 33796 25078 33916 25106
rect 33612 24942 33824 24970
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33600 24064 33652 24070
rect 33520 24024 33600 24052
rect 33600 24006 33652 24012
rect 33612 23662 33640 24006
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 33232 23588 33284 23594
rect 33232 23530 33284 23536
rect 33416 23588 33468 23594
rect 33416 23530 33468 23536
rect 33244 23322 33272 23530
rect 33232 23316 33284 23322
rect 33232 23258 33284 23264
rect 33244 22642 33272 23258
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 33508 22432 33560 22438
rect 33508 22374 33560 22380
rect 33140 22228 33192 22234
rect 33140 22170 33192 22176
rect 33416 21412 33468 21418
rect 33416 21354 33468 21360
rect 33428 21146 33456 21354
rect 33416 21140 33468 21146
rect 33416 21082 33468 21088
rect 33416 21004 33468 21010
rect 33416 20946 33468 20952
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 33152 20330 33180 20810
rect 33244 20534 33272 20878
rect 33322 20632 33378 20641
rect 33322 20567 33378 20576
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 33230 20360 33286 20369
rect 33140 20324 33192 20330
rect 33230 20295 33286 20304
rect 33140 20266 33192 20272
rect 32954 20088 33010 20097
rect 32954 20023 33010 20032
rect 33048 19236 33100 19242
rect 33048 19178 33100 19184
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 32956 18964 33008 18970
rect 32956 18906 33008 18912
rect 32588 16992 32640 16998
rect 32588 16934 32640 16940
rect 32680 16992 32732 16998
rect 32680 16934 32732 16940
rect 32772 16992 32824 16998
rect 32772 16934 32824 16940
rect 32600 16794 32628 16934
rect 32588 16788 32640 16794
rect 32588 16730 32640 16736
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32586 16280 32642 16289
rect 32586 16215 32642 16224
rect 32600 15026 32628 16215
rect 32496 15020 32548 15026
rect 32496 14962 32548 14968
rect 32588 15020 32640 15026
rect 32588 14962 32640 14968
rect 32404 14816 32456 14822
rect 32140 14776 32260 14804
rect 32128 14272 32180 14278
rect 32128 14214 32180 14220
rect 32140 14006 32168 14214
rect 32128 14000 32180 14006
rect 32128 13942 32180 13948
rect 32128 13184 32180 13190
rect 32128 13126 32180 13132
rect 32140 12238 32168 13126
rect 32232 12442 32260 14776
rect 32404 14758 32456 14764
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32220 12436 32272 12442
rect 32220 12378 32272 12384
rect 32128 12232 32180 12238
rect 32128 12174 32180 12180
rect 32036 12096 32088 12102
rect 32036 12038 32088 12044
rect 32036 11892 32088 11898
rect 32036 11834 32088 11840
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 31668 10056 31720 10062
rect 31772 10033 31800 11698
rect 31668 9998 31720 10004
rect 31758 10024 31814 10033
rect 31758 9959 31814 9968
rect 32048 9722 32076 11834
rect 32324 10470 32352 12922
rect 32416 11694 32444 14758
rect 32508 14618 32536 14962
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32508 12986 32536 13262
rect 32496 12980 32548 12986
rect 32496 12922 32548 12928
rect 32692 12238 32720 16934
rect 32968 16590 32996 18906
rect 32956 16584 33008 16590
rect 32956 16526 33008 16532
rect 32956 16448 33008 16454
rect 33060 16436 33088 19178
rect 33244 17338 33272 20295
rect 33232 17332 33284 17338
rect 33232 17274 33284 17280
rect 33232 16516 33284 16522
rect 33232 16458 33284 16464
rect 33008 16408 33088 16436
rect 32956 16390 33008 16396
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 32784 12434 32812 16186
rect 32864 15428 32916 15434
rect 32864 15370 32916 15376
rect 32876 12646 32904 15370
rect 32968 15162 32996 16390
rect 33244 15502 33272 16458
rect 33336 16046 33364 20567
rect 33428 17610 33456 20946
rect 33520 18834 33548 22374
rect 33704 21078 33732 24754
rect 33796 24410 33824 24942
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33888 24313 33916 25078
rect 33980 24818 34008 25774
rect 34060 25696 34112 25702
rect 34060 25638 34112 25644
rect 34072 25362 34100 25638
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 34164 24818 34192 29038
rect 34336 28416 34388 28422
rect 34334 28384 34336 28393
rect 34388 28384 34390 28393
rect 34334 28319 34390 28328
rect 34336 27872 34388 27878
rect 34336 27814 34388 27820
rect 34348 27690 34376 27814
rect 34256 27674 34376 27690
rect 34440 27674 34468 29038
rect 34624 28626 34652 29582
rect 34612 28620 34664 28626
rect 34612 28562 34664 28568
rect 34624 28082 34652 28562
rect 34716 28558 34744 29718
rect 35624 29640 35676 29646
rect 35622 29608 35624 29617
rect 35676 29608 35678 29617
rect 35622 29543 35678 29552
rect 36096 29510 36124 30194
rect 36084 29504 36136 29510
rect 36084 29446 36136 29452
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35348 29300 35400 29306
rect 35348 29242 35400 29248
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 34808 28558 34836 28902
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34704 28552 34756 28558
rect 34704 28494 34756 28500
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 34980 28552 35032 28558
rect 34980 28494 35032 28500
rect 35072 28552 35124 28558
rect 35072 28494 35124 28500
rect 35256 28552 35308 28558
rect 35360 28540 35388 29242
rect 36096 29238 36124 29446
rect 36084 29232 36136 29238
rect 36084 29174 36136 29180
rect 36176 29096 36228 29102
rect 36176 29038 36228 29044
rect 36188 28994 36216 29038
rect 35308 28512 35388 28540
rect 36096 28966 36216 28994
rect 35256 28494 35308 28500
rect 34612 28076 34664 28082
rect 34612 28018 34664 28024
rect 34256 27668 34388 27674
rect 34256 27662 34336 27668
rect 34256 27062 34284 27662
rect 34336 27610 34388 27616
rect 34428 27668 34480 27674
rect 34428 27610 34480 27616
rect 34336 27532 34388 27538
rect 34336 27474 34388 27480
rect 34348 27334 34376 27474
rect 34336 27328 34388 27334
rect 34336 27270 34388 27276
rect 34244 27056 34296 27062
rect 34244 26998 34296 27004
rect 34256 26382 34284 26998
rect 34336 26988 34388 26994
rect 34336 26930 34388 26936
rect 34428 26988 34480 26994
rect 34428 26930 34480 26936
rect 34348 26586 34376 26930
rect 34336 26580 34388 26586
rect 34336 26522 34388 26528
rect 34244 26376 34296 26382
rect 34244 26318 34296 26324
rect 34334 26072 34390 26081
rect 34334 26007 34390 26016
rect 34244 25900 34296 25906
rect 34244 25842 34296 25848
rect 34256 25809 34284 25842
rect 34242 25800 34298 25809
rect 34242 25735 34298 25744
rect 34244 25696 34296 25702
rect 34244 25638 34296 25644
rect 34256 25498 34284 25638
rect 34348 25498 34376 26007
rect 34440 25770 34468 26930
rect 34518 26888 34574 26897
rect 34518 26823 34574 26832
rect 34532 26518 34560 26823
rect 34520 26512 34572 26518
rect 34520 26454 34572 26460
rect 34532 26042 34560 26454
rect 34612 26308 34664 26314
rect 34612 26250 34664 26256
rect 34520 26036 34572 26042
rect 34520 25978 34572 25984
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34428 25764 34480 25770
rect 34428 25706 34480 25712
rect 34244 25492 34296 25498
rect 34244 25434 34296 25440
rect 34336 25492 34388 25498
rect 34336 25434 34388 25440
rect 34532 25430 34560 25842
rect 34520 25424 34572 25430
rect 34520 25366 34572 25372
rect 33968 24812 34020 24818
rect 33968 24754 34020 24760
rect 34152 24812 34204 24818
rect 34152 24754 34204 24760
rect 33874 24304 33930 24313
rect 33874 24239 33876 24248
rect 33928 24239 33930 24248
rect 33876 24210 33928 24216
rect 33784 24132 33836 24138
rect 33784 24074 33836 24080
rect 33876 24132 33928 24138
rect 33876 24074 33928 24080
rect 33796 23730 33824 24074
rect 33784 23724 33836 23730
rect 33784 23666 33836 23672
rect 33692 21072 33744 21078
rect 33692 21014 33744 21020
rect 33796 21010 33824 23666
rect 33888 23662 33916 24074
rect 33876 23656 33928 23662
rect 33876 23598 33928 23604
rect 33980 23594 34008 24754
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34060 24608 34112 24614
rect 34060 24550 34112 24556
rect 33968 23588 34020 23594
rect 33968 23530 34020 23536
rect 33876 23520 33928 23526
rect 34072 23497 34100 24550
rect 34440 24410 34468 24686
rect 34624 24614 34652 26250
rect 34612 24608 34664 24614
rect 34612 24550 34664 24556
rect 34428 24404 34480 24410
rect 34428 24346 34480 24352
rect 34624 24138 34652 24550
rect 34612 24132 34664 24138
rect 34612 24074 34664 24080
rect 34244 24064 34296 24070
rect 34244 24006 34296 24012
rect 33876 23462 33928 23468
rect 34058 23488 34114 23497
rect 33784 21004 33836 21010
rect 33784 20946 33836 20952
rect 33600 20800 33652 20806
rect 33600 20742 33652 20748
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 33416 17604 33468 17610
rect 33416 17546 33468 17552
rect 33508 17332 33560 17338
rect 33508 17274 33560 17280
rect 33416 17128 33468 17134
rect 33416 17070 33468 17076
rect 33428 16794 33456 17070
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 33324 16040 33376 16046
rect 33428 16017 33456 16730
rect 33324 15982 33376 15988
rect 33414 16008 33470 16017
rect 33414 15943 33470 15952
rect 33324 15700 33376 15706
rect 33324 15642 33376 15648
rect 33048 15496 33100 15502
rect 33232 15496 33284 15502
rect 33100 15444 33180 15450
rect 33048 15438 33180 15444
rect 33232 15438 33284 15444
rect 33060 15422 33180 15438
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 32956 15156 33008 15162
rect 32956 15098 33008 15104
rect 32956 14068 33008 14074
rect 32956 14010 33008 14016
rect 32864 12640 32916 12646
rect 32864 12582 32916 12588
rect 32784 12406 32904 12434
rect 32496 12232 32548 12238
rect 32496 12174 32548 12180
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32404 11688 32456 11694
rect 32404 11630 32456 11636
rect 32508 11558 32536 12174
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32772 12096 32824 12102
rect 32772 12038 32824 12044
rect 32496 11552 32548 11558
rect 32496 11494 32548 11500
rect 32404 11076 32456 11082
rect 32404 11018 32456 11024
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31680 8809 31708 8910
rect 31666 8800 31722 8809
rect 31666 8735 31722 8744
rect 31484 8424 31536 8430
rect 31484 8366 31536 8372
rect 31576 8356 31628 8362
rect 31576 8298 31628 8304
rect 31392 7948 31444 7954
rect 31392 7890 31444 7896
rect 31300 7472 31352 7478
rect 31300 7414 31352 7420
rect 31404 7410 31432 7890
rect 31588 7410 31616 8298
rect 31680 7750 31708 8735
rect 31760 8628 31812 8634
rect 31760 8570 31812 8576
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31576 7404 31628 7410
rect 31576 7346 31628 7352
rect 31024 7336 31076 7342
rect 31024 7278 31076 7284
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31022 6896 31078 6905
rect 30840 6860 30892 6866
rect 30840 6802 30892 6808
rect 30932 6860 30984 6866
rect 31312 6866 31340 7278
rect 31022 6831 31078 6840
rect 31300 6860 31352 6866
rect 30932 6802 30984 6808
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 29920 6248 29972 6254
rect 29920 6190 29972 6196
rect 29644 5908 29696 5914
rect 29644 5850 29696 5856
rect 28264 5772 28316 5778
rect 28264 5714 28316 5720
rect 29932 5710 29960 6190
rect 29920 5704 29972 5710
rect 29920 5646 29972 5652
rect 31036 5642 31064 6831
rect 31300 6802 31352 6808
rect 31772 6662 31800 8570
rect 31944 8016 31996 8022
rect 31944 7958 31996 7964
rect 31956 7886 31984 7958
rect 31944 7880 31996 7886
rect 31944 7822 31996 7828
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 32128 6656 32180 6662
rect 32128 6598 32180 6604
rect 32140 6118 32168 6598
rect 32128 6112 32180 6118
rect 32128 6054 32180 6060
rect 32416 5642 32444 11018
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 32508 8838 32536 8978
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 32600 7002 32628 12038
rect 32680 11552 32732 11558
rect 32680 11494 32732 11500
rect 32692 11150 32720 11494
rect 32680 11144 32732 11150
rect 32680 11086 32732 11092
rect 32678 9616 32734 9625
rect 32678 9551 32734 9560
rect 32692 9178 32720 9551
rect 32680 9172 32732 9178
rect 32680 9114 32732 9120
rect 32680 8832 32732 8838
rect 32680 8774 32732 8780
rect 32692 8498 32720 8774
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32692 7954 32720 8434
rect 32680 7948 32732 7954
rect 32680 7890 32732 7896
rect 32588 6996 32640 7002
rect 32588 6938 32640 6944
rect 32784 6254 32812 12038
rect 32876 9625 32904 12406
rect 32968 12238 32996 14010
rect 33060 13462 33088 15302
rect 33152 13462 33180 15422
rect 33244 15094 33272 15438
rect 33232 15088 33284 15094
rect 33232 15030 33284 15036
rect 33048 13456 33100 13462
rect 33048 13398 33100 13404
rect 33140 13456 33192 13462
rect 33140 13398 33192 13404
rect 33060 13258 33088 13398
rect 33048 13252 33100 13258
rect 33048 13194 33100 13200
rect 33140 12436 33192 12442
rect 33336 12434 33364 15642
rect 33428 15162 33456 15943
rect 33416 15156 33468 15162
rect 33416 15098 33468 15104
rect 33520 15042 33548 17274
rect 33428 15014 33548 15042
rect 33428 12986 33456 15014
rect 33508 14816 33560 14822
rect 33508 14758 33560 14764
rect 33416 12980 33468 12986
rect 33416 12922 33468 12928
rect 33520 12434 33548 14758
rect 33612 13938 33640 20742
rect 33888 20618 33916 23462
rect 34058 23423 34114 23432
rect 33968 22432 34020 22438
rect 33968 22374 34020 22380
rect 33796 20590 33916 20618
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33704 20330 33732 20402
rect 33692 20324 33744 20330
rect 33692 20266 33744 20272
rect 33704 15502 33732 20266
rect 33796 15570 33824 20590
rect 33876 20460 33928 20466
rect 33980 20448 34008 22374
rect 34256 22094 34284 24006
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34428 22976 34480 22982
rect 34428 22918 34480 22924
rect 34440 22778 34468 22918
rect 34428 22772 34480 22778
rect 34428 22714 34480 22720
rect 34336 22704 34388 22710
rect 34532 22658 34560 23802
rect 34388 22652 34560 22658
rect 34336 22646 34560 22652
rect 34348 22630 34560 22646
rect 34256 22066 34468 22094
rect 34244 21004 34296 21010
rect 34244 20946 34296 20952
rect 33928 20420 34008 20448
rect 33876 20402 33928 20408
rect 33784 15564 33836 15570
rect 33784 15506 33836 15512
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33796 15026 33824 15506
rect 33784 15020 33836 15026
rect 33784 14962 33836 14968
rect 33600 13932 33652 13938
rect 33600 13874 33652 13880
rect 33612 13138 33640 13874
rect 33888 13326 33916 20402
rect 34152 18828 34204 18834
rect 34152 18770 34204 18776
rect 33968 18624 34020 18630
rect 33968 18566 34020 18572
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 33612 13110 33916 13138
rect 33692 12980 33744 12986
rect 33692 12922 33744 12928
rect 33336 12406 33456 12434
rect 33520 12406 33640 12434
rect 33140 12378 33192 12384
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32968 11082 32996 12174
rect 33046 11792 33102 11801
rect 33046 11727 33102 11736
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32862 9616 32918 9625
rect 33060 9586 33088 11727
rect 33152 10810 33180 12378
rect 33322 11792 33378 11801
rect 33428 11762 33456 12406
rect 33612 11762 33640 12406
rect 33704 11898 33732 12922
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33322 11727 33324 11736
rect 33376 11727 33378 11736
rect 33416 11756 33468 11762
rect 33324 11698 33376 11704
rect 33416 11698 33468 11704
rect 33508 11756 33560 11762
rect 33508 11698 33560 11704
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 33692 11756 33744 11762
rect 33692 11698 33744 11704
rect 33232 11008 33284 11014
rect 33232 10950 33284 10956
rect 33140 10804 33192 10810
rect 33140 10746 33192 10752
rect 33244 9674 33272 10950
rect 33152 9646 33272 9674
rect 33152 9586 33180 9646
rect 32862 9551 32864 9560
rect 32916 9551 32918 9560
rect 33048 9580 33100 9586
rect 32864 9522 32916 9528
rect 33048 9522 33100 9528
rect 33140 9580 33192 9586
rect 33140 9522 33192 9528
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 33060 9058 33088 9522
rect 32876 9030 33088 9058
rect 32876 8906 32904 9030
rect 33152 8974 33180 9522
rect 33244 9450 33272 9522
rect 33232 9444 33284 9450
rect 33232 9386 33284 9392
rect 33244 9353 33272 9386
rect 33336 9382 33364 9522
rect 33324 9376 33376 9382
rect 33230 9344 33286 9353
rect 33324 9318 33376 9324
rect 33230 9279 33286 9288
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 32864 8900 32916 8906
rect 32864 8842 32916 8848
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33060 8362 33088 8774
rect 33428 8634 33456 11698
rect 33520 11014 33548 11698
rect 33508 11008 33560 11014
rect 33508 10950 33560 10956
rect 33612 10826 33640 11698
rect 33704 11354 33732 11698
rect 33888 11558 33916 13110
rect 33980 11762 34008 18566
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 34072 17270 34100 17478
rect 34060 17264 34112 17270
rect 34060 17206 34112 17212
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 33876 11552 33928 11558
rect 33876 11494 33928 11500
rect 33968 11552 34020 11558
rect 33968 11494 34020 11500
rect 33796 11354 33824 11494
rect 33692 11348 33744 11354
rect 33692 11290 33744 11296
rect 33784 11348 33836 11354
rect 33784 11290 33836 11296
rect 33692 11144 33744 11150
rect 33692 11086 33744 11092
rect 33520 10798 33640 10826
rect 33520 9586 33548 10798
rect 33704 10674 33732 11086
rect 33692 10668 33744 10674
rect 33692 10610 33744 10616
rect 33704 9722 33732 10610
rect 33692 9716 33744 9722
rect 33692 9658 33744 9664
rect 33508 9580 33560 9586
rect 33508 9522 33560 9528
rect 33600 9580 33652 9586
rect 33600 9522 33652 9528
rect 33612 9178 33640 9522
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33876 9104 33928 9110
rect 33876 9046 33928 9052
rect 33508 8900 33560 8906
rect 33508 8842 33560 8848
rect 33416 8628 33468 8634
rect 33416 8570 33468 8576
rect 33520 8498 33548 8842
rect 33888 8634 33916 9046
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 33508 8492 33560 8498
rect 33508 8434 33560 8440
rect 32864 8356 32916 8362
rect 32864 8298 32916 8304
rect 33048 8356 33100 8362
rect 33048 8298 33100 8304
rect 32876 7886 32904 8298
rect 33060 8022 33088 8298
rect 33520 8294 33548 8434
rect 33508 8288 33560 8294
rect 33508 8230 33560 8236
rect 33048 8016 33100 8022
rect 33048 7958 33100 7964
rect 33520 7886 33548 8230
rect 33888 7954 33916 8570
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32864 7880 32916 7886
rect 32864 7822 32916 7828
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33980 7478 34008 11494
rect 34072 10577 34100 17206
rect 34164 17202 34192 18770
rect 34256 18086 34284 20946
rect 34440 20466 34468 22066
rect 34532 21010 34560 22630
rect 34612 22500 34664 22506
rect 34612 22442 34664 22448
rect 34624 22098 34652 22442
rect 34612 22092 34664 22098
rect 34612 22034 34664 22040
rect 34520 21004 34572 21010
rect 34520 20946 34572 20952
rect 34520 20868 34572 20874
rect 34520 20810 34572 20816
rect 34428 20460 34480 20466
rect 34348 20420 34428 20448
rect 34244 18080 34296 18086
rect 34244 18022 34296 18028
rect 34152 17196 34204 17202
rect 34152 17138 34204 17144
rect 34164 16522 34192 17138
rect 34152 16516 34204 16522
rect 34152 16458 34204 16464
rect 34256 16130 34284 18022
rect 34348 16726 34376 20420
rect 34428 20402 34480 20408
rect 34428 19712 34480 19718
rect 34428 19654 34480 19660
rect 34440 18834 34468 19654
rect 34532 19174 34560 20810
rect 34520 19168 34572 19174
rect 34520 19110 34572 19116
rect 34428 18828 34480 18834
rect 34428 18770 34480 18776
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34426 18184 34482 18193
rect 34426 18119 34482 18128
rect 34440 17898 34468 18119
rect 34532 18057 34560 18566
rect 34518 18048 34574 18057
rect 34518 17983 34574 17992
rect 34440 17870 34560 17898
rect 34532 17218 34560 17870
rect 34440 17190 34560 17218
rect 34336 16720 34388 16726
rect 34336 16662 34388 16668
rect 34440 16538 34468 17190
rect 34624 16590 34652 22034
rect 34716 20890 34744 28494
rect 34992 28082 35020 28494
rect 35084 28121 35112 28494
rect 35070 28112 35126 28121
rect 34980 28076 35032 28082
rect 35268 28082 35296 28494
rect 35440 28484 35492 28490
rect 35440 28426 35492 28432
rect 35070 28047 35072 28056
rect 34980 28018 35032 28024
rect 35124 28047 35126 28056
rect 35256 28076 35308 28082
rect 35072 28018 35124 28024
rect 35256 28018 35308 28024
rect 34992 27946 35020 28018
rect 34980 27940 35032 27946
rect 34980 27882 35032 27888
rect 35084 27860 35112 28018
rect 35452 27985 35480 28426
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35532 28076 35584 28082
rect 35532 28018 35584 28024
rect 35438 27976 35494 27985
rect 35438 27911 35494 27920
rect 35544 27860 35572 28018
rect 35084 27832 35388 27860
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35360 27674 35388 27832
rect 35452 27832 35572 27860
rect 35348 27668 35400 27674
rect 35348 27610 35400 27616
rect 35254 27568 35310 27577
rect 35254 27503 35310 27512
rect 35268 27470 35296 27503
rect 35256 27464 35308 27470
rect 35256 27406 35308 27412
rect 35348 27464 35400 27470
rect 35348 27406 35400 27412
rect 35256 27328 35308 27334
rect 35256 27270 35308 27276
rect 35072 27056 35124 27062
rect 35070 27024 35072 27033
rect 35124 27024 35126 27033
rect 34796 26988 34848 26994
rect 35070 26959 35126 26968
rect 34796 26930 34848 26936
rect 34808 26858 34836 26930
rect 34796 26852 34848 26858
rect 34796 26794 34848 26800
rect 34808 26450 34836 26794
rect 35268 26738 35296 27270
rect 35360 27062 35388 27406
rect 35452 27112 35480 27832
rect 36096 27577 36124 28966
rect 36176 28076 36228 28082
rect 36176 28018 36228 28024
rect 36082 27568 36138 27577
rect 36082 27503 36138 27512
rect 35992 27464 36044 27470
rect 35992 27406 36044 27412
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35452 27084 35664 27112
rect 35348 27056 35400 27062
rect 35348 26998 35400 27004
rect 35532 26988 35584 26994
rect 35532 26930 35584 26936
rect 35268 26710 35480 26738
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 35164 26444 35216 26450
rect 35164 26386 35216 26392
rect 35072 26240 35124 26246
rect 35176 26217 35204 26386
rect 35256 26376 35308 26382
rect 35256 26318 35308 26324
rect 35072 26182 35124 26188
rect 35162 26208 35218 26217
rect 35084 25974 35112 26182
rect 35162 26143 35218 26152
rect 35072 25968 35124 25974
rect 35072 25910 35124 25916
rect 35176 25770 35204 26143
rect 35268 25906 35296 26318
rect 35348 26240 35400 26246
rect 35348 26182 35400 26188
rect 35256 25900 35308 25906
rect 35256 25842 35308 25848
rect 35360 25838 35388 26182
rect 35348 25832 35400 25838
rect 35348 25774 35400 25780
rect 35164 25764 35216 25770
rect 35164 25706 35216 25712
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34808 25294 34836 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 25498 35388 25774
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 35162 25392 35218 25401
rect 35162 25327 35218 25336
rect 34796 25288 34848 25294
rect 34796 25230 34848 25236
rect 35176 24886 35204 25327
rect 35256 25288 35308 25294
rect 35256 25230 35308 25236
rect 35268 24954 35296 25230
rect 35348 25220 35400 25226
rect 35348 25162 35400 25168
rect 35256 24948 35308 24954
rect 35256 24890 35308 24896
rect 35164 24880 35216 24886
rect 35164 24822 35216 24828
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35164 24404 35216 24410
rect 35164 24346 35216 24352
rect 34796 24200 34848 24206
rect 34980 24200 35032 24206
rect 34796 24142 34848 24148
rect 34978 24168 34980 24177
rect 35032 24168 35034 24177
rect 34808 23322 34836 24142
rect 34978 24103 35034 24112
rect 35176 23526 35204 24346
rect 35256 24200 35308 24206
rect 35256 24142 35308 24148
rect 35268 23866 35296 24142
rect 35360 24070 35388 25162
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 35256 23860 35308 23866
rect 35256 23802 35308 23808
rect 35360 23730 35388 24006
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 35164 23520 35216 23526
rect 35164 23462 35216 23468
rect 35348 23520 35400 23526
rect 35348 23462 35400 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 23316 34848 23322
rect 34848 23276 34928 23304
rect 34796 23258 34848 23264
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34808 21010 34836 22918
rect 34900 22642 34928 23276
rect 35256 23112 35308 23118
rect 35254 23080 35256 23089
rect 35308 23080 35310 23089
rect 35072 23044 35124 23050
rect 35254 23015 35310 23024
rect 35072 22986 35124 22992
rect 34888 22636 34940 22642
rect 34888 22578 34940 22584
rect 35084 22545 35112 22986
rect 35360 22642 35388 23462
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 35070 22536 35126 22545
rect 35070 22471 35126 22480
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35360 21350 35388 22578
rect 35348 21344 35400 21350
rect 35348 21286 35400 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35452 21162 35480 26710
rect 35544 26246 35572 26930
rect 35636 26314 35664 27084
rect 35716 26988 35768 26994
rect 35716 26930 35768 26936
rect 35728 26353 35756 26930
rect 36004 26790 36032 27406
rect 36084 27396 36136 27402
rect 36084 27338 36136 27344
rect 36096 26994 36124 27338
rect 36188 27305 36216 28018
rect 36268 27464 36320 27470
rect 36268 27406 36320 27412
rect 36174 27296 36230 27305
rect 36174 27231 36230 27240
rect 36084 26988 36136 26994
rect 36084 26930 36136 26936
rect 35992 26784 36044 26790
rect 35992 26726 36044 26732
rect 36280 26625 36308 27406
rect 36266 26616 36322 26625
rect 36266 26551 36322 26560
rect 36176 26376 36228 26382
rect 35714 26344 35770 26353
rect 35624 26308 35676 26314
rect 36176 26318 36228 26324
rect 35714 26279 35770 26288
rect 35624 26250 35676 26256
rect 35532 26240 35584 26246
rect 35532 26182 35584 26188
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35624 25968 35676 25974
rect 36188 25945 36216 26318
rect 36360 26308 36412 26314
rect 36360 26250 36412 26256
rect 35624 25910 35676 25916
rect 36174 25936 36230 25945
rect 35532 25764 35584 25770
rect 35532 25706 35584 25712
rect 35544 25498 35572 25706
rect 35532 25492 35584 25498
rect 35532 25434 35584 25440
rect 35636 25294 35664 25910
rect 35716 25900 35768 25906
rect 36174 25871 36230 25880
rect 35716 25842 35768 25848
rect 35728 25430 35756 25842
rect 35806 25528 35862 25537
rect 35806 25463 35862 25472
rect 35820 25430 35848 25463
rect 35716 25424 35768 25430
rect 35716 25366 35768 25372
rect 35808 25424 35860 25430
rect 35808 25366 35860 25372
rect 35624 25288 35676 25294
rect 35716 25288 35768 25294
rect 35624 25230 35676 25236
rect 35714 25256 35716 25265
rect 35992 25288 36044 25294
rect 35768 25256 35770 25265
rect 35992 25230 36044 25236
rect 35714 25191 35770 25200
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35808 24948 35860 24954
rect 35808 24890 35860 24896
rect 35820 24410 35848 24890
rect 35808 24404 35860 24410
rect 35808 24346 35860 24352
rect 35530 24168 35586 24177
rect 35530 24103 35532 24112
rect 35584 24103 35586 24112
rect 35532 24074 35584 24080
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 36004 22094 36032 25230
rect 36266 24848 36322 24857
rect 36266 24783 36322 24792
rect 36176 24744 36228 24750
rect 36176 24686 36228 24692
rect 36082 24576 36138 24585
rect 36082 24511 36138 24520
rect 36096 24206 36124 24511
rect 36188 24274 36216 24686
rect 36176 24268 36228 24274
rect 36176 24210 36228 24216
rect 36084 24200 36136 24206
rect 36084 24142 36136 24148
rect 36176 23724 36228 23730
rect 36176 23666 36228 23672
rect 36188 23225 36216 23666
rect 36174 23216 36230 23225
rect 36174 23151 36230 23160
rect 36176 22568 36228 22574
rect 36174 22536 36176 22545
rect 36228 22536 36230 22545
rect 36174 22471 36230 22480
rect 36176 22228 36228 22234
rect 36176 22170 36228 22176
rect 36004 22066 36124 22094
rect 35992 22024 36044 22030
rect 35992 21966 36044 21972
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 35544 21185 35572 21490
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35268 21134 35480 21162
rect 35530 21176 35586 21185
rect 34796 21004 34848 21010
rect 34796 20946 34848 20952
rect 34980 20936 35032 20942
rect 34978 20904 34980 20913
rect 35032 20904 35034 20913
rect 34716 20862 34836 20890
rect 34704 20800 34756 20806
rect 34702 20768 34704 20777
rect 34756 20768 34758 20777
rect 34702 20703 34758 20712
rect 34808 20466 34836 20862
rect 34978 20839 35034 20848
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 34704 20256 34756 20262
rect 34704 20198 34756 20204
rect 34716 19854 34744 20198
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34716 18766 34744 18906
rect 34808 18850 34836 20402
rect 35268 20398 35296 21134
rect 35530 21111 35586 21120
rect 35348 21004 35400 21010
rect 35348 20946 35400 20952
rect 35256 20392 35308 20398
rect 35256 20334 35308 20340
rect 35360 20262 35388 20946
rect 35728 20942 35756 21286
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 35440 20800 35492 20806
rect 35440 20742 35492 20748
rect 35348 20256 35400 20262
rect 35348 20198 35400 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35348 20052 35400 20058
rect 35348 19994 35400 20000
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34808 18822 34928 18850
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34612 16584 34664 16590
rect 34440 16510 34560 16538
rect 34612 16526 34664 16532
rect 34532 16250 34560 16510
rect 34716 16402 34744 18702
rect 34808 17270 34836 18822
rect 34900 18766 34928 18822
rect 34888 18760 34940 18766
rect 34888 18702 34940 18708
rect 35072 18692 35124 18698
rect 35072 18634 35124 18640
rect 35084 18086 35112 18634
rect 35072 18080 35124 18086
rect 35072 18022 35124 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 35360 17082 35388 19994
rect 34624 16374 34744 16402
rect 34808 17054 35388 17082
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34256 16102 34560 16130
rect 34428 16040 34480 16046
rect 34428 15982 34480 15988
rect 34336 13320 34388 13326
rect 34336 13262 34388 13268
rect 34348 11626 34376 13262
rect 34440 11830 34468 15982
rect 34532 14550 34560 16102
rect 34520 14544 34572 14550
rect 34520 14486 34572 14492
rect 34520 13184 34572 13190
rect 34520 13126 34572 13132
rect 34532 12238 34560 13126
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 34428 11824 34480 11830
rect 34428 11766 34480 11772
rect 34624 11762 34652 16374
rect 34704 16244 34756 16250
rect 34704 16186 34756 16192
rect 34612 11756 34664 11762
rect 34612 11698 34664 11704
rect 34336 11620 34388 11626
rect 34336 11562 34388 11568
rect 34612 11620 34664 11626
rect 34612 11562 34664 11568
rect 34336 11280 34388 11286
rect 34336 11222 34388 11228
rect 34348 11121 34376 11222
rect 34624 11218 34652 11562
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 34334 11112 34390 11121
rect 34334 11047 34390 11056
rect 34348 10742 34376 11047
rect 34336 10736 34388 10742
rect 34336 10678 34388 10684
rect 34624 10674 34652 11154
rect 34716 10810 34744 16186
rect 34808 14958 34836 17054
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35254 16552 35310 16561
rect 35164 16516 35216 16522
rect 35254 16487 35256 16496
rect 35164 16458 35216 16464
rect 35308 16487 35310 16496
rect 35256 16458 35308 16464
rect 35176 15978 35204 16458
rect 35348 16448 35400 16454
rect 35348 16390 35400 16396
rect 35164 15972 35216 15978
rect 35164 15914 35216 15920
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35072 15020 35124 15026
rect 35072 14962 35124 14968
rect 34796 14952 34848 14958
rect 35084 14929 35112 14962
rect 34796 14894 34848 14900
rect 35070 14920 35126 14929
rect 35070 14855 35126 14864
rect 34796 14816 34848 14822
rect 34796 14758 34848 14764
rect 34808 13530 34836 14758
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 13524 34848 13530
rect 34796 13466 34848 13472
rect 35360 13394 35388 16390
rect 35452 13462 35480 20742
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35532 20392 35584 20398
rect 35532 20334 35584 20340
rect 35544 20058 35572 20334
rect 35532 20052 35584 20058
rect 35532 19994 35584 20000
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35440 13456 35492 13462
rect 35440 13398 35492 13404
rect 35348 13388 35400 13394
rect 35348 13330 35400 13336
rect 35360 13274 35388 13330
rect 35360 13246 35480 13274
rect 34796 13184 34848 13190
rect 34796 13126 34848 13132
rect 34808 11150 34836 13126
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35256 12164 35308 12170
rect 35256 12106 35308 12112
rect 34886 12064 34942 12073
rect 34886 11999 34942 12008
rect 34900 11830 34928 11999
rect 35268 11898 35296 12106
rect 35256 11892 35308 11898
rect 35256 11834 35308 11840
rect 34888 11824 34940 11830
rect 34888 11766 34940 11772
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34704 10804 34756 10810
rect 34704 10746 34756 10752
rect 34796 10736 34848 10742
rect 34796 10678 34848 10684
rect 34612 10668 34664 10674
rect 34612 10610 34664 10616
rect 34058 10568 34114 10577
rect 34058 10503 34114 10512
rect 34072 7818 34100 10503
rect 34336 9988 34388 9994
rect 34336 9930 34388 9936
rect 34348 9722 34376 9930
rect 34808 9722 34836 10678
rect 35452 10674 35480 13246
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35440 10668 35492 10674
rect 35440 10610 35492 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 34336 9716 34388 9722
rect 34336 9658 34388 9664
rect 34796 9716 34848 9722
rect 34796 9658 34848 9664
rect 34334 9616 34390 9625
rect 34334 9551 34336 9560
rect 34388 9551 34390 9560
rect 34336 9522 34388 9528
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 36004 8974 36032 21966
rect 35992 8968 36044 8974
rect 35992 8910 36044 8916
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34992 8634 35020 8774
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 34520 8560 34572 8566
rect 34520 8502 34572 8508
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34060 7812 34112 7818
rect 34060 7754 34112 7760
rect 34164 7546 34192 8434
rect 34244 8356 34296 8362
rect 34244 8298 34296 8304
rect 34256 8022 34284 8298
rect 34244 8016 34296 8022
rect 34244 7958 34296 7964
rect 34336 7880 34388 7886
rect 34336 7822 34388 7828
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 33968 7472 34020 7478
rect 33968 7414 34020 7420
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 33152 6866 33180 7278
rect 33140 6860 33192 6866
rect 33140 6802 33192 6808
rect 33152 6458 33180 6802
rect 33784 6724 33836 6730
rect 33784 6666 33836 6672
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 32772 6248 32824 6254
rect 32772 6190 32824 6196
rect 33152 5778 33180 6394
rect 33796 6390 33824 6666
rect 33784 6384 33836 6390
rect 33784 6326 33836 6332
rect 33796 6118 33824 6326
rect 33784 6112 33836 6118
rect 33784 6054 33836 6060
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33796 5642 33824 6054
rect 34164 5914 34192 7482
rect 34348 7478 34376 7822
rect 34428 7812 34480 7818
rect 34428 7754 34480 7760
rect 34336 7472 34388 7478
rect 34336 7414 34388 7420
rect 34348 6730 34376 7414
rect 34440 7002 34468 7754
rect 34428 6996 34480 7002
rect 34428 6938 34480 6944
rect 34336 6724 34388 6730
rect 34336 6666 34388 6672
rect 34532 6458 34560 8502
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 34808 7546 34836 8434
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 36096 7886 36124 22066
rect 36188 15638 36216 22170
rect 36176 15632 36228 15638
rect 36176 15574 36228 15580
rect 36176 15020 36228 15026
rect 36176 14962 36228 14968
rect 36188 12753 36216 14962
rect 36174 12744 36230 12753
rect 36174 12679 36230 12688
rect 36188 10470 36216 12679
rect 36176 10464 36228 10470
rect 36176 10406 36228 10412
rect 36280 9926 36308 24783
rect 36372 24342 36400 26250
rect 36544 25492 36596 25498
rect 36544 25434 36596 25440
rect 36360 24336 36412 24342
rect 36360 24278 36412 24284
rect 36450 23624 36506 23633
rect 36450 23559 36506 23568
rect 36464 17542 36492 23559
rect 36452 17536 36504 17542
rect 36452 17478 36504 17484
rect 36556 17354 36584 25434
rect 36726 21584 36782 21593
rect 36726 21519 36782 21528
rect 36634 18320 36690 18329
rect 36634 18255 36690 18264
rect 36372 17326 36584 17354
rect 36268 9920 36320 9926
rect 36268 9862 36320 9868
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 34520 6452 34572 6458
rect 34520 6394 34572 6400
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34152 5908 34204 5914
rect 34152 5850 34204 5856
rect 31024 5636 31076 5642
rect 31024 5578 31076 5584
rect 32404 5636 32456 5642
rect 32404 5578 32456 5584
rect 33784 5636 33836 5642
rect 33784 5578 33836 5584
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 26700 4820 26752 4826
rect 26700 4762 26752 4768
rect 27344 4480 27396 4486
rect 27344 4422 27396 4428
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26620 3602 26648 3878
rect 26712 3670 26740 3878
rect 27356 3738 27384 4422
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 36096 3738 36124 7822
rect 36372 6662 36400 17326
rect 36452 17196 36504 17202
rect 36452 17138 36504 17144
rect 36360 6656 36412 6662
rect 36360 6598 36412 6604
rect 36464 4146 36492 17138
rect 36648 17082 36676 18255
rect 36556 17054 36676 17082
rect 36556 8090 36584 17054
rect 36544 8084 36596 8090
rect 36544 8026 36596 8032
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 36740 3942 36768 21519
rect 36728 3936 36780 3942
rect 36728 3878 36780 3884
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 36084 3732 36136 3738
rect 36084 3674 36136 3680
rect 26700 3664 26752 3670
rect 26700 3606 26752 3612
rect 26608 3596 26660 3602
rect 26608 3538 26660 3544
rect 27356 3534 27384 3674
rect 27344 3528 27396 3534
rect 27344 3470 27396 3476
rect 36082 3496 36138 3505
rect 36082 3431 36084 3440
rect 36136 3431 36138 3440
rect 36084 3402 36136 3408
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 24952 2440 25004 2446
rect 24952 2382 25004 2388
rect 24504 800 24532 2382
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25148 800 25176 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 18 0 74 800
rect 662 0 718 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 2686 31320 2742 31376
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 8298 34604 8354 34640
rect 8298 34584 8300 34604
rect 8300 34584 8352 34604
rect 8352 34584 8354 34604
rect 8666 34468 8722 34504
rect 8666 34448 8668 34468
rect 8668 34448 8720 34468
rect 8720 34448 8722 34468
rect 10230 35264 10286 35320
rect 9770 34312 9826 34368
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 5170 30676 5172 30696
rect 5172 30676 5224 30696
rect 5224 30676 5226 30696
rect 5170 30640 5226 30676
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 3698 29280 3754 29336
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4342 29144 4398 29200
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4158 28076 4214 28112
rect 4158 28056 4160 28076
rect 4160 28056 4212 28076
rect 4212 28056 4214 28076
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4710 29144 4766 29200
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4986 28076 5042 28112
rect 4986 28056 4988 28076
rect 4988 28056 5040 28076
rect 5040 28056 5042 28076
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 3146 26968 3202 27024
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4066 22072 4122 22128
rect 4342 22092 4398 22128
rect 4342 22072 4344 22092
rect 4344 22072 4396 22092
rect 4396 22072 4398 22092
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 5078 21972 5080 21992
rect 5080 21972 5132 21992
rect 5132 21972 5134 21992
rect 5078 21936 5134 21972
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 5998 25916 6000 25936
rect 6000 25916 6052 25936
rect 6052 25916 6054 25936
rect 5998 25880 6054 25916
rect 6826 26868 6828 26888
rect 6828 26868 6880 26888
rect 6880 26868 6882 26888
rect 6826 26832 6882 26868
rect 5998 23704 6054 23760
rect 5722 21972 5724 21992
rect 5724 21972 5776 21992
rect 5776 21972 5778 21992
rect 5722 21936 5778 21972
rect 6458 23568 6514 23624
rect 4894 20848 4950 20904
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4526 19896 4582 19952
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 5722 21140 5778 21176
rect 5722 21120 5724 21140
rect 5724 21120 5776 21140
rect 5776 21120 5778 21140
rect 5722 20576 5778 20632
rect 5998 19896 6054 19952
rect 5262 16632 5318 16688
rect 4894 16496 4950 16552
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 5538 16496 5594 16552
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4802 13948 4804 13968
rect 4804 13948 4856 13968
rect 4856 13948 4858 13968
rect 4802 13912 4858 13948
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 6918 24248 6974 24304
rect 6826 24148 6828 24168
rect 6828 24148 6880 24168
rect 6880 24148 6882 24168
rect 6826 24112 6882 24148
rect 7286 22208 7342 22264
rect 8298 29280 8354 29336
rect 7838 25880 7894 25936
rect 9310 32292 9366 32328
rect 9310 32272 9312 32292
rect 9312 32272 9364 32292
rect 9364 32272 9366 32292
rect 10138 33224 10194 33280
rect 9310 31456 9366 31512
rect 9126 31320 9182 31376
rect 9494 31592 9550 31648
rect 9034 30776 9090 30832
rect 9770 31592 9826 31648
rect 9862 30640 9918 30696
rect 9126 29280 9182 29336
rect 8942 28872 8998 28928
rect 8850 26832 8906 26888
rect 7746 25100 7748 25120
rect 7748 25100 7800 25120
rect 7800 25100 7802 25120
rect 7746 25064 7802 25100
rect 7654 22652 7656 22672
rect 7656 22652 7708 22672
rect 7708 22652 7710 22672
rect 7654 22616 7710 22652
rect 7378 20848 7434 20904
rect 7470 20576 7526 20632
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 5906 10104 5962 10160
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 938 4120 994 4176
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 8482 25472 8538 25528
rect 8390 24792 8446 24848
rect 8758 26016 8814 26072
rect 8574 24112 8630 24168
rect 9218 25744 9274 25800
rect 8022 21140 8078 21176
rect 8022 21120 8024 21140
rect 8024 21120 8076 21140
rect 8076 21120 8078 21140
rect 8022 14900 8024 14920
rect 8024 14900 8076 14920
rect 8076 14900 8078 14920
rect 8022 14864 8078 14900
rect 9218 23604 9220 23624
rect 9220 23604 9272 23624
rect 9272 23604 9274 23624
rect 9218 23568 9274 23604
rect 9218 21548 9274 21584
rect 9586 29008 9642 29064
rect 9770 29552 9826 29608
rect 9678 28600 9734 28656
rect 9770 27512 9826 27568
rect 10690 34992 10746 35048
rect 12162 34992 12218 35048
rect 10598 31728 10654 31784
rect 10322 29588 10324 29608
rect 10324 29588 10376 29608
rect 10376 29588 10378 29608
rect 10322 29552 10378 29588
rect 10046 29008 10102 29064
rect 10230 28872 10286 28928
rect 10230 28636 10232 28656
rect 10232 28636 10284 28656
rect 10284 28636 10286 28656
rect 10230 28600 10286 28636
rect 10046 27240 10102 27296
rect 10046 27104 10102 27160
rect 9678 24812 9734 24848
rect 9954 26152 10010 26208
rect 9678 24792 9680 24812
rect 9680 24792 9732 24812
rect 9732 24792 9734 24812
rect 9678 23316 9734 23352
rect 9678 23296 9680 23316
rect 9680 23296 9732 23316
rect 9732 23296 9734 23316
rect 9218 21528 9220 21548
rect 9220 21528 9272 21548
rect 9272 21528 9274 21548
rect 10322 27648 10378 27704
rect 10506 31340 10562 31376
rect 10506 31320 10508 31340
rect 10508 31320 10560 31340
rect 10560 31320 10562 31340
rect 10874 32952 10930 33008
rect 12898 35828 12954 35864
rect 12898 35808 12900 35828
rect 12900 35808 12952 35828
rect 12952 35808 12954 35828
rect 12714 35400 12770 35456
rect 12622 35028 12624 35048
rect 12624 35028 12676 35048
rect 12676 35028 12678 35048
rect 12622 34992 12678 35028
rect 10782 31456 10838 31512
rect 10966 31728 11022 31784
rect 11242 30540 11244 30560
rect 11244 30540 11296 30560
rect 11296 30540 11298 30560
rect 11242 30504 11298 30540
rect 11702 30368 11758 30424
rect 11426 30232 11482 30288
rect 10138 26832 10194 26888
rect 10322 26832 10378 26888
rect 10138 24284 10140 24304
rect 10140 24284 10192 24304
rect 10192 24284 10194 24304
rect 10138 24248 10194 24284
rect 10046 23180 10102 23216
rect 10046 23160 10048 23180
rect 10048 23160 10100 23180
rect 10100 23160 10102 23180
rect 10322 23704 10378 23760
rect 10046 23044 10102 23080
rect 10046 23024 10048 23044
rect 10048 23024 10100 23044
rect 10100 23024 10102 23044
rect 9862 21392 9918 21448
rect 10046 20984 10102 21040
rect 9678 20032 9734 20088
rect 10690 29028 10746 29064
rect 10690 29008 10692 29028
rect 10692 29008 10744 29028
rect 10744 29008 10746 29028
rect 11518 28620 11574 28656
rect 11518 28600 11520 28620
rect 11520 28600 11572 28620
rect 11572 28600 11574 28620
rect 11794 29008 11850 29064
rect 10690 26832 10746 26888
rect 10966 27104 11022 27160
rect 11150 26832 11206 26888
rect 10966 26696 11022 26752
rect 10782 25472 10838 25528
rect 10782 23160 10838 23216
rect 11150 26696 11206 26752
rect 11058 26424 11114 26480
rect 10598 21548 10654 21584
rect 10598 21528 10600 21548
rect 10600 21528 10652 21548
rect 10652 21528 10654 21548
rect 10414 20868 10470 20904
rect 10414 20848 10416 20868
rect 10416 20848 10468 20868
rect 10468 20848 10470 20868
rect 10414 18844 10416 18864
rect 10416 18844 10468 18864
rect 10468 18844 10470 18864
rect 10414 18808 10470 18844
rect 9770 17992 9826 18048
rect 6090 10140 6092 10160
rect 6092 10140 6144 10160
rect 6144 10140 6146 10160
rect 6090 10104 6146 10140
rect 6734 10104 6790 10160
rect 6182 9444 6238 9480
rect 6182 9424 6184 9444
rect 6184 9424 6236 9444
rect 6236 9424 6238 9444
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 8942 16532 8944 16552
rect 8944 16532 8996 16552
rect 8996 16532 8998 16552
rect 8942 16496 8998 16532
rect 8758 15564 8814 15600
rect 8758 15544 8760 15564
rect 8760 15544 8812 15564
rect 8812 15544 8814 15564
rect 8942 12824 8998 12880
rect 8666 12708 8722 12744
rect 8666 12688 8668 12708
rect 8668 12688 8720 12708
rect 8720 12688 8722 12708
rect 8666 12416 8722 12472
rect 8574 12280 8630 12336
rect 9402 15564 9458 15600
rect 9402 15544 9404 15564
rect 9404 15544 9456 15564
rect 9456 15544 9458 15564
rect 9494 14864 9550 14920
rect 9770 13932 9826 13968
rect 9770 13912 9772 13932
rect 9772 13912 9824 13932
rect 9824 13912 9826 13932
rect 9218 12280 9274 12336
rect 11242 23060 11244 23080
rect 11244 23060 11296 23080
rect 11296 23060 11298 23080
rect 11242 23024 11298 23060
rect 11518 25472 11574 25528
rect 11610 25372 11612 25392
rect 11612 25372 11664 25392
rect 11664 25372 11666 25392
rect 11610 25336 11666 25372
rect 12070 31764 12072 31784
rect 12072 31764 12124 31784
rect 12124 31764 12126 31784
rect 12070 31728 12126 31764
rect 13082 33088 13138 33144
rect 12070 29416 12126 29472
rect 12622 29280 12678 29336
rect 12530 29008 12586 29064
rect 12438 28872 12494 28928
rect 12530 28636 12532 28656
rect 12532 28636 12584 28656
rect 12584 28636 12586 28656
rect 12530 28600 12586 28636
rect 12898 29416 12954 29472
rect 12990 29008 13046 29064
rect 12530 27512 12586 27568
rect 12622 26832 12678 26888
rect 12530 26560 12586 26616
rect 13634 35400 13690 35456
rect 14186 35672 14242 35728
rect 13726 31728 13782 31784
rect 15658 35672 15714 35728
rect 14738 35264 14794 35320
rect 12990 27104 13046 27160
rect 12806 26424 12862 26480
rect 12530 26016 12586 26072
rect 12070 25608 12126 25664
rect 11518 24112 11574 24168
rect 12346 25608 12402 25664
rect 11978 23196 11980 23216
rect 11980 23196 12032 23216
rect 12032 23196 12034 23216
rect 11978 23160 12034 23196
rect 11058 18672 11114 18728
rect 10966 18420 11022 18456
rect 10966 18400 10968 18420
rect 10968 18400 11020 18420
rect 11020 18400 11022 18420
rect 11150 17856 11206 17912
rect 10138 12844 10194 12880
rect 10138 12824 10140 12844
rect 10140 12824 10192 12844
rect 10192 12824 10194 12844
rect 8666 10124 8722 10160
rect 8666 10104 8668 10124
rect 8668 10104 8720 10124
rect 8720 10104 8722 10124
rect 9678 10124 9734 10160
rect 9678 10104 9680 10124
rect 9680 10104 9732 10124
rect 9732 10104 9734 10124
rect 10230 12316 10232 12336
rect 10232 12316 10284 12336
rect 10284 12316 10286 12336
rect 10230 12280 10286 12316
rect 12530 24520 12586 24576
rect 12346 23704 12402 23760
rect 11702 20304 11758 20360
rect 13266 27104 13322 27160
rect 13266 26324 13268 26344
rect 13268 26324 13320 26344
rect 13320 26324 13322 26344
rect 13266 26288 13322 26324
rect 13266 26188 13268 26208
rect 13268 26188 13320 26208
rect 13320 26188 13322 26208
rect 13266 26152 13322 26188
rect 12622 24248 12678 24304
rect 13634 27376 13690 27432
rect 13542 26988 13598 27024
rect 13542 26968 13544 26988
rect 13544 26968 13596 26988
rect 13596 26968 13598 26988
rect 13726 26560 13782 26616
rect 12530 19896 12586 19952
rect 11518 18672 11574 18728
rect 11334 16224 11390 16280
rect 11150 12552 11206 12608
rect 10230 10124 10286 10160
rect 10230 10104 10232 10124
rect 10232 10104 10284 10124
rect 10284 10104 10286 10124
rect 10782 10668 10838 10704
rect 11150 12316 11152 12336
rect 11152 12316 11204 12336
rect 11204 12316 11206 12336
rect 11150 12280 11206 12316
rect 11426 12552 11482 12608
rect 10782 10648 10784 10668
rect 10784 10648 10836 10668
rect 10836 10648 10838 10668
rect 11242 10004 11244 10024
rect 11244 10004 11296 10024
rect 11296 10004 11298 10024
rect 11242 9968 11298 10004
rect 11242 8084 11298 8120
rect 11242 8064 11244 8084
rect 11244 8064 11296 8084
rect 11296 8064 11298 8084
rect 11150 7928 11206 7984
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 11610 14864 11666 14920
rect 12254 19216 12310 19272
rect 13910 26988 13966 27024
rect 13910 26968 13912 26988
rect 13912 26968 13964 26988
rect 13964 26968 13966 26988
rect 13910 26324 13912 26344
rect 13912 26324 13964 26344
rect 13964 26324 13966 26344
rect 13910 26288 13966 26324
rect 14094 29164 14150 29200
rect 14094 29144 14096 29164
rect 14096 29144 14148 29164
rect 14148 29144 14150 29164
rect 14554 30796 14610 30832
rect 14554 30776 14556 30796
rect 14556 30776 14608 30796
rect 14608 30776 14610 30796
rect 14462 29008 14518 29064
rect 14094 27240 14150 27296
rect 13910 24520 13966 24576
rect 13818 23840 13874 23896
rect 12254 14884 12310 14920
rect 12254 14864 12256 14884
rect 12256 14864 12308 14884
rect 12308 14864 12310 14884
rect 12254 13912 12310 13968
rect 12162 12824 12218 12880
rect 11978 12416 12034 12472
rect 11610 10004 11612 10024
rect 11612 10004 11664 10024
rect 11664 10004 11666 10024
rect 11610 9968 11666 10004
rect 14370 26324 14372 26344
rect 14372 26324 14424 26344
rect 14424 26324 14426 26344
rect 14370 26288 14426 26324
rect 18234 35808 18290 35864
rect 14738 29552 14794 29608
rect 15014 29280 15070 29336
rect 14646 26424 14702 26480
rect 14646 24928 14702 24984
rect 14094 23568 14150 23624
rect 14646 23432 14702 23488
rect 14186 23160 14242 23216
rect 13634 17332 13690 17368
rect 13634 17312 13636 17332
rect 13636 17312 13688 17332
rect 13688 17312 13690 17332
rect 13634 17040 13690 17096
rect 13726 16632 13782 16688
rect 14186 19216 14242 19272
rect 14094 18708 14096 18728
rect 14096 18708 14148 18728
rect 14148 18708 14150 18728
rect 14094 18672 14150 18708
rect 13910 16224 13966 16280
rect 13726 16088 13782 16144
rect 11610 7384 11666 7440
rect 11794 7148 11796 7168
rect 11796 7148 11848 7168
rect 11848 7148 11850 7168
rect 11794 7112 11850 7148
rect 12070 7248 12126 7304
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 13174 13368 13230 13424
rect 12530 7404 12586 7440
rect 13818 14900 13820 14920
rect 13820 14900 13872 14920
rect 13872 14900 13874 14920
rect 13818 14864 13874 14900
rect 14094 14592 14150 14648
rect 12990 11192 13046 11248
rect 13726 11600 13782 11656
rect 13634 11328 13690 11384
rect 12898 10648 12954 10704
rect 12530 7384 12532 7404
rect 12532 7384 12584 7404
rect 12584 7384 12586 7404
rect 12254 7112 12310 7168
rect 13450 8084 13506 8120
rect 13450 8064 13452 8084
rect 13452 8064 13504 8084
rect 13504 8064 13506 8084
rect 14370 16088 14426 16144
rect 14278 14592 14334 14648
rect 14094 9560 14150 9616
rect 14002 9424 14058 9480
rect 14002 7248 14058 7304
rect 15014 27512 15070 27568
rect 15014 26696 15070 26752
rect 15014 21664 15070 21720
rect 15842 27648 15898 27704
rect 15658 24248 15714 24304
rect 16670 31884 16726 31920
rect 16670 31864 16672 31884
rect 16672 31864 16724 31884
rect 16724 31864 16726 31884
rect 16578 30368 16634 30424
rect 17314 32952 17370 33008
rect 17866 32852 17868 32872
rect 17868 32852 17920 32872
rect 17920 32852 17922 32872
rect 17866 32816 17922 32852
rect 17866 31900 17868 31920
rect 17868 31900 17920 31920
rect 17920 31900 17922 31920
rect 17866 31864 17922 31900
rect 18142 32716 18144 32736
rect 18144 32716 18196 32736
rect 18196 32716 18198 32736
rect 18142 32680 18198 32716
rect 18050 32272 18106 32328
rect 16118 28056 16174 28112
rect 16394 27276 16396 27296
rect 16396 27276 16448 27296
rect 16448 27276 16450 27296
rect 16394 27240 16450 27276
rect 16026 25744 16082 25800
rect 16394 25608 16450 25664
rect 15474 21528 15530 21584
rect 15198 19896 15254 19952
rect 14738 17992 14794 18048
rect 15382 17992 15438 18048
rect 14646 16224 14702 16280
rect 14646 14764 14648 14784
rect 14648 14764 14700 14784
rect 14700 14764 14702 14784
rect 14646 14728 14702 14764
rect 14738 13912 14794 13968
rect 16026 21256 16082 21312
rect 16210 21120 16266 21176
rect 16854 28620 16910 28656
rect 16854 28600 16856 28620
rect 16856 28600 16908 28620
rect 16908 28600 16910 28620
rect 16946 28484 17002 28520
rect 16946 28464 16948 28484
rect 16948 28464 17000 28484
rect 17000 28464 17002 28484
rect 16762 27648 16818 27704
rect 16854 27512 16910 27568
rect 16762 27412 16764 27432
rect 16764 27412 16816 27432
rect 16816 27412 16818 27432
rect 16762 27376 16818 27412
rect 16578 25472 16634 25528
rect 16854 25064 16910 25120
rect 17866 30368 17922 30424
rect 17498 30232 17554 30288
rect 17222 28328 17278 28384
rect 17222 27920 17278 27976
rect 17314 27240 17370 27296
rect 16762 23432 16818 23488
rect 17406 26152 17462 26208
rect 19062 34312 19118 34368
rect 19338 33804 19340 33824
rect 19340 33804 19392 33824
rect 19392 33804 19394 33824
rect 19338 33768 19394 33804
rect 19798 33768 19854 33824
rect 19430 33360 19486 33416
rect 19154 33088 19210 33144
rect 18694 32836 18750 32872
rect 18694 32816 18696 32836
rect 18696 32816 18748 32836
rect 18748 32816 18750 32836
rect 18878 32716 18880 32736
rect 18880 32716 18932 32736
rect 18932 32716 18934 32736
rect 18878 32680 18934 32716
rect 17774 28500 17776 28520
rect 17776 28500 17828 28520
rect 17828 28500 17830 28520
rect 17774 28464 17830 28500
rect 17682 28056 17738 28112
rect 18142 28192 18198 28248
rect 17958 28056 18014 28112
rect 17774 26152 17830 26208
rect 17958 23704 18014 23760
rect 18142 26696 18198 26752
rect 18142 25336 18198 25392
rect 17222 21548 17278 21584
rect 17222 21528 17224 21548
rect 17224 21528 17276 21548
rect 17276 21528 17278 21548
rect 17498 20868 17554 20904
rect 17498 20848 17500 20868
rect 17500 20848 17552 20868
rect 17552 20848 17554 20868
rect 17406 20168 17462 20224
rect 17590 19760 17646 19816
rect 15566 15136 15622 15192
rect 15750 15136 15806 15192
rect 15750 14048 15806 14104
rect 15014 9560 15070 9616
rect 14830 8472 14886 8528
rect 14830 7112 14886 7168
rect 15198 9172 15254 9208
rect 15198 9152 15200 9172
rect 15200 9152 15252 9172
rect 15252 9152 15254 9172
rect 15106 7656 15162 7712
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 16210 16496 16266 16552
rect 16762 17312 16818 17368
rect 17130 18828 17186 18864
rect 17130 18808 17132 18828
rect 17132 18808 17184 18828
rect 17184 18808 17186 18828
rect 16394 14728 16450 14784
rect 16578 13776 16634 13832
rect 16394 13640 16450 13696
rect 16210 10104 16266 10160
rect 15842 7928 15898 7984
rect 16486 11736 16542 11792
rect 16762 11192 16818 11248
rect 17222 16396 17224 16416
rect 17224 16396 17276 16416
rect 17276 16396 17278 16416
rect 17222 16360 17278 16396
rect 17590 16768 17646 16824
rect 17866 20848 17922 20904
rect 18970 27956 18972 27976
rect 18972 27956 19024 27976
rect 19024 27956 19026 27976
rect 18970 27920 19026 27956
rect 19706 28192 19762 28248
rect 19430 27240 19486 27296
rect 18234 21664 18290 21720
rect 18418 21800 18474 21856
rect 17958 20712 18014 20768
rect 17866 19080 17922 19136
rect 17958 18400 18014 18456
rect 17958 16516 18014 16552
rect 17958 16496 17960 16516
rect 17960 16496 18012 16516
rect 18012 16496 18014 16516
rect 16946 13640 17002 13696
rect 17038 12280 17094 12336
rect 16762 9968 16818 10024
rect 16762 9444 16818 9480
rect 16762 9424 16764 9444
rect 16764 9424 16816 9444
rect 16816 9424 16818 9444
rect 17130 11192 17186 11248
rect 17590 15544 17646 15600
rect 17314 13776 17370 13832
rect 17406 13504 17462 13560
rect 17590 14728 17646 14784
rect 17590 14356 17592 14376
rect 17592 14356 17644 14376
rect 17644 14356 17646 14376
rect 17590 14320 17646 14356
rect 18510 20304 18566 20360
rect 18142 19236 18198 19272
rect 18142 19216 18144 19236
rect 18144 19216 18196 19236
rect 18196 19216 18198 19236
rect 18142 16768 18198 16824
rect 18142 15564 18198 15600
rect 18142 15544 18144 15564
rect 18144 15544 18196 15564
rect 18196 15544 18198 15564
rect 18142 15272 18198 15328
rect 18050 15000 18106 15056
rect 18510 17040 18566 17096
rect 18234 15020 18290 15056
rect 18234 15000 18236 15020
rect 18236 15000 18288 15020
rect 18288 15000 18290 15020
rect 18418 15000 18474 15056
rect 18326 14356 18328 14376
rect 18328 14356 18380 14376
rect 18380 14356 18382 14376
rect 18326 14320 18382 14356
rect 17958 14184 18014 14240
rect 17406 12960 17462 13016
rect 17314 12008 17370 12064
rect 17222 10124 17278 10160
rect 17774 12688 17830 12744
rect 17222 10104 17224 10124
rect 17224 10104 17276 10124
rect 17276 10104 17278 10124
rect 17314 10004 17316 10024
rect 17316 10004 17368 10024
rect 17368 10004 17370 10024
rect 17314 9968 17370 10004
rect 18050 13524 18106 13560
rect 18050 13504 18052 13524
rect 18052 13504 18104 13524
rect 18104 13504 18106 13524
rect 18050 13388 18106 13424
rect 18050 13368 18052 13388
rect 18052 13368 18104 13388
rect 18104 13368 18106 13388
rect 18418 14048 18474 14104
rect 18326 13368 18382 13424
rect 18786 21120 18842 21176
rect 18970 24248 19026 24304
rect 19062 23976 19118 24032
rect 19522 24792 19578 24848
rect 19706 24792 19762 24848
rect 19982 26424 20038 26480
rect 19982 25780 19984 25800
rect 19984 25780 20036 25800
rect 20036 25780 20038 25800
rect 19982 25744 20038 25780
rect 19338 23468 19340 23488
rect 19340 23468 19392 23488
rect 19392 23468 19394 23488
rect 19338 23432 19394 23468
rect 19154 23160 19210 23216
rect 19246 23024 19302 23080
rect 19246 22208 19302 22264
rect 19614 23704 19670 23760
rect 19614 23568 19670 23624
rect 19430 23060 19432 23080
rect 19432 23060 19484 23080
rect 19484 23060 19486 23080
rect 19430 23024 19486 23060
rect 19430 21972 19432 21992
rect 19432 21972 19484 21992
rect 19484 21972 19486 21992
rect 19430 21936 19486 21972
rect 19430 21684 19486 21720
rect 19430 21664 19432 21684
rect 19432 21664 19484 21684
rect 19484 21664 19486 21684
rect 18786 20476 18788 20496
rect 18788 20476 18840 20496
rect 18840 20476 18842 20496
rect 18786 20440 18842 20476
rect 19246 21004 19302 21040
rect 19246 20984 19248 21004
rect 19248 20984 19300 21004
rect 19300 20984 19302 21004
rect 19430 21120 19486 21176
rect 19246 20848 19302 20904
rect 19154 20032 19210 20088
rect 19614 20984 19670 21040
rect 19338 19624 19394 19680
rect 18878 17720 18934 17776
rect 18878 17448 18934 17504
rect 19246 19252 19248 19272
rect 19248 19252 19300 19272
rect 19300 19252 19302 19272
rect 19246 19216 19302 19252
rect 19154 18400 19210 18456
rect 19614 20576 19670 20632
rect 19706 20168 19762 20224
rect 19798 19780 19854 19816
rect 19798 19760 19800 19780
rect 19800 19760 19852 19780
rect 19852 19760 19854 19780
rect 19430 18572 19432 18592
rect 19432 18572 19484 18592
rect 19484 18572 19486 18592
rect 19430 18536 19486 18572
rect 19246 16088 19302 16144
rect 18970 15544 19026 15600
rect 19062 15156 19118 15192
rect 19798 17720 19854 17776
rect 19062 15136 19064 15156
rect 19064 15136 19116 15156
rect 19116 15136 19118 15156
rect 18878 14456 18934 14512
rect 19062 14612 19118 14648
rect 19062 14592 19064 14612
rect 19064 14592 19116 14612
rect 19116 14592 19118 14612
rect 18786 14356 18788 14376
rect 18788 14356 18840 14376
rect 18840 14356 18842 14376
rect 18786 14320 18842 14356
rect 18786 14220 18788 14240
rect 18788 14220 18840 14240
rect 18840 14220 18842 14240
rect 18786 14184 18842 14220
rect 19338 14592 19394 14648
rect 19338 13912 19394 13968
rect 18878 13640 18934 13696
rect 18326 11464 18382 11520
rect 17682 10260 17738 10296
rect 17682 10240 17684 10260
rect 17684 10240 17736 10260
rect 17736 10240 17738 10260
rect 17866 9152 17922 9208
rect 17314 7404 17370 7440
rect 18142 9152 18198 9208
rect 19522 13232 19578 13288
rect 19430 13096 19486 13152
rect 19062 11872 19118 11928
rect 18602 9172 18658 9208
rect 18602 9152 18604 9172
rect 18604 9152 18656 9172
rect 18656 9152 18658 9172
rect 18878 10648 18934 10704
rect 18878 9288 18934 9344
rect 19246 11464 19302 11520
rect 19338 11212 19394 11248
rect 19338 11192 19340 11212
rect 19340 11192 19392 11212
rect 19392 11192 19394 11212
rect 19338 10376 19394 10432
rect 19706 16108 19762 16144
rect 19706 16088 19708 16108
rect 19708 16088 19760 16108
rect 19760 16088 19762 16108
rect 20166 24248 20222 24304
rect 20258 23432 20314 23488
rect 20166 21664 20222 21720
rect 20074 20204 20076 20224
rect 20076 20204 20128 20224
rect 20128 20204 20130 20224
rect 20074 20168 20130 20204
rect 20350 21800 20406 21856
rect 20626 26152 20682 26208
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 21362 33360 21418 33416
rect 21822 33380 21878 33416
rect 21822 33360 21824 33380
rect 21824 33360 21876 33380
rect 21876 33360 21878 33380
rect 22190 34448 22246 34504
rect 21362 30232 21418 30288
rect 21086 29008 21142 29064
rect 20902 28872 20958 28928
rect 21086 28192 21142 28248
rect 20810 27240 20866 27296
rect 20626 24928 20682 24984
rect 20902 24928 20958 24984
rect 20534 23976 20590 24032
rect 20442 21664 20498 21720
rect 20442 21292 20444 21312
rect 20444 21292 20496 21312
rect 20496 21292 20498 21312
rect 20442 21256 20498 21292
rect 21546 25880 21602 25936
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 22466 35692 22522 35728
rect 22466 35672 22468 35692
rect 22468 35672 22520 35692
rect 22520 35672 22522 35692
rect 23018 35692 23074 35728
rect 23018 35672 23020 35692
rect 23020 35672 23072 35692
rect 23072 35672 23074 35692
rect 22282 32000 22338 32056
rect 22466 32000 22522 32056
rect 22190 31728 22246 31784
rect 22834 33360 22890 33416
rect 23018 32428 23074 32464
rect 23018 32408 23020 32428
rect 23020 32408 23072 32428
rect 23072 32408 23074 32428
rect 22926 32000 22982 32056
rect 21822 29960 21878 30016
rect 21914 29008 21970 29064
rect 21730 28620 21786 28656
rect 21730 28600 21732 28620
rect 21732 28600 21784 28620
rect 21784 28600 21786 28620
rect 22190 29044 22192 29064
rect 22192 29044 22244 29064
rect 22244 29044 22246 29064
rect 22190 29008 22246 29044
rect 21914 26696 21970 26752
rect 21730 24828 21732 24848
rect 21732 24828 21784 24848
rect 21784 24828 21786 24848
rect 21730 24792 21786 24828
rect 21730 24692 21732 24712
rect 21732 24692 21784 24712
rect 21784 24692 21786 24712
rect 21730 24656 21786 24692
rect 21362 23568 21418 23624
rect 20626 20304 20682 20360
rect 20074 17176 20130 17232
rect 20534 18400 20590 18456
rect 20534 17312 20590 17368
rect 20166 16532 20168 16552
rect 20168 16532 20220 16552
rect 20220 16532 20222 16552
rect 20166 16496 20222 16532
rect 20166 16088 20222 16144
rect 19798 15444 19800 15464
rect 19800 15444 19852 15464
rect 19852 15444 19854 15464
rect 19798 15408 19854 15444
rect 20534 16396 20536 16416
rect 20536 16396 20588 16416
rect 20588 16396 20590 16416
rect 20534 16360 20590 16396
rect 20534 15816 20590 15872
rect 20258 15544 20314 15600
rect 19982 14612 20038 14648
rect 19982 14592 19984 14612
rect 19984 14592 20036 14612
rect 20036 14592 20038 14612
rect 19798 14184 19854 14240
rect 20074 14184 20130 14240
rect 19890 13676 19935 13696
rect 19935 13676 19946 13696
rect 19890 13640 19946 13676
rect 20258 14456 20314 14512
rect 20258 14184 20314 14240
rect 19706 12688 19762 12744
rect 19798 12164 19854 12200
rect 19798 12144 19800 12164
rect 19800 12144 19852 12164
rect 19852 12144 19854 12164
rect 19522 9696 19578 9752
rect 19246 9016 19302 9072
rect 19154 8200 19210 8256
rect 17314 7384 17316 7404
rect 17316 7384 17368 7404
rect 17368 7384 17370 7404
rect 19338 8492 19394 8528
rect 19338 8472 19340 8492
rect 19340 8472 19392 8492
rect 19392 8472 19394 8492
rect 20166 13096 20222 13152
rect 19890 11192 19946 11248
rect 20350 11464 20406 11520
rect 20350 11056 20406 11112
rect 20074 10240 20130 10296
rect 20258 10376 20314 10432
rect 19522 8356 19578 8392
rect 19522 8336 19524 8356
rect 19524 8336 19576 8356
rect 19576 8336 19578 8356
rect 19338 7948 19394 7984
rect 19338 7928 19340 7948
rect 19340 7928 19392 7948
rect 19392 7928 19394 7948
rect 20166 9988 20222 10024
rect 20166 9968 20168 9988
rect 20168 9968 20220 9988
rect 20220 9968 20222 9988
rect 20258 9016 20314 9072
rect 20258 8744 20314 8800
rect 19890 7928 19946 7984
rect 19430 7792 19486 7848
rect 19706 7828 19708 7848
rect 19708 7828 19760 7848
rect 19760 7828 19762 7848
rect 19706 7792 19762 7828
rect 19338 7404 19394 7440
rect 19338 7384 19340 7404
rect 19340 7384 19392 7404
rect 19392 7384 19394 7404
rect 17774 6840 17830 6896
rect 19614 7384 19670 7440
rect 20166 7792 20222 7848
rect 21086 19216 21142 19272
rect 21086 18708 21088 18728
rect 21088 18708 21140 18728
rect 21140 18708 21142 18728
rect 21086 18672 21142 18708
rect 21454 22480 21510 22536
rect 21454 20440 21510 20496
rect 22650 29008 22706 29064
rect 22558 26968 22614 27024
rect 22374 24112 22430 24168
rect 22006 23568 22062 23624
rect 22558 23568 22614 23624
rect 22006 22888 22062 22944
rect 22466 22888 22522 22944
rect 21178 18536 21234 18592
rect 21822 18944 21878 19000
rect 21546 18536 21602 18592
rect 21822 18400 21878 18456
rect 21638 18128 21694 18184
rect 21454 17448 21510 17504
rect 20902 15000 20958 15056
rect 20810 13912 20866 13968
rect 20718 11872 20774 11928
rect 21546 17312 21602 17368
rect 21086 13368 21142 13424
rect 21454 13912 21510 13968
rect 21362 12960 21418 13016
rect 21730 15952 21786 16008
rect 21638 15680 21694 15736
rect 22006 19352 22062 19408
rect 22098 19216 22154 19272
rect 22098 18536 22154 18592
rect 21914 15136 21970 15192
rect 22282 18400 22338 18456
rect 23018 29416 23074 29472
rect 23110 29044 23112 29064
rect 23112 29044 23164 29064
rect 23164 29044 23166 29064
rect 23110 29008 23166 29044
rect 23110 28464 23166 28520
rect 22926 27648 22982 27704
rect 24214 31728 24270 31784
rect 24214 31184 24270 31240
rect 23018 27412 23020 27432
rect 23020 27412 23072 27432
rect 23072 27412 23074 27432
rect 23018 27376 23074 27412
rect 22926 25064 22982 25120
rect 22650 22636 22706 22672
rect 22650 22616 22652 22636
rect 22652 22616 22704 22636
rect 22704 22616 22706 22636
rect 22742 22516 22744 22536
rect 22744 22516 22796 22536
rect 22796 22516 22798 22536
rect 22742 22480 22798 22516
rect 23386 28364 23388 28384
rect 23388 28364 23440 28384
rect 23440 28364 23442 28384
rect 23386 28328 23442 28364
rect 24214 29996 24216 30016
rect 24216 29996 24268 30016
rect 24268 29996 24270 30016
rect 24214 29960 24270 29996
rect 23754 29144 23810 29200
rect 23662 25880 23718 25936
rect 24306 28076 24362 28112
rect 24306 28056 24308 28076
rect 24308 28056 24360 28076
rect 24360 28056 24362 28076
rect 23846 26696 23902 26752
rect 23202 23296 23258 23352
rect 23202 22072 23258 22128
rect 22282 16108 22338 16144
rect 22282 16088 22284 16108
rect 22284 16088 22336 16108
rect 22336 16088 22338 16108
rect 22190 14456 22246 14512
rect 21546 12300 21602 12336
rect 21546 12280 21548 12300
rect 21548 12280 21600 12300
rect 21600 12280 21602 12300
rect 20626 11772 20628 11792
rect 20628 11772 20680 11792
rect 20680 11772 20682 11792
rect 20626 11736 20682 11772
rect 20442 8880 20498 8936
rect 20626 8200 20682 8256
rect 17866 5364 17922 5400
rect 17866 5344 17868 5364
rect 17868 5344 17920 5364
rect 17920 5344 17922 5364
rect 17590 3984 17646 4040
rect 16762 1808 16818 1864
rect 18602 1808 18658 1864
rect 19522 4020 19524 4040
rect 19524 4020 19576 4040
rect 19576 4020 19578 4040
rect 19522 3984 19578 4020
rect 20534 6432 20590 6488
rect 20350 5244 20352 5264
rect 20352 5244 20404 5264
rect 20404 5244 20406 5264
rect 20350 5208 20406 5244
rect 20902 10920 20958 10976
rect 21270 11500 21272 11520
rect 21272 11500 21324 11520
rect 21324 11500 21326 11520
rect 21270 11464 21326 11500
rect 21178 11228 21180 11248
rect 21180 11228 21232 11248
rect 21232 11228 21234 11248
rect 21178 11192 21234 11228
rect 21178 10920 21234 10976
rect 20994 9968 21050 10024
rect 20994 9288 21050 9344
rect 21086 9152 21142 9208
rect 21546 11736 21602 11792
rect 21362 11192 21418 11248
rect 21454 9172 21510 9208
rect 21454 9152 21456 9172
rect 21456 9152 21508 9172
rect 21508 9152 21510 9172
rect 21638 10104 21694 10160
rect 21086 8336 21142 8392
rect 21270 8472 21326 8528
rect 21178 8200 21234 8256
rect 21914 12164 21970 12200
rect 21914 12144 21916 12164
rect 21916 12144 21968 12164
rect 21968 12144 21970 12164
rect 22282 12416 22338 12472
rect 22558 17076 22560 17096
rect 22560 17076 22612 17096
rect 22612 17076 22614 17096
rect 22558 17040 22614 17076
rect 22558 15680 22614 15736
rect 22466 14456 22522 14512
rect 22558 12844 22614 12880
rect 22558 12824 22560 12844
rect 22560 12824 22612 12844
rect 22612 12824 22614 12844
rect 22282 11076 22338 11112
rect 22282 11056 22284 11076
rect 22284 11056 22336 11076
rect 22336 11056 22338 11076
rect 21730 7964 21732 7984
rect 21732 7964 21784 7984
rect 21784 7964 21786 7984
rect 21730 7928 21786 7964
rect 22006 8236 22008 8256
rect 22008 8236 22060 8256
rect 22060 8236 22062 8256
rect 22006 8200 22062 8236
rect 21638 6976 21694 7032
rect 22098 7792 22154 7848
rect 21914 6568 21970 6624
rect 22098 5752 22154 5808
rect 22558 12008 22614 12064
rect 23110 18672 23166 18728
rect 23018 16496 23074 16552
rect 23294 21120 23350 21176
rect 23570 21936 23626 21992
rect 23386 20712 23442 20768
rect 23018 15156 23074 15192
rect 23018 15136 23020 15156
rect 23020 15136 23072 15156
rect 23072 15136 23074 15156
rect 23294 17332 23350 17368
rect 23294 17312 23296 17332
rect 23296 17312 23348 17332
rect 23348 17312 23350 17332
rect 23846 21428 23848 21448
rect 23848 21428 23900 21448
rect 23900 21428 23902 21448
rect 23846 21392 23902 21428
rect 24214 27648 24270 27704
rect 24306 26988 24362 27024
rect 24306 26968 24308 26988
rect 24308 26968 24360 26988
rect 24360 26968 24362 26988
rect 24306 26288 24362 26344
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 25962 32428 26018 32464
rect 25962 32408 25964 32428
rect 25964 32408 26016 32428
rect 26016 32408 26018 32428
rect 25318 30912 25374 30968
rect 24674 30676 24676 30696
rect 24676 30676 24728 30696
rect 24728 30676 24730 30696
rect 24674 30640 24730 30676
rect 25226 30232 25282 30288
rect 24766 29008 24822 29064
rect 24674 26288 24730 26344
rect 24766 24928 24822 24984
rect 25502 29960 25558 30016
rect 25318 29008 25374 29064
rect 25226 26968 25282 27024
rect 25778 27396 25834 27432
rect 25778 27376 25780 27396
rect 25780 27376 25832 27396
rect 25832 27376 25834 27396
rect 25594 27240 25650 27296
rect 25134 25764 25190 25800
rect 25134 25744 25136 25764
rect 25136 25744 25188 25764
rect 25188 25744 25190 25764
rect 25226 24656 25282 24712
rect 24582 23976 24638 24032
rect 24490 23740 24492 23760
rect 24492 23740 24544 23760
rect 24544 23740 24546 23760
rect 24490 23704 24546 23740
rect 24950 23724 25006 23760
rect 24950 23704 24952 23724
rect 24952 23704 25004 23724
rect 25004 23704 25006 23724
rect 24306 21836 24308 21856
rect 24308 21836 24360 21856
rect 24360 21836 24362 21856
rect 24306 21800 24362 21836
rect 23938 19216 23994 19272
rect 23662 16532 23664 16552
rect 23664 16532 23716 16552
rect 23716 16532 23718 16552
rect 22926 15020 22982 15056
rect 22926 15000 22928 15020
rect 22928 15000 22980 15020
rect 22980 15000 22982 15020
rect 22926 13912 22982 13968
rect 22834 11348 22890 11384
rect 22834 11328 22836 11348
rect 22836 11328 22888 11348
rect 22888 11328 22890 11348
rect 22650 9560 22706 9616
rect 22558 9152 22614 9208
rect 23662 16496 23718 16532
rect 24214 20576 24270 20632
rect 24122 16768 24178 16824
rect 24582 21936 24638 21992
rect 24674 21392 24730 21448
rect 24490 21292 24492 21312
rect 24492 21292 24544 21312
rect 24544 21292 24546 21312
rect 24490 21256 24546 21292
rect 24490 19624 24546 19680
rect 24398 19372 24454 19408
rect 24398 19352 24400 19372
rect 24400 19352 24452 19372
rect 24452 19352 24454 19372
rect 25042 22072 25098 22128
rect 24950 21664 25006 21720
rect 24950 21528 25006 21584
rect 24766 19624 24822 19680
rect 24674 19080 24730 19136
rect 24582 17992 24638 18048
rect 24398 17040 24454 17096
rect 27526 30252 27582 30288
rect 27526 30232 27528 30252
rect 27528 30232 27580 30252
rect 27580 30232 27582 30252
rect 28538 31864 28594 31920
rect 27802 29960 27858 30016
rect 26514 28464 26570 28520
rect 26330 28192 26386 28248
rect 26054 26968 26110 27024
rect 25686 26288 25742 26344
rect 25962 25900 26018 25936
rect 25962 25880 25964 25900
rect 25964 25880 26016 25900
rect 26016 25880 26018 25900
rect 25686 23724 25742 23760
rect 25686 23704 25688 23724
rect 25688 23704 25740 23724
rect 25740 23704 25742 23724
rect 25686 21972 25688 21992
rect 25688 21972 25740 21992
rect 25740 21972 25742 21992
rect 25686 21936 25742 21972
rect 25410 21528 25466 21584
rect 25594 21528 25650 21584
rect 25410 19916 25466 19952
rect 25410 19896 25412 19916
rect 25412 19896 25464 19916
rect 25464 19896 25466 19916
rect 24766 18164 24768 18184
rect 24768 18164 24820 18184
rect 24820 18164 24822 18184
rect 24766 18128 24822 18164
rect 24398 16632 24454 16688
rect 25318 18300 25320 18320
rect 25320 18300 25372 18320
rect 25372 18300 25374 18320
rect 25318 18264 25374 18300
rect 25226 17720 25282 17776
rect 25042 17604 25098 17640
rect 25042 17584 25044 17604
rect 25044 17584 25096 17604
rect 25096 17584 25098 17604
rect 24950 17176 25006 17232
rect 24490 15952 24546 16008
rect 24122 15816 24178 15872
rect 23754 14048 23810 14104
rect 23386 12164 23442 12200
rect 23386 12144 23388 12164
rect 23388 12144 23440 12164
rect 23440 12144 23442 12164
rect 23018 10376 23074 10432
rect 22834 9324 22836 9344
rect 22836 9324 22888 9344
rect 22888 9324 22890 9344
rect 22834 9288 22890 9324
rect 22742 8628 22798 8664
rect 22742 8608 22744 8628
rect 22744 8608 22796 8628
rect 22796 8608 22798 8628
rect 23018 8608 23074 8664
rect 22558 5244 22560 5264
rect 22560 5244 22612 5264
rect 22612 5244 22614 5264
rect 22558 5208 22614 5244
rect 23386 11600 23442 11656
rect 23754 11872 23810 11928
rect 23662 11464 23718 11520
rect 23938 14456 23994 14512
rect 24030 12416 24086 12472
rect 23938 11872 23994 11928
rect 23938 11328 23994 11384
rect 23846 11056 23902 11112
rect 23846 10784 23902 10840
rect 23570 9444 23626 9480
rect 23570 9424 23572 9444
rect 23572 9424 23624 9444
rect 23624 9424 23626 9444
rect 23938 10412 23940 10432
rect 23940 10412 23992 10432
rect 23992 10412 23994 10432
rect 23938 10376 23994 10412
rect 23754 7384 23810 7440
rect 24582 15544 24638 15600
rect 24214 15036 24216 15056
rect 24216 15036 24268 15056
rect 24268 15036 24270 15056
rect 24214 15000 24270 15036
rect 24214 11464 24270 11520
rect 24858 14864 24914 14920
rect 24766 14764 24768 14784
rect 24768 14764 24820 14784
rect 24820 14764 24822 14784
rect 24766 14728 24822 14764
rect 25042 15136 25098 15192
rect 24674 13640 24730 13696
rect 24490 11192 24546 11248
rect 24490 10784 24546 10840
rect 23386 5752 23442 5808
rect 24950 13640 25006 13696
rect 24398 7656 24454 7712
rect 24674 5752 24730 5808
rect 25686 18300 25688 18320
rect 25688 18300 25740 18320
rect 25740 18300 25742 18320
rect 25686 18264 25742 18300
rect 25594 16904 25650 16960
rect 25870 18944 25926 19000
rect 26054 23724 26110 23760
rect 26054 23704 26056 23724
rect 26056 23704 26108 23724
rect 26108 23704 26110 23724
rect 26146 23060 26148 23080
rect 26148 23060 26200 23080
rect 26200 23060 26202 23080
rect 26146 23024 26202 23060
rect 26422 24384 26478 24440
rect 26790 29028 26846 29064
rect 27434 29688 27490 29744
rect 26790 29008 26792 29028
rect 26792 29008 26844 29028
rect 26844 29008 26846 29028
rect 26698 26968 26754 27024
rect 26606 23296 26662 23352
rect 26514 22888 26570 22944
rect 27066 25336 27122 25392
rect 27250 29008 27306 29064
rect 26606 20984 26662 21040
rect 26606 20596 26662 20632
rect 26606 20576 26608 20596
rect 26608 20576 26660 20596
rect 26660 20576 26662 20596
rect 26514 19660 26516 19680
rect 26516 19660 26568 19680
rect 26568 19660 26570 19680
rect 26514 19624 26570 19660
rect 25962 16668 25964 16688
rect 25964 16668 26016 16688
rect 26016 16668 26018 16688
rect 25962 16632 26018 16668
rect 25778 16244 25834 16280
rect 25778 16224 25780 16244
rect 25780 16224 25832 16244
rect 25832 16224 25834 16244
rect 25318 14728 25374 14784
rect 25134 12280 25190 12336
rect 26238 17856 26294 17912
rect 26422 18420 26478 18456
rect 26422 18400 26424 18420
rect 26424 18400 26476 18420
rect 26476 18400 26478 18420
rect 26054 14320 26110 14376
rect 25962 13368 26018 13424
rect 25778 12688 25834 12744
rect 25686 12280 25742 12336
rect 25686 8608 25742 8664
rect 25502 8200 25558 8256
rect 26330 15156 26386 15192
rect 26330 15136 26332 15156
rect 26332 15136 26384 15156
rect 26384 15136 26386 15156
rect 26606 18536 26662 18592
rect 27158 23840 27214 23896
rect 27710 29552 27766 29608
rect 27342 23316 27398 23352
rect 27342 23296 27344 23316
rect 27344 23296 27396 23316
rect 27396 23296 27398 23316
rect 27250 23024 27306 23080
rect 26882 22480 26938 22536
rect 26882 21800 26938 21856
rect 26882 21664 26938 21720
rect 28170 30504 28226 30560
rect 28262 27532 28318 27568
rect 28262 27512 28264 27532
rect 28264 27512 28316 27532
rect 28316 27512 28318 27532
rect 28262 26424 28318 26480
rect 27894 24656 27950 24712
rect 28078 23568 28134 23624
rect 28170 22752 28226 22808
rect 26882 20712 26938 20768
rect 26882 19796 26884 19816
rect 26884 19796 26936 19816
rect 26936 19796 26938 19816
rect 26882 19760 26938 19796
rect 26606 15308 26608 15328
rect 26608 15308 26660 15328
rect 26660 15308 26662 15328
rect 26606 15272 26662 15308
rect 26606 14864 26662 14920
rect 26514 14320 26570 14376
rect 26606 14184 26662 14240
rect 26974 18708 26976 18728
rect 26976 18708 27028 18728
rect 27028 18708 27030 18728
rect 26974 18672 27030 18708
rect 27066 17856 27122 17912
rect 26974 15272 27030 15328
rect 26974 14340 27030 14376
rect 26974 14320 26976 14340
rect 26976 14320 27028 14340
rect 27028 14320 27030 14340
rect 26974 14068 27030 14104
rect 26974 14048 26976 14068
rect 26976 14048 27028 14068
rect 27028 14048 27030 14068
rect 26238 10920 26294 10976
rect 26790 12280 26846 12336
rect 26422 10668 26478 10704
rect 26422 10648 26424 10668
rect 26424 10648 26476 10668
rect 26476 10648 26478 10668
rect 26422 10240 26478 10296
rect 26422 10124 26478 10160
rect 26422 10104 26424 10124
rect 26424 10104 26476 10124
rect 26476 10104 26478 10124
rect 26330 9288 26386 9344
rect 25962 8472 26018 8528
rect 26698 10512 26754 10568
rect 27158 13776 27214 13832
rect 27894 20304 27950 20360
rect 27342 17448 27398 17504
rect 27434 17176 27490 17232
rect 27618 15680 27674 15736
rect 28170 21392 28226 21448
rect 28446 24792 28502 24848
rect 29550 31764 29552 31784
rect 29552 31764 29604 31784
rect 29604 31764 29606 31784
rect 29550 31728 29606 31764
rect 28906 30116 28962 30152
rect 28906 30096 28908 30116
rect 28908 30096 28960 30116
rect 28960 30096 28962 30116
rect 28906 29164 28962 29200
rect 28906 29144 28908 29164
rect 28908 29144 28960 29164
rect 28960 29144 28962 29164
rect 29458 30232 29514 30288
rect 29182 28192 29238 28248
rect 28998 27396 29054 27432
rect 28998 27376 29000 27396
rect 29000 27376 29052 27396
rect 29052 27376 29054 27396
rect 28354 24248 28410 24304
rect 28354 24148 28356 24168
rect 28356 24148 28408 24168
rect 28408 24148 28410 24168
rect 28354 24112 28410 24148
rect 28446 22752 28502 22808
rect 28906 25608 28962 25664
rect 28814 24112 28870 24168
rect 28722 24012 28724 24032
rect 28724 24012 28776 24032
rect 28776 24012 28778 24032
rect 28722 23976 28778 24012
rect 28446 21392 28502 21448
rect 28354 21120 28410 21176
rect 28354 19372 28410 19408
rect 28630 21392 28686 21448
rect 28722 21140 28778 21176
rect 28722 21120 28724 21140
rect 28724 21120 28776 21140
rect 28776 21120 28778 21140
rect 29274 27104 29330 27160
rect 29458 27512 29514 27568
rect 29182 26152 29238 26208
rect 29826 29008 29882 29064
rect 30010 28192 30066 28248
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 31206 31864 31262 31920
rect 30286 29824 30342 29880
rect 30378 29552 30434 29608
rect 30194 29300 30250 29336
rect 30194 29280 30196 29300
rect 30196 29280 30248 29300
rect 30248 29280 30250 29300
rect 30102 28056 30158 28112
rect 30010 27920 30066 27976
rect 29918 27784 29974 27840
rect 29918 27396 29974 27432
rect 29918 27376 29920 27396
rect 29920 27376 29972 27396
rect 29972 27376 29974 27396
rect 29642 27104 29698 27160
rect 29274 24928 29330 24984
rect 28354 19352 28356 19372
rect 28356 19352 28408 19372
rect 28408 19352 28410 19372
rect 27986 15272 28042 15328
rect 27158 11872 27214 11928
rect 27158 11636 27160 11656
rect 27160 11636 27212 11656
rect 27212 11636 27214 11656
rect 25778 6316 25834 6352
rect 25778 6296 25780 6316
rect 25780 6296 25832 6316
rect 25832 6296 25834 6316
rect 27158 11600 27214 11636
rect 26974 10376 27030 10432
rect 27158 9832 27214 9888
rect 27158 9580 27214 9616
rect 27158 9560 27160 9580
rect 27160 9560 27212 9580
rect 27212 9560 27214 9580
rect 27066 6568 27122 6624
rect 27618 14612 27674 14648
rect 27618 14592 27620 14612
rect 27620 14592 27672 14612
rect 27672 14592 27674 14612
rect 27618 13932 27674 13968
rect 27618 13912 27620 13932
rect 27620 13912 27672 13932
rect 27672 13912 27674 13932
rect 27618 12824 27674 12880
rect 27618 12164 27674 12200
rect 27618 12144 27620 12164
rect 27620 12144 27672 12164
rect 27672 12144 27674 12164
rect 27986 13912 28042 13968
rect 27986 13812 27988 13832
rect 27988 13812 28040 13832
rect 28040 13812 28042 13832
rect 27986 13776 28042 13812
rect 27894 12688 27950 12744
rect 28722 18844 28724 18864
rect 28724 18844 28776 18864
rect 28776 18844 28778 18864
rect 28722 18808 28778 18844
rect 29366 22636 29422 22672
rect 29366 22616 29368 22636
rect 29368 22616 29420 22636
rect 29420 22616 29422 22636
rect 29366 21800 29422 21856
rect 29918 26016 29974 26072
rect 30102 26832 30158 26888
rect 30378 27648 30434 27704
rect 29918 24112 29974 24168
rect 29734 22072 29790 22128
rect 30010 22072 30066 22128
rect 31114 30540 31116 30560
rect 31116 30540 31168 30560
rect 31168 30540 31170 30560
rect 30838 30096 30894 30152
rect 30746 29588 30748 29608
rect 30748 29588 30800 29608
rect 30800 29588 30802 29608
rect 30746 29552 30802 29588
rect 30654 27784 30710 27840
rect 30930 29552 30986 29608
rect 31114 30504 31170 30540
rect 31114 29008 31170 29064
rect 30930 27956 30932 27976
rect 30932 27956 30984 27976
rect 30984 27956 30986 27976
rect 30930 27920 30986 27956
rect 29550 19488 29606 19544
rect 29182 16108 29238 16144
rect 29182 16088 29184 16108
rect 29184 16088 29236 16108
rect 29236 16088 29238 16108
rect 29366 16108 29422 16144
rect 29366 16088 29368 16108
rect 29368 16088 29420 16108
rect 29420 16088 29422 16108
rect 28906 14728 28962 14784
rect 28170 12280 28226 12336
rect 27802 10920 27858 10976
rect 28170 11328 28226 11384
rect 27894 10004 27896 10024
rect 27896 10004 27948 10024
rect 27948 10004 27950 10024
rect 27894 9968 27950 10004
rect 27802 9560 27858 9616
rect 28170 10412 28172 10432
rect 28172 10412 28224 10432
rect 28224 10412 28226 10432
rect 28170 10376 28226 10412
rect 28078 10104 28134 10160
rect 27618 8200 27674 8256
rect 27894 8336 27950 8392
rect 28906 13796 28962 13832
rect 28906 13776 28908 13796
rect 28908 13776 28960 13796
rect 28960 13776 28962 13796
rect 29274 15136 29330 15192
rect 29826 19352 29882 19408
rect 30286 19488 30342 19544
rect 30654 25472 30710 25528
rect 30562 22072 30618 22128
rect 30562 20712 30618 20768
rect 31022 26308 31078 26344
rect 31022 26288 31024 26308
rect 31024 26288 31076 26308
rect 31076 26288 31078 26308
rect 30930 26016 30986 26072
rect 30930 25472 30986 25528
rect 30930 23024 30986 23080
rect 30838 22888 30894 22944
rect 31390 29688 31446 29744
rect 31390 28872 31446 28928
rect 31390 28328 31446 28384
rect 31298 28192 31354 28248
rect 31758 30096 31814 30152
rect 32126 30096 32182 30152
rect 32402 29688 32458 29744
rect 32310 29552 32366 29608
rect 31574 29044 31576 29064
rect 31576 29044 31628 29064
rect 31628 29044 31630 29064
rect 31574 29008 31630 29044
rect 31850 28736 31906 28792
rect 31574 28464 31630 28520
rect 31298 24828 31300 24848
rect 31300 24828 31352 24848
rect 31352 24828 31354 24848
rect 31298 24792 31354 24828
rect 31298 24384 31354 24440
rect 31942 28636 31944 28656
rect 31944 28636 31996 28656
rect 31996 28636 31998 28656
rect 31942 28600 31998 28636
rect 31666 28056 31722 28112
rect 31574 27784 31630 27840
rect 32494 29280 32550 29336
rect 32402 29164 32458 29200
rect 32402 29144 32404 29164
rect 32404 29144 32456 29164
rect 32456 29144 32458 29164
rect 32402 29008 32458 29064
rect 32310 28328 32366 28384
rect 32034 26036 32090 26072
rect 32034 26016 32036 26036
rect 32036 26016 32088 26036
rect 32088 26016 32090 26036
rect 32678 28500 32680 28520
rect 32680 28500 32732 28520
rect 32732 28500 32734 28520
rect 32678 28464 32734 28500
rect 32678 28056 32734 28112
rect 32494 27376 32550 27432
rect 32862 28872 32918 28928
rect 31758 25236 31760 25256
rect 31760 25236 31812 25256
rect 31812 25236 31814 25256
rect 31758 25200 31814 25236
rect 30838 19624 30894 19680
rect 28354 11092 28356 11112
rect 28356 11092 28408 11112
rect 28408 11092 28410 11112
rect 28354 11056 28410 11092
rect 28814 12416 28870 12472
rect 28722 12044 28724 12064
rect 28724 12044 28776 12064
rect 28776 12044 28778 12064
rect 28722 12008 28778 12044
rect 28538 10240 28594 10296
rect 28354 8916 28356 8936
rect 28356 8916 28408 8936
rect 28408 8916 28410 8936
rect 28354 8880 28410 8916
rect 29182 11600 29238 11656
rect 29274 10920 29330 10976
rect 28722 9696 28778 9752
rect 28722 9152 28778 9208
rect 29090 10376 29146 10432
rect 29274 10104 29330 10160
rect 28906 9982 28908 10024
rect 28908 9982 28960 10024
rect 28960 9982 28962 10024
rect 28906 9968 28962 9982
rect 29274 9832 29330 9888
rect 29550 13776 29606 13832
rect 29550 13504 29606 13560
rect 29550 11636 29552 11656
rect 29552 11636 29604 11656
rect 29604 11636 29606 11656
rect 29550 11600 29606 11636
rect 29550 11056 29606 11112
rect 29918 10668 29974 10704
rect 29918 10648 29920 10668
rect 29920 10648 29972 10668
rect 29972 10648 29974 10668
rect 29826 9868 29828 9888
rect 29828 9868 29880 9888
rect 29880 9868 29882 9888
rect 29826 9832 29882 9868
rect 29458 8200 29514 8256
rect 28998 7540 29054 7576
rect 28998 7520 29000 7540
rect 29000 7520 29052 7540
rect 29052 7520 29054 7540
rect 28722 6568 28778 6624
rect 30194 15988 30196 16008
rect 30196 15988 30248 16008
rect 30248 15988 30250 16008
rect 30194 15952 30250 15988
rect 30194 15408 30250 15464
rect 30562 13368 30618 13424
rect 30746 12708 30802 12744
rect 30746 12688 30748 12708
rect 30748 12688 30800 12708
rect 30800 12688 30802 12708
rect 30746 12416 30802 12472
rect 30930 17856 30986 17912
rect 31666 23024 31722 23080
rect 32034 25200 32090 25256
rect 31482 22480 31538 22536
rect 31850 22888 31906 22944
rect 31758 20984 31814 21040
rect 31482 20576 31538 20632
rect 31298 20440 31354 20496
rect 31390 19760 31446 19816
rect 31390 19624 31446 19680
rect 31206 16224 31262 16280
rect 31666 20440 31722 20496
rect 31666 20340 31668 20360
rect 31668 20340 31720 20360
rect 31720 20340 31722 20360
rect 31666 20304 31722 20340
rect 31574 16108 31630 16144
rect 31574 16088 31576 16108
rect 31576 16088 31628 16108
rect 31628 16088 31630 16108
rect 31298 15308 31300 15328
rect 31300 15308 31352 15328
rect 31352 15308 31354 15328
rect 31298 15272 31354 15308
rect 29826 8372 29828 8392
rect 29828 8372 29880 8392
rect 29880 8372 29882 8392
rect 29826 8336 29882 8372
rect 30562 7928 30618 7984
rect 30562 7248 30618 7304
rect 30194 6976 30250 7032
rect 31114 11464 31170 11520
rect 31206 10004 31208 10024
rect 31208 10004 31260 10024
rect 31260 10004 31262 10024
rect 31206 9968 31262 10004
rect 31850 20204 31852 20224
rect 31852 20204 31904 20224
rect 31904 20204 31906 20224
rect 31850 20168 31906 20204
rect 32218 25064 32274 25120
rect 32034 23296 32090 23352
rect 33230 30232 33286 30288
rect 33506 29824 33562 29880
rect 33414 29280 33470 29336
rect 33138 28736 33194 28792
rect 33598 29416 33654 29472
rect 33138 28328 33194 28384
rect 33046 28056 33102 28112
rect 32402 24928 32458 24984
rect 32586 25200 32642 25256
rect 32494 24792 32550 24848
rect 32310 22616 32366 22672
rect 32310 22072 32366 22128
rect 31666 12280 31722 12336
rect 32402 19352 32458 19408
rect 33414 28192 33470 28248
rect 33690 28600 33746 28656
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 33690 27648 33746 27704
rect 33046 25880 33102 25936
rect 33138 25744 33194 25800
rect 32770 24248 32826 24304
rect 33322 25608 33378 25664
rect 33414 25472 33470 25528
rect 33414 25064 33470 25120
rect 32954 22752 33010 22808
rect 32402 18128 32458 18184
rect 32310 17856 32366 17912
rect 32862 20748 32864 20768
rect 32864 20748 32916 20768
rect 32916 20748 32918 20768
rect 32862 20712 32918 20748
rect 33690 26968 33746 27024
rect 33874 28328 33930 28384
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 33874 27784 33930 27840
rect 33782 26288 33838 26344
rect 33690 25608 33746 25664
rect 33690 25236 33692 25256
rect 33692 25236 33744 25256
rect 33744 25236 33746 25256
rect 33690 25200 33746 25236
rect 33322 20576 33378 20632
rect 33230 20304 33286 20360
rect 32954 20032 33010 20088
rect 32586 16224 32642 16280
rect 31758 9968 31814 10024
rect 34334 28364 34336 28384
rect 34336 28364 34388 28384
rect 34388 28364 34390 28384
rect 34334 28328 34390 28364
rect 35622 29588 35624 29608
rect 35624 29588 35676 29608
rect 35676 29588 35678 29608
rect 35622 29552 35678 29588
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34334 26016 34390 26072
rect 34242 25744 34298 25800
rect 34518 26832 34574 26888
rect 33874 24268 33930 24304
rect 33874 24248 33876 24268
rect 33876 24248 33928 24268
rect 33928 24248 33930 24268
rect 33414 15952 33470 16008
rect 31666 8744 31722 8800
rect 31022 6840 31078 6896
rect 32678 9560 32734 9616
rect 34058 23432 34114 23488
rect 33046 11736 33102 11792
rect 32862 9580 32918 9616
rect 33322 11756 33378 11792
rect 33322 11736 33324 11756
rect 33324 11736 33376 11756
rect 33376 11736 33378 11756
rect 32862 9560 32864 9580
rect 32864 9560 32916 9580
rect 32916 9560 32918 9580
rect 33230 9288 33286 9344
rect 34426 18128 34482 18184
rect 34518 17992 34574 18048
rect 35070 28076 35126 28112
rect 35070 28056 35072 28076
rect 35072 28056 35124 28076
rect 35124 28056 35126 28076
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35438 27920 35494 27976
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35254 27512 35310 27568
rect 35070 27004 35072 27024
rect 35072 27004 35124 27024
rect 35124 27004 35126 27024
rect 35070 26968 35126 27004
rect 36082 27512 36138 27568
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35162 26152 35218 26208
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35162 25336 35218 25392
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34978 24148 34980 24168
rect 34980 24148 35032 24168
rect 35032 24148 35034 24168
rect 34978 24112 35034 24148
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35254 23060 35256 23080
rect 35256 23060 35308 23080
rect 35308 23060 35310 23080
rect 35254 23024 35310 23060
rect 35070 22480 35126 22536
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 36174 27240 36230 27296
rect 36266 26560 36322 26616
rect 35714 26288 35770 26344
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 36174 25880 36230 25936
rect 35806 25472 35862 25528
rect 35714 25236 35716 25256
rect 35716 25236 35768 25256
rect 35768 25236 35770 25256
rect 35714 25200 35770 25236
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35530 24132 35586 24168
rect 35530 24112 35532 24132
rect 35532 24112 35584 24132
rect 35584 24112 35586 24132
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 36266 24792 36322 24848
rect 36082 24520 36138 24576
rect 36174 23160 36230 23216
rect 36174 22516 36176 22536
rect 36176 22516 36228 22536
rect 36228 22516 36230 22536
rect 36174 22480 36230 22516
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34702 20748 34704 20768
rect 34704 20748 34756 20768
rect 34756 20748 34758 20768
rect 34702 20712 34758 20748
rect 34978 20884 34980 20904
rect 34980 20884 35032 20904
rect 35032 20884 35034 20904
rect 34978 20848 35034 20884
rect 35530 21120 35586 21176
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34334 11056 34390 11112
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35254 16516 35310 16552
rect 35254 16496 35256 16516
rect 35256 16496 35308 16516
rect 35308 16496 35310 16516
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35070 14864 35126 14920
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34886 12008 34942 12064
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34058 10512 34114 10568
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34334 9580 34390 9616
rect 34334 9560 34336 9580
rect 34336 9560 34388 9580
rect 34388 9560 34390 9580
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 36174 12688 36230 12744
rect 36450 23568 36506 23624
rect 36726 21528 36782 21584
rect 36634 18264 36690 18320
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 36082 3460 36138 3496
rect 36082 3440 36084 3460
rect 36084 3440 36136 3460
rect 36136 3440 36138 3460
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36138 800 36168
rect 0 36078 1042 36138
rect 0 36048 800 36078
rect 982 35910 1042 36078
rect 614 35850 1042 35910
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 12893 35866 12959 35869
rect 18229 35866 18295 35869
rect 12893 35864 18295 35866
rect 614 35594 674 35850
rect 12893 35808 12898 35864
rect 12954 35808 18234 35864
rect 18290 35808 18295 35864
rect 12893 35806 18295 35808
rect 12893 35803 12959 35806
rect 18229 35803 18295 35806
rect 14181 35730 14247 35733
rect 15653 35730 15719 35733
rect 14181 35728 15719 35730
rect 14181 35672 14186 35728
rect 14242 35672 15658 35728
rect 15714 35672 15719 35728
rect 14181 35670 15719 35672
rect 14181 35667 14247 35670
rect 15653 35667 15719 35670
rect 22461 35730 22527 35733
rect 23013 35730 23079 35733
rect 22461 35728 23079 35730
rect 22461 35672 22466 35728
rect 22522 35672 23018 35728
rect 23074 35672 23079 35728
rect 22461 35670 23079 35672
rect 22461 35667 22527 35670
rect 23013 35667 23079 35670
rect 8886 35594 8892 35596
rect 614 35534 8892 35594
rect 8886 35532 8892 35534
rect 8956 35532 8962 35596
rect 12709 35458 12775 35461
rect 13629 35458 13695 35461
rect 12709 35456 13695 35458
rect 12709 35400 12714 35456
rect 12770 35400 13634 35456
rect 13690 35400 13695 35456
rect 12709 35398 13695 35400
rect 12709 35395 12775 35398
rect 13629 35395 13695 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 10225 35322 10291 35325
rect 14733 35322 14799 35325
rect 10225 35320 14799 35322
rect 10225 35264 10230 35320
rect 10286 35264 14738 35320
rect 14794 35264 14799 35320
rect 10225 35262 14799 35264
rect 10225 35259 10291 35262
rect 14733 35259 14799 35262
rect 10685 35050 10751 35053
rect 12157 35050 12223 35053
rect 12617 35050 12683 35053
rect 10685 35048 12683 35050
rect 10685 34992 10690 35048
rect 10746 34992 12162 35048
rect 12218 34992 12622 35048
rect 12678 34992 12683 35048
rect 10685 34990 12683 34992
rect 10685 34987 10751 34990
rect 12157 34987 12223 34990
rect 12617 34987 12683 34990
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 8293 34644 8359 34645
rect 8293 34642 8340 34644
rect 8248 34640 8340 34642
rect 8248 34584 8298 34640
rect 8248 34582 8340 34584
rect 8293 34580 8340 34582
rect 8404 34580 8410 34644
rect 8293 34579 8359 34580
rect 8661 34506 8727 34509
rect 22185 34506 22251 34509
rect 8661 34504 22251 34506
rect 8661 34448 8666 34504
rect 8722 34448 22190 34504
rect 22246 34448 22251 34504
rect 8661 34446 22251 34448
rect 8661 34443 8727 34446
rect 22185 34443 22251 34446
rect 9765 34370 9831 34373
rect 9990 34370 9996 34372
rect 9765 34368 9996 34370
rect 9765 34312 9770 34368
rect 9826 34312 9996 34368
rect 9765 34310 9996 34312
rect 9765 34307 9831 34310
rect 9990 34308 9996 34310
rect 10060 34308 10066 34372
rect 13670 34308 13676 34372
rect 13740 34370 13746 34372
rect 19057 34370 19123 34373
rect 13740 34368 19123 34370
rect 13740 34312 19062 34368
rect 19118 34312 19123 34368
rect 13740 34310 19123 34312
rect 13740 34308 13746 34310
rect 19057 34307 19123 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19333 33826 19399 33829
rect 19793 33826 19859 33829
rect 19333 33824 19859 33826
rect 19333 33768 19338 33824
rect 19394 33768 19798 33824
rect 19854 33768 19859 33824
rect 19333 33766 19859 33768
rect 19333 33763 19399 33766
rect 19793 33763 19859 33766
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 19425 33418 19491 33421
rect 21357 33418 21423 33421
rect 21817 33418 21883 33421
rect 22829 33418 22895 33421
rect 19425 33416 22895 33418
rect 19425 33360 19430 33416
rect 19486 33360 21362 33416
rect 21418 33360 21822 33416
rect 21878 33360 22834 33416
rect 22890 33360 22895 33416
rect 19425 33358 22895 33360
rect 19425 33355 19491 33358
rect 21357 33355 21423 33358
rect 21817 33355 21883 33358
rect 22829 33355 22895 33358
rect 9806 33220 9812 33284
rect 9876 33282 9882 33284
rect 10133 33282 10199 33285
rect 9876 33280 10199 33282
rect 9876 33224 10138 33280
rect 10194 33224 10199 33280
rect 9876 33222 10199 33224
rect 9876 33220 9882 33222
rect 10133 33219 10199 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 13077 33146 13143 33149
rect 19149 33146 19215 33149
rect 13077 33144 19215 33146
rect 13077 33088 13082 33144
rect 13138 33088 19154 33144
rect 19210 33088 19215 33144
rect 13077 33086 19215 33088
rect 13077 33083 13143 33086
rect 19149 33083 19215 33086
rect 10869 33010 10935 33013
rect 17309 33010 17375 33013
rect 10869 33008 17375 33010
rect 10869 32952 10874 33008
rect 10930 32952 17314 33008
rect 17370 32952 17375 33008
rect 10869 32950 17375 32952
rect 10869 32947 10935 32950
rect 17309 32947 17375 32950
rect 17861 32874 17927 32877
rect 18689 32874 18755 32877
rect 17861 32872 18755 32874
rect 17861 32816 17866 32872
rect 17922 32816 18694 32872
rect 18750 32816 18755 32872
rect 17861 32814 18755 32816
rect 17861 32811 17927 32814
rect 18689 32811 18755 32814
rect 18137 32738 18203 32741
rect 18873 32738 18939 32741
rect 18137 32736 18939 32738
rect 18137 32680 18142 32736
rect 18198 32680 18878 32736
rect 18934 32680 18939 32736
rect 18137 32678 18939 32680
rect 18137 32675 18203 32678
rect 18873 32675 18939 32678
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 23013 32466 23079 32469
rect 25957 32466 26023 32469
rect 23013 32464 26023 32466
rect 23013 32408 23018 32464
rect 23074 32408 25962 32464
rect 26018 32408 26023 32464
rect 23013 32406 26023 32408
rect 23013 32403 23079 32406
rect 25957 32403 26023 32406
rect 9305 32330 9371 32333
rect 18045 32330 18111 32333
rect 9305 32328 18111 32330
rect 9305 32272 9310 32328
rect 9366 32272 18050 32328
rect 18106 32272 18111 32328
rect 9305 32270 18111 32272
rect 9305 32267 9371 32270
rect 18045 32267 18111 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 22277 32058 22343 32061
rect 22142 32056 22343 32058
rect 22142 32000 22282 32056
rect 22338 32000 22343 32056
rect 22142 31998 22343 32000
rect 16665 31922 16731 31925
rect 17861 31922 17927 31925
rect 16665 31920 17927 31922
rect 16665 31864 16670 31920
rect 16726 31864 17866 31920
rect 17922 31864 17927 31920
rect 16665 31862 17927 31864
rect 16665 31859 16731 31862
rect 17861 31859 17927 31862
rect 22142 31789 22202 31998
rect 22277 31995 22343 31998
rect 22461 32058 22527 32061
rect 22921 32058 22987 32061
rect 22461 32056 22987 32058
rect 22461 32000 22466 32056
rect 22522 32000 22926 32056
rect 22982 32000 22987 32056
rect 22461 31998 22987 32000
rect 22461 31995 22527 31998
rect 22921 31995 22987 31998
rect 28533 31922 28599 31925
rect 31201 31922 31267 31925
rect 28533 31920 31267 31922
rect 28533 31864 28538 31920
rect 28594 31864 31206 31920
rect 31262 31864 31267 31920
rect 28533 31862 31267 31864
rect 28533 31859 28599 31862
rect 31201 31859 31267 31862
rect 10593 31786 10659 31789
rect 10961 31786 11027 31789
rect 12065 31786 12131 31789
rect 13721 31786 13787 31789
rect 10593 31784 13787 31786
rect 10593 31728 10598 31784
rect 10654 31728 10966 31784
rect 11022 31728 12070 31784
rect 12126 31728 13726 31784
rect 13782 31728 13787 31784
rect 10593 31726 13787 31728
rect 22142 31784 22251 31789
rect 22142 31728 22190 31784
rect 22246 31728 22251 31784
rect 22142 31726 22251 31728
rect 10593 31723 10659 31726
rect 10961 31723 11027 31726
rect 12065 31723 12131 31726
rect 13721 31723 13787 31726
rect 22185 31723 22251 31726
rect 24209 31786 24275 31789
rect 29545 31786 29611 31789
rect 24209 31784 29611 31786
rect 24209 31728 24214 31784
rect 24270 31728 29550 31784
rect 29606 31728 29611 31784
rect 24209 31726 29611 31728
rect 24209 31723 24275 31726
rect 29545 31723 29611 31726
rect 9489 31650 9555 31653
rect 9765 31650 9831 31653
rect 9489 31648 9831 31650
rect 9489 31592 9494 31648
rect 9550 31592 9770 31648
rect 9826 31592 9831 31648
rect 9489 31590 9831 31592
rect 9489 31587 9555 31590
rect 9765 31587 9831 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 9305 31514 9371 31517
rect 10777 31514 10843 31517
rect 9305 31512 10843 31514
rect 9305 31456 9310 31512
rect 9366 31456 10782 31512
rect 10838 31456 10843 31512
rect 9305 31454 10843 31456
rect 9305 31451 9371 31454
rect 10777 31451 10843 31454
rect 0 31378 800 31408
rect 2681 31378 2747 31381
rect 0 31376 2747 31378
rect 0 31320 2686 31376
rect 2742 31320 2747 31376
rect 0 31318 2747 31320
rect 0 31288 800 31318
rect 2681 31315 2747 31318
rect 9121 31378 9187 31381
rect 10501 31378 10567 31381
rect 9121 31376 10567 31378
rect 9121 31320 9126 31376
rect 9182 31320 10506 31376
rect 10562 31320 10567 31376
rect 9121 31318 10567 31320
rect 9121 31315 9187 31318
rect 10501 31315 10567 31318
rect 24209 31244 24275 31245
rect 24158 31180 24164 31244
rect 24228 31242 24275 31244
rect 24228 31240 24320 31242
rect 24270 31184 24320 31240
rect 24228 31182 24320 31184
rect 24228 31180 24275 31182
rect 24209 31179 24275 31180
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 13486 30908 13492 30972
rect 13556 30970 13562 30972
rect 25313 30970 25379 30973
rect 13556 30968 25379 30970
rect 13556 30912 25318 30968
rect 25374 30912 25379 30968
rect 13556 30910 25379 30912
rect 13556 30908 13562 30910
rect 25313 30907 25379 30910
rect 9029 30834 9095 30837
rect 14549 30834 14615 30837
rect 9029 30832 14615 30834
rect 9029 30776 9034 30832
rect 9090 30776 14554 30832
rect 14610 30776 14615 30832
rect 9029 30774 14615 30776
rect 9029 30771 9095 30774
rect 14549 30771 14615 30774
rect 0 30698 800 30728
rect 5165 30698 5231 30701
rect 0 30696 5231 30698
rect 0 30640 5170 30696
rect 5226 30640 5231 30696
rect 0 30638 5231 30640
rect 0 30608 800 30638
rect 5165 30635 5231 30638
rect 9857 30698 9923 30701
rect 9990 30698 9996 30700
rect 9857 30696 9996 30698
rect 9857 30640 9862 30696
rect 9918 30640 9996 30696
rect 9857 30638 9996 30640
rect 9857 30635 9923 30638
rect 9990 30636 9996 30638
rect 10060 30636 10066 30700
rect 21950 30636 21956 30700
rect 22020 30698 22026 30700
rect 24669 30698 24735 30701
rect 22020 30696 24735 30698
rect 22020 30640 24674 30696
rect 24730 30640 24735 30696
rect 22020 30638 24735 30640
rect 22020 30636 22026 30638
rect 24669 30635 24735 30638
rect 11237 30562 11303 30565
rect 11830 30562 11836 30564
rect 11237 30560 11836 30562
rect 11237 30504 11242 30560
rect 11298 30504 11836 30560
rect 11237 30502 11836 30504
rect 11237 30499 11303 30502
rect 11830 30500 11836 30502
rect 11900 30500 11906 30564
rect 28165 30562 28231 30565
rect 31109 30562 31175 30565
rect 28165 30560 31175 30562
rect 28165 30504 28170 30560
rect 28226 30504 31114 30560
rect 31170 30504 31175 30560
rect 28165 30502 31175 30504
rect 28165 30499 28231 30502
rect 31109 30499 31175 30502
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 10910 30364 10916 30428
rect 10980 30426 10986 30428
rect 11697 30426 11763 30429
rect 16573 30428 16639 30429
rect 16573 30426 16620 30428
rect 10980 30424 11763 30426
rect 10980 30368 11702 30424
rect 11758 30368 11763 30424
rect 10980 30366 11763 30368
rect 16528 30424 16620 30426
rect 16684 30426 16690 30428
rect 17861 30426 17927 30429
rect 16684 30424 17927 30426
rect 16528 30368 16578 30424
rect 16684 30368 17866 30424
rect 17922 30368 17927 30424
rect 16528 30366 16620 30368
rect 10980 30364 10986 30366
rect 11697 30363 11763 30366
rect 16573 30364 16620 30366
rect 16684 30366 17927 30368
rect 16684 30364 16690 30366
rect 16573 30363 16639 30364
rect 17861 30363 17927 30366
rect 11421 30290 11487 30293
rect 13854 30290 13860 30292
rect 11421 30288 13860 30290
rect 11421 30232 11426 30288
rect 11482 30232 13860 30288
rect 11421 30230 13860 30232
rect 11421 30227 11487 30230
rect 13854 30228 13860 30230
rect 13924 30290 13930 30292
rect 17493 30290 17559 30293
rect 21357 30290 21423 30293
rect 13924 30288 21423 30290
rect 13924 30232 17498 30288
rect 17554 30232 21362 30288
rect 21418 30232 21423 30288
rect 13924 30230 21423 30232
rect 13924 30228 13930 30230
rect 17493 30227 17559 30230
rect 21357 30227 21423 30230
rect 25221 30290 25287 30293
rect 25446 30290 25452 30292
rect 25221 30288 25452 30290
rect 25221 30232 25226 30288
rect 25282 30232 25452 30288
rect 25221 30230 25452 30232
rect 25221 30227 25287 30230
rect 25446 30228 25452 30230
rect 25516 30290 25522 30292
rect 27521 30290 27587 30293
rect 25516 30288 27587 30290
rect 25516 30232 27526 30288
rect 27582 30232 27587 30288
rect 25516 30230 27587 30232
rect 25516 30228 25522 30230
rect 27521 30227 27587 30230
rect 29453 30290 29519 30293
rect 33225 30290 33291 30293
rect 29453 30288 33291 30290
rect 29453 30232 29458 30288
rect 29514 30232 33230 30288
rect 33286 30232 33291 30288
rect 29453 30230 33291 30232
rect 29453 30227 29519 30230
rect 33225 30227 33291 30230
rect 28901 30154 28967 30157
rect 30833 30154 30899 30157
rect 28901 30152 30899 30154
rect 28901 30096 28906 30152
rect 28962 30096 30838 30152
rect 30894 30096 30899 30152
rect 28901 30094 30899 30096
rect 28901 30091 28967 30094
rect 30833 30091 30899 30094
rect 31753 30154 31819 30157
rect 31886 30154 31892 30156
rect 31753 30152 31892 30154
rect 31753 30096 31758 30152
rect 31814 30096 31892 30152
rect 31753 30094 31892 30096
rect 31753 30091 31819 30094
rect 31886 30092 31892 30094
rect 31956 30092 31962 30156
rect 32121 30154 32187 30157
rect 32254 30154 32260 30156
rect 32078 30152 32260 30154
rect 32078 30096 32126 30152
rect 32182 30096 32260 30152
rect 32078 30094 32260 30096
rect 32078 30091 32187 30094
rect 32254 30092 32260 30094
rect 32324 30092 32330 30156
rect 21817 30018 21883 30021
rect 24209 30018 24275 30021
rect 25497 30018 25563 30021
rect 21817 30016 25563 30018
rect 21817 29960 21822 30016
rect 21878 29960 24214 30016
rect 24270 29960 25502 30016
rect 25558 29960 25563 30016
rect 21817 29958 25563 29960
rect 21817 29955 21883 29958
rect 24209 29955 24275 29958
rect 25497 29955 25563 29958
rect 27797 30018 27863 30021
rect 32078 30018 32138 30091
rect 27797 30016 32138 30018
rect 27797 29960 27802 30016
rect 27858 29960 32138 30016
rect 27797 29958 32138 29960
rect 27797 29955 27863 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 30281 29882 30347 29885
rect 33501 29882 33567 29885
rect 30281 29880 33567 29882
rect 30281 29824 30286 29880
rect 30342 29824 33506 29880
rect 33562 29824 33567 29880
rect 30281 29822 33567 29824
rect 30281 29819 30347 29822
rect 33501 29819 33567 29822
rect 27429 29746 27495 29749
rect 31385 29746 31451 29749
rect 32397 29748 32463 29749
rect 32397 29746 32444 29748
rect 27429 29744 32444 29746
rect 32508 29746 32514 29748
rect 27429 29688 27434 29744
rect 27490 29688 31390 29744
rect 31446 29688 32402 29744
rect 27429 29686 32444 29688
rect 27429 29683 27495 29686
rect 31385 29683 31451 29686
rect 32397 29684 32444 29686
rect 32508 29686 32590 29746
rect 32508 29684 32514 29686
rect 32397 29683 32463 29684
rect 9765 29610 9831 29613
rect 10317 29610 10383 29613
rect 14733 29610 14799 29613
rect 27705 29610 27771 29613
rect 9765 29608 14799 29610
rect 9765 29552 9770 29608
rect 9826 29552 10322 29608
rect 10378 29552 14738 29608
rect 14794 29552 14799 29608
rect 9765 29550 14799 29552
rect 9765 29547 9831 29550
rect 10317 29547 10383 29550
rect 14733 29547 14799 29550
rect 22050 29608 27771 29610
rect 22050 29552 27710 29608
rect 27766 29552 27771 29608
rect 22050 29550 27771 29552
rect 12065 29474 12131 29477
rect 12893 29474 12959 29477
rect 12065 29472 12959 29474
rect 12065 29416 12070 29472
rect 12126 29416 12898 29472
rect 12954 29416 12959 29472
rect 12065 29414 12959 29416
rect 12065 29411 12131 29414
rect 12893 29411 12959 29414
rect 4870 29408 5186 29409
rect 0 29338 800 29368
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 3693 29338 3759 29341
rect 0 29336 3759 29338
rect 0 29280 3698 29336
rect 3754 29280 3759 29336
rect 0 29278 3759 29280
rect 0 29248 800 29278
rect 3693 29275 3759 29278
rect 8293 29338 8359 29341
rect 9121 29338 9187 29341
rect 8293 29336 9187 29338
rect 8293 29280 8298 29336
rect 8354 29280 9126 29336
rect 9182 29280 9187 29336
rect 8293 29278 9187 29280
rect 8293 29275 8359 29278
rect 9121 29275 9187 29278
rect 12617 29338 12683 29341
rect 15009 29338 15075 29341
rect 22050 29338 22110 29550
rect 27705 29547 27771 29550
rect 30373 29610 30439 29613
rect 30741 29610 30807 29613
rect 30373 29608 30807 29610
rect 30373 29552 30378 29608
rect 30434 29552 30746 29608
rect 30802 29552 30807 29608
rect 30373 29550 30807 29552
rect 30373 29547 30439 29550
rect 30741 29547 30807 29550
rect 30925 29610 30991 29613
rect 32305 29610 32371 29613
rect 30925 29608 32371 29610
rect 30925 29552 30930 29608
rect 30986 29552 32310 29608
rect 32366 29552 32371 29608
rect 30925 29550 32371 29552
rect 30925 29547 30991 29550
rect 32305 29547 32371 29550
rect 35382 29548 35388 29612
rect 35452 29610 35458 29612
rect 35617 29610 35683 29613
rect 35452 29608 35683 29610
rect 35452 29552 35622 29608
rect 35678 29552 35683 29608
rect 35452 29550 35683 29552
rect 35452 29548 35458 29550
rect 35617 29547 35683 29550
rect 23013 29474 23079 29477
rect 33593 29474 33659 29477
rect 12617 29336 22110 29338
rect 12617 29280 12622 29336
rect 12678 29280 15014 29336
rect 15070 29280 22110 29336
rect 12617 29278 22110 29280
rect 22188 29472 33659 29474
rect 22188 29416 23018 29472
rect 23074 29416 33598 29472
rect 33654 29416 33659 29472
rect 22188 29414 33659 29416
rect 12617 29275 12683 29278
rect 15009 29275 15075 29278
rect 4337 29202 4403 29205
rect 4705 29202 4771 29205
rect 14089 29202 14155 29205
rect 22188 29202 22248 29414
rect 23013 29411 23079 29414
rect 33593 29411 33659 29414
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 30189 29338 30255 29341
rect 30414 29338 30420 29340
rect 30189 29336 30420 29338
rect 30189 29280 30194 29336
rect 30250 29280 30420 29336
rect 30189 29278 30420 29280
rect 30189 29275 30255 29278
rect 30414 29276 30420 29278
rect 30484 29276 30490 29340
rect 32489 29338 32555 29341
rect 33409 29338 33475 29341
rect 30652 29336 33475 29338
rect 30652 29280 32494 29336
rect 32550 29280 33414 29336
rect 33470 29280 33475 29336
rect 30652 29278 33475 29280
rect 4337 29200 14155 29202
rect 4337 29144 4342 29200
rect 4398 29144 4710 29200
rect 4766 29144 14094 29200
rect 14150 29144 14155 29200
rect 4337 29142 14155 29144
rect 4337 29139 4403 29142
rect 4705 29139 4771 29142
rect 14089 29139 14155 29142
rect 22050 29142 22248 29202
rect 23749 29202 23815 29205
rect 28901 29202 28967 29205
rect 30652 29202 30712 29278
rect 32489 29275 32555 29278
rect 33409 29275 33475 29278
rect 32397 29202 32463 29205
rect 23749 29200 30712 29202
rect 23749 29144 23754 29200
rect 23810 29144 28906 29200
rect 28962 29144 30712 29200
rect 23749 29142 30712 29144
rect 30790 29200 32463 29202
rect 30790 29144 32402 29200
rect 32458 29144 32463 29200
rect 30790 29142 32463 29144
rect 5758 29004 5764 29068
rect 5828 29066 5834 29068
rect 9581 29066 9647 29069
rect 5828 29064 9647 29066
rect 5828 29008 9586 29064
rect 9642 29008 9647 29064
rect 5828 29006 9647 29008
rect 5828 29004 5834 29006
rect 9581 29003 9647 29006
rect 10041 29066 10107 29069
rect 10685 29066 10751 29069
rect 10041 29064 10751 29066
rect 10041 29008 10046 29064
rect 10102 29008 10690 29064
rect 10746 29008 10751 29064
rect 10041 29006 10751 29008
rect 10041 29003 10107 29006
rect 10685 29003 10751 29006
rect 11789 29066 11855 29069
rect 12525 29068 12591 29069
rect 12198 29066 12204 29068
rect 11789 29064 12204 29066
rect 11789 29008 11794 29064
rect 11850 29008 12204 29064
rect 11789 29006 12204 29008
rect 11789 29003 11855 29006
rect 12198 29004 12204 29006
rect 12268 29004 12274 29068
rect 12525 29064 12572 29068
rect 12636 29066 12642 29068
rect 12985 29066 13051 29069
rect 14457 29066 14523 29069
rect 12525 29008 12530 29064
rect 12525 29004 12572 29008
rect 12636 29006 12682 29066
rect 12985 29064 14523 29066
rect 12985 29008 12990 29064
rect 13046 29008 14462 29064
rect 14518 29008 14523 29064
rect 12985 29006 14523 29008
rect 12636 29004 12642 29006
rect 12525 29003 12591 29004
rect 12985 29003 13051 29006
rect 14457 29003 14523 29006
rect 21081 29066 21147 29069
rect 21909 29066 21975 29069
rect 21081 29064 21975 29066
rect 21081 29008 21086 29064
rect 21142 29008 21914 29064
rect 21970 29008 21975 29064
rect 21081 29006 21975 29008
rect 21081 29003 21147 29006
rect 21909 29003 21975 29006
rect 7598 28868 7604 28932
rect 7668 28930 7674 28932
rect 8937 28930 9003 28933
rect 7668 28928 9003 28930
rect 7668 28872 8942 28928
rect 8998 28872 9003 28928
rect 7668 28870 9003 28872
rect 7668 28868 7674 28870
rect 8937 28867 9003 28870
rect 10225 28930 10291 28933
rect 12433 28930 12499 28933
rect 10225 28928 12499 28930
rect 10225 28872 10230 28928
rect 10286 28872 12438 28928
rect 12494 28872 12499 28928
rect 10225 28870 12499 28872
rect 10225 28867 10291 28870
rect 12433 28867 12499 28870
rect 20897 28930 20963 28933
rect 22050 28930 22110 29142
rect 23749 29139 23815 29142
rect 28901 29139 28967 29142
rect 22185 29066 22251 29069
rect 22645 29066 22711 29069
rect 22185 29064 22711 29066
rect 22185 29008 22190 29064
rect 22246 29008 22650 29064
rect 22706 29008 22711 29064
rect 22185 29006 22711 29008
rect 22185 29003 22251 29006
rect 22645 29003 22711 29006
rect 23105 29066 23171 29069
rect 24761 29066 24827 29069
rect 25313 29066 25379 29069
rect 23105 29064 25379 29066
rect 23105 29008 23110 29064
rect 23166 29008 24766 29064
rect 24822 29008 25318 29064
rect 25374 29008 25379 29064
rect 23105 29006 25379 29008
rect 23105 29003 23171 29006
rect 24761 29003 24827 29006
rect 25313 29003 25379 29006
rect 26785 29066 26851 29069
rect 27245 29066 27311 29069
rect 26785 29064 27311 29066
rect 26785 29008 26790 29064
rect 26846 29008 27250 29064
rect 27306 29008 27311 29064
rect 26785 29006 27311 29008
rect 26785 29003 26851 29006
rect 27245 29003 27311 29006
rect 29821 29066 29887 29069
rect 30790 29066 30850 29142
rect 32397 29139 32463 29142
rect 29821 29064 30850 29066
rect 29821 29008 29826 29064
rect 29882 29008 30850 29064
rect 29821 29006 30850 29008
rect 31109 29066 31175 29069
rect 31569 29068 31635 29069
rect 31518 29066 31524 29068
rect 31109 29064 31524 29066
rect 31588 29066 31635 29068
rect 32397 29068 32463 29069
rect 32397 29066 32444 29068
rect 31588 29064 31680 29066
rect 31109 29008 31114 29064
rect 31170 29008 31524 29064
rect 31630 29008 31680 29064
rect 31109 29006 31524 29008
rect 29821 29003 29887 29006
rect 31109 29003 31175 29006
rect 31518 29004 31524 29006
rect 31588 29006 31680 29008
rect 32352 29064 32444 29066
rect 32352 29008 32402 29064
rect 32352 29006 32444 29008
rect 31588 29004 31635 29006
rect 31569 29003 31635 29004
rect 32397 29004 32444 29006
rect 32508 29004 32514 29068
rect 32397 29003 32463 29004
rect 20897 28928 22110 28930
rect 20897 28872 20902 28928
rect 20958 28872 22110 28928
rect 20897 28870 22110 28872
rect 31385 28930 31451 28933
rect 32857 28930 32923 28933
rect 31385 28928 32923 28930
rect 31385 28872 31390 28928
rect 31446 28872 32862 28928
rect 32918 28872 32923 28928
rect 31385 28870 32923 28872
rect 20897 28867 20963 28870
rect 31385 28867 31451 28870
rect 32857 28867 32923 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 31845 28794 31911 28797
rect 33133 28794 33199 28797
rect 31845 28792 33199 28794
rect 31845 28736 31850 28792
rect 31906 28736 33138 28792
rect 33194 28736 33199 28792
rect 31845 28734 33199 28736
rect 31845 28731 31911 28734
rect 33133 28731 33199 28734
rect 9673 28658 9739 28661
rect 10225 28658 10291 28661
rect 10358 28658 10364 28660
rect 9673 28656 10364 28658
rect 9673 28600 9678 28656
rect 9734 28600 10230 28656
rect 10286 28600 10364 28656
rect 9673 28598 10364 28600
rect 9673 28595 9739 28598
rect 10225 28595 10291 28598
rect 10358 28596 10364 28598
rect 10428 28596 10434 28660
rect 11513 28658 11579 28661
rect 12525 28658 12591 28661
rect 11513 28656 12591 28658
rect 11513 28600 11518 28656
rect 11574 28600 12530 28656
rect 12586 28600 12591 28656
rect 11513 28598 12591 28600
rect 11513 28595 11579 28598
rect 12525 28595 12591 28598
rect 16849 28658 16915 28661
rect 21725 28658 21791 28661
rect 16849 28656 21791 28658
rect 16849 28600 16854 28656
rect 16910 28600 21730 28656
rect 21786 28600 21791 28656
rect 16849 28598 21791 28600
rect 16849 28595 16915 28598
rect 21725 28595 21791 28598
rect 31937 28658 32003 28661
rect 33685 28658 33751 28661
rect 31937 28656 33751 28658
rect 31937 28600 31942 28656
rect 31998 28600 33690 28656
rect 33746 28600 33751 28656
rect 31937 28598 33751 28600
rect 31937 28595 32003 28598
rect 33685 28595 33751 28598
rect 16941 28522 17007 28525
rect 17769 28522 17835 28525
rect 16941 28520 17835 28522
rect 16941 28464 16946 28520
rect 17002 28464 17774 28520
rect 17830 28464 17835 28520
rect 16941 28462 17835 28464
rect 16941 28459 17007 28462
rect 17769 28459 17835 28462
rect 23105 28522 23171 28525
rect 23105 28520 23306 28522
rect 23105 28464 23110 28520
rect 23166 28464 23306 28520
rect 23105 28462 23306 28464
rect 23105 28459 23171 28462
rect 17217 28388 17283 28389
rect 23246 28388 23306 28462
rect 23422 28460 23428 28524
rect 23492 28522 23498 28524
rect 26509 28522 26575 28525
rect 23492 28520 26575 28522
rect 23492 28464 26514 28520
rect 26570 28464 26575 28520
rect 23492 28462 26575 28464
rect 23492 28460 23498 28462
rect 26509 28459 26575 28462
rect 31569 28522 31635 28525
rect 32673 28522 32739 28525
rect 31569 28520 32739 28522
rect 31569 28464 31574 28520
rect 31630 28464 32678 28520
rect 32734 28464 32739 28520
rect 31569 28462 32739 28464
rect 31569 28459 31635 28462
rect 32673 28459 32739 28462
rect 17166 28324 17172 28388
rect 17236 28386 17283 28388
rect 17236 28384 17328 28386
rect 17278 28328 17328 28384
rect 17236 28326 17328 28328
rect 17236 28324 17283 28326
rect 23238 28324 23244 28388
rect 23308 28386 23314 28388
rect 23381 28386 23447 28389
rect 23308 28384 23447 28386
rect 23308 28328 23386 28384
rect 23442 28328 23447 28384
rect 23308 28326 23447 28328
rect 23308 28324 23314 28326
rect 17217 28323 17283 28324
rect 23381 28323 23447 28326
rect 31385 28386 31451 28389
rect 32070 28386 32076 28388
rect 31385 28384 32076 28386
rect 31385 28328 31390 28384
rect 31446 28328 32076 28384
rect 31385 28326 32076 28328
rect 31385 28323 31451 28326
rect 32070 28324 32076 28326
rect 32140 28324 32146 28388
rect 32305 28386 32371 28389
rect 33133 28386 33199 28389
rect 32305 28384 33199 28386
rect 32305 28328 32310 28384
rect 32366 28328 33138 28384
rect 33194 28328 33199 28384
rect 32305 28326 33199 28328
rect 32305 28323 32371 28326
rect 33133 28323 33199 28326
rect 33358 28324 33364 28388
rect 33428 28386 33434 28388
rect 33869 28386 33935 28389
rect 34329 28386 34395 28389
rect 33428 28384 34395 28386
rect 33428 28328 33874 28384
rect 33930 28328 34334 28384
rect 34390 28328 34395 28384
rect 33428 28326 34395 28328
rect 33428 28324 33434 28326
rect 33869 28323 33935 28326
rect 34329 28323 34395 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 8518 28188 8524 28252
rect 8588 28250 8594 28252
rect 18137 28250 18203 28253
rect 8588 28248 18203 28250
rect 8588 28192 18142 28248
rect 18198 28192 18203 28248
rect 8588 28190 18203 28192
rect 8588 28188 8594 28190
rect 18137 28187 18203 28190
rect 19701 28250 19767 28253
rect 21081 28250 21147 28253
rect 26325 28250 26391 28253
rect 26550 28250 26556 28252
rect 19701 28248 26556 28250
rect 19701 28192 19706 28248
rect 19762 28192 21086 28248
rect 21142 28192 26330 28248
rect 26386 28192 26556 28248
rect 19701 28190 26556 28192
rect 19701 28187 19767 28190
rect 21081 28187 21147 28190
rect 26325 28187 26391 28190
rect 26550 28188 26556 28190
rect 26620 28188 26626 28252
rect 29177 28250 29243 28253
rect 30005 28250 30071 28253
rect 31293 28250 31359 28253
rect 33409 28250 33475 28253
rect 29177 28248 31218 28250
rect 29177 28192 29182 28248
rect 29238 28192 30010 28248
rect 30066 28192 31218 28248
rect 29177 28190 31218 28192
rect 29177 28187 29243 28190
rect 30005 28187 30071 28190
rect 4153 28114 4219 28117
rect 4981 28114 5047 28117
rect 4153 28112 5047 28114
rect 4153 28056 4158 28112
rect 4214 28056 4986 28112
rect 5042 28056 5047 28112
rect 4153 28054 5047 28056
rect 4153 28051 4219 28054
rect 4981 28051 5047 28054
rect 16113 28114 16179 28117
rect 17677 28114 17743 28117
rect 17953 28114 18019 28117
rect 16113 28112 18019 28114
rect 16113 28056 16118 28112
rect 16174 28056 17682 28112
rect 17738 28056 17958 28112
rect 18014 28056 18019 28112
rect 16113 28054 18019 28056
rect 16113 28051 16179 28054
rect 17677 28051 17743 28054
rect 17953 28051 18019 28054
rect 24301 28114 24367 28117
rect 26182 28114 26188 28116
rect 24301 28112 26188 28114
rect 24301 28056 24306 28112
rect 24362 28056 26188 28112
rect 24301 28054 26188 28056
rect 24301 28051 24367 28054
rect 26182 28052 26188 28054
rect 26252 28114 26258 28116
rect 30097 28114 30163 28117
rect 26252 28112 30163 28114
rect 26252 28056 30102 28112
rect 30158 28056 30163 28112
rect 26252 28054 30163 28056
rect 31158 28114 31218 28190
rect 31293 28248 33475 28250
rect 31293 28192 31298 28248
rect 31354 28192 33414 28248
rect 33470 28192 33475 28248
rect 31293 28190 33475 28192
rect 31293 28187 31359 28190
rect 33409 28187 33475 28190
rect 31661 28114 31727 28117
rect 31158 28112 31727 28114
rect 31158 28056 31666 28112
rect 31722 28056 31727 28112
rect 31158 28054 31727 28056
rect 26252 28052 26258 28054
rect 30097 28051 30163 28054
rect 31661 28051 31727 28054
rect 32070 28052 32076 28116
rect 32140 28114 32146 28116
rect 32673 28114 32739 28117
rect 33041 28114 33107 28117
rect 35065 28114 35131 28117
rect 32140 28112 35131 28114
rect 32140 28056 32678 28112
rect 32734 28056 33046 28112
rect 33102 28056 35070 28112
rect 35126 28056 35131 28112
rect 32140 28054 35131 28056
rect 32140 28052 32146 28054
rect 32673 28051 32739 28054
rect 33041 28051 33107 28054
rect 35065 28051 35131 28054
rect 17217 27978 17283 27981
rect 17350 27978 17356 27980
rect 17217 27976 17356 27978
rect 17217 27920 17222 27976
rect 17278 27920 17356 27976
rect 17217 27918 17356 27920
rect 17217 27915 17283 27918
rect 17350 27916 17356 27918
rect 17420 27978 17426 27980
rect 18965 27978 19031 27981
rect 17420 27976 19031 27978
rect 17420 27920 18970 27976
rect 19026 27920 19031 27976
rect 17420 27918 19031 27920
rect 17420 27916 17426 27918
rect 18965 27915 19031 27918
rect 30005 27978 30071 27981
rect 30925 27978 30991 27981
rect 35433 27978 35499 27981
rect 30005 27976 35499 27978
rect 30005 27920 30010 27976
rect 30066 27920 30930 27976
rect 30986 27920 35438 27976
rect 35494 27920 35499 27976
rect 30005 27918 35499 27920
rect 30005 27915 30071 27918
rect 30925 27915 30991 27918
rect 35433 27915 35499 27918
rect 29913 27842 29979 27845
rect 30649 27842 30715 27845
rect 29913 27840 30715 27842
rect 29913 27784 29918 27840
rect 29974 27784 30654 27840
rect 30710 27784 30715 27840
rect 29913 27782 30715 27784
rect 29913 27779 29979 27782
rect 30649 27779 30715 27782
rect 31569 27842 31635 27845
rect 33869 27842 33935 27845
rect 31569 27840 33935 27842
rect 31569 27784 31574 27840
rect 31630 27784 33874 27840
rect 33930 27784 33935 27840
rect 31569 27782 33935 27784
rect 31569 27779 31635 27782
rect 33869 27779 33935 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 10317 27706 10383 27709
rect 15837 27706 15903 27709
rect 16757 27706 16823 27709
rect 10317 27704 16823 27706
rect 10317 27648 10322 27704
rect 10378 27648 15842 27704
rect 15898 27648 16762 27704
rect 16818 27648 16823 27704
rect 10317 27646 16823 27648
rect 10317 27643 10383 27646
rect 15837 27643 15903 27646
rect 16757 27643 16823 27646
rect 22921 27706 22987 27709
rect 24209 27706 24275 27709
rect 22921 27704 24275 27706
rect 22921 27648 22926 27704
rect 22982 27648 24214 27704
rect 24270 27648 24275 27704
rect 22921 27646 24275 27648
rect 22921 27643 22987 27646
rect 24209 27643 24275 27646
rect 30373 27706 30439 27709
rect 33685 27706 33751 27709
rect 30373 27704 33751 27706
rect 30373 27648 30378 27704
rect 30434 27648 33690 27704
rect 33746 27648 33751 27704
rect 30373 27646 33751 27648
rect 30373 27643 30439 27646
rect 33685 27643 33751 27646
rect 9765 27570 9831 27573
rect 12525 27570 12591 27573
rect 15009 27570 15075 27573
rect 16849 27570 16915 27573
rect 28257 27570 28323 27573
rect 9765 27568 13922 27570
rect 9765 27512 9770 27568
rect 9826 27512 12530 27568
rect 12586 27512 13922 27568
rect 9765 27510 13922 27512
rect 9765 27507 9831 27510
rect 12525 27507 12591 27510
rect 13629 27436 13695 27437
rect 13629 27434 13676 27436
rect 13584 27432 13676 27434
rect 13584 27376 13634 27432
rect 13584 27374 13676 27376
rect 13629 27372 13676 27374
rect 13740 27372 13746 27436
rect 13862 27434 13922 27510
rect 15009 27568 16915 27570
rect 15009 27512 15014 27568
rect 15070 27512 16854 27568
rect 16910 27512 16915 27568
rect 15009 27510 16915 27512
rect 15009 27507 15075 27510
rect 16849 27507 16915 27510
rect 22050 27568 28323 27570
rect 22050 27512 28262 27568
rect 28318 27512 28323 27568
rect 22050 27510 28323 27512
rect 16757 27434 16823 27437
rect 22050 27434 22110 27510
rect 28257 27507 28323 27510
rect 29453 27570 29519 27573
rect 35249 27570 35315 27573
rect 36077 27570 36143 27573
rect 29453 27568 36143 27570
rect 29453 27512 29458 27568
rect 29514 27512 35254 27568
rect 35310 27512 36082 27568
rect 36138 27512 36143 27568
rect 29453 27510 36143 27512
rect 29453 27507 29519 27510
rect 35249 27507 35315 27510
rect 36077 27507 36143 27510
rect 13862 27432 22110 27434
rect 13862 27376 16762 27432
rect 16818 27376 22110 27432
rect 13862 27374 22110 27376
rect 23013 27434 23079 27437
rect 25773 27434 25839 27437
rect 23013 27432 25839 27434
rect 23013 27376 23018 27432
rect 23074 27376 25778 27432
rect 25834 27376 25839 27432
rect 23013 27374 25839 27376
rect 13629 27371 13695 27372
rect 16757 27371 16823 27374
rect 23013 27371 23079 27374
rect 25773 27371 25839 27374
rect 28993 27434 29059 27437
rect 29913 27434 29979 27437
rect 28993 27432 29979 27434
rect 28993 27376 28998 27432
rect 29054 27376 29918 27432
rect 29974 27376 29979 27432
rect 28993 27374 29979 27376
rect 28993 27371 29059 27374
rect 29913 27371 29979 27374
rect 30414 27372 30420 27436
rect 30484 27434 30490 27436
rect 32489 27434 32555 27437
rect 30484 27432 32555 27434
rect 30484 27376 32494 27432
rect 32550 27376 32555 27432
rect 30484 27374 32555 27376
rect 30484 27372 30490 27374
rect 32489 27371 32555 27374
rect 10041 27298 10107 27301
rect 14089 27298 14155 27301
rect 10041 27296 14155 27298
rect 10041 27240 10046 27296
rect 10102 27240 14094 27296
rect 14150 27240 14155 27296
rect 10041 27238 14155 27240
rect 10041 27235 10107 27238
rect 14089 27235 14155 27238
rect 16389 27298 16455 27301
rect 17309 27298 17375 27301
rect 16389 27296 17375 27298
rect 16389 27240 16394 27296
rect 16450 27240 17314 27296
rect 17370 27240 17375 27296
rect 16389 27238 17375 27240
rect 16389 27235 16455 27238
rect 17309 27235 17375 27238
rect 19425 27298 19491 27301
rect 20805 27298 20871 27301
rect 25589 27298 25655 27301
rect 19425 27296 25655 27298
rect 19425 27240 19430 27296
rect 19486 27240 20810 27296
rect 20866 27240 25594 27296
rect 25650 27240 25655 27296
rect 19425 27238 25655 27240
rect 19425 27235 19491 27238
rect 20805 27235 20871 27238
rect 25589 27235 25655 27238
rect 36169 27298 36235 27301
rect 36895 27298 37695 27328
rect 36169 27296 37695 27298
rect 36169 27240 36174 27296
rect 36230 27240 37695 27296
rect 36169 27238 37695 27240
rect 36169 27235 36235 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 36895 27208 37695 27238
rect 35590 27167 35906 27168
rect 10041 27162 10107 27165
rect 10961 27162 11027 27165
rect 10041 27160 11027 27162
rect 10041 27104 10046 27160
rect 10102 27104 10966 27160
rect 11022 27104 11027 27160
rect 10041 27102 11027 27104
rect 10041 27099 10107 27102
rect 10961 27099 11027 27102
rect 12985 27162 13051 27165
rect 13261 27162 13327 27165
rect 29269 27162 29335 27165
rect 29637 27162 29703 27165
rect 12985 27160 13968 27162
rect 12985 27104 12990 27160
rect 13046 27104 13266 27160
rect 13322 27104 13968 27160
rect 12985 27102 13968 27104
rect 12985 27099 13051 27102
rect 13261 27099 13327 27102
rect 13908 27029 13968 27102
rect 29269 27160 29703 27162
rect 29269 27104 29274 27160
rect 29330 27104 29642 27160
rect 29698 27104 29703 27160
rect 29269 27102 29703 27104
rect 29269 27099 29335 27102
rect 29637 27099 29703 27102
rect 3141 27026 3207 27029
rect 13537 27026 13603 27029
rect 3141 27024 13603 27026
rect 3141 26968 3146 27024
rect 3202 26968 13542 27024
rect 13598 26968 13603 27024
rect 3141 26966 13603 26968
rect 3141 26963 3207 26966
rect 13537 26963 13603 26966
rect 13905 27024 13971 27029
rect 13905 26968 13910 27024
rect 13966 26968 13971 27024
rect 13905 26963 13971 26968
rect 22553 27026 22619 27029
rect 24301 27026 24367 27029
rect 25221 27026 25287 27029
rect 26049 27026 26115 27029
rect 26693 27026 26759 27029
rect 22553 27024 26759 27026
rect 22553 26968 22558 27024
rect 22614 26968 24306 27024
rect 24362 26968 25226 27024
rect 25282 26968 26054 27024
rect 26110 26968 26698 27024
rect 26754 26968 26759 27024
rect 22553 26966 26759 26968
rect 22553 26963 22619 26966
rect 24301 26963 24367 26966
rect 25221 26963 25287 26966
rect 26049 26963 26115 26966
rect 26693 26963 26759 26966
rect 33685 27026 33751 27029
rect 35065 27026 35131 27029
rect 33685 27024 35131 27026
rect 33685 26968 33690 27024
rect 33746 26968 35070 27024
rect 35126 26968 35131 27024
rect 33685 26966 35131 26968
rect 33685 26963 33751 26966
rect 35065 26963 35131 26966
rect 6821 26890 6887 26893
rect 8845 26890 8911 26893
rect 6821 26888 8911 26890
rect 6821 26832 6826 26888
rect 6882 26832 8850 26888
rect 8906 26832 8911 26888
rect 6821 26830 8911 26832
rect 6821 26827 6887 26830
rect 8845 26827 8911 26830
rect 10133 26890 10199 26893
rect 10317 26890 10383 26893
rect 10685 26890 10751 26893
rect 11145 26890 11211 26893
rect 10133 26888 10751 26890
rect 10133 26832 10138 26888
rect 10194 26832 10322 26888
rect 10378 26832 10690 26888
rect 10746 26832 10751 26888
rect 10133 26830 10751 26832
rect 10133 26827 10199 26830
rect 10317 26827 10383 26830
rect 10685 26827 10751 26830
rect 10964 26888 11211 26890
rect 10964 26832 11150 26888
rect 11206 26832 11211 26888
rect 10964 26830 11211 26832
rect 10964 26757 11024 26830
rect 11145 26827 11211 26830
rect 12617 26890 12683 26893
rect 13486 26890 13492 26892
rect 12617 26888 13492 26890
rect 12617 26832 12622 26888
rect 12678 26832 13492 26888
rect 12617 26830 13492 26832
rect 12617 26827 12683 26830
rect 13486 26828 13492 26830
rect 13556 26828 13562 26892
rect 30097 26890 30163 26893
rect 34513 26890 34579 26893
rect 30097 26888 34579 26890
rect 30097 26832 30102 26888
rect 30158 26832 34518 26888
rect 34574 26832 34579 26888
rect 30097 26830 34579 26832
rect 30097 26827 30163 26830
rect 34513 26827 34579 26830
rect 10961 26752 11027 26757
rect 10961 26696 10966 26752
rect 11022 26696 11027 26752
rect 10961 26691 11027 26696
rect 11145 26754 11211 26757
rect 15009 26754 15075 26757
rect 18137 26756 18203 26757
rect 11145 26752 15075 26754
rect 11145 26696 11150 26752
rect 11206 26696 15014 26752
rect 15070 26696 15075 26752
rect 11145 26694 15075 26696
rect 11145 26691 11211 26694
rect 15009 26691 15075 26694
rect 18086 26692 18092 26756
rect 18156 26754 18203 26756
rect 21909 26754 21975 26757
rect 23841 26754 23907 26757
rect 18156 26752 18248 26754
rect 18198 26696 18248 26752
rect 18156 26694 18248 26696
rect 21909 26752 23907 26754
rect 21909 26696 21914 26752
rect 21970 26696 23846 26752
rect 23902 26696 23907 26752
rect 21909 26694 23907 26696
rect 18156 26692 18203 26694
rect 18137 26691 18203 26692
rect 21909 26691 21975 26694
rect 23841 26691 23907 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 12525 26618 12591 26621
rect 13721 26618 13787 26621
rect 36261 26618 36327 26621
rect 36895 26618 37695 26648
rect 12525 26616 20178 26618
rect 12525 26560 12530 26616
rect 12586 26560 13726 26616
rect 13782 26560 20178 26616
rect 12525 26558 20178 26560
rect 12525 26555 12591 26558
rect 13721 26555 13787 26558
rect 11053 26482 11119 26485
rect 12801 26482 12867 26485
rect 14641 26482 14707 26485
rect 11053 26480 14707 26482
rect 11053 26424 11058 26480
rect 11114 26424 12806 26480
rect 12862 26424 14646 26480
rect 14702 26424 14707 26480
rect 11053 26422 14707 26424
rect 11053 26419 11119 26422
rect 12801 26419 12867 26422
rect 14641 26419 14707 26422
rect 19006 26420 19012 26484
rect 19076 26482 19082 26484
rect 19977 26482 20043 26485
rect 19076 26480 20043 26482
rect 19076 26424 19982 26480
rect 20038 26424 20043 26480
rect 19076 26422 20043 26424
rect 20118 26482 20178 26558
rect 36261 26616 37695 26618
rect 36261 26560 36266 26616
rect 36322 26560 37695 26616
rect 36261 26558 37695 26560
rect 36261 26555 36327 26558
rect 36895 26528 37695 26558
rect 28257 26482 28323 26485
rect 20118 26480 28323 26482
rect 20118 26424 28262 26480
rect 28318 26424 28323 26480
rect 20118 26422 28323 26424
rect 19076 26420 19082 26422
rect 19977 26419 20043 26422
rect 28257 26419 28323 26422
rect 13261 26346 13327 26349
rect 13905 26346 13971 26349
rect 14365 26346 14431 26349
rect 24301 26346 24367 26349
rect 13261 26344 13784 26346
rect 13261 26288 13266 26344
rect 13322 26288 13784 26344
rect 13261 26286 13784 26288
rect 13261 26283 13327 26286
rect 9949 26210 10015 26213
rect 13261 26210 13327 26213
rect 9949 26208 13327 26210
rect 9949 26152 9954 26208
rect 10010 26152 13266 26208
rect 13322 26152 13327 26208
rect 9949 26150 13327 26152
rect 13724 26210 13784 26286
rect 13905 26344 24367 26346
rect 13905 26288 13910 26344
rect 13966 26288 14370 26344
rect 14426 26288 24306 26344
rect 24362 26288 24367 26344
rect 13905 26286 24367 26288
rect 13905 26283 13971 26286
rect 14365 26283 14431 26286
rect 24301 26283 24367 26286
rect 24526 26284 24532 26348
rect 24596 26346 24602 26348
rect 24669 26346 24735 26349
rect 24596 26344 24735 26346
rect 24596 26288 24674 26344
rect 24730 26288 24735 26344
rect 24596 26286 24735 26288
rect 24596 26284 24602 26286
rect 24669 26283 24735 26286
rect 24894 26284 24900 26348
rect 24964 26346 24970 26348
rect 25681 26346 25747 26349
rect 24964 26344 25747 26346
rect 24964 26288 25686 26344
rect 25742 26288 25747 26344
rect 24964 26286 25747 26288
rect 24964 26284 24970 26286
rect 25681 26283 25747 26286
rect 31017 26346 31083 26349
rect 33777 26346 33843 26349
rect 35709 26346 35775 26349
rect 31017 26344 35775 26346
rect 31017 26288 31022 26344
rect 31078 26288 33782 26344
rect 33838 26288 35714 26344
rect 35770 26288 35775 26344
rect 31017 26286 35775 26288
rect 31017 26283 31083 26286
rect 33777 26283 33843 26286
rect 35709 26283 35775 26286
rect 17401 26210 17467 26213
rect 17769 26210 17835 26213
rect 13724 26208 17835 26210
rect 13724 26152 17406 26208
rect 17462 26152 17774 26208
rect 17830 26152 17835 26208
rect 13724 26150 17835 26152
rect 9949 26147 10015 26150
rect 13261 26147 13327 26150
rect 17401 26147 17467 26150
rect 17769 26147 17835 26150
rect 20110 26148 20116 26212
rect 20180 26210 20186 26212
rect 20621 26210 20687 26213
rect 20180 26208 20687 26210
rect 20180 26152 20626 26208
rect 20682 26152 20687 26208
rect 20180 26150 20687 26152
rect 20180 26148 20186 26150
rect 20621 26147 20687 26150
rect 28942 26148 28948 26212
rect 29012 26210 29018 26212
rect 29177 26210 29243 26213
rect 35157 26210 35223 26213
rect 29012 26208 35223 26210
rect 29012 26152 29182 26208
rect 29238 26152 35162 26208
rect 35218 26152 35223 26208
rect 29012 26150 35223 26152
rect 29012 26148 29018 26150
rect 29177 26147 29243 26150
rect 35157 26147 35223 26150
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 8753 26074 8819 26077
rect 12525 26074 12591 26077
rect 8753 26072 12591 26074
rect 8753 26016 8758 26072
rect 8814 26016 12530 26072
rect 12586 26016 12591 26072
rect 8753 26014 12591 26016
rect 8753 26011 8819 26014
rect 12525 26011 12591 26014
rect 29913 26074 29979 26077
rect 30925 26074 30991 26077
rect 29913 26072 30991 26074
rect 29913 26016 29918 26072
rect 29974 26016 30930 26072
rect 30986 26016 30991 26072
rect 29913 26014 30991 26016
rect 29913 26011 29979 26014
rect 30925 26011 30991 26014
rect 32029 26074 32095 26077
rect 34329 26074 34395 26077
rect 32029 26072 34395 26074
rect 32029 26016 32034 26072
rect 32090 26016 34334 26072
rect 34390 26016 34395 26072
rect 32029 26014 34395 26016
rect 32029 26011 32095 26014
rect 34329 26011 34395 26014
rect 5993 25938 6059 25941
rect 7833 25938 7899 25941
rect 20110 25938 20116 25940
rect 5993 25936 20116 25938
rect 5993 25880 5998 25936
rect 6054 25880 7838 25936
rect 7894 25880 20116 25936
rect 5993 25878 20116 25880
rect 5993 25875 6059 25878
rect 7833 25875 7899 25878
rect 20110 25876 20116 25878
rect 20180 25876 20186 25940
rect 21541 25938 21607 25941
rect 23657 25938 23723 25941
rect 21541 25936 23723 25938
rect 21541 25880 21546 25936
rect 21602 25880 23662 25936
rect 23718 25880 23723 25936
rect 21541 25878 23723 25880
rect 21541 25875 21607 25878
rect 23657 25875 23723 25878
rect 25957 25938 26023 25941
rect 31518 25938 31524 25940
rect 25957 25936 31524 25938
rect 25957 25880 25962 25936
rect 26018 25880 31524 25936
rect 25957 25878 31524 25880
rect 25957 25875 26023 25878
rect 31518 25876 31524 25878
rect 31588 25876 31594 25940
rect 32254 25876 32260 25940
rect 32324 25938 32330 25940
rect 33041 25938 33107 25941
rect 32324 25936 33107 25938
rect 32324 25880 33046 25936
rect 33102 25880 33107 25936
rect 32324 25878 33107 25880
rect 32324 25876 32330 25878
rect 33041 25875 33107 25878
rect 36169 25938 36235 25941
rect 36895 25938 37695 25968
rect 36169 25936 37695 25938
rect 36169 25880 36174 25936
rect 36230 25880 37695 25936
rect 36169 25878 37695 25880
rect 36169 25875 36235 25878
rect 36895 25848 37695 25878
rect 9213 25802 9279 25805
rect 16021 25802 16087 25805
rect 9213 25800 16087 25802
rect 9213 25744 9218 25800
rect 9274 25744 16026 25800
rect 16082 25744 16087 25800
rect 9213 25742 16087 25744
rect 9213 25739 9279 25742
rect 16021 25739 16087 25742
rect 19977 25802 20043 25805
rect 25129 25802 25195 25805
rect 19977 25800 25195 25802
rect 19977 25744 19982 25800
rect 20038 25744 25134 25800
rect 25190 25744 25195 25800
rect 19977 25742 25195 25744
rect 19977 25739 20043 25742
rect 25129 25739 25195 25742
rect 33133 25802 33199 25805
rect 34237 25802 34303 25805
rect 33133 25800 34303 25802
rect 33133 25744 33138 25800
rect 33194 25744 34242 25800
rect 34298 25744 34303 25800
rect 33133 25742 34303 25744
rect 33133 25739 33199 25742
rect 34237 25739 34303 25742
rect 12065 25666 12131 25669
rect 12341 25666 12407 25669
rect 16389 25666 16455 25669
rect 12065 25664 16455 25666
rect 12065 25608 12070 25664
rect 12126 25608 12346 25664
rect 12402 25608 16394 25664
rect 16450 25608 16455 25664
rect 12065 25606 16455 25608
rect 12065 25603 12131 25606
rect 12341 25603 12407 25606
rect 16389 25603 16455 25606
rect 28901 25666 28967 25669
rect 33317 25666 33383 25669
rect 33685 25666 33751 25669
rect 28901 25664 33751 25666
rect 28901 25608 28906 25664
rect 28962 25608 33322 25664
rect 33378 25608 33690 25664
rect 33746 25608 33751 25664
rect 28901 25606 33751 25608
rect 28901 25603 28967 25606
rect 33317 25603 33383 25606
rect 33685 25603 33751 25606
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 8477 25532 8543 25533
rect 8477 25530 8524 25532
rect 8432 25528 8524 25530
rect 8432 25472 8482 25528
rect 8432 25470 8524 25472
rect 8477 25468 8524 25470
rect 8588 25468 8594 25532
rect 10777 25530 10843 25533
rect 11513 25530 11579 25533
rect 10777 25528 11579 25530
rect 10777 25472 10782 25528
rect 10838 25472 11518 25528
rect 11574 25472 11579 25528
rect 10777 25470 11579 25472
rect 8477 25467 8543 25468
rect 10777 25467 10843 25470
rect 11513 25467 11579 25470
rect 16573 25532 16639 25533
rect 16573 25528 16620 25532
rect 16684 25530 16690 25532
rect 30649 25530 30715 25533
rect 30925 25530 30991 25533
rect 33409 25530 33475 25533
rect 16573 25472 16578 25528
rect 16573 25468 16620 25472
rect 16684 25470 16730 25530
rect 30649 25528 33475 25530
rect 30649 25472 30654 25528
rect 30710 25472 30930 25528
rect 30986 25472 33414 25528
rect 33470 25472 33475 25528
rect 30649 25470 33475 25472
rect 16684 25468 16690 25470
rect 16573 25467 16639 25468
rect 30649 25467 30715 25470
rect 30925 25467 30991 25470
rect 33409 25467 33475 25470
rect 35382 25468 35388 25532
rect 35452 25530 35458 25532
rect 35801 25530 35867 25533
rect 35452 25528 35867 25530
rect 35452 25472 35806 25528
rect 35862 25472 35867 25528
rect 35452 25470 35867 25472
rect 35452 25468 35458 25470
rect 11605 25394 11671 25397
rect 18137 25394 18203 25397
rect 27061 25394 27127 25397
rect 35157 25394 35223 25397
rect 35390 25394 35450 25468
rect 35801 25467 35867 25470
rect 11605 25392 18203 25394
rect 11605 25336 11610 25392
rect 11666 25336 18142 25392
rect 18198 25336 18203 25392
rect 11605 25334 18203 25336
rect 11605 25331 11671 25334
rect 18137 25331 18203 25334
rect 22050 25392 35450 25394
rect 22050 25336 27066 25392
rect 27122 25336 35162 25392
rect 35218 25336 35450 25392
rect 22050 25334 35450 25336
rect 16062 25196 16068 25260
rect 16132 25258 16138 25260
rect 22050 25258 22110 25334
rect 27061 25331 27127 25334
rect 35157 25331 35223 25334
rect 16132 25198 22110 25258
rect 31753 25258 31819 25261
rect 32029 25258 32095 25261
rect 31753 25256 32095 25258
rect 31753 25200 31758 25256
rect 31814 25200 32034 25256
rect 32090 25200 32095 25256
rect 31753 25198 32095 25200
rect 16132 25196 16138 25198
rect 31753 25195 31819 25198
rect 32029 25195 32095 25198
rect 32581 25258 32647 25261
rect 33685 25258 33751 25261
rect 32581 25256 33751 25258
rect 32581 25200 32586 25256
rect 32642 25200 33690 25256
rect 33746 25200 33751 25256
rect 32581 25198 33751 25200
rect 32581 25195 32647 25198
rect 33685 25195 33751 25198
rect 35709 25258 35775 25261
rect 36895 25258 37695 25288
rect 35709 25256 37695 25258
rect 35709 25200 35714 25256
rect 35770 25200 37695 25256
rect 35709 25198 37695 25200
rect 35709 25195 35775 25198
rect 36895 25168 37695 25198
rect 7741 25122 7807 25125
rect 16849 25122 16915 25125
rect 7741 25120 16915 25122
rect 7741 25064 7746 25120
rect 7802 25064 16854 25120
rect 16910 25064 16915 25120
rect 7741 25062 16915 25064
rect 7741 25059 7807 25062
rect 16849 25059 16915 25062
rect 22921 25122 22987 25125
rect 23054 25122 23060 25124
rect 22921 25120 23060 25122
rect 22921 25064 22926 25120
rect 22982 25064 23060 25120
rect 22921 25062 23060 25064
rect 22921 25059 22987 25062
rect 23054 25060 23060 25062
rect 23124 25060 23130 25124
rect 32213 25122 32279 25125
rect 33409 25122 33475 25125
rect 32213 25120 33475 25122
rect 32213 25064 32218 25120
rect 32274 25064 33414 25120
rect 33470 25064 33475 25120
rect 32213 25062 33475 25064
rect 32213 25059 32279 25062
rect 33409 25059 33475 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 14641 24986 14707 24989
rect 14774 24986 14780 24988
rect 14641 24984 14780 24986
rect 14641 24928 14646 24984
rect 14702 24928 14780 24984
rect 14641 24926 14780 24928
rect 14641 24923 14707 24926
rect 14774 24924 14780 24926
rect 14844 24924 14850 24988
rect 20621 24986 20687 24989
rect 20897 24986 20963 24989
rect 24761 24986 24827 24989
rect 20621 24984 24827 24986
rect 20621 24928 20626 24984
rect 20682 24928 20902 24984
rect 20958 24928 24766 24984
rect 24822 24928 24827 24984
rect 20621 24926 24827 24928
rect 20621 24923 20687 24926
rect 20897 24923 20963 24926
rect 24761 24923 24827 24926
rect 29269 24988 29335 24989
rect 29269 24984 29316 24988
rect 29380 24986 29386 24988
rect 32397 24986 32463 24989
rect 29269 24928 29274 24984
rect 29269 24924 29316 24928
rect 29380 24926 29426 24986
rect 32397 24984 32690 24986
rect 32397 24928 32402 24984
rect 32458 24928 32690 24984
rect 32397 24926 32690 24928
rect 29380 24924 29386 24926
rect 29269 24923 29335 24924
rect 32397 24923 32463 24926
rect 8385 24852 8451 24853
rect 8334 24850 8340 24852
rect 8294 24790 8340 24850
rect 8404 24848 8451 24852
rect 8446 24792 8451 24848
rect 8334 24788 8340 24790
rect 8404 24788 8451 24792
rect 8385 24787 8451 24788
rect 9673 24850 9739 24853
rect 12566 24850 12572 24852
rect 9673 24848 12572 24850
rect 9673 24792 9678 24848
rect 9734 24792 12572 24848
rect 9673 24790 12572 24792
rect 9673 24787 9739 24790
rect 12566 24788 12572 24790
rect 12636 24788 12642 24852
rect 19517 24850 19583 24853
rect 19701 24850 19767 24853
rect 21725 24850 21791 24853
rect 28441 24850 28507 24853
rect 31293 24852 31359 24853
rect 31293 24850 31340 24852
rect 19517 24848 28507 24850
rect 19517 24792 19522 24848
rect 19578 24792 19706 24848
rect 19762 24792 21730 24848
rect 21786 24792 28446 24848
rect 28502 24792 28507 24848
rect 19517 24790 28507 24792
rect 31248 24848 31340 24850
rect 31248 24792 31298 24848
rect 31248 24790 31340 24792
rect 19517 24787 19583 24790
rect 19701 24787 19767 24790
rect 21725 24787 21791 24790
rect 28441 24787 28507 24790
rect 31293 24788 31340 24790
rect 31404 24788 31410 24852
rect 31518 24788 31524 24852
rect 31588 24850 31594 24852
rect 32489 24850 32555 24853
rect 31588 24848 32555 24850
rect 31588 24792 32494 24848
rect 32550 24792 32555 24848
rect 31588 24790 32555 24792
rect 31588 24788 31594 24790
rect 31293 24787 31359 24788
rect 32489 24787 32555 24790
rect 32630 24850 32690 24926
rect 36261 24850 36327 24853
rect 32630 24848 36327 24850
rect 32630 24792 36266 24848
rect 36322 24792 36327 24848
rect 32630 24790 36327 24792
rect 21725 24714 21791 24717
rect 25221 24714 25287 24717
rect 21725 24712 25287 24714
rect 21725 24656 21730 24712
rect 21786 24656 25226 24712
rect 25282 24656 25287 24712
rect 21725 24654 25287 24656
rect 21725 24651 21791 24654
rect 25221 24651 25287 24654
rect 27889 24714 27955 24717
rect 32630 24714 32690 24790
rect 36261 24787 36327 24790
rect 27889 24712 32690 24714
rect 27889 24656 27894 24712
rect 27950 24656 32690 24712
rect 27889 24654 32690 24656
rect 27889 24651 27955 24654
rect 12525 24578 12591 24581
rect 13905 24578 13971 24581
rect 12525 24576 13971 24578
rect 12525 24520 12530 24576
rect 12586 24520 13910 24576
rect 13966 24520 13971 24576
rect 12525 24518 13971 24520
rect 12525 24515 12591 24518
rect 13905 24515 13971 24518
rect 36077 24578 36143 24581
rect 36895 24578 37695 24608
rect 36077 24576 37695 24578
rect 36077 24520 36082 24576
rect 36138 24520 37695 24576
rect 36077 24518 37695 24520
rect 36077 24515 36143 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 36895 24488 37695 24518
rect 34930 24447 35246 24448
rect 26417 24442 26483 24445
rect 31293 24442 31359 24445
rect 32070 24442 32076 24444
rect 26417 24440 32076 24442
rect 26417 24384 26422 24440
rect 26478 24384 31298 24440
rect 31354 24384 32076 24440
rect 26417 24382 32076 24384
rect 26417 24379 26483 24382
rect 31293 24379 31359 24382
rect 32070 24380 32076 24382
rect 32140 24380 32146 24444
rect 6913 24306 6979 24309
rect 10133 24308 10199 24309
rect 10133 24306 10180 24308
rect 6913 24304 10180 24306
rect 6913 24248 6918 24304
rect 6974 24248 10138 24304
rect 6913 24246 10180 24248
rect 6913 24243 6979 24246
rect 10133 24244 10180 24246
rect 10244 24244 10250 24308
rect 12617 24306 12683 24309
rect 15653 24306 15719 24309
rect 12617 24304 15719 24306
rect 12617 24248 12622 24304
rect 12678 24248 15658 24304
rect 15714 24248 15719 24304
rect 12617 24246 15719 24248
rect 10133 24243 10199 24244
rect 12617 24243 12683 24246
rect 15653 24243 15719 24246
rect 18965 24306 19031 24309
rect 20161 24306 20227 24309
rect 18965 24304 20227 24306
rect 18965 24248 18970 24304
rect 19026 24248 20166 24304
rect 20222 24248 20227 24304
rect 18965 24246 20227 24248
rect 18965 24243 19031 24246
rect 20161 24243 20227 24246
rect 28349 24306 28415 24309
rect 28758 24306 28764 24308
rect 28349 24304 28764 24306
rect 28349 24248 28354 24304
rect 28410 24248 28764 24304
rect 28349 24246 28764 24248
rect 28349 24243 28415 24246
rect 28758 24244 28764 24246
rect 28828 24244 28834 24308
rect 32765 24306 32831 24309
rect 33869 24306 33935 24309
rect 32765 24304 33935 24306
rect 32765 24248 32770 24304
rect 32826 24248 33874 24304
rect 33930 24248 33935 24304
rect 32765 24246 33935 24248
rect 32765 24243 32831 24246
rect 33869 24243 33935 24246
rect 6310 24108 6316 24172
rect 6380 24170 6386 24172
rect 6821 24170 6887 24173
rect 8569 24170 8635 24173
rect 6380 24168 8635 24170
rect 6380 24112 6826 24168
rect 6882 24112 8574 24168
rect 8630 24112 8635 24168
rect 6380 24110 8635 24112
rect 6380 24108 6386 24110
rect 6821 24107 6887 24110
rect 8569 24107 8635 24110
rect 11513 24170 11579 24173
rect 22369 24170 22435 24173
rect 11513 24168 22435 24170
rect 11513 24112 11518 24168
rect 11574 24112 22374 24168
rect 22430 24112 22435 24168
rect 11513 24110 22435 24112
rect 11513 24107 11579 24110
rect 22369 24107 22435 24110
rect 28349 24170 28415 24173
rect 28809 24170 28875 24173
rect 28349 24168 28875 24170
rect 28349 24112 28354 24168
rect 28410 24112 28814 24168
rect 28870 24112 28875 24168
rect 28349 24110 28875 24112
rect 28349 24107 28415 24110
rect 28809 24107 28875 24110
rect 29913 24170 29979 24173
rect 34973 24170 35039 24173
rect 29913 24168 35039 24170
rect 29913 24112 29918 24168
rect 29974 24112 34978 24168
rect 35034 24112 35039 24168
rect 29913 24110 35039 24112
rect 29913 24107 29979 24110
rect 34973 24107 35039 24110
rect 35525 24170 35591 24173
rect 35525 24168 36370 24170
rect 35525 24112 35530 24168
rect 35586 24112 36370 24168
rect 35525 24110 36370 24112
rect 35525 24107 35591 24110
rect 19057 24034 19123 24037
rect 20529 24034 20595 24037
rect 19057 24032 20595 24034
rect 19057 23976 19062 24032
rect 19118 23976 20534 24032
rect 20590 23976 20595 24032
rect 19057 23974 20595 23976
rect 19057 23971 19123 23974
rect 20529 23971 20595 23974
rect 24577 24034 24643 24037
rect 28717 24034 28783 24037
rect 24577 24032 28783 24034
rect 24577 23976 24582 24032
rect 24638 23976 28722 24032
rect 28778 23976 28783 24032
rect 24577 23974 28783 23976
rect 24577 23971 24643 23974
rect 28717 23971 28783 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 13813 23898 13879 23901
rect 17166 23898 17172 23900
rect 13813 23896 17172 23898
rect 13813 23840 13818 23896
rect 13874 23840 17172 23896
rect 13813 23838 17172 23840
rect 13813 23835 13879 23838
rect 17166 23836 17172 23838
rect 17236 23898 17242 23900
rect 27153 23898 27219 23901
rect 28942 23898 28948 23900
rect 17236 23896 28948 23898
rect 17236 23840 27158 23896
rect 27214 23840 28948 23896
rect 17236 23838 28948 23840
rect 17236 23836 17242 23838
rect 27153 23835 27219 23838
rect 28942 23836 28948 23838
rect 29012 23836 29018 23900
rect 36310 23898 36370 24110
rect 36895 23898 37695 23928
rect 36310 23838 37695 23898
rect 36895 23808 37695 23838
rect 5993 23764 6059 23765
rect 5942 23762 5948 23764
rect 5902 23702 5948 23762
rect 6012 23760 6059 23764
rect 6054 23704 6059 23760
rect 5942 23700 5948 23702
rect 6012 23700 6059 23704
rect 5993 23699 6059 23700
rect 10317 23762 10383 23765
rect 12341 23762 12407 23765
rect 10317 23760 12407 23762
rect 10317 23704 10322 23760
rect 10378 23704 12346 23760
rect 12402 23704 12407 23760
rect 10317 23702 12407 23704
rect 10317 23699 10383 23702
rect 12341 23699 12407 23702
rect 13670 23700 13676 23764
rect 13740 23762 13746 23764
rect 17953 23762 18019 23765
rect 13740 23760 18019 23762
rect 13740 23704 17958 23760
rect 18014 23704 18019 23760
rect 13740 23702 18019 23704
rect 13740 23700 13746 23702
rect 17953 23699 18019 23702
rect 19609 23762 19675 23765
rect 24485 23762 24551 23765
rect 19609 23760 24551 23762
rect 19609 23704 19614 23760
rect 19670 23704 24490 23760
rect 24546 23704 24551 23760
rect 19609 23702 24551 23704
rect 19609 23699 19675 23702
rect 24485 23699 24551 23702
rect 24945 23762 25011 23765
rect 25681 23762 25747 23765
rect 26049 23762 26115 23765
rect 24945 23760 31770 23762
rect 24945 23704 24950 23760
rect 25006 23704 25686 23760
rect 25742 23704 26054 23760
rect 26110 23704 31770 23760
rect 24945 23702 31770 23704
rect 24945 23699 25011 23702
rect 25681 23699 25747 23702
rect 26049 23699 26115 23702
rect 6453 23626 6519 23629
rect 9213 23626 9279 23629
rect 14089 23628 14155 23629
rect 6453 23624 9279 23626
rect 6453 23568 6458 23624
rect 6514 23568 9218 23624
rect 9274 23568 9279 23624
rect 6453 23566 9279 23568
rect 6453 23563 6519 23566
rect 9213 23563 9279 23566
rect 14038 23564 14044 23628
rect 14108 23626 14155 23628
rect 14108 23624 14200 23626
rect 14150 23568 14200 23624
rect 14108 23566 14200 23568
rect 14108 23564 14155 23566
rect 15326 23564 15332 23628
rect 15396 23626 15402 23628
rect 19609 23626 19675 23629
rect 15396 23624 19675 23626
rect 15396 23568 19614 23624
rect 19670 23568 19675 23624
rect 15396 23566 19675 23568
rect 15396 23564 15402 23566
rect 14089 23563 14155 23564
rect 19609 23563 19675 23566
rect 21357 23626 21423 23629
rect 22001 23626 22067 23629
rect 21357 23624 22067 23626
rect 21357 23568 21362 23624
rect 21418 23568 22006 23624
rect 22062 23568 22067 23624
rect 21357 23566 22067 23568
rect 21357 23563 21423 23566
rect 22001 23563 22067 23566
rect 22134 23564 22140 23628
rect 22204 23626 22210 23628
rect 22553 23626 22619 23629
rect 22204 23624 22619 23626
rect 22204 23568 22558 23624
rect 22614 23568 22619 23624
rect 22204 23566 22619 23568
rect 22204 23564 22210 23566
rect 22553 23563 22619 23566
rect 27838 23564 27844 23628
rect 27908 23626 27914 23628
rect 28073 23626 28139 23629
rect 27908 23624 28139 23626
rect 27908 23568 28078 23624
rect 28134 23568 28139 23624
rect 27908 23566 28139 23568
rect 31710 23626 31770 23702
rect 36445 23626 36511 23629
rect 31710 23624 36511 23626
rect 31710 23568 36450 23624
rect 36506 23568 36511 23624
rect 31710 23566 36511 23568
rect 27908 23564 27914 23566
rect 28073 23563 28139 23566
rect 36445 23563 36511 23566
rect 14641 23490 14707 23493
rect 16757 23492 16823 23493
rect 14958 23490 14964 23492
rect 14641 23488 14964 23490
rect 14641 23432 14646 23488
rect 14702 23432 14964 23488
rect 14641 23430 14964 23432
rect 14641 23427 14707 23430
rect 14958 23428 14964 23430
rect 15028 23428 15034 23492
rect 16757 23488 16804 23492
rect 16868 23490 16874 23492
rect 19333 23490 19399 23493
rect 20253 23490 20319 23493
rect 34053 23492 34119 23493
rect 16757 23432 16762 23488
rect 16757 23428 16804 23432
rect 16868 23430 16914 23490
rect 19333 23488 20319 23490
rect 19333 23432 19338 23488
rect 19394 23432 20258 23488
rect 20314 23432 20319 23488
rect 19333 23430 20319 23432
rect 16868 23428 16874 23430
rect 16757 23427 16823 23428
rect 19333 23427 19399 23430
rect 20253 23427 20319 23430
rect 28758 23428 28764 23492
rect 28828 23490 28834 23492
rect 29126 23490 29132 23492
rect 28828 23430 29132 23490
rect 28828 23428 28834 23430
rect 29126 23428 29132 23430
rect 29196 23428 29202 23492
rect 34053 23488 34100 23492
rect 34164 23490 34170 23492
rect 34053 23432 34058 23488
rect 34053 23428 34100 23432
rect 34164 23430 34210 23490
rect 34164 23428 34170 23430
rect 34053 23427 34119 23428
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 9673 23354 9739 23357
rect 9806 23354 9812 23356
rect 9673 23352 9812 23354
rect 9673 23296 9678 23352
rect 9734 23296 9812 23352
rect 9673 23294 9812 23296
rect 9673 23291 9739 23294
rect 9806 23292 9812 23294
rect 9876 23292 9882 23356
rect 16430 23292 16436 23356
rect 16500 23354 16506 23356
rect 18086 23354 18092 23356
rect 16500 23294 18092 23354
rect 16500 23292 16506 23294
rect 18086 23292 18092 23294
rect 18156 23292 18162 23356
rect 23197 23354 23263 23357
rect 26601 23354 26667 23357
rect 27337 23354 27403 23357
rect 23197 23352 27403 23354
rect 23197 23296 23202 23352
rect 23258 23296 26606 23352
rect 26662 23296 27342 23352
rect 27398 23296 27403 23352
rect 23197 23294 27403 23296
rect 23197 23291 23263 23294
rect 26601 23291 26667 23294
rect 27337 23291 27403 23294
rect 31334 23292 31340 23356
rect 31404 23354 31410 23356
rect 32029 23354 32095 23357
rect 31404 23352 32095 23354
rect 31404 23296 32034 23352
rect 32090 23296 32095 23352
rect 31404 23294 32095 23296
rect 31404 23292 31410 23294
rect 32029 23291 32095 23294
rect 10041 23218 10107 23221
rect 10777 23218 10843 23221
rect 11973 23218 12039 23221
rect 10041 23216 12039 23218
rect 10041 23160 10046 23216
rect 10102 23160 10782 23216
rect 10838 23160 11978 23216
rect 12034 23160 12039 23216
rect 10041 23158 12039 23160
rect 10041 23155 10107 23158
rect 10777 23155 10843 23158
rect 11973 23155 12039 23158
rect 14181 23218 14247 23221
rect 19149 23218 19215 23221
rect 14181 23216 19215 23218
rect 14181 23160 14186 23216
rect 14242 23160 19154 23216
rect 19210 23160 19215 23216
rect 14181 23158 19215 23160
rect 14181 23155 14247 23158
rect 19149 23155 19215 23158
rect 36169 23218 36235 23221
rect 36895 23218 37695 23248
rect 36169 23216 37695 23218
rect 36169 23160 36174 23216
rect 36230 23160 37695 23216
rect 36169 23158 37695 23160
rect 36169 23155 36235 23158
rect 36895 23128 37695 23158
rect 10041 23082 10107 23085
rect 11237 23082 11303 23085
rect 10041 23080 11303 23082
rect 10041 23024 10046 23080
rect 10102 23024 11242 23080
rect 11298 23024 11303 23080
rect 10041 23022 11303 23024
rect 10041 23019 10107 23022
rect 11237 23019 11303 23022
rect 13302 23020 13308 23084
rect 13372 23082 13378 23084
rect 19241 23082 19307 23085
rect 13372 23080 19307 23082
rect 13372 23024 19246 23080
rect 19302 23024 19307 23080
rect 13372 23022 19307 23024
rect 13372 23020 13378 23022
rect 19241 23019 19307 23022
rect 19425 23082 19491 23085
rect 23422 23082 23428 23084
rect 19425 23080 23428 23082
rect 19425 23024 19430 23080
rect 19486 23024 23428 23080
rect 19425 23022 23428 23024
rect 19425 23019 19491 23022
rect 23422 23020 23428 23022
rect 23492 23020 23498 23084
rect 26141 23082 26207 23085
rect 26366 23082 26372 23084
rect 26141 23080 26372 23082
rect 26141 23024 26146 23080
rect 26202 23024 26372 23080
rect 26141 23022 26372 23024
rect 26141 23019 26207 23022
rect 26366 23020 26372 23022
rect 26436 23082 26442 23084
rect 27245 23082 27311 23085
rect 26436 23080 27311 23082
rect 26436 23024 27250 23080
rect 27306 23024 27311 23080
rect 26436 23022 27311 23024
rect 26436 23020 26442 23022
rect 27245 23019 27311 23022
rect 30925 23082 30991 23085
rect 31661 23082 31727 23085
rect 35249 23082 35315 23085
rect 30925 23080 35315 23082
rect 30925 23024 30930 23080
rect 30986 23024 31666 23080
rect 31722 23024 35254 23080
rect 35310 23024 35315 23080
rect 30925 23022 35315 23024
rect 30925 23019 30991 23022
rect 31661 23019 31727 23022
rect 35249 23019 35315 23022
rect 22001 22946 22067 22949
rect 22461 22946 22527 22949
rect 26509 22946 26575 22949
rect 22001 22944 26575 22946
rect 22001 22888 22006 22944
rect 22062 22888 22466 22944
rect 22522 22888 26514 22944
rect 26570 22888 26575 22944
rect 22001 22886 26575 22888
rect 22001 22883 22067 22886
rect 22461 22883 22527 22886
rect 26509 22883 26575 22886
rect 30833 22946 30899 22949
rect 31845 22946 31911 22949
rect 30833 22944 31911 22946
rect 30833 22888 30838 22944
rect 30894 22888 31850 22944
rect 31906 22888 31911 22944
rect 30833 22886 31911 22888
rect 30833 22883 30899 22886
rect 31845 22883 31911 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 16614 22748 16620 22812
rect 16684 22810 16690 22812
rect 28165 22810 28231 22813
rect 16684 22808 28231 22810
rect 16684 22752 28170 22808
rect 28226 22752 28231 22808
rect 16684 22750 28231 22752
rect 16684 22748 16690 22750
rect 28165 22747 28231 22750
rect 28441 22810 28507 22813
rect 32949 22810 33015 22813
rect 28441 22808 33015 22810
rect 28441 22752 28446 22808
rect 28502 22752 32954 22808
rect 33010 22752 33015 22808
rect 28441 22750 33015 22752
rect 28441 22747 28507 22750
rect 32949 22747 33015 22750
rect 7414 22612 7420 22676
rect 7484 22674 7490 22676
rect 7649 22674 7715 22677
rect 7484 22672 7715 22674
rect 7484 22616 7654 22672
rect 7710 22616 7715 22672
rect 7484 22614 7715 22616
rect 7484 22612 7490 22614
rect 7649 22611 7715 22614
rect 22645 22674 22711 22677
rect 29361 22674 29427 22677
rect 29494 22674 29500 22676
rect 22645 22672 29500 22674
rect 22645 22616 22650 22672
rect 22706 22616 29366 22672
rect 29422 22616 29500 22672
rect 22645 22614 29500 22616
rect 22645 22611 22711 22614
rect 29361 22611 29427 22614
rect 29494 22612 29500 22614
rect 29564 22612 29570 22676
rect 32305 22674 32371 22677
rect 32438 22674 32444 22676
rect 32305 22672 32444 22674
rect 32305 22616 32310 22672
rect 32366 22616 32444 22672
rect 32305 22614 32444 22616
rect 32305 22611 32371 22614
rect 32438 22612 32444 22614
rect 32508 22612 32514 22676
rect 21449 22538 21515 22541
rect 21582 22538 21588 22540
rect 21449 22536 21588 22538
rect 21449 22480 21454 22536
rect 21510 22480 21588 22536
rect 21449 22478 21588 22480
rect 21449 22475 21515 22478
rect 21582 22476 21588 22478
rect 21652 22476 21658 22540
rect 22737 22538 22803 22541
rect 22870 22538 22876 22540
rect 22737 22536 22876 22538
rect 22737 22480 22742 22536
rect 22798 22480 22876 22536
rect 22737 22478 22876 22480
rect 22737 22475 22803 22478
rect 22870 22476 22876 22478
rect 22940 22476 22946 22540
rect 26877 22538 26943 22541
rect 31477 22538 31543 22541
rect 26877 22536 31543 22538
rect 26877 22480 26882 22536
rect 26938 22480 31482 22536
rect 31538 22480 31543 22536
rect 26877 22478 31543 22480
rect 26877 22475 26943 22478
rect 31477 22475 31543 22478
rect 33726 22476 33732 22540
rect 33796 22538 33802 22540
rect 35065 22538 35131 22541
rect 33796 22536 35131 22538
rect 33796 22480 35070 22536
rect 35126 22480 35131 22536
rect 33796 22478 35131 22480
rect 33796 22476 33802 22478
rect 35065 22475 35131 22478
rect 36169 22538 36235 22541
rect 36895 22538 37695 22568
rect 36169 22536 37695 22538
rect 36169 22480 36174 22536
rect 36230 22480 37695 22536
rect 36169 22478 37695 22480
rect 36169 22475 36235 22478
rect 36895 22448 37695 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 7281 22266 7347 22269
rect 4616 22264 7347 22266
rect 4616 22208 7286 22264
rect 7342 22208 7347 22264
rect 4616 22206 7347 22208
rect 4061 22130 4127 22133
rect 4337 22130 4403 22133
rect 4616 22130 4676 22206
rect 7281 22203 7347 22206
rect 17534 22204 17540 22268
rect 17604 22266 17610 22268
rect 19241 22266 19307 22269
rect 17604 22264 19307 22266
rect 17604 22208 19246 22264
rect 19302 22208 19307 22264
rect 17604 22206 19307 22208
rect 17604 22204 17610 22206
rect 19241 22203 19307 22206
rect 4061 22128 4676 22130
rect 4061 22072 4066 22128
rect 4122 22072 4342 22128
rect 4398 22072 4676 22128
rect 4061 22070 4676 22072
rect 23197 22130 23263 22133
rect 25037 22130 25103 22133
rect 23197 22128 25103 22130
rect 23197 22072 23202 22128
rect 23258 22072 25042 22128
rect 25098 22072 25103 22128
rect 23197 22070 25103 22072
rect 4061 22067 4127 22070
rect 4337 22067 4403 22070
rect 23197 22067 23263 22070
rect 25037 22067 25103 22070
rect 29729 22130 29795 22133
rect 30005 22130 30071 22133
rect 29729 22128 30071 22130
rect 29729 22072 29734 22128
rect 29790 22072 30010 22128
rect 30066 22072 30071 22128
rect 29729 22070 30071 22072
rect 29729 22067 29795 22070
rect 30005 22067 30071 22070
rect 30557 22130 30623 22133
rect 32305 22130 32371 22133
rect 30557 22128 32371 22130
rect 30557 22072 30562 22128
rect 30618 22072 32310 22128
rect 32366 22072 32371 22128
rect 30557 22070 32371 22072
rect 30557 22067 30623 22070
rect 32305 22067 32371 22070
rect 5073 21994 5139 21997
rect 5717 21994 5783 21997
rect 19425 21996 19491 21997
rect 5073 21992 5783 21994
rect 5073 21936 5078 21992
rect 5134 21936 5722 21992
rect 5778 21936 5783 21992
rect 5073 21934 5783 21936
rect 5073 21931 5139 21934
rect 5717 21931 5783 21934
rect 19374 21932 19380 21996
rect 19444 21994 19491 21996
rect 23565 21994 23631 21997
rect 24342 21994 24348 21996
rect 19444 21992 19536 21994
rect 19486 21936 19536 21992
rect 19444 21934 19536 21936
rect 23565 21992 24348 21994
rect 23565 21936 23570 21992
rect 23626 21936 24348 21992
rect 23565 21934 24348 21936
rect 19444 21932 19491 21934
rect 19425 21931 19491 21932
rect 23565 21931 23631 21934
rect 24342 21932 24348 21934
rect 24412 21994 24418 21996
rect 24577 21994 24643 21997
rect 24412 21992 24643 21994
rect 24412 21936 24582 21992
rect 24638 21936 24643 21992
rect 24412 21934 24643 21936
rect 24412 21932 24418 21934
rect 24577 21931 24643 21934
rect 25681 21994 25747 21997
rect 25681 21992 30114 21994
rect 25681 21936 25686 21992
rect 25742 21936 30114 21992
rect 25681 21934 30114 21936
rect 25681 21931 25747 21934
rect 18413 21858 18479 21861
rect 20345 21858 20411 21861
rect 18413 21856 20411 21858
rect 18413 21800 18418 21856
rect 18474 21800 20350 21856
rect 20406 21800 20411 21856
rect 18413 21798 20411 21800
rect 18413 21795 18479 21798
rect 20345 21795 20411 21798
rect 23054 21796 23060 21860
rect 23124 21858 23130 21860
rect 24301 21858 24367 21861
rect 24710 21858 24716 21860
rect 23124 21856 24716 21858
rect 23124 21800 24306 21856
rect 24362 21800 24716 21856
rect 23124 21798 24716 21800
rect 23124 21796 23130 21798
rect 24301 21795 24367 21798
rect 24710 21796 24716 21798
rect 24780 21796 24786 21860
rect 26182 21796 26188 21860
rect 26252 21858 26258 21860
rect 26877 21858 26943 21861
rect 26252 21856 26943 21858
rect 26252 21800 26882 21856
rect 26938 21800 26943 21856
rect 26252 21798 26943 21800
rect 26252 21796 26258 21798
rect 26877 21795 26943 21798
rect 29361 21858 29427 21861
rect 29862 21858 29868 21860
rect 29361 21856 29868 21858
rect 29361 21800 29366 21856
rect 29422 21800 29868 21856
rect 29361 21798 29868 21800
rect 29361 21795 29427 21798
rect 29862 21796 29868 21798
rect 29932 21796 29938 21860
rect 30054 21858 30114 21934
rect 31710 21934 36186 21994
rect 31710 21858 31770 21934
rect 30054 21798 31770 21858
rect 36126 21858 36186 21934
rect 36895 21858 37695 21888
rect 36126 21798 37695 21858
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 36895 21768 37695 21798
rect 35590 21727 35906 21728
rect 15009 21722 15075 21725
rect 18229 21722 18295 21725
rect 15009 21720 18295 21722
rect 15009 21664 15014 21720
rect 15070 21664 18234 21720
rect 18290 21664 18295 21720
rect 15009 21662 18295 21664
rect 15009 21659 15075 21662
rect 18229 21659 18295 21662
rect 19425 21722 19491 21725
rect 20161 21722 20227 21725
rect 20437 21722 20503 21725
rect 19425 21720 20503 21722
rect 19425 21664 19430 21720
rect 19486 21664 20166 21720
rect 20222 21664 20442 21720
rect 20498 21664 20503 21720
rect 19425 21662 20503 21664
rect 19425 21659 19491 21662
rect 20161 21659 20227 21662
rect 20437 21659 20503 21662
rect 24945 21722 25011 21725
rect 26877 21722 26943 21725
rect 24945 21720 26943 21722
rect 24945 21664 24950 21720
rect 25006 21664 26882 21720
rect 26938 21664 26943 21720
rect 24945 21662 26943 21664
rect 24945 21659 25011 21662
rect 26877 21659 26943 21662
rect 9213 21586 9279 21589
rect 10593 21586 10659 21589
rect 9213 21584 10659 21586
rect 9213 21528 9218 21584
rect 9274 21528 10598 21584
rect 10654 21528 10659 21584
rect 9213 21526 10659 21528
rect 9213 21523 9279 21526
rect 10593 21523 10659 21526
rect 15469 21586 15535 21589
rect 16062 21586 16068 21588
rect 15469 21584 16068 21586
rect 15469 21528 15474 21584
rect 15530 21528 16068 21584
rect 15469 21526 16068 21528
rect 15469 21523 15535 21526
rect 16062 21524 16068 21526
rect 16132 21524 16138 21588
rect 17217 21586 17283 21589
rect 24945 21586 25011 21589
rect 25405 21586 25471 21589
rect 17217 21584 25471 21586
rect 17217 21528 17222 21584
rect 17278 21528 24950 21584
rect 25006 21528 25410 21584
rect 25466 21528 25471 21584
rect 17217 21526 25471 21528
rect 17217 21523 17283 21526
rect 24945 21523 25011 21526
rect 25405 21523 25471 21526
rect 25589 21586 25655 21589
rect 36721 21586 36787 21589
rect 25589 21584 36787 21586
rect 25589 21528 25594 21584
rect 25650 21528 36726 21584
rect 36782 21528 36787 21584
rect 25589 21526 36787 21528
rect 25589 21523 25655 21526
rect 36721 21523 36787 21526
rect 9857 21450 9923 21453
rect 23841 21450 23907 21453
rect 9857 21448 23907 21450
rect 9857 21392 9862 21448
rect 9918 21392 23846 21448
rect 23902 21392 23907 21448
rect 9857 21390 23907 21392
rect 9857 21387 9923 21390
rect 23841 21387 23907 21390
rect 24526 21388 24532 21452
rect 24596 21450 24602 21452
rect 24669 21450 24735 21453
rect 24596 21448 24735 21450
rect 24596 21392 24674 21448
rect 24730 21392 24735 21448
rect 24596 21390 24735 21392
rect 24596 21388 24602 21390
rect 24669 21387 24735 21390
rect 28165 21450 28231 21453
rect 28441 21450 28507 21453
rect 28625 21452 28691 21453
rect 28165 21448 28507 21450
rect 28165 21392 28170 21448
rect 28226 21392 28446 21448
rect 28502 21392 28507 21448
rect 28165 21390 28507 21392
rect 28165 21387 28231 21390
rect 28441 21387 28507 21390
rect 28574 21388 28580 21452
rect 28644 21450 28691 21452
rect 28644 21448 28736 21450
rect 28686 21392 28736 21448
rect 28644 21390 28736 21392
rect 28644 21388 28691 21390
rect 28625 21387 28691 21388
rect 16021 21314 16087 21317
rect 20437 21314 20503 21317
rect 24485 21316 24551 21317
rect 24485 21314 24532 21316
rect 16021 21312 20503 21314
rect 16021 21256 16026 21312
rect 16082 21256 20442 21312
rect 20498 21256 20503 21312
rect 16021 21254 20503 21256
rect 24440 21312 24532 21314
rect 24440 21256 24490 21312
rect 24440 21254 24532 21256
rect 16021 21251 16087 21254
rect 20437 21251 20503 21254
rect 24485 21252 24532 21254
rect 24596 21252 24602 21316
rect 24485 21251 24551 21252
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 5717 21178 5783 21181
rect 8017 21178 8083 21181
rect 5717 21176 8083 21178
rect 5717 21120 5722 21176
rect 5778 21120 8022 21176
rect 8078 21120 8083 21176
rect 5717 21118 8083 21120
rect 5717 21115 5783 21118
rect 8017 21115 8083 21118
rect 16205 21178 16271 21181
rect 18781 21178 18847 21181
rect 16205 21176 18847 21178
rect 16205 21120 16210 21176
rect 16266 21120 18786 21176
rect 18842 21120 18847 21176
rect 16205 21118 18847 21120
rect 16205 21115 16271 21118
rect 18781 21115 18847 21118
rect 19425 21178 19491 21181
rect 23289 21178 23355 21181
rect 19425 21176 23355 21178
rect 19425 21120 19430 21176
rect 19486 21120 23294 21176
rect 23350 21120 23355 21176
rect 19425 21118 23355 21120
rect 19425 21115 19491 21118
rect 23289 21115 23355 21118
rect 28349 21178 28415 21181
rect 28717 21178 28783 21181
rect 28349 21176 28783 21178
rect 28349 21120 28354 21176
rect 28410 21120 28722 21176
rect 28778 21120 28783 21176
rect 28349 21118 28783 21120
rect 28349 21115 28415 21118
rect 28717 21115 28783 21118
rect 35525 21178 35591 21181
rect 36895 21178 37695 21208
rect 35525 21176 37695 21178
rect 35525 21120 35530 21176
rect 35586 21120 37695 21176
rect 35525 21118 37695 21120
rect 35525 21115 35591 21118
rect 36895 21088 37695 21118
rect 10041 21042 10107 21045
rect 19241 21042 19307 21045
rect 19609 21044 19675 21045
rect 10041 21040 19307 21042
rect 10041 20984 10046 21040
rect 10102 20984 19246 21040
rect 19302 20984 19307 21040
rect 10041 20982 19307 20984
rect 10041 20979 10107 20982
rect 19241 20979 19307 20982
rect 19558 20980 19564 21044
rect 19628 21042 19675 21044
rect 26601 21042 26667 21045
rect 31753 21042 31819 21045
rect 31886 21042 31892 21044
rect 19628 21040 19720 21042
rect 19670 20984 19720 21040
rect 19628 20982 19720 20984
rect 26601 21040 31632 21042
rect 26601 20984 26606 21040
rect 26662 20984 31632 21040
rect 26601 20982 31632 20984
rect 19628 20980 19675 20982
rect 19609 20979 19675 20980
rect 26601 20979 26667 20982
rect 4654 20844 4660 20908
rect 4724 20906 4730 20908
rect 4889 20906 4955 20909
rect 4724 20904 4955 20906
rect 4724 20848 4894 20904
rect 4950 20848 4955 20904
rect 4724 20846 4955 20848
rect 4724 20844 4730 20846
rect 4889 20843 4955 20846
rect 7373 20906 7439 20909
rect 10409 20906 10475 20909
rect 7373 20904 10475 20906
rect 7373 20848 7378 20904
rect 7434 20848 10414 20904
rect 10470 20848 10475 20904
rect 7373 20846 10475 20848
rect 7373 20843 7439 20846
rect 10409 20843 10475 20846
rect 17493 20906 17559 20909
rect 17861 20906 17927 20909
rect 19241 20906 19307 20909
rect 17493 20904 19307 20906
rect 17493 20848 17498 20904
rect 17554 20848 17866 20904
rect 17922 20848 19246 20904
rect 19302 20848 19307 20904
rect 17493 20846 19307 20848
rect 31572 20906 31632 20982
rect 31753 21040 31892 21042
rect 31753 20984 31758 21040
rect 31814 20984 31892 21040
rect 31753 20982 31892 20984
rect 31753 20979 31819 20982
rect 31886 20980 31892 20982
rect 31956 20980 31962 21044
rect 31572 20846 31770 20906
rect 17493 20843 17559 20846
rect 17861 20843 17927 20846
rect 19241 20843 19307 20846
rect 17953 20768 18019 20773
rect 17953 20712 17958 20768
rect 18014 20712 18019 20768
rect 17953 20707 18019 20712
rect 23381 20770 23447 20773
rect 24158 20770 24164 20772
rect 23381 20768 24164 20770
rect 23381 20712 23386 20768
rect 23442 20712 24164 20768
rect 23381 20710 24164 20712
rect 23381 20707 23447 20710
rect 24158 20708 24164 20710
rect 24228 20708 24234 20772
rect 26877 20770 26943 20773
rect 30557 20770 30623 20773
rect 31518 20770 31524 20772
rect 26877 20768 31524 20770
rect 26877 20712 26882 20768
rect 26938 20712 30562 20768
rect 30618 20712 31524 20768
rect 26877 20710 31524 20712
rect 26877 20707 26943 20710
rect 30557 20707 30623 20710
rect 31518 20708 31524 20710
rect 31588 20708 31594 20772
rect 31710 20770 31770 20846
rect 31886 20844 31892 20908
rect 31956 20906 31962 20908
rect 34973 20906 35039 20909
rect 31956 20904 35039 20906
rect 31956 20848 34978 20904
rect 35034 20848 35039 20904
rect 31956 20846 35039 20848
rect 31956 20844 31962 20846
rect 34973 20843 35039 20846
rect 32857 20770 32923 20773
rect 34697 20772 34763 20773
rect 34646 20770 34652 20772
rect 31710 20768 32923 20770
rect 31710 20712 32862 20768
rect 32918 20712 32923 20768
rect 31710 20710 32923 20712
rect 34606 20710 34652 20770
rect 34716 20768 34763 20772
rect 34758 20712 34763 20768
rect 32857 20707 32923 20710
rect 34646 20708 34652 20710
rect 34716 20708 34763 20712
rect 34697 20707 34763 20708
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 5717 20636 5783 20637
rect 5717 20632 5764 20636
rect 5828 20634 5834 20636
rect 7465 20634 7531 20637
rect 7598 20634 7604 20636
rect 5717 20576 5722 20632
rect 5717 20572 5764 20576
rect 5828 20574 5874 20634
rect 7465 20632 7604 20634
rect 7465 20576 7470 20632
rect 7526 20576 7604 20632
rect 7465 20574 7604 20576
rect 5828 20572 5834 20574
rect 5717 20571 5783 20572
rect 7465 20571 7531 20574
rect 7598 20572 7604 20574
rect 7668 20572 7674 20636
rect 17718 20572 17724 20636
rect 17788 20634 17794 20636
rect 17956 20634 18016 20707
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 17788 20574 18016 20634
rect 17788 20572 17794 20574
rect 18638 20572 18644 20636
rect 18708 20634 18714 20636
rect 19609 20634 19675 20637
rect 18708 20632 19675 20634
rect 18708 20576 19614 20632
rect 19670 20576 19675 20632
rect 18708 20574 19675 20576
rect 18708 20572 18714 20574
rect 19609 20571 19675 20574
rect 24209 20634 24275 20637
rect 26601 20636 26667 20637
rect 26550 20634 26556 20636
rect 24209 20632 26556 20634
rect 26620 20634 26667 20636
rect 31477 20634 31543 20637
rect 33317 20634 33383 20637
rect 26620 20632 26712 20634
rect 24209 20576 24214 20632
rect 24270 20576 26556 20632
rect 26662 20576 26712 20632
rect 24209 20574 26556 20576
rect 24209 20571 24275 20574
rect 26550 20572 26556 20574
rect 26620 20574 26712 20576
rect 31477 20632 33383 20634
rect 31477 20576 31482 20632
rect 31538 20576 33322 20632
rect 33378 20576 33383 20632
rect 31477 20574 33383 20576
rect 26620 20572 26667 20574
rect 26601 20571 26667 20572
rect 31477 20571 31543 20574
rect 33317 20571 33383 20574
rect 8886 20436 8892 20500
rect 8956 20498 8962 20500
rect 18781 20498 18847 20501
rect 8956 20496 18847 20498
rect 8956 20440 18786 20496
rect 18842 20440 18847 20496
rect 8956 20438 18847 20440
rect 8956 20436 8962 20438
rect 18781 20435 18847 20438
rect 19374 20436 19380 20500
rect 19444 20498 19450 20500
rect 21449 20498 21515 20501
rect 19444 20496 21515 20498
rect 19444 20440 21454 20496
rect 21510 20440 21515 20496
rect 19444 20438 21515 20440
rect 19444 20436 19450 20438
rect 21449 20435 21515 20438
rect 31293 20498 31359 20501
rect 31661 20498 31727 20501
rect 31293 20496 31727 20498
rect 31293 20440 31298 20496
rect 31354 20440 31666 20496
rect 31722 20440 31727 20496
rect 31293 20438 31727 20440
rect 31293 20435 31359 20438
rect 31661 20435 31727 20438
rect 36895 20500 37695 20528
rect 36895 20436 37044 20500
rect 37108 20436 37695 20500
rect 36895 20408 37695 20436
rect 11697 20362 11763 20365
rect 11830 20362 11836 20364
rect 11697 20360 11836 20362
rect 11697 20304 11702 20360
rect 11758 20304 11836 20360
rect 11697 20302 11836 20304
rect 11697 20299 11763 20302
rect 11830 20300 11836 20302
rect 11900 20300 11906 20364
rect 18505 20362 18571 20365
rect 19558 20362 19564 20364
rect 18505 20360 19564 20362
rect 18505 20304 18510 20360
rect 18566 20304 19564 20360
rect 18505 20302 19564 20304
rect 18505 20299 18571 20302
rect 19558 20300 19564 20302
rect 19628 20362 19634 20364
rect 20478 20362 20484 20364
rect 19628 20302 20484 20362
rect 19628 20300 19634 20302
rect 20478 20300 20484 20302
rect 20548 20300 20554 20364
rect 20621 20362 20687 20365
rect 20846 20362 20852 20364
rect 20621 20360 20852 20362
rect 20621 20304 20626 20360
rect 20682 20304 20852 20360
rect 20621 20302 20852 20304
rect 20621 20299 20687 20302
rect 20846 20300 20852 20302
rect 20916 20300 20922 20364
rect 27889 20362 27955 20365
rect 31661 20362 31727 20365
rect 33225 20362 33291 20365
rect 27889 20360 33291 20362
rect 27889 20304 27894 20360
rect 27950 20304 31666 20360
rect 31722 20304 33230 20360
rect 33286 20304 33291 20360
rect 27889 20302 33291 20304
rect 27889 20299 27955 20302
rect 31661 20299 31727 20302
rect 33225 20299 33291 20302
rect 17401 20226 17467 20229
rect 19701 20226 19767 20229
rect 20069 20228 20135 20229
rect 31845 20228 31911 20229
rect 20069 20226 20116 20228
rect 17401 20224 19767 20226
rect 17401 20168 17406 20224
rect 17462 20168 19706 20224
rect 19762 20168 19767 20224
rect 17401 20166 19767 20168
rect 20024 20224 20116 20226
rect 20024 20168 20074 20224
rect 20024 20166 20116 20168
rect 17401 20163 17467 20166
rect 19701 20163 19767 20166
rect 20069 20164 20116 20166
rect 20180 20164 20186 20228
rect 31845 20226 31892 20228
rect 31800 20224 31892 20226
rect 31800 20168 31850 20224
rect 31800 20166 31892 20168
rect 31845 20164 31892 20166
rect 31956 20164 31962 20228
rect 20069 20163 20135 20164
rect 31845 20163 31911 20164
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 9673 20090 9739 20093
rect 10174 20090 10180 20092
rect 9673 20088 10180 20090
rect 9673 20032 9678 20088
rect 9734 20032 10180 20088
rect 9673 20030 10180 20032
rect 9673 20027 9739 20030
rect 10174 20028 10180 20030
rect 10244 20028 10250 20092
rect 18270 20028 18276 20092
rect 18340 20090 18346 20092
rect 19149 20090 19215 20093
rect 32949 20090 33015 20093
rect 18340 20088 33015 20090
rect 18340 20032 19154 20088
rect 19210 20032 32954 20088
rect 33010 20032 33015 20088
rect 18340 20030 33015 20032
rect 18340 20028 18346 20030
rect 19149 20027 19215 20030
rect 32949 20027 33015 20030
rect 4521 19954 4587 19957
rect 5993 19954 6059 19957
rect 4521 19952 6059 19954
rect 4521 19896 4526 19952
rect 4582 19896 5998 19952
rect 6054 19896 6059 19952
rect 4521 19894 6059 19896
rect 4521 19891 4587 19894
rect 5993 19891 6059 19894
rect 12525 19954 12591 19957
rect 15193 19954 15259 19957
rect 25405 19956 25471 19957
rect 25405 19954 25452 19956
rect 12525 19952 15259 19954
rect 12525 19896 12530 19952
rect 12586 19896 15198 19952
rect 15254 19896 15259 19952
rect 12525 19894 15259 19896
rect 25364 19952 25452 19954
rect 25516 19954 25522 19956
rect 37038 19954 37044 19956
rect 25364 19896 25410 19952
rect 25364 19894 25452 19896
rect 12525 19891 12591 19894
rect 15193 19891 15259 19894
rect 25405 19892 25452 19894
rect 25516 19894 37044 19954
rect 25516 19892 25522 19894
rect 37038 19892 37044 19894
rect 37108 19892 37114 19956
rect 25405 19891 25471 19892
rect 17585 19818 17651 19821
rect 19793 19818 19859 19821
rect 17585 19816 19859 19818
rect 17585 19760 17590 19816
rect 17646 19760 19798 19816
rect 19854 19760 19859 19816
rect 17585 19758 19859 19760
rect 17585 19755 17651 19758
rect 19793 19755 19859 19758
rect 26877 19818 26943 19821
rect 27102 19818 27108 19820
rect 26877 19816 27108 19818
rect 26877 19760 26882 19816
rect 26938 19760 27108 19816
rect 26877 19758 27108 19760
rect 26877 19755 26943 19758
rect 27102 19756 27108 19758
rect 27172 19756 27178 19820
rect 31385 19818 31451 19821
rect 33358 19818 33364 19820
rect 31385 19816 33364 19818
rect 31385 19760 31390 19816
rect 31446 19760 33364 19816
rect 31385 19758 33364 19760
rect 31385 19755 31451 19758
rect 33358 19756 33364 19758
rect 33428 19756 33434 19820
rect 19333 19682 19399 19685
rect 23238 19682 23244 19684
rect 19333 19680 23244 19682
rect 19333 19624 19338 19680
rect 19394 19624 23244 19680
rect 19333 19622 23244 19624
rect 19333 19619 19399 19622
rect 23238 19620 23244 19622
rect 23308 19620 23314 19684
rect 24485 19682 24551 19685
rect 24761 19682 24827 19685
rect 24485 19680 24827 19682
rect 24485 19624 24490 19680
rect 24546 19624 24766 19680
rect 24822 19624 24827 19680
rect 24485 19622 24827 19624
rect 24485 19619 24551 19622
rect 24761 19619 24827 19622
rect 25630 19620 25636 19684
rect 25700 19682 25706 19684
rect 26509 19682 26575 19685
rect 25700 19680 26575 19682
rect 25700 19624 26514 19680
rect 26570 19624 26575 19680
rect 25700 19622 26575 19624
rect 25700 19620 25706 19622
rect 26509 19619 26575 19622
rect 30833 19682 30899 19685
rect 31385 19682 31451 19685
rect 30833 19680 31451 19682
rect 30833 19624 30838 19680
rect 30894 19624 31390 19680
rect 31446 19624 31451 19680
rect 30833 19622 31451 19624
rect 30833 19619 30899 19622
rect 31385 19619 31451 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 29545 19546 29611 19549
rect 30281 19546 30347 19549
rect 29545 19544 30347 19546
rect 29545 19488 29550 19544
rect 29606 19488 30286 19544
rect 30342 19488 30347 19544
rect 29545 19486 30347 19488
rect 29545 19483 29611 19486
rect 30281 19483 30347 19486
rect 16246 19348 16252 19412
rect 16316 19410 16322 19412
rect 17534 19410 17540 19412
rect 16316 19350 17540 19410
rect 16316 19348 16322 19350
rect 17534 19348 17540 19350
rect 17604 19348 17610 19412
rect 22001 19410 22067 19413
rect 24393 19410 24459 19413
rect 22001 19408 24459 19410
rect 22001 19352 22006 19408
rect 22062 19352 24398 19408
rect 24454 19352 24459 19408
rect 22001 19350 24459 19352
rect 22001 19347 22067 19350
rect 24393 19347 24459 19350
rect 28206 19348 28212 19412
rect 28276 19410 28282 19412
rect 28349 19410 28415 19413
rect 28276 19408 28415 19410
rect 28276 19352 28354 19408
rect 28410 19352 28415 19408
rect 28276 19350 28415 19352
rect 28276 19348 28282 19350
rect 28349 19347 28415 19350
rect 29821 19410 29887 19413
rect 30414 19410 30420 19412
rect 29821 19408 30420 19410
rect 29821 19352 29826 19408
rect 29882 19352 30420 19408
rect 29821 19350 30420 19352
rect 29821 19347 29887 19350
rect 30414 19348 30420 19350
rect 30484 19348 30490 19412
rect 32254 19348 32260 19412
rect 32324 19410 32330 19412
rect 32397 19410 32463 19413
rect 32324 19408 32463 19410
rect 32324 19352 32402 19408
rect 32458 19352 32463 19408
rect 32324 19350 32463 19352
rect 32324 19348 32330 19350
rect 32397 19347 32463 19350
rect 12249 19276 12315 19277
rect 12198 19274 12204 19276
rect 12158 19214 12204 19274
rect 12268 19272 12315 19276
rect 12310 19216 12315 19272
rect 12198 19212 12204 19214
rect 12268 19212 12315 19216
rect 12249 19211 12315 19212
rect 14181 19274 14247 19277
rect 15326 19274 15332 19276
rect 14181 19272 15332 19274
rect 14181 19216 14186 19272
rect 14242 19216 15332 19272
rect 14181 19214 15332 19216
rect 14181 19211 14247 19214
rect 15326 19212 15332 19214
rect 15396 19212 15402 19276
rect 18137 19274 18203 19277
rect 19241 19274 19307 19277
rect 18137 19272 19307 19274
rect 18137 19216 18142 19272
rect 18198 19216 19246 19272
rect 19302 19216 19307 19272
rect 18137 19214 19307 19216
rect 18137 19211 18203 19214
rect 19241 19211 19307 19214
rect 21081 19274 21147 19277
rect 22093 19274 22159 19277
rect 21081 19272 22159 19274
rect 21081 19216 21086 19272
rect 21142 19216 22098 19272
rect 22154 19216 22159 19272
rect 21081 19214 22159 19216
rect 21081 19211 21147 19214
rect 22093 19211 22159 19214
rect 23933 19274 23999 19277
rect 25998 19274 26004 19276
rect 23933 19272 26004 19274
rect 23933 19216 23938 19272
rect 23994 19216 26004 19272
rect 23933 19214 26004 19216
rect 23933 19211 23999 19214
rect 25998 19212 26004 19214
rect 26068 19212 26074 19276
rect 17861 19138 17927 19141
rect 24669 19138 24735 19141
rect 17861 19136 24735 19138
rect 17861 19080 17866 19136
rect 17922 19080 24674 19136
rect 24730 19080 24735 19136
rect 17861 19078 24735 19080
rect 17861 19075 17927 19078
rect 24669 19075 24735 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 21817 19002 21883 19005
rect 25865 19002 25931 19005
rect 21817 19000 25931 19002
rect 21817 18944 21822 19000
rect 21878 18944 25870 19000
rect 25926 18944 25931 19000
rect 21817 18942 25931 18944
rect 21817 18939 21883 18942
rect 25865 18939 25931 18942
rect 10409 18866 10475 18869
rect 17125 18866 17191 18869
rect 28717 18868 28783 18869
rect 28717 18866 28764 18868
rect 10409 18864 17191 18866
rect 10409 18808 10414 18864
rect 10470 18808 17130 18864
rect 17186 18808 17191 18864
rect 10409 18806 17191 18808
rect 28672 18864 28764 18866
rect 28672 18808 28722 18864
rect 28672 18806 28764 18808
rect 10409 18803 10475 18806
rect 17125 18803 17191 18806
rect 28717 18804 28764 18806
rect 28828 18804 28834 18868
rect 28717 18803 28783 18804
rect 11053 18730 11119 18733
rect 11513 18732 11579 18733
rect 11278 18730 11284 18732
rect 11053 18728 11284 18730
rect 11053 18672 11058 18728
rect 11114 18672 11284 18728
rect 11053 18670 11284 18672
rect 11053 18667 11119 18670
rect 11278 18668 11284 18670
rect 11348 18668 11354 18732
rect 11462 18668 11468 18732
rect 11532 18730 11579 18732
rect 14089 18730 14155 18733
rect 20662 18730 20668 18732
rect 11532 18728 11624 18730
rect 11574 18672 11624 18728
rect 11532 18670 11624 18672
rect 14089 18728 20668 18730
rect 14089 18672 14094 18728
rect 14150 18672 20668 18728
rect 14089 18670 20668 18672
rect 11532 18668 11579 18670
rect 11513 18667 11579 18668
rect 14089 18667 14155 18670
rect 20662 18668 20668 18670
rect 20732 18668 20738 18732
rect 21081 18730 21147 18733
rect 23105 18730 23171 18733
rect 26969 18730 27035 18733
rect 21081 18728 27035 18730
rect 21081 18672 21086 18728
rect 21142 18672 23110 18728
rect 23166 18672 26974 18728
rect 27030 18672 27035 18728
rect 21081 18670 27035 18672
rect 21081 18667 21147 18670
rect 23105 18667 23171 18670
rect 26969 18667 27035 18670
rect 19425 18594 19491 18597
rect 21173 18594 21239 18597
rect 19425 18592 21239 18594
rect 19425 18536 19430 18592
rect 19486 18536 21178 18592
rect 21234 18536 21239 18592
rect 19425 18534 21239 18536
rect 19425 18531 19491 18534
rect 21173 18531 21239 18534
rect 21541 18594 21607 18597
rect 21766 18594 21772 18596
rect 21541 18592 21772 18594
rect 21541 18536 21546 18592
rect 21602 18536 21772 18592
rect 21541 18534 21772 18536
rect 21541 18531 21607 18534
rect 21766 18532 21772 18534
rect 21836 18532 21842 18596
rect 22093 18594 22159 18597
rect 26601 18594 26667 18597
rect 22093 18592 26667 18594
rect 22093 18536 22098 18592
rect 22154 18536 26606 18592
rect 26662 18536 26667 18592
rect 22093 18534 26667 18536
rect 22093 18531 22159 18534
rect 26601 18531 26667 18534
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 10961 18460 11027 18461
rect 10910 18396 10916 18460
rect 10980 18458 11027 18460
rect 17953 18458 18019 18461
rect 19149 18458 19215 18461
rect 10980 18456 11072 18458
rect 11022 18400 11072 18456
rect 10980 18398 11072 18400
rect 17953 18456 19215 18458
rect 17953 18400 17958 18456
rect 18014 18400 19154 18456
rect 19210 18400 19215 18456
rect 17953 18398 19215 18400
rect 10980 18396 11027 18398
rect 10961 18395 11027 18396
rect 17953 18395 18019 18398
rect 19149 18395 19215 18398
rect 20529 18458 20595 18461
rect 21817 18458 21883 18461
rect 20529 18456 21883 18458
rect 20529 18400 20534 18456
rect 20590 18400 21822 18456
rect 21878 18400 21883 18456
rect 20529 18398 21883 18400
rect 20529 18395 20595 18398
rect 21817 18395 21883 18398
rect 22277 18458 22343 18461
rect 26417 18458 26483 18461
rect 22277 18456 26483 18458
rect 22277 18400 22282 18456
rect 22338 18400 26422 18456
rect 26478 18400 26483 18456
rect 22277 18398 26483 18400
rect 22277 18395 22343 18398
rect 26417 18395 26483 18398
rect 14038 18260 14044 18324
rect 14108 18322 14114 18324
rect 25313 18322 25379 18325
rect 14108 18320 25379 18322
rect 14108 18264 25318 18320
rect 25374 18264 25379 18320
rect 14108 18262 25379 18264
rect 14108 18260 14114 18262
rect 25313 18259 25379 18262
rect 25681 18322 25747 18325
rect 26182 18322 26188 18324
rect 25681 18320 26188 18322
rect 25681 18264 25686 18320
rect 25742 18264 26188 18320
rect 25681 18262 26188 18264
rect 25681 18259 25747 18262
rect 26182 18260 26188 18262
rect 26252 18260 26258 18324
rect 36629 18322 36695 18325
rect 31710 18320 36695 18322
rect 31710 18264 36634 18320
rect 36690 18264 36695 18320
rect 31710 18262 36695 18264
rect 21633 18188 21699 18189
rect 21582 18186 21588 18188
rect 21542 18126 21588 18186
rect 21652 18184 21699 18188
rect 21694 18128 21699 18184
rect 21582 18124 21588 18126
rect 21652 18124 21699 18128
rect 21633 18123 21699 18124
rect 24761 18186 24827 18189
rect 31710 18186 31770 18262
rect 36629 18259 36695 18262
rect 24761 18184 31770 18186
rect 24761 18128 24766 18184
rect 24822 18128 31770 18184
rect 24761 18126 31770 18128
rect 32397 18186 32463 18189
rect 34421 18186 34487 18189
rect 32397 18184 34487 18186
rect 32397 18128 32402 18184
rect 32458 18128 34426 18184
rect 34482 18128 34487 18184
rect 32397 18126 34487 18128
rect 24761 18123 24827 18126
rect 32397 18123 32463 18126
rect 34421 18123 34487 18126
rect 9765 18050 9831 18053
rect 10358 18050 10364 18052
rect 9765 18048 10364 18050
rect 9765 17992 9770 18048
rect 9826 17992 10364 18048
rect 9765 17990 10364 17992
rect 9765 17987 9831 17990
rect 10358 17988 10364 17990
rect 10428 17988 10434 18052
rect 13118 17988 13124 18052
rect 13188 18050 13194 18052
rect 14733 18050 14799 18053
rect 13188 18048 14799 18050
rect 13188 17992 14738 18048
rect 14794 17992 14799 18048
rect 13188 17990 14799 17992
rect 13188 17988 13194 17990
rect 14733 17987 14799 17990
rect 15142 17988 15148 18052
rect 15212 18050 15218 18052
rect 15377 18050 15443 18053
rect 15212 18048 15443 18050
rect 15212 17992 15382 18048
rect 15438 17992 15443 18048
rect 15212 17990 15443 17992
rect 15212 17988 15218 17990
rect 15377 17987 15443 17990
rect 23054 17988 23060 18052
rect 23124 18050 23130 18052
rect 24577 18050 24643 18053
rect 34513 18050 34579 18053
rect 23124 18048 24643 18050
rect 23124 17992 24582 18048
rect 24638 17992 24643 18048
rect 23124 17990 24643 17992
rect 23124 17988 23130 17990
rect 24577 17987 24643 17990
rect 30422 18048 34579 18050
rect 30422 17992 34518 18048
rect 34574 17992 34579 18048
rect 30422 17990 34579 17992
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 11145 17914 11211 17917
rect 13854 17914 13860 17916
rect 11145 17912 13860 17914
rect 11145 17856 11150 17912
rect 11206 17856 13860 17912
rect 11145 17854 13860 17856
rect 11145 17851 11211 17854
rect 13854 17852 13860 17854
rect 13924 17852 13930 17916
rect 14774 17852 14780 17916
rect 14844 17914 14850 17916
rect 26233 17914 26299 17917
rect 14844 17912 26299 17914
rect 14844 17856 26238 17912
rect 26294 17856 26299 17912
rect 14844 17854 26299 17856
rect 14844 17852 14850 17854
rect 26233 17851 26299 17854
rect 27061 17914 27127 17917
rect 30422 17914 30482 17990
rect 34513 17987 34579 17990
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 27061 17912 30482 17914
rect 27061 17856 27066 17912
rect 27122 17856 30482 17912
rect 27061 17854 30482 17856
rect 30925 17914 30991 17917
rect 32305 17914 32371 17917
rect 30925 17912 32371 17914
rect 30925 17856 30930 17912
rect 30986 17856 32310 17912
rect 32366 17856 32371 17912
rect 30925 17854 32371 17856
rect 27061 17851 27127 17854
rect 30925 17851 30991 17854
rect 32305 17851 32371 17854
rect 18873 17778 18939 17781
rect 19006 17778 19012 17780
rect 18873 17776 19012 17778
rect 18873 17720 18878 17776
rect 18934 17720 19012 17776
rect 18873 17718 19012 17720
rect 18873 17715 18939 17718
rect 19006 17716 19012 17718
rect 19076 17716 19082 17780
rect 19793 17778 19859 17781
rect 25221 17778 25287 17781
rect 19793 17776 25287 17778
rect 19793 17720 19798 17776
rect 19854 17720 25226 17776
rect 25282 17720 25287 17776
rect 19793 17718 25287 17720
rect 19793 17715 19859 17718
rect 25221 17715 25287 17718
rect 14958 17580 14964 17644
rect 15028 17642 15034 17644
rect 25037 17642 25103 17645
rect 15028 17640 25103 17642
rect 15028 17584 25042 17640
rect 25098 17584 25103 17640
rect 15028 17582 25103 17584
rect 15028 17580 15034 17582
rect 25037 17579 25103 17582
rect 18873 17506 18939 17509
rect 19374 17506 19380 17508
rect 18873 17504 19380 17506
rect 18873 17448 18878 17504
rect 18934 17448 19380 17504
rect 18873 17446 19380 17448
rect 18873 17443 18939 17446
rect 19374 17444 19380 17446
rect 19444 17444 19450 17508
rect 21449 17506 21515 17509
rect 27337 17506 27403 17509
rect 21449 17504 27403 17506
rect 21449 17448 21454 17504
rect 21510 17448 27342 17504
rect 27398 17448 27403 17504
rect 21449 17446 27403 17448
rect 21449 17443 21515 17446
rect 27337 17443 27403 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 13629 17370 13695 17373
rect 16614 17370 16620 17372
rect 13629 17368 16620 17370
rect 13629 17312 13634 17368
rect 13690 17312 16620 17368
rect 13629 17310 16620 17312
rect 13629 17307 13695 17310
rect 16614 17308 16620 17310
rect 16684 17308 16690 17372
rect 16757 17370 16823 17373
rect 20529 17370 20595 17373
rect 16757 17368 20595 17370
rect 16757 17312 16762 17368
rect 16818 17312 20534 17368
rect 20590 17312 20595 17368
rect 16757 17310 20595 17312
rect 16757 17307 16823 17310
rect 20529 17307 20595 17310
rect 21541 17370 21607 17373
rect 23289 17370 23355 17373
rect 21541 17368 23355 17370
rect 21541 17312 21546 17368
rect 21602 17312 23294 17368
rect 23350 17312 23355 17368
rect 21541 17310 23355 17312
rect 21541 17307 21607 17310
rect 23289 17307 23355 17310
rect 16430 17172 16436 17236
rect 16500 17234 16506 17236
rect 17902 17234 17908 17236
rect 16500 17174 17908 17234
rect 16500 17172 16506 17174
rect 17902 17172 17908 17174
rect 17972 17172 17978 17236
rect 20069 17234 20135 17237
rect 24945 17234 25011 17237
rect 27429 17234 27495 17237
rect 20069 17232 27495 17234
rect 20069 17176 20074 17232
rect 20130 17176 24950 17232
rect 25006 17176 27434 17232
rect 27490 17176 27495 17232
rect 20069 17174 27495 17176
rect 20069 17171 20135 17174
rect 24945 17171 25011 17174
rect 27429 17171 27495 17174
rect 13629 17098 13695 17101
rect 18505 17098 18571 17101
rect 13629 17096 18571 17098
rect 13629 17040 13634 17096
rect 13690 17040 18510 17096
rect 18566 17040 18571 17096
rect 13629 17038 18571 17040
rect 13629 17035 13695 17038
rect 18505 17035 18571 17038
rect 21766 17036 21772 17100
rect 21836 17098 21842 17100
rect 22553 17098 22619 17101
rect 21836 17096 22619 17098
rect 21836 17040 22558 17096
rect 22614 17040 22619 17096
rect 21836 17038 22619 17040
rect 21836 17036 21842 17038
rect 22553 17035 22619 17038
rect 24393 17098 24459 17101
rect 24710 17098 24716 17100
rect 24393 17096 24716 17098
rect 24393 17040 24398 17096
rect 24454 17040 24716 17096
rect 24393 17038 24716 17040
rect 24393 17035 24459 17038
rect 24710 17036 24716 17038
rect 24780 17098 24786 17100
rect 25814 17098 25820 17100
rect 24780 17038 25820 17098
rect 24780 17036 24786 17038
rect 25814 17036 25820 17038
rect 25884 17036 25890 17100
rect 16798 16900 16804 16964
rect 16868 16962 16874 16964
rect 19742 16962 19748 16964
rect 16868 16902 19748 16962
rect 16868 16900 16874 16902
rect 19742 16900 19748 16902
rect 19812 16962 19818 16964
rect 25589 16962 25655 16965
rect 19812 16960 25655 16962
rect 19812 16904 25594 16960
rect 25650 16904 25655 16960
rect 19812 16902 25655 16904
rect 19812 16900 19818 16902
rect 25589 16899 25655 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 17585 16828 17651 16829
rect 18137 16828 18203 16829
rect 17534 16764 17540 16828
rect 17604 16826 17651 16828
rect 18086 16826 18092 16828
rect 17604 16824 17696 16826
rect 17646 16768 17696 16824
rect 17604 16766 17696 16768
rect 18046 16766 18092 16826
rect 18156 16824 18203 16828
rect 18198 16768 18203 16824
rect 17604 16764 17651 16766
rect 18086 16764 18092 16766
rect 18156 16764 18203 16768
rect 22502 16764 22508 16828
rect 22572 16826 22578 16828
rect 24117 16826 24183 16829
rect 22572 16824 24183 16826
rect 22572 16768 24122 16824
rect 24178 16768 24183 16824
rect 22572 16766 24183 16768
rect 22572 16764 22578 16766
rect 17585 16763 17651 16764
rect 18137 16763 18203 16764
rect 24117 16763 24183 16766
rect 5257 16690 5323 16693
rect 7414 16690 7420 16692
rect 5257 16688 7420 16690
rect 5257 16632 5262 16688
rect 5318 16632 7420 16688
rect 5257 16630 7420 16632
rect 5257 16627 5323 16630
rect 7414 16628 7420 16630
rect 7484 16628 7490 16692
rect 13721 16690 13787 16693
rect 24393 16690 24459 16693
rect 13721 16688 24459 16690
rect 13721 16632 13726 16688
rect 13782 16632 24398 16688
rect 24454 16632 24459 16688
rect 13721 16630 24459 16632
rect 13721 16627 13787 16630
rect 24393 16627 24459 16630
rect 25446 16628 25452 16692
rect 25516 16690 25522 16692
rect 25957 16690 26023 16693
rect 25516 16688 26023 16690
rect 25516 16632 25962 16688
rect 26018 16632 26023 16688
rect 25516 16630 26023 16632
rect 25516 16628 25522 16630
rect 25957 16627 26023 16630
rect 4889 16554 4955 16557
rect 5533 16554 5599 16557
rect 8937 16554 9003 16557
rect 4889 16552 9003 16554
rect 4889 16496 4894 16552
rect 4950 16496 5538 16552
rect 5594 16496 8942 16552
rect 8998 16496 9003 16552
rect 4889 16494 9003 16496
rect 4889 16491 4955 16494
rect 5533 16491 5599 16494
rect 8937 16491 9003 16494
rect 13486 16492 13492 16556
rect 13556 16554 13562 16556
rect 14038 16554 14044 16556
rect 13556 16494 14044 16554
rect 13556 16492 13562 16494
rect 14038 16492 14044 16494
rect 14108 16492 14114 16556
rect 16205 16554 16271 16557
rect 17953 16554 18019 16557
rect 16205 16552 18019 16554
rect 16205 16496 16210 16552
rect 16266 16496 17958 16552
rect 18014 16496 18019 16552
rect 16205 16494 18019 16496
rect 16205 16491 16271 16494
rect 17953 16491 18019 16494
rect 20161 16554 20227 16557
rect 23013 16554 23079 16557
rect 23422 16554 23428 16556
rect 20161 16552 22938 16554
rect 20161 16496 20166 16552
rect 20222 16496 22938 16552
rect 20161 16494 22938 16496
rect 20161 16491 20227 16494
rect 17217 16418 17283 16421
rect 20529 16418 20595 16421
rect 17217 16416 20595 16418
rect 17217 16360 17222 16416
rect 17278 16360 20534 16416
rect 20590 16360 20595 16416
rect 17217 16358 20595 16360
rect 22878 16418 22938 16494
rect 23013 16552 23428 16554
rect 23013 16496 23018 16552
rect 23074 16496 23428 16552
rect 23013 16494 23428 16496
rect 23013 16491 23079 16494
rect 23422 16492 23428 16494
rect 23492 16492 23498 16556
rect 23657 16554 23723 16557
rect 28758 16554 28764 16556
rect 23657 16552 28764 16554
rect 23657 16496 23662 16552
rect 23718 16496 28764 16552
rect 23657 16494 28764 16496
rect 23657 16491 23723 16494
rect 28758 16492 28764 16494
rect 28828 16492 28834 16556
rect 35249 16554 35315 16557
rect 31710 16552 35315 16554
rect 31710 16496 35254 16552
rect 35310 16496 35315 16552
rect 31710 16494 35315 16496
rect 26918 16418 26924 16420
rect 22878 16358 26924 16418
rect 17217 16355 17283 16358
rect 20529 16355 20595 16358
rect 26918 16356 26924 16358
rect 26988 16418 26994 16420
rect 31710 16418 31770 16494
rect 35249 16491 35315 16494
rect 26988 16358 31770 16418
rect 26988 16356 26994 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 11329 16282 11395 16285
rect 13905 16282 13971 16285
rect 11329 16280 13971 16282
rect 11329 16224 11334 16280
rect 11390 16224 13910 16280
rect 13966 16224 13971 16280
rect 11329 16222 13971 16224
rect 11329 16219 11395 16222
rect 13905 16219 13971 16222
rect 14641 16282 14707 16285
rect 25773 16282 25839 16285
rect 14641 16280 25839 16282
rect 14641 16224 14646 16280
rect 14702 16224 25778 16280
rect 25834 16224 25839 16280
rect 14641 16222 25839 16224
rect 14641 16219 14707 16222
rect 25773 16219 25839 16222
rect 31201 16282 31267 16285
rect 32581 16282 32647 16285
rect 31201 16280 32647 16282
rect 31201 16224 31206 16280
rect 31262 16224 32586 16280
rect 32642 16224 32647 16280
rect 31201 16222 32647 16224
rect 31201 16219 31267 16222
rect 32581 16219 32647 16222
rect 13721 16146 13787 16149
rect 14365 16146 14431 16149
rect 19241 16146 19307 16149
rect 13721 16144 19307 16146
rect 13721 16088 13726 16144
rect 13782 16088 14370 16144
rect 14426 16088 19246 16144
rect 19302 16088 19307 16144
rect 13721 16086 19307 16088
rect 13721 16083 13787 16086
rect 14365 16083 14431 16086
rect 19241 16083 19307 16086
rect 19701 16146 19767 16149
rect 20161 16146 20227 16149
rect 19701 16144 20227 16146
rect 19701 16088 19706 16144
rect 19762 16088 20166 16144
rect 20222 16088 20227 16144
rect 19701 16086 20227 16088
rect 19701 16083 19767 16086
rect 20161 16083 20227 16086
rect 22277 16146 22343 16149
rect 28390 16146 28396 16148
rect 22277 16144 28396 16146
rect 22277 16088 22282 16144
rect 22338 16088 28396 16144
rect 22277 16086 28396 16088
rect 22277 16083 22343 16086
rect 28390 16084 28396 16086
rect 28460 16146 28466 16148
rect 29177 16146 29243 16149
rect 28460 16144 29243 16146
rect 28460 16088 29182 16144
rect 29238 16088 29243 16144
rect 28460 16086 29243 16088
rect 28460 16084 28466 16086
rect 29177 16083 29243 16086
rect 29361 16146 29427 16149
rect 31569 16146 31635 16149
rect 29361 16144 31635 16146
rect 29361 16088 29366 16144
rect 29422 16088 31574 16144
rect 31630 16088 31635 16144
rect 29361 16086 31635 16088
rect 29361 16083 29427 16086
rect 31569 16083 31635 16086
rect 21725 16010 21791 16013
rect 24485 16010 24551 16013
rect 21725 16008 24551 16010
rect 21725 15952 21730 16008
rect 21786 15952 24490 16008
rect 24546 15952 24551 16008
rect 21725 15950 24551 15952
rect 21725 15947 21791 15950
rect 24485 15947 24551 15950
rect 30189 16010 30255 16013
rect 33409 16010 33475 16013
rect 30189 16008 33475 16010
rect 30189 15952 30194 16008
rect 30250 15952 33414 16008
rect 33470 15952 33475 16008
rect 30189 15950 33475 15952
rect 30189 15947 30255 15950
rect 33409 15947 33475 15950
rect 20529 15874 20595 15877
rect 24117 15874 24183 15877
rect 20529 15872 24183 15874
rect 20529 15816 20534 15872
rect 20590 15816 24122 15872
rect 24178 15816 24183 15872
rect 20529 15814 24183 15816
rect 20529 15811 20595 15814
rect 24117 15811 24183 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 21633 15738 21699 15741
rect 22553 15738 22619 15741
rect 27613 15738 27679 15741
rect 21633 15736 27679 15738
rect 21633 15680 21638 15736
rect 21694 15680 22558 15736
rect 22614 15680 27618 15736
rect 27674 15680 27679 15736
rect 21633 15678 27679 15680
rect 21633 15675 21699 15678
rect 22553 15675 22619 15678
rect 27613 15675 27679 15678
rect 8753 15602 8819 15605
rect 9397 15602 9463 15605
rect 8753 15600 9463 15602
rect 8753 15544 8758 15600
rect 8814 15544 9402 15600
rect 9458 15544 9463 15600
rect 8753 15542 9463 15544
rect 8753 15539 8819 15542
rect 9397 15539 9463 15542
rect 17585 15602 17651 15605
rect 18137 15602 18203 15605
rect 18965 15604 19031 15605
rect 18270 15602 18276 15604
rect 17585 15600 18276 15602
rect 17585 15544 17590 15600
rect 17646 15544 18142 15600
rect 18198 15544 18276 15600
rect 17585 15542 18276 15544
rect 17585 15539 17651 15542
rect 18137 15539 18203 15542
rect 18270 15540 18276 15542
rect 18340 15540 18346 15604
rect 18965 15600 19012 15604
rect 19076 15602 19082 15604
rect 20253 15602 20319 15605
rect 21398 15602 21404 15604
rect 18965 15544 18970 15600
rect 18965 15540 19012 15544
rect 19076 15542 19122 15602
rect 20253 15600 21404 15602
rect 20253 15544 20258 15600
rect 20314 15544 21404 15600
rect 20253 15542 21404 15544
rect 19076 15540 19082 15542
rect 18965 15539 19031 15540
rect 20253 15539 20319 15542
rect 21398 15540 21404 15542
rect 21468 15540 21474 15604
rect 21950 15540 21956 15604
rect 22020 15602 22026 15604
rect 24577 15602 24643 15605
rect 22020 15600 24643 15602
rect 22020 15544 24582 15600
rect 24638 15544 24643 15600
rect 22020 15542 24643 15544
rect 22020 15540 22026 15542
rect 24577 15539 24643 15542
rect 19793 15466 19859 15469
rect 20478 15466 20484 15468
rect 19793 15464 20484 15466
rect 19793 15408 19798 15464
rect 19854 15408 20484 15464
rect 19793 15406 20484 15408
rect 19793 15403 19859 15406
rect 20478 15404 20484 15406
rect 20548 15404 20554 15468
rect 30189 15466 30255 15469
rect 33726 15466 33732 15468
rect 30189 15464 33732 15466
rect 30189 15408 30194 15464
rect 30250 15408 33732 15464
rect 30189 15406 33732 15408
rect 30189 15403 30255 15406
rect 33726 15404 33732 15406
rect 33796 15404 33802 15468
rect 18137 15330 18203 15333
rect 26601 15330 26667 15333
rect 18137 15328 26667 15330
rect 18137 15272 18142 15328
rect 18198 15272 26606 15328
rect 26662 15272 26667 15328
rect 18137 15270 26667 15272
rect 18137 15267 18203 15270
rect 26601 15267 26667 15270
rect 26969 15330 27035 15333
rect 27286 15330 27292 15332
rect 26969 15328 27292 15330
rect 26969 15272 26974 15328
rect 27030 15272 27292 15328
rect 26969 15270 27292 15272
rect 26969 15267 27035 15270
rect 27286 15268 27292 15270
rect 27356 15268 27362 15332
rect 27838 15268 27844 15332
rect 27908 15330 27914 15332
rect 27981 15330 28047 15333
rect 27908 15328 28047 15330
rect 27908 15272 27986 15328
rect 28042 15272 28047 15328
rect 27908 15270 28047 15272
rect 27908 15268 27914 15270
rect 27981 15267 28047 15270
rect 31150 15268 31156 15332
rect 31220 15330 31226 15332
rect 31293 15330 31359 15333
rect 31220 15328 31359 15330
rect 31220 15272 31298 15328
rect 31354 15272 31359 15328
rect 31220 15270 31359 15272
rect 31220 15268 31226 15270
rect 31293 15267 31359 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 15561 15194 15627 15197
rect 15745 15194 15811 15197
rect 15561 15192 15811 15194
rect 15561 15136 15566 15192
rect 15622 15136 15750 15192
rect 15806 15136 15811 15192
rect 15561 15134 15811 15136
rect 15561 15131 15627 15134
rect 15745 15131 15811 15134
rect 19057 15194 19123 15197
rect 21909 15194 21975 15197
rect 23013 15194 23079 15197
rect 19057 15192 23079 15194
rect 19057 15136 19062 15192
rect 19118 15136 21914 15192
rect 21970 15136 23018 15192
rect 23074 15136 23079 15192
rect 19057 15134 23079 15136
rect 19057 15131 19123 15134
rect 21909 15131 21975 15134
rect 23013 15131 23079 15134
rect 24894 15132 24900 15196
rect 24964 15194 24970 15196
rect 25037 15194 25103 15197
rect 24964 15192 25103 15194
rect 24964 15136 25042 15192
rect 25098 15136 25103 15192
rect 24964 15134 25103 15136
rect 24964 15132 24970 15134
rect 25037 15131 25103 15134
rect 26325 15196 26391 15197
rect 29269 15196 29335 15197
rect 26325 15192 26372 15196
rect 26436 15194 26442 15196
rect 29269 15194 29316 15196
rect 26325 15136 26330 15192
rect 26325 15132 26372 15136
rect 26436 15134 26482 15194
rect 29224 15192 29316 15194
rect 29224 15136 29274 15192
rect 29224 15134 29316 15136
rect 26436 15132 26442 15134
rect 29269 15132 29316 15134
rect 29380 15132 29386 15196
rect 26325 15131 26391 15132
rect 29269 15131 29335 15132
rect 18045 15058 18111 15061
rect 18229 15060 18295 15061
rect 18229 15058 18276 15060
rect 18045 15056 18276 15058
rect 18045 15000 18050 15056
rect 18106 15000 18234 15056
rect 18045 14998 18276 15000
rect 18045 14995 18111 14998
rect 18229 14996 18276 14998
rect 18340 14996 18346 15060
rect 18413 15058 18479 15061
rect 19190 15058 19196 15060
rect 18413 15056 19196 15058
rect 18413 15000 18418 15056
rect 18474 15000 19196 15056
rect 18413 14998 19196 15000
rect 18229 14995 18295 14996
rect 18413 14995 18479 14998
rect 19190 14996 19196 14998
rect 19260 14996 19266 15060
rect 19558 14996 19564 15060
rect 19628 15058 19634 15060
rect 20897 15058 20963 15061
rect 22921 15058 22987 15061
rect 19628 15056 22987 15058
rect 19628 15000 20902 15056
rect 20958 15000 22926 15056
rect 22982 15000 22987 15056
rect 19628 14998 22987 15000
rect 19628 14996 19634 14998
rect 20897 14995 20963 14998
rect 22921 14995 22987 14998
rect 24209 15058 24275 15061
rect 28574 15058 28580 15060
rect 24209 15056 28580 15058
rect 24209 15000 24214 15056
rect 24270 15000 28580 15056
rect 24209 14998 28580 15000
rect 24209 14995 24275 14998
rect 28574 14996 28580 14998
rect 28644 14996 28650 15060
rect 8017 14922 8083 14925
rect 9489 14922 9555 14925
rect 8017 14920 9555 14922
rect 8017 14864 8022 14920
rect 8078 14864 9494 14920
rect 9550 14864 9555 14920
rect 8017 14862 9555 14864
rect 8017 14859 8083 14862
rect 9489 14859 9555 14862
rect 11605 14922 11671 14925
rect 12249 14922 12315 14925
rect 11605 14920 12315 14922
rect 11605 14864 11610 14920
rect 11666 14864 12254 14920
rect 12310 14864 12315 14920
rect 11605 14862 12315 14864
rect 11605 14859 11671 14862
rect 12249 14859 12315 14862
rect 13813 14922 13879 14925
rect 24853 14922 24919 14925
rect 13813 14920 24919 14922
rect 13813 14864 13818 14920
rect 13874 14864 24858 14920
rect 24914 14864 24919 14920
rect 13813 14862 24919 14864
rect 13813 14859 13879 14862
rect 24853 14859 24919 14862
rect 26601 14922 26667 14925
rect 35065 14922 35131 14925
rect 26601 14920 35131 14922
rect 26601 14864 26606 14920
rect 26662 14864 35070 14920
rect 35126 14864 35131 14920
rect 26601 14862 35131 14864
rect 26601 14859 26667 14862
rect 35065 14859 35131 14862
rect 14641 14786 14707 14789
rect 16389 14786 16455 14789
rect 14641 14784 16455 14786
rect 14641 14728 14646 14784
rect 14702 14728 16394 14784
rect 16450 14728 16455 14784
rect 14641 14726 16455 14728
rect 14641 14723 14707 14726
rect 16389 14723 16455 14726
rect 17585 14786 17651 14789
rect 24761 14786 24827 14789
rect 17585 14784 24827 14786
rect 17585 14728 17590 14784
rect 17646 14728 24766 14784
rect 24822 14728 24827 14784
rect 17585 14726 24827 14728
rect 17585 14723 17651 14726
rect 24761 14723 24827 14726
rect 25313 14786 25379 14789
rect 28901 14786 28967 14789
rect 25313 14784 28967 14786
rect 25313 14728 25318 14784
rect 25374 14728 28906 14784
rect 28962 14728 28967 14784
rect 25313 14726 28967 14728
rect 25313 14723 25379 14726
rect 28901 14723 28967 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 14089 14650 14155 14653
rect 14273 14650 14339 14653
rect 19057 14650 19123 14653
rect 14089 14648 14339 14650
rect 14089 14592 14094 14648
rect 14150 14592 14278 14648
rect 14334 14592 14339 14648
rect 14089 14590 14339 14592
rect 14089 14587 14155 14590
rect 14273 14587 14339 14590
rect 17910 14648 19123 14650
rect 17910 14592 19062 14648
rect 19118 14592 19123 14648
rect 17910 14590 19123 14592
rect 13302 14452 13308 14516
rect 13372 14514 13378 14516
rect 17910 14514 17970 14590
rect 19057 14587 19123 14590
rect 19333 14650 19399 14653
rect 19977 14650 20043 14653
rect 27613 14650 27679 14653
rect 19333 14648 20043 14650
rect 19333 14592 19338 14648
rect 19394 14592 19982 14648
rect 20038 14592 20043 14648
rect 19333 14590 20043 14592
rect 19333 14587 19399 14590
rect 19977 14587 20043 14590
rect 26328 14648 27679 14650
rect 26328 14592 27618 14648
rect 27674 14592 27679 14648
rect 26328 14590 27679 14592
rect 18873 14514 18939 14517
rect 13372 14454 17970 14514
rect 18462 14512 18939 14514
rect 18462 14456 18878 14512
rect 18934 14456 18939 14512
rect 18462 14454 18939 14456
rect 13372 14452 13378 14454
rect 17585 14378 17651 14381
rect 18321 14378 18387 14381
rect 17585 14376 18387 14378
rect 17585 14320 17590 14376
rect 17646 14320 18326 14376
rect 18382 14320 18387 14376
rect 17585 14318 18387 14320
rect 17585 14315 17651 14318
rect 18321 14315 18387 14318
rect 17953 14242 18019 14245
rect 18462 14242 18522 14454
rect 18873 14451 18939 14454
rect 20253 14516 20319 14517
rect 20253 14512 20300 14516
rect 20364 14514 20370 14516
rect 22185 14514 22251 14517
rect 22461 14514 22527 14517
rect 20253 14456 20258 14512
rect 20253 14452 20300 14456
rect 20364 14454 20410 14514
rect 22185 14512 22527 14514
rect 22185 14456 22190 14512
rect 22246 14456 22466 14512
rect 22522 14456 22527 14512
rect 22185 14454 22527 14456
rect 20364 14452 20370 14454
rect 20253 14451 20319 14452
rect 22185 14451 22251 14454
rect 22461 14451 22527 14454
rect 23933 14514 23999 14517
rect 26328 14514 26388 14590
rect 27613 14587 27679 14590
rect 23933 14512 26388 14514
rect 23933 14456 23938 14512
rect 23994 14456 26388 14512
rect 23933 14454 26388 14456
rect 23933 14451 23999 14454
rect 18781 14378 18847 14381
rect 21214 14378 21220 14380
rect 18781 14376 21220 14378
rect 18781 14320 18786 14376
rect 18842 14320 21220 14376
rect 18781 14318 21220 14320
rect 18781 14315 18847 14318
rect 21214 14316 21220 14318
rect 21284 14316 21290 14380
rect 26049 14378 26115 14381
rect 26366 14378 26372 14380
rect 26049 14376 26372 14378
rect 26049 14320 26054 14376
rect 26110 14320 26372 14376
rect 26049 14318 26372 14320
rect 26049 14315 26115 14318
rect 26366 14316 26372 14318
rect 26436 14316 26442 14380
rect 26509 14378 26575 14381
rect 26969 14378 27035 14381
rect 26509 14376 27035 14378
rect 26509 14320 26514 14376
rect 26570 14320 26974 14376
rect 27030 14320 27035 14376
rect 26509 14318 27035 14320
rect 26509 14315 26575 14318
rect 26969 14315 27035 14318
rect 17953 14240 18522 14242
rect 17953 14184 17958 14240
rect 18014 14184 18522 14240
rect 17953 14182 18522 14184
rect 18781 14240 18847 14245
rect 18781 14184 18786 14240
rect 18842 14184 18847 14240
rect 17953 14179 18019 14182
rect 18781 14179 18847 14184
rect 19793 14242 19859 14245
rect 20069 14242 20135 14245
rect 19793 14240 20135 14242
rect 19793 14184 19798 14240
rect 19854 14184 20074 14240
rect 20130 14184 20135 14240
rect 19793 14182 20135 14184
rect 19793 14179 19859 14182
rect 20069 14179 20135 14182
rect 20253 14242 20319 14245
rect 26601 14242 26667 14245
rect 20253 14240 26667 14242
rect 20253 14184 20258 14240
rect 20314 14184 26606 14240
rect 26662 14184 26667 14240
rect 20253 14182 26667 14184
rect 20253 14179 20319 14182
rect 26601 14179 26667 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 15745 14106 15811 14109
rect 18413 14106 18479 14109
rect 18784 14106 18844 14179
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 23749 14106 23815 14109
rect 26969 14108 27035 14109
rect 15745 14104 23815 14106
rect 15745 14048 15750 14104
rect 15806 14048 18418 14104
rect 18474 14048 23754 14104
rect 23810 14048 23815 14104
rect 15745 14046 23815 14048
rect 15745 14043 15811 14046
rect 18413 14043 18479 14046
rect 23749 14043 23815 14046
rect 26918 14044 26924 14108
rect 26988 14106 27035 14108
rect 26988 14104 27080 14106
rect 27030 14048 27080 14104
rect 26988 14046 27080 14048
rect 26988 14044 27035 14046
rect 26969 14043 27035 14044
rect 4654 13908 4660 13972
rect 4724 13970 4730 13972
rect 4797 13970 4863 13973
rect 4724 13968 4863 13970
rect 4724 13912 4802 13968
rect 4858 13912 4863 13968
rect 4724 13910 4863 13912
rect 4724 13908 4730 13910
rect 4797 13907 4863 13910
rect 9765 13970 9831 13973
rect 12249 13970 12315 13973
rect 14733 13970 14799 13973
rect 9765 13968 14799 13970
rect 9765 13912 9770 13968
rect 9826 13912 12254 13968
rect 12310 13912 14738 13968
rect 14794 13912 14799 13968
rect 9765 13910 14799 13912
rect 9765 13907 9831 13910
rect 12249 13907 12315 13910
rect 14733 13907 14799 13910
rect 19333 13970 19399 13973
rect 20805 13970 20871 13973
rect 21449 13970 21515 13973
rect 19333 13968 21515 13970
rect 19333 13912 19338 13968
rect 19394 13912 20810 13968
rect 20866 13912 21454 13968
rect 21510 13912 21515 13968
rect 19333 13910 21515 13912
rect 19333 13907 19399 13910
rect 20805 13907 20871 13910
rect 21449 13907 21515 13910
rect 22921 13970 22987 13973
rect 26182 13970 26188 13972
rect 22921 13968 26188 13970
rect 22921 13912 22926 13968
rect 22982 13912 26188 13968
rect 22921 13910 26188 13912
rect 22921 13907 22987 13910
rect 26182 13908 26188 13910
rect 26252 13970 26258 13972
rect 27613 13970 27679 13973
rect 27981 13970 28047 13973
rect 26252 13968 27679 13970
rect 26252 13912 27618 13968
rect 27674 13912 27679 13968
rect 26252 13910 27679 13912
rect 26252 13908 26258 13910
rect 27613 13907 27679 13910
rect 27846 13968 28047 13970
rect 27846 13912 27986 13968
rect 28042 13912 28047 13968
rect 27846 13910 28047 13912
rect 16573 13834 16639 13837
rect 17309 13834 17375 13837
rect 16573 13832 17375 13834
rect 16573 13776 16578 13832
rect 16634 13776 17314 13832
rect 17370 13776 17375 13832
rect 16573 13774 17375 13776
rect 16573 13771 16639 13774
rect 17309 13771 17375 13774
rect 27153 13834 27219 13837
rect 27846 13834 27906 13910
rect 27981 13907 28047 13910
rect 27153 13832 27906 13834
rect 27153 13776 27158 13832
rect 27214 13776 27906 13832
rect 27153 13774 27906 13776
rect 27981 13834 28047 13837
rect 28901 13834 28967 13837
rect 27981 13832 28967 13834
rect 27981 13776 27986 13832
rect 28042 13776 28906 13832
rect 28962 13776 28967 13832
rect 27981 13774 28967 13776
rect 27153 13771 27219 13774
rect 27981 13771 28047 13774
rect 28901 13771 28967 13774
rect 29545 13832 29611 13837
rect 29545 13776 29550 13832
rect 29606 13776 29611 13832
rect 29545 13771 29611 13776
rect 16389 13698 16455 13701
rect 16941 13698 17007 13701
rect 16389 13696 17007 13698
rect 16389 13640 16394 13696
rect 16450 13640 16946 13696
rect 17002 13640 17007 13696
rect 16389 13638 17007 13640
rect 16389 13635 16455 13638
rect 16941 13635 17007 13638
rect 18873 13698 18939 13701
rect 19558 13698 19564 13700
rect 18873 13696 19564 13698
rect 18873 13640 18878 13696
rect 18934 13640 19564 13696
rect 18873 13638 19564 13640
rect 18873 13635 18939 13638
rect 19558 13636 19564 13638
rect 19628 13636 19634 13700
rect 19885 13698 19951 13701
rect 20478 13698 20484 13700
rect 19885 13696 20484 13698
rect 19885 13640 19890 13696
rect 19946 13640 20484 13696
rect 19885 13638 20484 13640
rect 19885 13635 19951 13638
rect 20478 13636 20484 13638
rect 20548 13636 20554 13700
rect 24526 13636 24532 13700
rect 24596 13698 24602 13700
rect 24669 13698 24735 13701
rect 24596 13696 24735 13698
rect 24596 13640 24674 13696
rect 24730 13640 24735 13696
rect 24596 13638 24735 13640
rect 24596 13636 24602 13638
rect 24669 13635 24735 13638
rect 24945 13698 25011 13701
rect 26734 13698 26740 13700
rect 24945 13696 26740 13698
rect 24945 13640 24950 13696
rect 25006 13640 26740 13696
rect 24945 13638 26740 13640
rect 24945 13635 25011 13638
rect 26734 13636 26740 13638
rect 26804 13636 26810 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 29548 13565 29608 13771
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 17401 13562 17467 13565
rect 18045 13562 18111 13565
rect 17401 13560 22110 13562
rect 17401 13504 17406 13560
rect 17462 13504 18050 13560
rect 18106 13504 22110 13560
rect 17401 13502 22110 13504
rect 17401 13499 17467 13502
rect 18045 13499 18111 13502
rect 13169 13426 13235 13429
rect 18045 13426 18111 13429
rect 13169 13424 18111 13426
rect 13169 13368 13174 13424
rect 13230 13368 18050 13424
rect 18106 13368 18111 13424
rect 13169 13366 18111 13368
rect 13169 13363 13235 13366
rect 18045 13363 18111 13366
rect 18321 13426 18387 13429
rect 18454 13426 18460 13428
rect 18321 13424 18460 13426
rect 18321 13368 18326 13424
rect 18382 13368 18460 13424
rect 18321 13366 18460 13368
rect 18321 13363 18387 13366
rect 18454 13364 18460 13366
rect 18524 13426 18530 13428
rect 21081 13426 21147 13429
rect 18524 13424 21147 13426
rect 18524 13368 21086 13424
rect 21142 13368 21147 13424
rect 18524 13366 21147 13368
rect 22050 13426 22110 13502
rect 23974 13500 23980 13564
rect 24044 13562 24050 13564
rect 25630 13562 25636 13564
rect 24044 13502 25636 13562
rect 24044 13500 24050 13502
rect 25630 13500 25636 13502
rect 25700 13500 25706 13564
rect 29545 13560 29611 13565
rect 29545 13504 29550 13560
rect 29606 13504 29611 13560
rect 29545 13499 29611 13504
rect 25957 13426 26023 13429
rect 30557 13426 30623 13429
rect 22050 13424 30623 13426
rect 22050 13368 25962 13424
rect 26018 13368 30562 13424
rect 30618 13368 30623 13424
rect 22050 13366 30623 13368
rect 18524 13364 18530 13366
rect 21081 13363 21147 13366
rect 25957 13363 26023 13366
rect 30557 13363 30623 13366
rect 19517 13292 19583 13293
rect 19517 13288 19564 13292
rect 19628 13290 19634 13292
rect 19517 13232 19522 13288
rect 19517 13228 19564 13232
rect 19628 13230 19674 13290
rect 19628 13228 19634 13230
rect 19517 13227 19583 13228
rect 19425 13154 19491 13157
rect 20161 13154 20227 13157
rect 23238 13154 23244 13156
rect 19425 13152 23244 13154
rect 19425 13096 19430 13152
rect 19486 13096 20166 13152
rect 20222 13096 23244 13152
rect 19425 13094 23244 13096
rect 19425 13091 19491 13094
rect 20161 13091 20227 13094
rect 23238 13092 23244 13094
rect 23308 13092 23314 13156
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 17401 13018 17467 13021
rect 21357 13018 21423 13021
rect 17401 13016 21423 13018
rect 17401 12960 17406 13016
rect 17462 12960 21362 13016
rect 21418 12960 21423 13016
rect 17401 12958 21423 12960
rect 17401 12955 17467 12958
rect 21357 12955 21423 12958
rect 8937 12880 9003 12885
rect 10133 12884 10199 12885
rect 10133 12882 10180 12884
rect 8937 12824 8942 12880
rect 8998 12824 9003 12880
rect 8937 12819 9003 12824
rect 10088 12880 10180 12882
rect 10088 12824 10138 12880
rect 10088 12822 10180 12824
rect 10133 12820 10180 12822
rect 10244 12820 10250 12884
rect 12157 12882 12223 12885
rect 12022 12880 12223 12882
rect 12022 12824 12162 12880
rect 12218 12824 12223 12880
rect 12022 12822 12223 12824
rect 10133 12819 10199 12820
rect 8661 12744 8727 12749
rect 8661 12688 8666 12744
rect 8722 12688 8727 12744
rect 8661 12683 8727 12688
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 8664 12477 8724 12683
rect 8661 12472 8727 12477
rect 8661 12416 8666 12472
rect 8722 12416 8727 12472
rect 8661 12411 8727 12416
rect 8569 12338 8635 12341
rect 8940 12338 9000 12819
rect 11145 12610 11211 12613
rect 11421 12610 11487 12613
rect 11145 12608 11487 12610
rect 11145 12552 11150 12608
rect 11206 12552 11426 12608
rect 11482 12552 11487 12608
rect 11145 12550 11487 12552
rect 11145 12547 11211 12550
rect 11421 12547 11487 12550
rect 12022 12477 12082 12822
rect 12157 12819 12223 12822
rect 20662 12820 20668 12884
rect 20732 12882 20738 12884
rect 22553 12882 22619 12885
rect 20732 12880 22619 12882
rect 20732 12824 22558 12880
rect 22614 12824 22619 12880
rect 20732 12822 22619 12824
rect 20732 12820 20738 12822
rect 22553 12819 22619 12822
rect 27613 12882 27679 12885
rect 27838 12882 27844 12884
rect 27613 12880 27844 12882
rect 27613 12824 27618 12880
rect 27674 12824 27844 12880
rect 27613 12822 27844 12824
rect 27613 12819 27679 12822
rect 27838 12820 27844 12822
rect 27908 12820 27914 12884
rect 17769 12746 17835 12749
rect 18086 12746 18092 12748
rect 17769 12744 18092 12746
rect 17769 12688 17774 12744
rect 17830 12688 18092 12744
rect 17769 12686 18092 12688
rect 17769 12683 17835 12686
rect 18086 12684 18092 12686
rect 18156 12684 18162 12748
rect 19701 12746 19767 12749
rect 25773 12746 25839 12749
rect 19701 12744 25839 12746
rect 19701 12688 19706 12744
rect 19762 12688 25778 12744
rect 25834 12688 25839 12744
rect 19701 12686 25839 12688
rect 19701 12683 19767 12686
rect 25773 12683 25839 12686
rect 27889 12746 27955 12749
rect 28022 12746 28028 12748
rect 27889 12744 28028 12746
rect 27889 12688 27894 12744
rect 27950 12688 28028 12744
rect 27889 12686 28028 12688
rect 27889 12683 27955 12686
rect 28022 12684 28028 12686
rect 28092 12684 28098 12748
rect 30741 12746 30807 12749
rect 36169 12746 36235 12749
rect 30741 12744 36235 12746
rect 30741 12688 30746 12744
rect 30802 12688 36174 12744
rect 36230 12688 36235 12744
rect 30741 12686 36235 12688
rect 30741 12683 30807 12686
rect 36169 12683 36235 12686
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 11973 12472 12082 12477
rect 11973 12416 11978 12472
rect 12034 12416 12082 12472
rect 11973 12414 12082 12416
rect 22277 12474 22343 12477
rect 24025 12474 24091 12477
rect 28809 12474 28875 12477
rect 22277 12472 22616 12474
rect 22277 12416 22282 12472
rect 22338 12416 22616 12472
rect 22277 12414 22616 12416
rect 11973 12411 12039 12414
rect 22277 12411 22343 12414
rect 9213 12338 9279 12341
rect 8569 12336 9279 12338
rect 8569 12280 8574 12336
rect 8630 12280 9218 12336
rect 9274 12280 9279 12336
rect 8569 12278 9279 12280
rect 8569 12275 8635 12278
rect 9213 12275 9279 12278
rect 10225 12338 10291 12341
rect 11145 12338 11211 12341
rect 10225 12336 11211 12338
rect 10225 12280 10230 12336
rect 10286 12280 11150 12336
rect 11206 12280 11211 12336
rect 10225 12278 11211 12280
rect 10225 12275 10291 12278
rect 11145 12275 11211 12278
rect 17033 12338 17099 12341
rect 21541 12338 21607 12341
rect 17033 12336 21607 12338
rect 17033 12280 17038 12336
rect 17094 12280 21546 12336
rect 21602 12280 21607 12336
rect 17033 12278 21607 12280
rect 17033 12275 17099 12278
rect 21541 12275 21607 12278
rect 19793 12202 19859 12205
rect 21909 12202 21975 12205
rect 19793 12200 21975 12202
rect 19793 12144 19798 12200
rect 19854 12144 21914 12200
rect 21970 12144 21975 12200
rect 19793 12142 21975 12144
rect 19793 12139 19859 12142
rect 21909 12139 21975 12142
rect 22556 12069 22616 12414
rect 24025 12472 28875 12474
rect 24025 12416 24030 12472
rect 24086 12416 28814 12472
rect 28870 12416 28875 12472
rect 24025 12414 28875 12416
rect 24025 12411 24091 12414
rect 28809 12411 28875 12414
rect 30741 12474 30807 12477
rect 32070 12474 32076 12476
rect 30741 12472 32076 12474
rect 30741 12416 30746 12472
rect 30802 12416 32076 12472
rect 30741 12414 32076 12416
rect 30741 12411 30807 12414
rect 32070 12412 32076 12414
rect 32140 12412 32146 12476
rect 25129 12338 25195 12341
rect 25681 12338 25747 12341
rect 25129 12336 25747 12338
rect 25129 12280 25134 12336
rect 25190 12280 25686 12336
rect 25742 12280 25747 12336
rect 25129 12278 25747 12280
rect 25129 12275 25195 12278
rect 25681 12275 25747 12278
rect 26785 12338 26851 12341
rect 27102 12338 27108 12340
rect 26785 12336 27108 12338
rect 26785 12280 26790 12336
rect 26846 12280 27108 12336
rect 26785 12278 27108 12280
rect 26785 12275 26851 12278
rect 27102 12276 27108 12278
rect 27172 12338 27178 12340
rect 28165 12338 28231 12341
rect 27172 12336 28231 12338
rect 27172 12280 28170 12336
rect 28226 12280 28231 12336
rect 27172 12278 28231 12280
rect 27172 12276 27178 12278
rect 28165 12275 28231 12278
rect 31661 12338 31727 12341
rect 31886 12338 31892 12340
rect 31661 12336 31892 12338
rect 31661 12280 31666 12336
rect 31722 12280 31892 12336
rect 31661 12278 31892 12280
rect 31661 12275 31727 12278
rect 31886 12276 31892 12278
rect 31956 12276 31962 12340
rect 23381 12202 23447 12205
rect 27613 12202 27679 12205
rect 23381 12200 27679 12202
rect 23381 12144 23386 12200
rect 23442 12144 27618 12200
rect 27674 12144 27679 12200
rect 23381 12142 27679 12144
rect 23381 12139 23447 12142
rect 27613 12139 27679 12142
rect 17309 12066 17375 12069
rect 17534 12066 17540 12068
rect 17309 12064 17540 12066
rect 17309 12008 17314 12064
rect 17370 12008 17540 12064
rect 17309 12006 17540 12008
rect 17309 12003 17375 12006
rect 17534 12004 17540 12006
rect 17604 12066 17610 12068
rect 22318 12066 22324 12068
rect 17604 12006 22324 12066
rect 17604 12004 17610 12006
rect 22318 12004 22324 12006
rect 22388 12004 22394 12068
rect 22553 12066 22619 12069
rect 28717 12066 28783 12069
rect 22553 12064 28783 12066
rect 22553 12008 22558 12064
rect 22614 12008 28722 12064
rect 28778 12008 28783 12064
rect 22553 12006 28783 12008
rect 22553 12003 22619 12006
rect 28717 12003 28783 12006
rect 34646 12004 34652 12068
rect 34716 12066 34722 12068
rect 34881 12066 34947 12069
rect 34716 12064 34947 12066
rect 34716 12008 34886 12064
rect 34942 12008 34947 12064
rect 34716 12006 34947 12008
rect 34716 12004 34722 12006
rect 34881 12003 34947 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 19057 11932 19123 11933
rect 19006 11868 19012 11932
rect 19076 11930 19123 11932
rect 20713 11930 20779 11933
rect 23749 11930 23815 11933
rect 23933 11930 23999 11933
rect 27153 11930 27219 11933
rect 19076 11928 19168 11930
rect 19118 11872 19168 11928
rect 19076 11870 19168 11872
rect 20713 11928 21788 11930
rect 20713 11872 20718 11928
rect 20774 11872 21788 11928
rect 20713 11870 21788 11872
rect 19076 11868 19123 11870
rect 19057 11867 19123 11868
rect 20713 11867 20779 11870
rect 16246 11732 16252 11796
rect 16316 11794 16322 11796
rect 16481 11794 16547 11797
rect 16316 11792 16547 11794
rect 16316 11736 16486 11792
rect 16542 11736 16547 11792
rect 16316 11734 16547 11736
rect 16316 11732 16322 11734
rect 16481 11731 16547 11734
rect 20621 11794 20687 11797
rect 21541 11794 21607 11797
rect 20621 11792 21607 11794
rect 20621 11736 20626 11792
rect 20682 11736 21546 11792
rect 21602 11736 21607 11792
rect 20621 11734 21607 11736
rect 21728 11794 21788 11870
rect 23749 11928 27219 11930
rect 23749 11872 23754 11928
rect 23810 11872 23938 11928
rect 23994 11872 27158 11928
rect 27214 11872 27219 11928
rect 23749 11870 27219 11872
rect 23749 11867 23815 11870
rect 23933 11867 23999 11870
rect 27153 11867 27219 11870
rect 33041 11794 33107 11797
rect 33317 11796 33383 11797
rect 33317 11794 33364 11796
rect 21728 11734 29010 11794
rect 20621 11731 20687 11734
rect 21541 11731 21607 11734
rect 13721 11658 13787 11661
rect 20110 11658 20116 11660
rect 13721 11656 20116 11658
rect 13721 11600 13726 11656
rect 13782 11600 20116 11656
rect 13721 11598 20116 11600
rect 13721 11595 13787 11598
rect 20110 11596 20116 11598
rect 20180 11658 20186 11660
rect 23381 11658 23447 11661
rect 20180 11656 23447 11658
rect 20180 11600 23386 11656
rect 23442 11600 23447 11656
rect 20180 11598 23447 11600
rect 20180 11596 20186 11598
rect 23381 11595 23447 11598
rect 27153 11658 27219 11661
rect 27286 11658 27292 11660
rect 27153 11656 27292 11658
rect 27153 11600 27158 11656
rect 27214 11600 27292 11656
rect 27153 11598 27292 11600
rect 27153 11595 27219 11598
rect 27286 11596 27292 11598
rect 27356 11596 27362 11660
rect 18321 11524 18387 11525
rect 19241 11524 19307 11525
rect 20345 11524 20411 11525
rect 21265 11524 21331 11525
rect 18270 11460 18276 11524
rect 18340 11522 18387 11524
rect 18340 11520 18432 11522
rect 18382 11464 18432 11520
rect 18340 11462 18432 11464
rect 18340 11460 18387 11462
rect 19190 11460 19196 11524
rect 19260 11522 19307 11524
rect 19260 11520 19352 11522
rect 19302 11464 19352 11520
rect 19260 11462 19352 11464
rect 19260 11460 19307 11462
rect 20294 11460 20300 11524
rect 20364 11522 20411 11524
rect 20364 11520 20456 11522
rect 20406 11464 20456 11520
rect 20364 11462 20456 11464
rect 20364 11460 20411 11462
rect 21214 11460 21220 11524
rect 21284 11522 21331 11524
rect 21284 11520 21376 11522
rect 21326 11464 21376 11520
rect 21284 11462 21376 11464
rect 21284 11460 21331 11462
rect 21950 11460 21956 11524
rect 22020 11522 22026 11524
rect 22502 11522 22508 11524
rect 22020 11462 22508 11522
rect 22020 11460 22026 11462
rect 22502 11460 22508 11462
rect 22572 11460 22578 11524
rect 23238 11460 23244 11524
rect 23308 11522 23314 11524
rect 23657 11522 23723 11525
rect 24209 11522 24275 11525
rect 23308 11520 23723 11522
rect 23308 11464 23662 11520
rect 23718 11464 23723 11520
rect 23308 11462 23723 11464
rect 23308 11460 23314 11462
rect 18321 11459 18387 11460
rect 19241 11459 19307 11460
rect 20345 11459 20411 11460
rect 21265 11459 21331 11460
rect 23657 11459 23723 11462
rect 23982 11520 24275 11522
rect 23982 11464 24214 11520
rect 24270 11464 24275 11520
rect 23982 11462 24275 11464
rect 28950 11522 29010 11734
rect 33041 11792 33364 11794
rect 33041 11736 33046 11792
rect 33102 11736 33322 11792
rect 33041 11734 33364 11736
rect 33041 11731 33107 11734
rect 33317 11732 33364 11734
rect 33428 11732 33434 11796
rect 33317 11731 33383 11732
rect 29177 11660 29243 11661
rect 29545 11660 29611 11661
rect 29126 11596 29132 11660
rect 29196 11658 29243 11660
rect 29196 11656 29288 11658
rect 29238 11600 29288 11656
rect 29196 11598 29288 11600
rect 29196 11596 29243 11598
rect 29494 11596 29500 11660
rect 29564 11658 29611 11660
rect 29564 11656 29656 11658
rect 29606 11600 29656 11656
rect 29564 11598 29656 11600
rect 29564 11596 29611 11598
rect 29177 11595 29243 11596
rect 29545 11595 29611 11596
rect 31109 11522 31175 11525
rect 28950 11520 31175 11522
rect 28950 11464 31114 11520
rect 31170 11464 31175 11520
rect 28950 11462 31175 11464
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 23982 11389 24042 11462
rect 24209 11459 24275 11462
rect 31109 11459 31175 11462
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 13629 11386 13695 11389
rect 22829 11386 22895 11389
rect 23054 11386 23060 11388
rect 13629 11384 22570 11386
rect 13629 11328 13634 11384
rect 13690 11328 22570 11384
rect 13629 11326 22570 11328
rect 13629 11323 13695 11326
rect 12985 11250 13051 11253
rect 13118 11250 13124 11252
rect 12985 11248 13124 11250
rect 12985 11192 12990 11248
rect 13046 11192 13124 11248
rect 12985 11190 13124 11192
rect 12985 11187 13051 11190
rect 13118 11188 13124 11190
rect 13188 11188 13194 11252
rect 16614 11188 16620 11252
rect 16684 11250 16690 11252
rect 16757 11250 16823 11253
rect 16684 11248 16823 11250
rect 16684 11192 16762 11248
rect 16818 11192 16823 11248
rect 16684 11190 16823 11192
rect 16684 11188 16690 11190
rect 16757 11187 16823 11190
rect 17125 11250 17191 11253
rect 19333 11250 19399 11253
rect 19742 11250 19748 11252
rect 17125 11248 19748 11250
rect 17125 11192 17130 11248
rect 17186 11192 19338 11248
rect 19394 11192 19748 11248
rect 17125 11190 19748 11192
rect 17125 11187 17191 11190
rect 19333 11187 19399 11190
rect 19742 11188 19748 11190
rect 19812 11188 19818 11252
rect 19885 11250 19951 11253
rect 21173 11250 21239 11253
rect 19885 11248 21239 11250
rect 19885 11192 19890 11248
rect 19946 11192 21178 11248
rect 21234 11192 21239 11248
rect 19885 11190 21239 11192
rect 19885 11187 19951 11190
rect 21173 11187 21239 11190
rect 21357 11250 21423 11253
rect 21582 11250 21588 11252
rect 21357 11248 21588 11250
rect 21357 11192 21362 11248
rect 21418 11192 21588 11248
rect 21357 11190 21588 11192
rect 21357 11187 21423 11190
rect 21582 11188 21588 11190
rect 21652 11188 21658 11252
rect 22510 11250 22570 11326
rect 22829 11384 23060 11386
rect 22829 11328 22834 11384
rect 22890 11328 23060 11384
rect 22829 11326 23060 11328
rect 22829 11323 22895 11326
rect 23054 11324 23060 11326
rect 23124 11324 23130 11388
rect 23933 11384 24042 11389
rect 28165 11388 28231 11389
rect 28165 11386 28212 11388
rect 23933 11328 23938 11384
rect 23994 11328 24042 11384
rect 23933 11326 24042 11328
rect 28120 11384 28212 11386
rect 28120 11328 28170 11384
rect 28120 11326 28212 11328
rect 23933 11323 23999 11326
rect 28165 11324 28212 11326
rect 28276 11324 28282 11388
rect 28165 11323 28231 11324
rect 24485 11250 24551 11253
rect 22510 11248 27722 11250
rect 22510 11192 24490 11248
rect 24546 11192 27722 11248
rect 22510 11190 27722 11192
rect 24485 11187 24551 11190
rect 20345 11114 20411 11117
rect 20846 11114 20852 11116
rect 20345 11112 20852 11114
rect 20345 11056 20350 11112
rect 20406 11056 20852 11112
rect 20345 11054 20852 11056
rect 20345 11051 20411 11054
rect 20846 11052 20852 11054
rect 20916 11052 20922 11116
rect 22277 11114 22343 11117
rect 23841 11114 23907 11117
rect 22277 11112 23907 11114
rect 22277 11056 22282 11112
rect 22338 11056 23846 11112
rect 23902 11056 23907 11112
rect 22277 11054 23907 11056
rect 22277 11051 22343 11054
rect 23841 11051 23907 11054
rect 20897 10978 20963 10981
rect 21173 10978 21239 10981
rect 26233 10978 26299 10981
rect 20897 10976 26299 10978
rect 20897 10920 20902 10976
rect 20958 10920 21178 10976
rect 21234 10920 26238 10976
rect 26294 10920 26299 10976
rect 20897 10918 26299 10920
rect 27662 10978 27722 11190
rect 28349 11114 28415 11117
rect 29545 11114 29611 11117
rect 28349 11112 29611 11114
rect 28349 11056 28354 11112
rect 28410 11056 29550 11112
rect 29606 11056 29611 11112
rect 28349 11054 29611 11056
rect 28349 11051 28415 11054
rect 29545 11051 29611 11054
rect 34094 11052 34100 11116
rect 34164 11114 34170 11116
rect 34329 11114 34395 11117
rect 34164 11112 34395 11114
rect 34164 11056 34334 11112
rect 34390 11056 34395 11112
rect 34164 11054 34395 11056
rect 34164 11052 34170 11054
rect 34329 11051 34395 11054
rect 27797 10978 27863 10981
rect 27662 10976 27863 10978
rect 27662 10920 27802 10976
rect 27858 10920 27863 10976
rect 27662 10918 27863 10920
rect 20897 10915 20963 10918
rect 21173 10915 21239 10918
rect 26233 10915 26299 10918
rect 27797 10915 27863 10918
rect 29269 10978 29335 10981
rect 30414 10978 30420 10980
rect 29269 10976 30420 10978
rect 29269 10920 29274 10976
rect 29330 10920 30420 10976
rect 29269 10918 30420 10920
rect 29269 10915 29335 10918
rect 30414 10916 30420 10918
rect 30484 10916 30490 10980
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 23841 10842 23907 10845
rect 23974 10842 23980 10844
rect 22050 10840 23980 10842
rect 22050 10784 23846 10840
rect 23902 10784 23980 10840
rect 22050 10782 23980 10784
rect 10777 10706 10843 10709
rect 12893 10706 12959 10709
rect 10777 10704 12959 10706
rect 10777 10648 10782 10704
rect 10838 10648 12898 10704
rect 12954 10648 12959 10704
rect 10777 10646 12959 10648
rect 10777 10643 10843 10646
rect 12893 10643 12959 10646
rect 18873 10706 18939 10709
rect 22050 10706 22110 10782
rect 23841 10779 23907 10782
rect 23974 10780 23980 10782
rect 24044 10780 24050 10844
rect 24342 10780 24348 10844
rect 24412 10842 24418 10844
rect 24485 10842 24551 10845
rect 24412 10840 24551 10842
rect 24412 10784 24490 10840
rect 24546 10784 24551 10840
rect 24412 10782 24551 10784
rect 24412 10780 24418 10782
rect 24485 10779 24551 10782
rect 18873 10704 22110 10706
rect 18873 10648 18878 10704
rect 18934 10648 22110 10704
rect 18873 10646 22110 10648
rect 26417 10706 26483 10709
rect 29913 10706 29979 10709
rect 26417 10704 29979 10706
rect 26417 10648 26422 10704
rect 26478 10648 29918 10704
rect 29974 10648 29979 10704
rect 26417 10646 29979 10648
rect 18873 10643 18939 10646
rect 26417 10643 26483 10646
rect 29913 10643 29979 10646
rect 19558 10508 19564 10572
rect 19628 10570 19634 10572
rect 26693 10570 26759 10573
rect 34053 10570 34119 10573
rect 19628 10568 34119 10570
rect 19628 10512 26698 10568
rect 26754 10512 34058 10568
rect 34114 10512 34119 10568
rect 19628 10510 34119 10512
rect 19628 10508 19634 10510
rect 26693 10507 26759 10510
rect 34053 10507 34119 10510
rect 19333 10434 19399 10437
rect 20253 10434 20319 10437
rect 23013 10434 23079 10437
rect 23933 10434 23999 10437
rect 26969 10434 27035 10437
rect 19333 10432 27035 10434
rect 19333 10376 19338 10432
rect 19394 10376 20258 10432
rect 20314 10376 23018 10432
rect 23074 10376 23938 10432
rect 23994 10376 26974 10432
rect 27030 10376 27035 10432
rect 19333 10374 27035 10376
rect 19333 10371 19399 10374
rect 20253 10371 20319 10374
rect 23013 10371 23079 10374
rect 23933 10371 23999 10374
rect 26969 10371 27035 10374
rect 28165 10434 28231 10437
rect 29085 10434 29151 10437
rect 28165 10432 29151 10434
rect 28165 10376 28170 10432
rect 28226 10376 29090 10432
rect 29146 10376 29151 10432
rect 28165 10374 29151 10376
rect 28165 10371 28231 10374
rect 29085 10371 29151 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 17677 10300 17743 10301
rect 17677 10298 17724 10300
rect 17632 10296 17724 10298
rect 17632 10240 17682 10296
rect 17632 10238 17724 10240
rect 17677 10236 17724 10238
rect 17788 10236 17794 10300
rect 20069 10298 20135 10301
rect 26417 10298 26483 10301
rect 20069 10296 26483 10298
rect 20069 10240 20074 10296
rect 20130 10240 26422 10296
rect 26478 10240 26483 10296
rect 20069 10238 26483 10240
rect 17677 10235 17743 10236
rect 20069 10235 20135 10238
rect 26417 10235 26483 10238
rect 28022 10236 28028 10300
rect 28092 10298 28098 10300
rect 28533 10298 28599 10301
rect 28092 10296 28599 10298
rect 28092 10240 28538 10296
rect 28594 10240 28599 10296
rect 28092 10238 28599 10240
rect 28092 10236 28098 10238
rect 28533 10235 28599 10238
rect 5901 10164 5967 10165
rect 5901 10162 5948 10164
rect 5856 10160 5948 10162
rect 5856 10104 5906 10160
rect 5856 10102 5948 10104
rect 5901 10100 5948 10102
rect 6012 10100 6018 10164
rect 6085 10162 6151 10165
rect 6729 10162 6795 10165
rect 8661 10162 8727 10165
rect 6085 10160 8727 10162
rect 6085 10104 6090 10160
rect 6146 10104 6734 10160
rect 6790 10104 8666 10160
rect 8722 10104 8727 10160
rect 6085 10102 8727 10104
rect 5901 10099 5967 10100
rect 6085 10099 6151 10102
rect 6729 10099 6795 10102
rect 8661 10099 8727 10102
rect 9673 10162 9739 10165
rect 10225 10162 10291 10165
rect 9673 10160 10291 10162
rect 9673 10104 9678 10160
rect 9734 10104 10230 10160
rect 10286 10104 10291 10160
rect 9673 10102 10291 10104
rect 9673 10099 9739 10102
rect 10225 10099 10291 10102
rect 16205 10162 16271 10165
rect 17217 10162 17283 10165
rect 16205 10160 17283 10162
rect 16205 10104 16210 10160
rect 16266 10104 17222 10160
rect 17278 10104 17283 10160
rect 16205 10102 17283 10104
rect 16205 10099 16271 10102
rect 17217 10099 17283 10102
rect 21633 10162 21699 10165
rect 26417 10164 26483 10165
rect 21950 10162 21956 10164
rect 21633 10160 21956 10162
rect 21633 10104 21638 10160
rect 21694 10104 21956 10160
rect 21633 10102 21956 10104
rect 21633 10099 21699 10102
rect 21950 10100 21956 10102
rect 22020 10100 22026 10164
rect 26366 10100 26372 10164
rect 26436 10162 26483 10164
rect 28073 10162 28139 10165
rect 29269 10162 29335 10165
rect 26436 10160 26528 10162
rect 26478 10104 26528 10160
rect 26436 10102 26528 10104
rect 28073 10160 29335 10162
rect 28073 10104 28078 10160
rect 28134 10104 29274 10160
rect 29330 10104 29335 10160
rect 28073 10102 29335 10104
rect 26436 10100 26483 10102
rect 26417 10099 26483 10100
rect 28073 10099 28139 10102
rect 29269 10099 29335 10102
rect 11237 10026 11303 10029
rect 11605 10026 11671 10029
rect 11237 10024 11671 10026
rect 11237 9968 11242 10024
rect 11298 9968 11610 10024
rect 11666 9968 11671 10024
rect 11237 9966 11671 9968
rect 11237 9963 11303 9966
rect 11605 9963 11671 9966
rect 16757 10026 16823 10029
rect 17309 10026 17375 10029
rect 16757 10024 17375 10026
rect 16757 9968 16762 10024
rect 16818 9968 17314 10024
rect 17370 9968 17375 10024
rect 16757 9966 17375 9968
rect 16757 9963 16823 9966
rect 17309 9963 17375 9966
rect 20161 10026 20227 10029
rect 20989 10026 21055 10029
rect 27889 10028 27955 10029
rect 20161 10024 21055 10026
rect 20161 9968 20166 10024
rect 20222 9968 20994 10024
rect 21050 9968 21055 10024
rect 20161 9966 21055 9968
rect 20161 9963 20227 9966
rect 20989 9963 21055 9966
rect 27838 9964 27844 10028
rect 27908 10026 27955 10028
rect 27908 10024 28000 10026
rect 27950 9968 28000 10024
rect 27908 9966 28000 9968
rect 27908 9964 27955 9966
rect 28758 9964 28764 10028
rect 28828 10026 28834 10028
rect 28901 10026 28967 10029
rect 28828 10024 28967 10026
rect 28828 9968 28906 10024
rect 28962 9968 28967 10024
rect 28828 9966 28967 9968
rect 28828 9964 28834 9966
rect 27889 9963 27955 9964
rect 28901 9963 28967 9966
rect 31201 10026 31267 10029
rect 31753 10026 31819 10029
rect 31201 10024 31819 10026
rect 31201 9968 31206 10024
rect 31262 9968 31758 10024
rect 31814 9968 31819 10024
rect 31201 9966 31819 9968
rect 31201 9963 31267 9966
rect 31753 9963 31819 9966
rect 27153 9890 27219 9893
rect 29269 9890 29335 9893
rect 29821 9890 29887 9893
rect 27153 9888 29887 9890
rect 27153 9832 27158 9888
rect 27214 9832 29274 9888
rect 29330 9832 29826 9888
rect 29882 9832 29887 9888
rect 27153 9830 29887 9832
rect 27153 9827 27219 9830
rect 29269 9827 29335 9830
rect 29821 9827 29887 9830
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 19517 9754 19583 9757
rect 28717 9754 28783 9757
rect 19517 9752 28783 9754
rect 19517 9696 19522 9752
rect 19578 9696 28722 9752
rect 28778 9696 28783 9752
rect 19517 9694 28783 9696
rect 19517 9691 19583 9694
rect 28717 9691 28783 9694
rect 14089 9618 14155 9621
rect 14774 9618 14780 9620
rect 14089 9616 14780 9618
rect 14089 9560 14094 9616
rect 14150 9560 14780 9616
rect 14089 9558 14780 9560
rect 14089 9555 14155 9558
rect 14774 9556 14780 9558
rect 14844 9618 14850 9620
rect 15009 9618 15075 9621
rect 14844 9616 15075 9618
rect 14844 9560 15014 9616
rect 15070 9560 15075 9616
rect 14844 9558 15075 9560
rect 14844 9556 14850 9558
rect 15009 9555 15075 9558
rect 15150 9558 22110 9618
rect 6177 9482 6243 9485
rect 6310 9482 6316 9484
rect 6177 9480 6316 9482
rect 6177 9424 6182 9480
rect 6238 9424 6316 9480
rect 6177 9422 6316 9424
rect 6177 9419 6243 9422
rect 6310 9420 6316 9422
rect 6380 9420 6386 9484
rect 13997 9482 14063 9485
rect 15150 9482 15210 9558
rect 13997 9480 15210 9482
rect 13997 9424 14002 9480
rect 14058 9424 15210 9480
rect 13997 9422 15210 9424
rect 16757 9480 16823 9485
rect 16757 9424 16762 9480
rect 16818 9424 16823 9480
rect 13997 9419 14063 9422
rect 16757 9419 16823 9424
rect 22050 9482 22110 9558
rect 22318 9556 22324 9620
rect 22388 9618 22394 9620
rect 22645 9618 22711 9621
rect 22388 9616 22711 9618
rect 22388 9560 22650 9616
rect 22706 9560 22711 9616
rect 22388 9558 22711 9560
rect 22388 9556 22394 9558
rect 22645 9555 22711 9558
rect 26734 9556 26740 9620
rect 26804 9618 26810 9620
rect 27153 9618 27219 9621
rect 26804 9616 27219 9618
rect 26804 9560 27158 9616
rect 27214 9560 27219 9616
rect 26804 9558 27219 9560
rect 26804 9556 26810 9558
rect 27153 9555 27219 9558
rect 27797 9618 27863 9621
rect 32673 9618 32739 9621
rect 27797 9616 32739 9618
rect 27797 9560 27802 9616
rect 27858 9560 32678 9616
rect 32734 9560 32739 9616
rect 27797 9558 32739 9560
rect 27797 9555 27863 9558
rect 32673 9555 32739 9558
rect 32857 9618 32923 9621
rect 34329 9618 34395 9621
rect 32857 9616 34395 9618
rect 32857 9560 32862 9616
rect 32918 9560 34334 9616
rect 34390 9560 34395 9616
rect 32857 9558 34395 9560
rect 32857 9555 32923 9558
rect 34329 9555 34395 9558
rect 22050 9422 22386 9482
rect 16760 9346 16820 9419
rect 18873 9346 18939 9349
rect 16760 9344 18939 9346
rect 16760 9288 18878 9344
rect 18934 9288 18939 9344
rect 16760 9286 18939 9288
rect 18873 9283 18939 9286
rect 20989 9346 21055 9349
rect 22326 9346 22386 9422
rect 23422 9420 23428 9484
rect 23492 9482 23498 9484
rect 23565 9482 23631 9485
rect 23492 9480 23631 9482
rect 23492 9424 23570 9480
rect 23626 9424 23631 9480
rect 23492 9422 23631 9424
rect 23492 9420 23498 9422
rect 23565 9419 23631 9422
rect 26182 9420 26188 9484
rect 26252 9482 26258 9484
rect 26252 9422 31770 9482
rect 26252 9420 26258 9422
rect 22829 9346 22895 9349
rect 26325 9346 26391 9349
rect 20989 9344 22110 9346
rect 20989 9288 20994 9344
rect 21050 9288 22110 9344
rect 20989 9286 22110 9288
rect 22326 9344 26391 9346
rect 22326 9288 22834 9344
rect 22890 9288 26330 9344
rect 26386 9288 26391 9344
rect 22326 9286 26391 9288
rect 31710 9346 31770 9422
rect 33225 9346 33291 9349
rect 31710 9344 33291 9346
rect 31710 9288 33230 9344
rect 33286 9288 33291 9344
rect 31710 9286 33291 9288
rect 20989 9283 21055 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 15193 9212 15259 9213
rect 15142 9148 15148 9212
rect 15212 9210 15259 9212
rect 17861 9210 17927 9213
rect 18137 9210 18203 9213
rect 18597 9212 18663 9213
rect 18597 9210 18644 9212
rect 15212 9208 15304 9210
rect 15254 9152 15304 9208
rect 15212 9150 15304 9152
rect 17861 9208 18203 9210
rect 17861 9152 17866 9208
rect 17922 9152 18142 9208
rect 18198 9152 18203 9208
rect 17861 9150 18203 9152
rect 18552 9208 18644 9210
rect 18552 9152 18602 9208
rect 18552 9150 18644 9152
rect 15212 9148 15259 9150
rect 15193 9147 15259 9148
rect 17861 9147 17927 9150
rect 18137 9147 18203 9150
rect 18597 9148 18644 9150
rect 18708 9148 18714 9212
rect 21081 9210 21147 9213
rect 21449 9210 21515 9213
rect 21081 9208 21515 9210
rect 21081 9152 21086 9208
rect 21142 9152 21454 9208
rect 21510 9152 21515 9208
rect 21081 9150 21515 9152
rect 22050 9210 22110 9286
rect 22829 9283 22895 9286
rect 26325 9283 26391 9286
rect 33225 9283 33291 9286
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 22553 9210 22619 9213
rect 28390 9210 28396 9212
rect 22050 9150 22386 9210
rect 18597 9147 18663 9148
rect 21081 9147 21147 9150
rect 21449 9147 21515 9150
rect 19241 9074 19307 9077
rect 20253 9074 20319 9077
rect 19241 9072 20319 9074
rect 19241 9016 19246 9072
rect 19302 9016 20258 9072
rect 20314 9016 20319 9072
rect 19241 9014 20319 9016
rect 22326 9074 22386 9150
rect 22553 9208 28396 9210
rect 22553 9152 22558 9208
rect 22614 9152 28396 9208
rect 22553 9150 28396 9152
rect 22553 9147 22619 9150
rect 28390 9148 28396 9150
rect 28460 9210 28466 9212
rect 28717 9210 28783 9213
rect 28460 9208 28783 9210
rect 28460 9152 28722 9208
rect 28778 9152 28783 9208
rect 28460 9150 28783 9152
rect 28460 9148 28466 9150
rect 28717 9147 28783 9150
rect 26182 9074 26188 9076
rect 22326 9014 26188 9074
rect 19241 9011 19307 9014
rect 20253 9011 20319 9014
rect 26182 9012 26188 9014
rect 26252 9012 26258 9076
rect 20437 8938 20503 8941
rect 28349 8938 28415 8941
rect 20437 8936 28415 8938
rect 20437 8880 20442 8936
rect 20498 8880 28354 8936
rect 28410 8880 28415 8936
rect 20437 8878 28415 8880
rect 20437 8875 20503 8878
rect 28349 8875 28415 8878
rect 20253 8802 20319 8805
rect 21398 8802 21404 8804
rect 20253 8800 21404 8802
rect 20253 8744 20258 8800
rect 20314 8744 21404 8800
rect 20253 8742 21404 8744
rect 20253 8739 20319 8742
rect 21398 8740 21404 8742
rect 21468 8802 21474 8804
rect 31518 8802 31524 8804
rect 21468 8742 31524 8802
rect 21468 8740 21474 8742
rect 31518 8740 31524 8742
rect 31588 8802 31594 8804
rect 31661 8802 31727 8805
rect 31588 8800 31727 8802
rect 31588 8744 31666 8800
rect 31722 8744 31727 8800
rect 31588 8742 31727 8744
rect 31588 8740 31594 8742
rect 31661 8739 31727 8742
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 22737 8666 22803 8669
rect 22870 8666 22876 8668
rect 22737 8664 22876 8666
rect 22737 8608 22742 8664
rect 22798 8608 22876 8664
rect 22737 8606 22876 8608
rect 22737 8603 22803 8606
rect 22870 8604 22876 8606
rect 22940 8604 22946 8668
rect 23013 8666 23079 8669
rect 25681 8666 25747 8669
rect 23013 8664 25747 8666
rect 23013 8608 23018 8664
rect 23074 8608 25686 8664
rect 25742 8608 25747 8664
rect 23013 8606 25747 8608
rect 23013 8603 23079 8606
rect 25681 8603 25747 8606
rect 14825 8530 14891 8533
rect 19333 8532 19399 8533
rect 14958 8530 14964 8532
rect 14825 8528 14964 8530
rect 14825 8472 14830 8528
rect 14886 8472 14964 8528
rect 14825 8470 14964 8472
rect 14825 8467 14891 8470
rect 14958 8468 14964 8470
rect 15028 8468 15034 8532
rect 19333 8528 19380 8532
rect 19444 8530 19450 8532
rect 21265 8530 21331 8533
rect 25957 8530 26023 8533
rect 19333 8472 19338 8528
rect 19333 8468 19380 8472
rect 19444 8470 19490 8530
rect 21265 8528 26023 8530
rect 21265 8472 21270 8528
rect 21326 8472 25962 8528
rect 26018 8472 26023 8528
rect 21265 8470 26023 8472
rect 19444 8468 19450 8470
rect 19333 8467 19399 8468
rect 21265 8467 21331 8470
rect 25957 8467 26023 8470
rect 19517 8396 19583 8397
rect 19517 8394 19564 8396
rect 19472 8392 19564 8394
rect 19472 8336 19522 8392
rect 19472 8334 19564 8336
rect 19517 8332 19564 8334
rect 19628 8332 19634 8396
rect 20478 8332 20484 8396
rect 20548 8394 20554 8396
rect 21081 8394 21147 8397
rect 27889 8394 27955 8397
rect 28574 8394 28580 8396
rect 20548 8392 21834 8394
rect 20548 8336 21086 8392
rect 21142 8336 21834 8392
rect 20548 8334 21834 8336
rect 20548 8332 20554 8334
rect 19517 8331 19583 8332
rect 21081 8331 21147 8334
rect 19149 8258 19215 8261
rect 20621 8258 20687 8261
rect 19149 8256 20687 8258
rect 19149 8200 19154 8256
rect 19210 8200 20626 8256
rect 20682 8200 20687 8256
rect 19149 8198 20687 8200
rect 19149 8195 19215 8198
rect 20621 8195 20687 8198
rect 21173 8260 21239 8261
rect 21173 8256 21220 8260
rect 21284 8258 21290 8260
rect 21173 8200 21178 8256
rect 21173 8196 21220 8200
rect 21284 8198 21330 8258
rect 21284 8196 21290 8198
rect 21173 8195 21239 8196
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 11237 8124 11303 8125
rect 13445 8124 13511 8125
rect 11237 8122 11284 8124
rect 11192 8120 11284 8122
rect 11192 8064 11242 8120
rect 11192 8062 11284 8064
rect 11237 8060 11284 8062
rect 11348 8060 11354 8124
rect 13445 8122 13492 8124
rect 13400 8120 13492 8122
rect 13400 8064 13450 8120
rect 13400 8062 13492 8064
rect 13445 8060 13492 8062
rect 13556 8060 13562 8124
rect 21774 8122 21834 8334
rect 22142 8392 28580 8394
rect 22142 8336 27894 8392
rect 27950 8336 28580 8392
rect 22142 8334 28580 8336
rect 22001 8260 22067 8261
rect 21950 8258 21956 8260
rect 21910 8198 21956 8258
rect 22020 8256 22067 8260
rect 22062 8200 22067 8256
rect 21950 8196 21956 8198
rect 22020 8196 22067 8200
rect 22001 8195 22067 8196
rect 22142 8122 22202 8334
rect 27889 8331 27955 8334
rect 28574 8332 28580 8334
rect 28644 8394 28650 8396
rect 29821 8394 29887 8397
rect 28644 8392 29887 8394
rect 28644 8336 29826 8392
rect 29882 8336 29887 8392
rect 28644 8334 29887 8336
rect 28644 8332 28650 8334
rect 29821 8331 29887 8334
rect 25497 8258 25563 8261
rect 27613 8258 27679 8261
rect 25497 8256 27679 8258
rect 25497 8200 25502 8256
rect 25558 8200 27618 8256
rect 27674 8200 27679 8256
rect 25497 8198 27679 8200
rect 25497 8195 25563 8198
rect 27613 8195 27679 8198
rect 29453 8260 29519 8261
rect 29453 8256 29500 8260
rect 29564 8258 29570 8260
rect 29453 8200 29458 8256
rect 29453 8196 29500 8200
rect 29564 8198 29610 8258
rect 29564 8196 29570 8198
rect 29453 8195 29519 8196
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 21774 8062 22202 8122
rect 11237 8059 11303 8060
rect 13445 8059 13511 8060
rect 11145 7986 11211 7989
rect 11462 7986 11468 7988
rect 11145 7984 11468 7986
rect 11145 7928 11150 7984
rect 11206 7928 11468 7984
rect 11145 7926 11468 7928
rect 11145 7923 11211 7926
rect 11462 7924 11468 7926
rect 11532 7986 11538 7988
rect 15837 7986 15903 7989
rect 11532 7984 15903 7986
rect 11532 7928 15842 7984
rect 15898 7928 15903 7984
rect 11532 7926 15903 7928
rect 11532 7924 11538 7926
rect 15837 7923 15903 7926
rect 19333 7986 19399 7989
rect 19885 7986 19951 7989
rect 19333 7984 19951 7986
rect 19333 7928 19338 7984
rect 19394 7928 19890 7984
rect 19946 7928 19951 7984
rect 19333 7926 19951 7928
rect 19333 7923 19399 7926
rect 19885 7923 19951 7926
rect 21725 7986 21791 7989
rect 30557 7986 30623 7989
rect 21725 7984 30623 7986
rect 21725 7928 21730 7984
rect 21786 7928 30562 7984
rect 30618 7928 30623 7984
rect 21725 7926 30623 7928
rect 21725 7923 21791 7926
rect 30557 7923 30623 7926
rect 19425 7850 19491 7853
rect 19701 7850 19767 7853
rect 20161 7850 20227 7853
rect 22093 7850 22159 7853
rect 19425 7848 22159 7850
rect 19425 7792 19430 7848
rect 19486 7792 19706 7848
rect 19762 7792 20166 7848
rect 20222 7792 22098 7848
rect 22154 7792 22159 7848
rect 19425 7790 22159 7792
rect 19425 7787 19491 7790
rect 19701 7787 19767 7790
rect 20161 7787 20227 7790
rect 22093 7787 22159 7790
rect 15101 7714 15167 7717
rect 24393 7714 24459 7717
rect 15101 7712 24459 7714
rect 15101 7656 15106 7712
rect 15162 7656 24398 7712
rect 24454 7656 24459 7712
rect 15101 7654 24459 7656
rect 15101 7651 15167 7654
rect 24393 7651 24459 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 28758 7516 28764 7580
rect 28828 7578 28834 7580
rect 28993 7578 29059 7581
rect 28828 7576 29059 7578
rect 28828 7520 28998 7576
rect 29054 7520 29059 7576
rect 28828 7518 29059 7520
rect 28828 7516 28834 7518
rect 28993 7515 29059 7518
rect 11605 7442 11671 7445
rect 12525 7442 12591 7445
rect 17309 7444 17375 7445
rect 19333 7444 19399 7445
rect 17309 7442 17356 7444
rect 11605 7440 12591 7442
rect 11605 7384 11610 7440
rect 11666 7384 12530 7440
rect 12586 7384 12591 7440
rect 11605 7382 12591 7384
rect 17264 7440 17356 7442
rect 17264 7384 17314 7440
rect 17264 7382 17356 7384
rect 11605 7379 11671 7382
rect 12525 7379 12591 7382
rect 17309 7380 17356 7382
rect 17420 7380 17426 7444
rect 19333 7440 19380 7444
rect 19444 7442 19450 7444
rect 19609 7442 19675 7445
rect 23749 7442 23815 7445
rect 19333 7384 19338 7440
rect 19333 7380 19380 7384
rect 19444 7382 19490 7442
rect 19609 7440 23815 7442
rect 19609 7384 19614 7440
rect 19670 7384 23754 7440
rect 23810 7384 23815 7440
rect 19609 7382 23815 7384
rect 19444 7380 19450 7382
rect 17309 7379 17375 7380
rect 19333 7379 19399 7380
rect 19609 7379 19675 7382
rect 23749 7379 23815 7382
rect 12065 7306 12131 7309
rect 13997 7306 14063 7309
rect 12065 7304 14063 7306
rect 12065 7248 12070 7304
rect 12126 7248 14002 7304
rect 14058 7248 14063 7304
rect 12065 7246 14063 7248
rect 12065 7243 12131 7246
rect 13997 7243 14063 7246
rect 30557 7306 30623 7309
rect 32438 7306 32444 7308
rect 30557 7304 32444 7306
rect 30557 7248 30562 7304
rect 30618 7248 32444 7304
rect 30557 7246 32444 7248
rect 30557 7243 30623 7246
rect 32438 7244 32444 7246
rect 32508 7244 32514 7308
rect 11789 7170 11855 7173
rect 12249 7170 12315 7173
rect 14825 7170 14891 7173
rect 11789 7168 14891 7170
rect 11789 7112 11794 7168
rect 11850 7112 12254 7168
rect 12310 7112 14830 7168
rect 14886 7112 14891 7168
rect 11789 7110 14891 7112
rect 11789 7107 11855 7110
rect 12249 7107 12315 7110
rect 14825 7107 14891 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 21633 7036 21699 7037
rect 21582 6972 21588 7036
rect 21652 7034 21699 7036
rect 21652 7032 21744 7034
rect 21694 6976 21744 7032
rect 21652 6974 21744 6976
rect 21652 6972 21699 6974
rect 29862 6972 29868 7036
rect 29932 7034 29938 7036
rect 30189 7034 30255 7037
rect 29932 7032 30255 7034
rect 29932 6976 30194 7032
rect 30250 6976 30255 7032
rect 29932 6974 30255 6976
rect 29932 6972 29938 6974
rect 21633 6971 21699 6972
rect 30189 6971 30255 6974
rect 13670 6836 13676 6900
rect 13740 6898 13746 6900
rect 17769 6898 17835 6901
rect 13740 6896 17835 6898
rect 13740 6840 17774 6896
rect 17830 6840 17835 6896
rect 13740 6838 17835 6840
rect 13740 6836 13746 6838
rect 17769 6835 17835 6838
rect 31017 6898 31083 6901
rect 31150 6898 31156 6900
rect 31017 6896 31156 6898
rect 31017 6840 31022 6896
rect 31078 6840 31156 6896
rect 31017 6838 31156 6840
rect 31017 6835 31083 6838
rect 31150 6836 31156 6838
rect 31220 6836 31226 6900
rect 21909 6626 21975 6629
rect 27061 6626 27127 6629
rect 21909 6624 27127 6626
rect 21909 6568 21914 6624
rect 21970 6568 27066 6624
rect 27122 6568 27127 6624
rect 21909 6566 27127 6568
rect 21909 6563 21975 6566
rect 27061 6563 27127 6566
rect 28717 6626 28783 6629
rect 32254 6626 32260 6628
rect 28717 6624 32260 6626
rect 28717 6568 28722 6624
rect 28778 6568 32260 6624
rect 28717 6566 32260 6568
rect 28717 6563 28783 6566
rect 32254 6564 32260 6566
rect 32324 6564 32330 6628
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 20529 6490 20595 6493
rect 22502 6490 22508 6492
rect 20529 6488 22508 6490
rect 20529 6432 20534 6488
rect 20590 6432 22508 6488
rect 20529 6430 22508 6432
rect 20529 6427 20595 6430
rect 22502 6428 22508 6430
rect 22572 6428 22578 6492
rect 25773 6356 25839 6357
rect 25773 6354 25820 6356
rect 25728 6352 25820 6354
rect 25728 6296 25778 6352
rect 25728 6294 25820 6296
rect 25773 6292 25820 6294
rect 25884 6292 25890 6356
rect 25773 6291 25839 6292
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 22093 5812 22159 5813
rect 22093 5810 22140 5812
rect 22048 5808 22140 5810
rect 22204 5810 22210 5812
rect 23381 5810 23447 5813
rect 22204 5808 23447 5810
rect 22048 5752 22098 5808
rect 22204 5752 23386 5808
rect 23442 5752 23447 5808
rect 22048 5750 22140 5752
rect 22093 5748 22140 5750
rect 22204 5750 23447 5752
rect 22204 5748 22210 5750
rect 22093 5747 22159 5748
rect 23381 5747 23447 5750
rect 24669 5810 24735 5813
rect 25446 5810 25452 5812
rect 24669 5808 25452 5810
rect 24669 5752 24674 5808
rect 24730 5752 25452 5808
rect 24669 5750 25452 5752
rect 24669 5747 24735 5750
rect 25446 5748 25452 5750
rect 25516 5748 25522 5812
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 17861 5404 17927 5405
rect 17861 5402 17908 5404
rect 17816 5400 17908 5402
rect 17816 5344 17866 5400
rect 17816 5342 17908 5344
rect 17861 5340 17908 5342
rect 17972 5340 17978 5404
rect 17861 5339 17927 5340
rect 20345 5266 20411 5269
rect 22553 5266 22619 5269
rect 20345 5264 22619 5266
rect 20345 5208 20350 5264
rect 20406 5208 22558 5264
rect 22614 5208 22619 5264
rect 20345 5206 22619 5208
rect 20345 5203 20411 5206
rect 22553 5203 22619 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 17585 4042 17651 4045
rect 19517 4042 19583 4045
rect 17585 4040 19583 4042
rect 17585 3984 17590 4040
rect 17646 3984 19522 4040
rect 19578 3984 19583 4040
rect 17585 3982 19583 3984
rect 17585 3979 17651 3982
rect 19517 3979 19583 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 36077 3498 36143 3501
rect 36895 3498 37695 3528
rect 36077 3496 37695 3498
rect 36077 3440 36082 3496
rect 36138 3440 37695 3496
rect 36077 3438 37695 3440
rect 36077 3435 36143 3438
rect 36895 3408 37695 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 16757 1866 16823 1869
rect 18597 1866 18663 1869
rect 16757 1864 18663 1866
rect 16757 1808 16762 1864
rect 16818 1808 18602 1864
rect 18658 1808 18663 1864
rect 16757 1806 18663 1808
rect 16757 1803 16823 1806
rect 18597 1803 18663 1806
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 8892 35532 8956 35596
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 8340 34640 8404 34644
rect 8340 34584 8354 34640
rect 8354 34584 8404 34640
rect 8340 34580 8404 34584
rect 9996 34308 10060 34372
rect 13676 34308 13740 34372
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 9812 33220 9876 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 24164 31240 24228 31244
rect 24164 31184 24214 31240
rect 24214 31184 24228 31240
rect 24164 31180 24228 31184
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 13492 30908 13556 30972
rect 9996 30636 10060 30700
rect 21956 30636 22020 30700
rect 11836 30500 11900 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 10916 30364 10980 30428
rect 16620 30424 16684 30428
rect 16620 30368 16634 30424
rect 16634 30368 16684 30424
rect 16620 30364 16684 30368
rect 13860 30228 13924 30292
rect 25452 30228 25516 30292
rect 31892 30092 31956 30156
rect 32260 30092 32324 30156
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 32444 29744 32508 29748
rect 32444 29688 32458 29744
rect 32458 29688 32508 29744
rect 32444 29684 32508 29688
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35388 29548 35452 29612
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 30420 29276 30484 29340
rect 5764 29004 5828 29068
rect 12204 29004 12268 29068
rect 12572 29064 12636 29068
rect 12572 29008 12586 29064
rect 12586 29008 12636 29064
rect 12572 29004 12636 29008
rect 7604 28868 7668 28932
rect 31524 29064 31588 29068
rect 31524 29008 31574 29064
rect 31574 29008 31588 29064
rect 31524 29004 31588 29008
rect 32444 29064 32508 29068
rect 32444 29008 32458 29064
rect 32458 29008 32508 29064
rect 32444 29004 32508 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 10364 28596 10428 28660
rect 23428 28460 23492 28524
rect 17172 28384 17236 28388
rect 17172 28328 17222 28384
rect 17222 28328 17236 28384
rect 17172 28324 17236 28328
rect 23244 28324 23308 28388
rect 32076 28324 32140 28388
rect 33364 28324 33428 28388
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 8524 28188 8588 28252
rect 26556 28188 26620 28252
rect 26188 28052 26252 28116
rect 32076 28052 32140 28116
rect 17356 27916 17420 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 13676 27432 13740 27436
rect 13676 27376 13690 27432
rect 13690 27376 13740 27432
rect 13676 27372 13740 27376
rect 30420 27372 30484 27436
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 13492 26828 13556 26892
rect 18092 26752 18156 26756
rect 18092 26696 18142 26752
rect 18142 26696 18156 26752
rect 18092 26692 18156 26696
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19012 26420 19076 26484
rect 24532 26284 24596 26348
rect 24900 26284 24964 26348
rect 20116 26148 20180 26212
rect 28948 26148 29012 26212
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 20116 25876 20180 25940
rect 31524 25876 31588 25940
rect 32260 25876 32324 25940
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 8524 25528 8588 25532
rect 8524 25472 8538 25528
rect 8538 25472 8588 25528
rect 8524 25468 8588 25472
rect 16620 25528 16684 25532
rect 16620 25472 16634 25528
rect 16634 25472 16684 25528
rect 16620 25468 16684 25472
rect 35388 25468 35452 25532
rect 16068 25196 16132 25260
rect 23060 25060 23124 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 14780 24924 14844 24988
rect 29316 24984 29380 24988
rect 29316 24928 29330 24984
rect 29330 24928 29380 24984
rect 29316 24924 29380 24928
rect 8340 24848 8404 24852
rect 8340 24792 8390 24848
rect 8390 24792 8404 24848
rect 8340 24788 8404 24792
rect 12572 24788 12636 24852
rect 31340 24848 31404 24852
rect 31340 24792 31354 24848
rect 31354 24792 31404 24848
rect 31340 24788 31404 24792
rect 31524 24788 31588 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 32076 24380 32140 24444
rect 10180 24304 10244 24308
rect 10180 24248 10194 24304
rect 10194 24248 10244 24304
rect 10180 24244 10244 24248
rect 28764 24244 28828 24308
rect 6316 24108 6380 24172
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 17172 23836 17236 23900
rect 28948 23836 29012 23900
rect 5948 23760 6012 23764
rect 5948 23704 5998 23760
rect 5998 23704 6012 23760
rect 5948 23700 6012 23704
rect 13676 23700 13740 23764
rect 14044 23624 14108 23628
rect 14044 23568 14094 23624
rect 14094 23568 14108 23624
rect 14044 23564 14108 23568
rect 15332 23564 15396 23628
rect 22140 23564 22204 23628
rect 27844 23564 27908 23628
rect 14964 23428 15028 23492
rect 16804 23488 16868 23492
rect 16804 23432 16818 23488
rect 16818 23432 16868 23488
rect 16804 23428 16868 23432
rect 28764 23428 28828 23492
rect 29132 23428 29196 23492
rect 34100 23488 34164 23492
rect 34100 23432 34114 23488
rect 34114 23432 34164 23488
rect 34100 23428 34164 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 9812 23292 9876 23356
rect 16436 23292 16500 23356
rect 18092 23292 18156 23356
rect 31340 23292 31404 23356
rect 13308 23020 13372 23084
rect 23428 23020 23492 23084
rect 26372 23020 26436 23084
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 16620 22748 16684 22812
rect 7420 22612 7484 22676
rect 29500 22612 29564 22676
rect 32444 22612 32508 22676
rect 21588 22476 21652 22540
rect 22876 22476 22940 22540
rect 33732 22476 33796 22540
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 17540 22204 17604 22268
rect 19380 21992 19444 21996
rect 19380 21936 19430 21992
rect 19430 21936 19444 21992
rect 19380 21932 19444 21936
rect 24348 21932 24412 21996
rect 23060 21796 23124 21860
rect 24716 21796 24780 21860
rect 26188 21796 26252 21860
rect 29868 21796 29932 21860
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 16068 21524 16132 21588
rect 24532 21388 24596 21452
rect 28580 21448 28644 21452
rect 28580 21392 28630 21448
rect 28630 21392 28644 21448
rect 28580 21388 28644 21392
rect 24532 21312 24596 21316
rect 24532 21256 24546 21312
rect 24546 21256 24596 21312
rect 24532 21252 24596 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19564 21040 19628 21044
rect 19564 20984 19614 21040
rect 19614 20984 19628 21040
rect 19564 20980 19628 20984
rect 4660 20844 4724 20908
rect 31892 20980 31956 21044
rect 24164 20708 24228 20772
rect 31524 20708 31588 20772
rect 31892 20844 31956 20908
rect 34652 20768 34716 20772
rect 34652 20712 34702 20768
rect 34702 20712 34716 20768
rect 34652 20708 34716 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 5764 20632 5828 20636
rect 5764 20576 5778 20632
rect 5778 20576 5828 20632
rect 5764 20572 5828 20576
rect 7604 20572 7668 20636
rect 17724 20572 17788 20636
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 18644 20572 18708 20636
rect 26556 20632 26620 20636
rect 26556 20576 26606 20632
rect 26606 20576 26620 20632
rect 26556 20572 26620 20576
rect 8892 20436 8956 20500
rect 19380 20436 19444 20500
rect 37044 20436 37108 20500
rect 11836 20300 11900 20364
rect 19564 20300 19628 20364
rect 20484 20300 20548 20364
rect 20852 20300 20916 20364
rect 20116 20224 20180 20228
rect 20116 20168 20130 20224
rect 20130 20168 20180 20224
rect 20116 20164 20180 20168
rect 31892 20224 31956 20228
rect 31892 20168 31906 20224
rect 31906 20168 31956 20224
rect 31892 20164 31956 20168
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 10180 20028 10244 20092
rect 18276 20028 18340 20092
rect 25452 19952 25516 19956
rect 25452 19896 25466 19952
rect 25466 19896 25516 19952
rect 25452 19892 25516 19896
rect 37044 19892 37108 19956
rect 27108 19756 27172 19820
rect 33364 19756 33428 19820
rect 23244 19620 23308 19684
rect 25636 19620 25700 19684
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 16252 19348 16316 19412
rect 17540 19348 17604 19412
rect 28212 19348 28276 19412
rect 30420 19348 30484 19412
rect 32260 19348 32324 19412
rect 12204 19272 12268 19276
rect 12204 19216 12254 19272
rect 12254 19216 12268 19272
rect 12204 19212 12268 19216
rect 15332 19212 15396 19276
rect 26004 19212 26068 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 28764 18864 28828 18868
rect 28764 18808 28778 18864
rect 28778 18808 28828 18864
rect 28764 18804 28828 18808
rect 11284 18668 11348 18732
rect 11468 18728 11532 18732
rect 11468 18672 11518 18728
rect 11518 18672 11532 18728
rect 11468 18668 11532 18672
rect 20668 18668 20732 18732
rect 21772 18532 21836 18596
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 10916 18456 10980 18460
rect 10916 18400 10966 18456
rect 10966 18400 10980 18456
rect 10916 18396 10980 18400
rect 14044 18260 14108 18324
rect 26188 18260 26252 18324
rect 21588 18184 21652 18188
rect 21588 18128 21638 18184
rect 21638 18128 21652 18184
rect 21588 18124 21652 18128
rect 10364 17988 10428 18052
rect 13124 17988 13188 18052
rect 15148 17988 15212 18052
rect 23060 17988 23124 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 13860 17852 13924 17916
rect 14780 17852 14844 17916
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19012 17716 19076 17780
rect 14964 17580 15028 17644
rect 19380 17444 19444 17508
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 16620 17308 16684 17372
rect 16436 17172 16500 17236
rect 17908 17172 17972 17236
rect 21772 17036 21836 17100
rect 24716 17036 24780 17100
rect 25820 17036 25884 17100
rect 16804 16900 16868 16964
rect 19748 16900 19812 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 17540 16824 17604 16828
rect 17540 16768 17590 16824
rect 17590 16768 17604 16824
rect 17540 16764 17604 16768
rect 18092 16824 18156 16828
rect 18092 16768 18142 16824
rect 18142 16768 18156 16824
rect 18092 16764 18156 16768
rect 22508 16764 22572 16828
rect 7420 16628 7484 16692
rect 25452 16628 25516 16692
rect 13492 16492 13556 16556
rect 14044 16492 14108 16556
rect 23428 16492 23492 16556
rect 28764 16492 28828 16556
rect 26924 16356 26988 16420
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 28396 16084 28460 16148
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 18276 15540 18340 15604
rect 19012 15600 19076 15604
rect 19012 15544 19026 15600
rect 19026 15544 19076 15600
rect 19012 15540 19076 15544
rect 21404 15540 21468 15604
rect 21956 15540 22020 15604
rect 20484 15404 20548 15468
rect 33732 15404 33796 15468
rect 27292 15268 27356 15332
rect 27844 15268 27908 15332
rect 31156 15268 31220 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 24900 15132 24964 15196
rect 26372 15192 26436 15196
rect 26372 15136 26386 15192
rect 26386 15136 26436 15192
rect 26372 15132 26436 15136
rect 29316 15192 29380 15196
rect 29316 15136 29330 15192
rect 29330 15136 29380 15192
rect 29316 15132 29380 15136
rect 18276 15056 18340 15060
rect 18276 15000 18290 15056
rect 18290 15000 18340 15056
rect 18276 14996 18340 15000
rect 19196 14996 19260 15060
rect 19564 14996 19628 15060
rect 28580 14996 28644 15060
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 13308 14452 13372 14516
rect 20300 14512 20364 14516
rect 20300 14456 20314 14512
rect 20314 14456 20364 14512
rect 20300 14452 20364 14456
rect 21220 14316 21284 14380
rect 26372 14316 26436 14380
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 26924 14104 26988 14108
rect 26924 14048 26974 14104
rect 26974 14048 26988 14104
rect 26924 14044 26988 14048
rect 4660 13908 4724 13972
rect 26188 13908 26252 13972
rect 19564 13636 19628 13700
rect 20484 13636 20548 13700
rect 24532 13636 24596 13700
rect 26740 13636 26804 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 18460 13364 18524 13428
rect 23980 13500 24044 13564
rect 25636 13500 25700 13564
rect 19564 13288 19628 13292
rect 19564 13232 19578 13288
rect 19578 13232 19628 13288
rect 19564 13228 19628 13232
rect 23244 13092 23308 13156
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 10180 12880 10244 12884
rect 10180 12824 10194 12880
rect 10194 12824 10244 12880
rect 10180 12820 10244 12824
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 20668 12820 20732 12884
rect 27844 12820 27908 12884
rect 18092 12684 18156 12748
rect 28028 12684 28092 12748
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 32076 12412 32140 12476
rect 27108 12276 27172 12340
rect 31892 12276 31956 12340
rect 17540 12004 17604 12068
rect 22324 12004 22388 12068
rect 34652 12004 34716 12068
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 19012 11928 19076 11932
rect 19012 11872 19062 11928
rect 19062 11872 19076 11928
rect 19012 11868 19076 11872
rect 16252 11732 16316 11796
rect 20116 11596 20180 11660
rect 27292 11596 27356 11660
rect 18276 11520 18340 11524
rect 18276 11464 18326 11520
rect 18326 11464 18340 11520
rect 18276 11460 18340 11464
rect 19196 11520 19260 11524
rect 19196 11464 19246 11520
rect 19246 11464 19260 11520
rect 19196 11460 19260 11464
rect 20300 11520 20364 11524
rect 20300 11464 20350 11520
rect 20350 11464 20364 11520
rect 20300 11460 20364 11464
rect 21220 11520 21284 11524
rect 21220 11464 21270 11520
rect 21270 11464 21284 11520
rect 21220 11460 21284 11464
rect 21956 11460 22020 11524
rect 22508 11460 22572 11524
rect 23244 11460 23308 11524
rect 33364 11792 33428 11796
rect 33364 11736 33378 11792
rect 33378 11736 33428 11792
rect 33364 11732 33428 11736
rect 29132 11656 29196 11660
rect 29132 11600 29182 11656
rect 29182 11600 29196 11656
rect 29132 11596 29196 11600
rect 29500 11656 29564 11660
rect 29500 11600 29550 11656
rect 29550 11600 29564 11656
rect 29500 11596 29564 11600
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 13124 11188 13188 11252
rect 16620 11188 16684 11252
rect 19748 11188 19812 11252
rect 21588 11188 21652 11252
rect 23060 11324 23124 11388
rect 28212 11384 28276 11388
rect 28212 11328 28226 11384
rect 28226 11328 28276 11384
rect 28212 11324 28276 11328
rect 20852 11052 20916 11116
rect 34100 11052 34164 11116
rect 30420 10916 30484 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 23980 10780 24044 10844
rect 24348 10780 24412 10844
rect 19564 10508 19628 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 17724 10296 17788 10300
rect 17724 10240 17738 10296
rect 17738 10240 17788 10296
rect 17724 10236 17788 10240
rect 28028 10236 28092 10300
rect 5948 10160 6012 10164
rect 5948 10104 5962 10160
rect 5962 10104 6012 10160
rect 5948 10100 6012 10104
rect 21956 10100 22020 10164
rect 26372 10160 26436 10164
rect 26372 10104 26422 10160
rect 26422 10104 26436 10160
rect 26372 10100 26436 10104
rect 27844 10024 27908 10028
rect 27844 9968 27894 10024
rect 27894 9968 27908 10024
rect 27844 9964 27908 9968
rect 28764 9964 28828 10028
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 14780 9556 14844 9620
rect 6316 9420 6380 9484
rect 22324 9556 22388 9620
rect 26740 9556 26804 9620
rect 23428 9420 23492 9484
rect 26188 9420 26252 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 15148 9208 15212 9212
rect 15148 9152 15198 9208
rect 15198 9152 15212 9208
rect 15148 9148 15212 9152
rect 18644 9208 18708 9212
rect 18644 9152 18658 9208
rect 18658 9152 18708 9208
rect 18644 9148 18708 9152
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 28396 9148 28460 9212
rect 26188 9012 26252 9076
rect 21404 8740 21468 8804
rect 31524 8740 31588 8804
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 22876 8604 22940 8668
rect 14964 8468 15028 8532
rect 19380 8528 19444 8532
rect 19380 8472 19394 8528
rect 19394 8472 19444 8528
rect 19380 8468 19444 8472
rect 19564 8392 19628 8396
rect 19564 8336 19578 8392
rect 19578 8336 19628 8392
rect 19564 8332 19628 8336
rect 20484 8332 20548 8396
rect 21220 8256 21284 8260
rect 21220 8200 21234 8256
rect 21234 8200 21284 8256
rect 21220 8196 21284 8200
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 11284 8120 11348 8124
rect 11284 8064 11298 8120
rect 11298 8064 11348 8120
rect 11284 8060 11348 8064
rect 13492 8120 13556 8124
rect 13492 8064 13506 8120
rect 13506 8064 13556 8120
rect 13492 8060 13556 8064
rect 21956 8256 22020 8260
rect 21956 8200 22006 8256
rect 22006 8200 22020 8256
rect 21956 8196 22020 8200
rect 28580 8332 28644 8396
rect 29500 8256 29564 8260
rect 29500 8200 29514 8256
rect 29514 8200 29564 8256
rect 29500 8196 29564 8200
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 11468 7924 11532 7988
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 28764 7516 28828 7580
rect 17356 7440 17420 7444
rect 17356 7384 17370 7440
rect 17370 7384 17420 7440
rect 17356 7380 17420 7384
rect 19380 7440 19444 7444
rect 19380 7384 19394 7440
rect 19394 7384 19444 7440
rect 19380 7380 19444 7384
rect 32444 7244 32508 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 21588 7032 21652 7036
rect 21588 6976 21638 7032
rect 21638 6976 21652 7032
rect 21588 6972 21652 6976
rect 29868 6972 29932 7036
rect 13676 6836 13740 6900
rect 31156 6836 31220 6900
rect 32260 6564 32324 6628
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 22508 6428 22572 6492
rect 25820 6352 25884 6356
rect 25820 6296 25834 6352
rect 25834 6296 25884 6352
rect 25820 6292 25884 6296
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 22140 5808 22204 5812
rect 22140 5752 22154 5808
rect 22154 5752 22204 5808
rect 22140 5748 22204 5752
rect 25452 5748 25516 5812
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 17908 5400 17972 5404
rect 17908 5344 17922 5400
rect 17922 5344 17972 5400
rect 17908 5340 17972 5344
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 8891 35596 8957 35597
rect 8891 35532 8892 35596
rect 8956 35532 8957 35596
rect 8891 35531 8957 35532
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 8339 34644 8405 34645
rect 8339 34580 8340 34644
rect 8404 34580 8405 34644
rect 8339 34579 8405 34580
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 5763 29068 5829 29069
rect 5763 29004 5764 29068
rect 5828 29004 5829 29068
rect 5763 29003 5829 29004
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4659 20908 4725 20909
rect 4659 20844 4660 20908
rect 4724 20844 4725 20908
rect 4659 20843 4725 20844
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4662 13973 4722 20843
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 5766 20637 5826 29003
rect 7603 28932 7669 28933
rect 7603 28868 7604 28932
rect 7668 28868 7669 28932
rect 7603 28867 7669 28868
rect 6315 24172 6381 24173
rect 6315 24108 6316 24172
rect 6380 24108 6381 24172
rect 6315 24107 6381 24108
rect 5947 23764 6013 23765
rect 5947 23700 5948 23764
rect 6012 23700 6013 23764
rect 5947 23699 6013 23700
rect 5763 20636 5829 20637
rect 5763 20572 5764 20636
rect 5828 20572 5829 20636
rect 5763 20571 5829 20572
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4659 13972 4725 13973
rect 4659 13908 4660 13972
rect 4724 13908 4725 13972
rect 4659 13907 4725 13908
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 5950 10165 6010 23699
rect 5947 10164 6013 10165
rect 5947 10100 5948 10164
rect 6012 10100 6013 10164
rect 5947 10099 6013 10100
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 6318 9485 6378 24107
rect 7419 22676 7485 22677
rect 7419 22612 7420 22676
rect 7484 22612 7485 22676
rect 7419 22611 7485 22612
rect 7422 16693 7482 22611
rect 7606 20637 7666 28867
rect 8342 24853 8402 34579
rect 8523 28252 8589 28253
rect 8523 28188 8524 28252
rect 8588 28188 8589 28252
rect 8523 28187 8589 28188
rect 8526 25533 8586 28187
rect 8523 25532 8589 25533
rect 8523 25468 8524 25532
rect 8588 25468 8589 25532
rect 8523 25467 8589 25468
rect 8339 24852 8405 24853
rect 8339 24788 8340 24852
rect 8404 24788 8405 24852
rect 8339 24787 8405 24788
rect 7603 20636 7669 20637
rect 7603 20572 7604 20636
rect 7668 20572 7669 20636
rect 7603 20571 7669 20572
rect 8894 20501 8954 35531
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 9995 34372 10061 34373
rect 9995 34308 9996 34372
rect 10060 34308 10061 34372
rect 9995 34307 10061 34308
rect 13675 34372 13741 34373
rect 13675 34308 13676 34372
rect 13740 34308 13741 34372
rect 13675 34307 13741 34308
rect 9811 33284 9877 33285
rect 9811 33220 9812 33284
rect 9876 33220 9877 33284
rect 9811 33219 9877 33220
rect 9814 23357 9874 33219
rect 9998 30701 10058 34307
rect 13491 30972 13557 30973
rect 13491 30908 13492 30972
rect 13556 30908 13557 30972
rect 13491 30907 13557 30908
rect 9995 30700 10061 30701
rect 9995 30636 9996 30700
rect 10060 30636 10061 30700
rect 9995 30635 10061 30636
rect 11835 30564 11901 30565
rect 11835 30500 11836 30564
rect 11900 30500 11901 30564
rect 11835 30499 11901 30500
rect 10915 30428 10981 30429
rect 10915 30364 10916 30428
rect 10980 30364 10981 30428
rect 10915 30363 10981 30364
rect 10363 28660 10429 28661
rect 10363 28596 10364 28660
rect 10428 28596 10429 28660
rect 10363 28595 10429 28596
rect 10179 24308 10245 24309
rect 10179 24244 10180 24308
rect 10244 24244 10245 24308
rect 10179 24243 10245 24244
rect 9811 23356 9877 23357
rect 9811 23292 9812 23356
rect 9876 23292 9877 23356
rect 9811 23291 9877 23292
rect 8891 20500 8957 20501
rect 8891 20436 8892 20500
rect 8956 20436 8957 20500
rect 8891 20435 8957 20436
rect 10182 20093 10242 24243
rect 10179 20092 10245 20093
rect 10179 20028 10180 20092
rect 10244 20028 10245 20092
rect 10179 20027 10245 20028
rect 7419 16692 7485 16693
rect 7419 16628 7420 16692
rect 7484 16628 7485 16692
rect 7419 16627 7485 16628
rect 10182 12885 10242 20027
rect 10366 18053 10426 28595
rect 10918 18461 10978 30363
rect 11838 20365 11898 30499
rect 12203 29068 12269 29069
rect 12203 29004 12204 29068
rect 12268 29004 12269 29068
rect 12203 29003 12269 29004
rect 12571 29068 12637 29069
rect 12571 29004 12572 29068
rect 12636 29004 12637 29068
rect 12571 29003 12637 29004
rect 11835 20364 11901 20365
rect 11835 20300 11836 20364
rect 11900 20300 11901 20364
rect 11835 20299 11901 20300
rect 12206 19277 12266 29003
rect 12574 24853 12634 29003
rect 13494 26893 13554 30907
rect 13678 27437 13738 34307
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 24163 31244 24229 31245
rect 24163 31180 24164 31244
rect 24228 31180 24229 31244
rect 24163 31179 24229 31180
rect 21955 30700 22021 30701
rect 21955 30636 21956 30700
rect 22020 30636 22021 30700
rect 21955 30635 22021 30636
rect 16619 30428 16685 30429
rect 16619 30364 16620 30428
rect 16684 30364 16685 30428
rect 16619 30363 16685 30364
rect 13859 30292 13925 30293
rect 13859 30228 13860 30292
rect 13924 30228 13925 30292
rect 13859 30227 13925 30228
rect 13675 27436 13741 27437
rect 13675 27372 13676 27436
rect 13740 27372 13741 27436
rect 13675 27371 13741 27372
rect 13491 26892 13557 26893
rect 13491 26828 13492 26892
rect 13556 26828 13557 26892
rect 13491 26827 13557 26828
rect 12571 24852 12637 24853
rect 12571 24788 12572 24852
rect 12636 24788 12637 24852
rect 12571 24787 12637 24788
rect 13675 23764 13741 23765
rect 13675 23700 13676 23764
rect 13740 23700 13741 23764
rect 13675 23699 13741 23700
rect 13307 23084 13373 23085
rect 13307 23020 13308 23084
rect 13372 23020 13373 23084
rect 13307 23019 13373 23020
rect 12203 19276 12269 19277
rect 12203 19212 12204 19276
rect 12268 19212 12269 19276
rect 12203 19211 12269 19212
rect 11283 18732 11349 18733
rect 11283 18668 11284 18732
rect 11348 18668 11349 18732
rect 11283 18667 11349 18668
rect 11467 18732 11533 18733
rect 11467 18668 11468 18732
rect 11532 18668 11533 18732
rect 11467 18667 11533 18668
rect 10915 18460 10981 18461
rect 10915 18396 10916 18460
rect 10980 18396 10981 18460
rect 10915 18395 10981 18396
rect 10363 18052 10429 18053
rect 10363 17988 10364 18052
rect 10428 17988 10429 18052
rect 10363 17987 10429 17988
rect 10179 12884 10245 12885
rect 10179 12820 10180 12884
rect 10244 12820 10245 12884
rect 10179 12819 10245 12820
rect 6315 9484 6381 9485
rect 6315 9420 6316 9484
rect 6380 9420 6381 9484
rect 6315 9419 6381 9420
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 11286 8125 11346 18667
rect 11283 8124 11349 8125
rect 11283 8060 11284 8124
rect 11348 8060 11349 8124
rect 11283 8059 11349 8060
rect 11470 7989 11530 18667
rect 13123 18052 13189 18053
rect 13123 17988 13124 18052
rect 13188 17988 13189 18052
rect 13123 17987 13189 17988
rect 13126 11253 13186 17987
rect 13310 14517 13370 23019
rect 13491 16556 13557 16557
rect 13491 16492 13492 16556
rect 13556 16492 13557 16556
rect 13491 16491 13557 16492
rect 13307 14516 13373 14517
rect 13307 14452 13308 14516
rect 13372 14452 13373 14516
rect 13307 14451 13373 14452
rect 13123 11252 13189 11253
rect 13123 11188 13124 11252
rect 13188 11188 13189 11252
rect 13123 11187 13189 11188
rect 13494 8125 13554 16491
rect 13491 8124 13557 8125
rect 13491 8060 13492 8124
rect 13556 8060 13557 8124
rect 13491 8059 13557 8060
rect 11467 7988 11533 7989
rect 11467 7924 11468 7988
rect 11532 7924 11533 7988
rect 11467 7923 11533 7924
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 13678 6901 13738 23699
rect 13862 17917 13922 30227
rect 16622 25533 16682 30363
rect 17171 28388 17237 28389
rect 17171 28324 17172 28388
rect 17236 28324 17237 28388
rect 17171 28323 17237 28324
rect 16619 25532 16685 25533
rect 16619 25468 16620 25532
rect 16684 25468 16685 25532
rect 16619 25467 16685 25468
rect 16067 25260 16133 25261
rect 16067 25196 16068 25260
rect 16132 25196 16133 25260
rect 16067 25195 16133 25196
rect 14779 24988 14845 24989
rect 14779 24924 14780 24988
rect 14844 24924 14845 24988
rect 14779 24923 14845 24924
rect 14043 23628 14109 23629
rect 14043 23564 14044 23628
rect 14108 23564 14109 23628
rect 14043 23563 14109 23564
rect 14046 18325 14106 23563
rect 14043 18324 14109 18325
rect 14043 18260 14044 18324
rect 14108 18260 14109 18324
rect 14043 18259 14109 18260
rect 13859 17916 13925 17917
rect 13859 17852 13860 17916
rect 13924 17852 13925 17916
rect 13859 17851 13925 17852
rect 14046 16557 14106 18259
rect 14782 17917 14842 24923
rect 15331 23628 15397 23629
rect 15331 23564 15332 23628
rect 15396 23564 15397 23628
rect 15331 23563 15397 23564
rect 14963 23492 15029 23493
rect 14963 23428 14964 23492
rect 15028 23428 15029 23492
rect 14963 23427 15029 23428
rect 14779 17916 14845 17917
rect 14779 17852 14780 17916
rect 14844 17852 14845 17916
rect 14779 17851 14845 17852
rect 14043 16556 14109 16557
rect 14043 16492 14044 16556
rect 14108 16492 14109 16556
rect 14043 16491 14109 16492
rect 14782 9621 14842 17851
rect 14966 17645 15026 23427
rect 15334 19277 15394 23563
rect 16070 21589 16130 25195
rect 17174 23901 17234 28323
rect 17355 27980 17421 27981
rect 17355 27916 17356 27980
rect 17420 27916 17421 27980
rect 17355 27915 17421 27916
rect 17171 23900 17237 23901
rect 17171 23836 17172 23900
rect 17236 23836 17237 23900
rect 17171 23835 17237 23836
rect 16803 23492 16869 23493
rect 16803 23428 16804 23492
rect 16868 23428 16869 23492
rect 16803 23427 16869 23428
rect 16435 23356 16501 23357
rect 16435 23292 16436 23356
rect 16500 23292 16501 23356
rect 16435 23291 16501 23292
rect 16067 21588 16133 21589
rect 16067 21524 16068 21588
rect 16132 21524 16133 21588
rect 16067 21523 16133 21524
rect 16251 19412 16317 19413
rect 16251 19348 16252 19412
rect 16316 19348 16317 19412
rect 16251 19347 16317 19348
rect 15331 19276 15397 19277
rect 15331 19212 15332 19276
rect 15396 19212 15397 19276
rect 15331 19211 15397 19212
rect 15147 18052 15213 18053
rect 15147 17988 15148 18052
rect 15212 17988 15213 18052
rect 15147 17987 15213 17988
rect 14963 17644 15029 17645
rect 14963 17580 14964 17644
rect 15028 17580 15029 17644
rect 14963 17579 15029 17580
rect 14779 9620 14845 9621
rect 14779 9556 14780 9620
rect 14844 9556 14845 9620
rect 14779 9555 14845 9556
rect 14966 8533 15026 17579
rect 15150 9213 15210 17987
rect 16254 11797 16314 19347
rect 16438 17237 16498 23291
rect 16619 22812 16685 22813
rect 16619 22748 16620 22812
rect 16684 22748 16685 22812
rect 16619 22747 16685 22748
rect 16622 17373 16682 22747
rect 16619 17372 16685 17373
rect 16619 17308 16620 17372
rect 16684 17308 16685 17372
rect 16619 17307 16685 17308
rect 16435 17236 16501 17237
rect 16435 17172 16436 17236
rect 16500 17172 16501 17236
rect 16435 17171 16501 17172
rect 16251 11796 16317 11797
rect 16251 11732 16252 11796
rect 16316 11732 16317 11796
rect 16251 11731 16317 11732
rect 16622 11253 16682 17307
rect 16806 16965 16866 23427
rect 16803 16964 16869 16965
rect 16803 16900 16804 16964
rect 16868 16900 16869 16964
rect 16803 16899 16869 16900
rect 16619 11252 16685 11253
rect 16619 11188 16620 11252
rect 16684 11188 16685 11252
rect 16619 11187 16685 11188
rect 15147 9212 15213 9213
rect 15147 9148 15148 9212
rect 15212 9148 15213 9212
rect 15147 9147 15213 9148
rect 14963 8532 15029 8533
rect 14963 8468 14964 8532
rect 15028 8468 15029 8532
rect 14963 8467 15029 8468
rect 17358 7445 17418 27915
rect 18091 26756 18157 26757
rect 18091 26692 18092 26756
rect 18156 26692 18157 26756
rect 18091 26691 18157 26692
rect 18094 23357 18154 26691
rect 19011 26484 19077 26485
rect 19011 26420 19012 26484
rect 19076 26420 19077 26484
rect 19011 26419 19077 26420
rect 18091 23356 18157 23357
rect 18091 23292 18092 23356
rect 18156 23292 18157 23356
rect 18091 23291 18157 23292
rect 17539 22268 17605 22269
rect 17539 22204 17540 22268
rect 17604 22204 17605 22268
rect 17539 22203 17605 22204
rect 17542 19413 17602 22203
rect 17723 20636 17789 20637
rect 17723 20572 17724 20636
rect 17788 20572 17789 20636
rect 17723 20571 17789 20572
rect 18643 20636 18709 20637
rect 18643 20572 18644 20636
rect 18708 20572 18709 20636
rect 18643 20571 18709 20572
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 17539 16828 17605 16829
rect 17539 16764 17540 16828
rect 17604 16764 17605 16828
rect 17539 16763 17605 16764
rect 17542 12069 17602 16763
rect 17539 12068 17605 12069
rect 17539 12004 17540 12068
rect 17604 12004 17605 12068
rect 17539 12003 17605 12004
rect 17726 10301 17786 20571
rect 18275 20092 18341 20093
rect 18275 20028 18276 20092
rect 18340 20028 18341 20092
rect 18275 20027 18341 20028
rect 17907 17236 17973 17237
rect 17907 17172 17908 17236
rect 17972 17172 17973 17236
rect 17907 17171 17973 17172
rect 17723 10300 17789 10301
rect 17723 10236 17724 10300
rect 17788 10236 17789 10300
rect 17723 10235 17789 10236
rect 17355 7444 17421 7445
rect 17355 7380 17356 7444
rect 17420 7380 17421 7444
rect 17355 7379 17421 7380
rect 13675 6900 13741 6901
rect 13675 6836 13676 6900
rect 13740 6836 13741 6900
rect 13675 6835 13741 6836
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 17910 5405 17970 17171
rect 18091 16828 18157 16829
rect 18091 16764 18092 16828
rect 18156 16764 18157 16828
rect 18091 16763 18157 16764
rect 18094 12749 18154 16763
rect 18278 15605 18338 20027
rect 18275 15604 18341 15605
rect 18275 15540 18276 15604
rect 18340 15602 18341 15604
rect 18340 15542 18522 15602
rect 18340 15540 18341 15542
rect 18275 15539 18341 15540
rect 18275 15060 18341 15061
rect 18275 14996 18276 15060
rect 18340 14996 18341 15060
rect 18275 14995 18341 14996
rect 18091 12748 18157 12749
rect 18091 12684 18092 12748
rect 18156 12684 18157 12748
rect 18091 12683 18157 12684
rect 18278 11525 18338 14995
rect 18462 13429 18522 15542
rect 18459 13428 18525 13429
rect 18459 13364 18460 13428
rect 18524 13364 18525 13428
rect 18459 13363 18525 13364
rect 18275 11524 18341 11525
rect 18275 11460 18276 11524
rect 18340 11460 18341 11524
rect 18275 11459 18341 11460
rect 18646 9213 18706 20571
rect 19014 17781 19074 26419
rect 20115 26212 20181 26213
rect 20115 26148 20116 26212
rect 20180 26148 20181 26212
rect 20115 26147 20181 26148
rect 20118 25941 20178 26147
rect 20115 25940 20181 25941
rect 20115 25876 20116 25940
rect 20180 25876 20181 25940
rect 20115 25875 20181 25876
rect 19379 21996 19445 21997
rect 19379 21932 19380 21996
rect 19444 21932 19445 21996
rect 19379 21931 19445 21932
rect 19382 20501 19442 21931
rect 19563 21044 19629 21045
rect 19563 20980 19564 21044
rect 19628 20980 19629 21044
rect 19563 20979 19629 20980
rect 19379 20500 19445 20501
rect 19379 20436 19380 20500
rect 19444 20436 19445 20500
rect 19379 20435 19445 20436
rect 19011 17780 19077 17781
rect 19011 17716 19012 17780
rect 19076 17716 19077 17780
rect 19011 17715 19077 17716
rect 19382 17509 19442 20435
rect 19566 20365 19626 20979
rect 19563 20364 19629 20365
rect 19563 20300 19564 20364
rect 19628 20300 19629 20364
rect 19563 20299 19629 20300
rect 20118 20229 20178 25875
rect 21587 22540 21653 22541
rect 21587 22476 21588 22540
rect 21652 22476 21653 22540
rect 21587 22475 21653 22476
rect 20483 20364 20549 20365
rect 20483 20300 20484 20364
rect 20548 20300 20549 20364
rect 20483 20299 20549 20300
rect 20851 20364 20917 20365
rect 20851 20300 20852 20364
rect 20916 20300 20917 20364
rect 20851 20299 20917 20300
rect 20115 20228 20181 20229
rect 20115 20164 20116 20228
rect 20180 20164 20181 20228
rect 20115 20163 20181 20164
rect 19379 17508 19445 17509
rect 19379 17444 19380 17508
rect 19444 17444 19445 17508
rect 19379 17443 19445 17444
rect 19747 16964 19813 16965
rect 19747 16900 19748 16964
rect 19812 16900 19813 16964
rect 19747 16899 19813 16900
rect 19011 15604 19077 15605
rect 19011 15540 19012 15604
rect 19076 15540 19077 15604
rect 19011 15539 19077 15540
rect 19014 11933 19074 15539
rect 19195 15060 19261 15061
rect 19195 14996 19196 15060
rect 19260 14996 19261 15060
rect 19195 14995 19261 14996
rect 19563 15060 19629 15061
rect 19563 14996 19564 15060
rect 19628 14996 19629 15060
rect 19563 14995 19629 14996
rect 19011 11932 19077 11933
rect 19011 11868 19012 11932
rect 19076 11868 19077 11932
rect 19011 11867 19077 11868
rect 19198 11525 19258 14995
rect 19566 13701 19626 14995
rect 19563 13700 19629 13701
rect 19563 13636 19564 13700
rect 19628 13636 19629 13700
rect 19563 13635 19629 13636
rect 19563 13292 19629 13293
rect 19563 13228 19564 13292
rect 19628 13228 19629 13292
rect 19563 13227 19629 13228
rect 19195 11524 19261 11525
rect 19195 11460 19196 11524
rect 19260 11460 19261 11524
rect 19195 11459 19261 11460
rect 19566 10573 19626 13227
rect 19750 11253 19810 16899
rect 20118 11661 20178 20163
rect 20486 15469 20546 20299
rect 20667 18732 20733 18733
rect 20667 18668 20668 18732
rect 20732 18668 20733 18732
rect 20667 18667 20733 18668
rect 20483 15468 20549 15469
rect 20483 15404 20484 15468
rect 20548 15404 20549 15468
rect 20483 15403 20549 15404
rect 20299 14516 20365 14517
rect 20299 14452 20300 14516
rect 20364 14452 20365 14516
rect 20299 14451 20365 14452
rect 20115 11660 20181 11661
rect 20115 11596 20116 11660
rect 20180 11596 20181 11660
rect 20115 11595 20181 11596
rect 20302 11525 20362 14451
rect 20486 13701 20546 15403
rect 20483 13700 20549 13701
rect 20483 13636 20484 13700
rect 20548 13636 20549 13700
rect 20483 13635 20549 13636
rect 20299 11524 20365 11525
rect 20299 11460 20300 11524
rect 20364 11460 20365 11524
rect 20299 11459 20365 11460
rect 19747 11252 19813 11253
rect 19747 11188 19748 11252
rect 19812 11188 19813 11252
rect 19747 11187 19813 11188
rect 19563 10572 19629 10573
rect 19563 10508 19564 10572
rect 19628 10508 19629 10572
rect 19563 10507 19629 10508
rect 18643 9212 18709 9213
rect 18643 9148 18644 9212
rect 18708 9148 18709 9212
rect 18643 9147 18709 9148
rect 19379 8532 19445 8533
rect 19379 8468 19380 8532
rect 19444 8468 19445 8532
rect 19379 8467 19445 8468
rect 19382 7445 19442 8467
rect 19566 8397 19626 10507
rect 20486 8397 20546 13635
rect 20670 12885 20730 18667
rect 20667 12884 20733 12885
rect 20667 12820 20668 12884
rect 20732 12820 20733 12884
rect 20667 12819 20733 12820
rect 20854 11117 20914 20299
rect 21590 18189 21650 22475
rect 21771 18596 21837 18597
rect 21771 18532 21772 18596
rect 21836 18532 21837 18596
rect 21771 18531 21837 18532
rect 21587 18188 21653 18189
rect 21587 18124 21588 18188
rect 21652 18124 21653 18188
rect 21587 18123 21653 18124
rect 21774 17101 21834 18531
rect 21771 17100 21837 17101
rect 21771 17036 21772 17100
rect 21836 17036 21837 17100
rect 21771 17035 21837 17036
rect 21958 15605 22018 30635
rect 23427 28524 23493 28525
rect 23427 28460 23428 28524
rect 23492 28460 23493 28524
rect 23427 28459 23493 28460
rect 23243 28388 23309 28389
rect 23243 28324 23244 28388
rect 23308 28324 23309 28388
rect 23243 28323 23309 28324
rect 23059 25124 23125 25125
rect 23059 25060 23060 25124
rect 23124 25060 23125 25124
rect 23059 25059 23125 25060
rect 22139 23628 22205 23629
rect 22139 23564 22140 23628
rect 22204 23564 22205 23628
rect 22139 23563 22205 23564
rect 21403 15604 21469 15605
rect 21403 15540 21404 15604
rect 21468 15540 21469 15604
rect 21403 15539 21469 15540
rect 21955 15604 22021 15605
rect 21955 15540 21956 15604
rect 22020 15540 22021 15604
rect 21955 15539 22021 15540
rect 21219 14380 21285 14381
rect 21219 14316 21220 14380
rect 21284 14316 21285 14380
rect 21219 14315 21285 14316
rect 21222 11525 21282 14315
rect 21219 11524 21285 11525
rect 21219 11460 21220 11524
rect 21284 11460 21285 11524
rect 21219 11459 21285 11460
rect 20851 11116 20917 11117
rect 20851 11052 20852 11116
rect 20916 11052 20917 11116
rect 20851 11051 20917 11052
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 20483 8396 20549 8397
rect 20483 8332 20484 8396
rect 20548 8332 20549 8396
rect 20483 8331 20549 8332
rect 21222 8261 21282 11459
rect 21406 8805 21466 15539
rect 21958 11525 22018 15539
rect 21955 11524 22021 11525
rect 21955 11460 21956 11524
rect 22020 11460 22021 11524
rect 21955 11459 22021 11460
rect 21587 11252 21653 11253
rect 21587 11188 21588 11252
rect 21652 11188 21653 11252
rect 21587 11187 21653 11188
rect 21403 8804 21469 8805
rect 21403 8740 21404 8804
rect 21468 8740 21469 8804
rect 21403 8739 21469 8740
rect 21219 8260 21285 8261
rect 21219 8196 21220 8260
rect 21284 8196 21285 8260
rect 21219 8195 21285 8196
rect 19379 7444 19445 7445
rect 19379 7380 19380 7444
rect 19444 7380 19445 7444
rect 19379 7379 19445 7380
rect 21590 7037 21650 11187
rect 21955 10164 22021 10165
rect 21955 10100 21956 10164
rect 22020 10100 22021 10164
rect 21955 10099 22021 10100
rect 21958 8261 22018 10099
rect 21955 8260 22021 8261
rect 21955 8196 21956 8260
rect 22020 8196 22021 8260
rect 21955 8195 22021 8196
rect 21587 7036 21653 7037
rect 21587 6972 21588 7036
rect 21652 6972 21653 7036
rect 21587 6971 21653 6972
rect 22142 5813 22202 23563
rect 22875 22540 22941 22541
rect 22875 22476 22876 22540
rect 22940 22476 22941 22540
rect 22875 22475 22941 22476
rect 22507 16828 22573 16829
rect 22507 16764 22508 16828
rect 22572 16764 22573 16828
rect 22507 16763 22573 16764
rect 22510 12450 22570 16763
rect 22326 12390 22570 12450
rect 22326 12069 22386 12390
rect 22323 12068 22389 12069
rect 22323 12004 22324 12068
rect 22388 12004 22389 12068
rect 22323 12003 22389 12004
rect 22326 9621 22386 12003
rect 22507 11524 22573 11525
rect 22507 11460 22508 11524
rect 22572 11460 22573 11524
rect 22507 11459 22573 11460
rect 22323 9620 22389 9621
rect 22323 9556 22324 9620
rect 22388 9556 22389 9620
rect 22323 9555 22389 9556
rect 22510 6493 22570 11459
rect 22878 8669 22938 22475
rect 23062 21861 23122 25059
rect 23059 21860 23125 21861
rect 23059 21796 23060 21860
rect 23124 21796 23125 21860
rect 23059 21795 23125 21796
rect 23246 19685 23306 28323
rect 23430 23085 23490 28459
rect 23427 23084 23493 23085
rect 23427 23020 23428 23084
rect 23492 23020 23493 23084
rect 23427 23019 23493 23020
rect 24166 20773 24226 31179
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 25451 30292 25517 30293
rect 25451 30228 25452 30292
rect 25516 30228 25517 30292
rect 25451 30227 25517 30228
rect 24531 26348 24597 26349
rect 24531 26284 24532 26348
rect 24596 26284 24597 26348
rect 24531 26283 24597 26284
rect 24899 26348 24965 26349
rect 24899 26284 24900 26348
rect 24964 26284 24965 26348
rect 24899 26283 24965 26284
rect 24347 21996 24413 21997
rect 24347 21932 24348 21996
rect 24412 21932 24413 21996
rect 24347 21931 24413 21932
rect 24163 20772 24229 20773
rect 24163 20708 24164 20772
rect 24228 20708 24229 20772
rect 24163 20707 24229 20708
rect 23243 19684 23309 19685
rect 23243 19620 23244 19684
rect 23308 19620 23309 19684
rect 23243 19619 23309 19620
rect 23059 18052 23125 18053
rect 23059 17988 23060 18052
rect 23124 17988 23125 18052
rect 23059 17987 23125 17988
rect 23062 11389 23122 17987
rect 23427 16556 23493 16557
rect 23427 16492 23428 16556
rect 23492 16492 23493 16556
rect 23427 16491 23493 16492
rect 23243 13156 23309 13157
rect 23243 13092 23244 13156
rect 23308 13092 23309 13156
rect 23243 13091 23309 13092
rect 23246 11525 23306 13091
rect 23243 11524 23309 11525
rect 23243 11460 23244 11524
rect 23308 11460 23309 11524
rect 23243 11459 23309 11460
rect 23059 11388 23125 11389
rect 23059 11324 23060 11388
rect 23124 11324 23125 11388
rect 23059 11323 23125 11324
rect 23430 9485 23490 16491
rect 23979 13564 24045 13565
rect 23979 13500 23980 13564
rect 24044 13500 24045 13564
rect 23979 13499 24045 13500
rect 23982 10845 24042 13499
rect 24350 10845 24410 21931
rect 24534 21453 24594 26283
rect 24715 21860 24781 21861
rect 24715 21796 24716 21860
rect 24780 21796 24781 21860
rect 24715 21795 24781 21796
rect 24531 21452 24597 21453
rect 24531 21388 24532 21452
rect 24596 21388 24597 21452
rect 24531 21387 24597 21388
rect 24531 21316 24597 21317
rect 24531 21252 24532 21316
rect 24596 21252 24597 21316
rect 24531 21251 24597 21252
rect 24534 13701 24594 21251
rect 24718 17101 24778 21795
rect 24715 17100 24781 17101
rect 24715 17036 24716 17100
rect 24780 17036 24781 17100
rect 24715 17035 24781 17036
rect 24902 15197 24962 26283
rect 25454 19957 25514 30227
rect 31891 30156 31957 30157
rect 31891 30092 31892 30156
rect 31956 30092 31957 30156
rect 31891 30091 31957 30092
rect 32259 30156 32325 30157
rect 32259 30092 32260 30156
rect 32324 30092 32325 30156
rect 32259 30091 32325 30092
rect 30419 29340 30485 29341
rect 30419 29276 30420 29340
rect 30484 29276 30485 29340
rect 30419 29275 30485 29276
rect 26555 28252 26621 28253
rect 26555 28188 26556 28252
rect 26620 28188 26621 28252
rect 26555 28187 26621 28188
rect 26187 28116 26253 28117
rect 26187 28052 26188 28116
rect 26252 28052 26253 28116
rect 26187 28051 26253 28052
rect 26190 22110 26250 28051
rect 26371 23084 26437 23085
rect 26371 23020 26372 23084
rect 26436 23020 26437 23084
rect 26371 23019 26437 23020
rect 26006 22050 26250 22110
rect 25451 19956 25517 19957
rect 25451 19892 25452 19956
rect 25516 19892 25517 19956
rect 25451 19891 25517 19892
rect 25635 19684 25701 19685
rect 25635 19620 25636 19684
rect 25700 19620 25701 19684
rect 25635 19619 25701 19620
rect 25451 16692 25517 16693
rect 25451 16628 25452 16692
rect 25516 16628 25517 16692
rect 25451 16627 25517 16628
rect 24899 15196 24965 15197
rect 24899 15132 24900 15196
rect 24964 15132 24965 15196
rect 24899 15131 24965 15132
rect 24531 13700 24597 13701
rect 24531 13636 24532 13700
rect 24596 13636 24597 13700
rect 24531 13635 24597 13636
rect 23979 10844 24045 10845
rect 23979 10780 23980 10844
rect 24044 10780 24045 10844
rect 23979 10779 24045 10780
rect 24347 10844 24413 10845
rect 24347 10780 24348 10844
rect 24412 10780 24413 10844
rect 24347 10779 24413 10780
rect 23427 9484 23493 9485
rect 23427 9420 23428 9484
rect 23492 9420 23493 9484
rect 23427 9419 23493 9420
rect 22875 8668 22941 8669
rect 22875 8604 22876 8668
rect 22940 8604 22941 8668
rect 22875 8603 22941 8604
rect 22507 6492 22573 6493
rect 22507 6428 22508 6492
rect 22572 6428 22573 6492
rect 22507 6427 22573 6428
rect 25454 5813 25514 16627
rect 25638 13565 25698 19619
rect 26006 19277 26066 22050
rect 26187 21860 26253 21861
rect 26187 21796 26188 21860
rect 26252 21796 26253 21860
rect 26187 21795 26253 21796
rect 26003 19276 26069 19277
rect 26003 19212 26004 19276
rect 26068 19212 26069 19276
rect 26003 19211 26069 19212
rect 26190 18325 26250 21795
rect 26187 18324 26253 18325
rect 26187 18260 26188 18324
rect 26252 18260 26253 18324
rect 26187 18259 26253 18260
rect 25819 17100 25885 17101
rect 25819 17036 25820 17100
rect 25884 17036 25885 17100
rect 25819 17035 25885 17036
rect 25635 13564 25701 13565
rect 25635 13500 25636 13564
rect 25700 13500 25701 13564
rect 25635 13499 25701 13500
rect 25822 6357 25882 17035
rect 26190 13973 26250 18259
rect 26374 15197 26434 23019
rect 26558 20637 26618 28187
rect 30422 27437 30482 29275
rect 31523 29068 31589 29069
rect 31523 29004 31524 29068
rect 31588 29004 31589 29068
rect 31523 29003 31589 29004
rect 30419 27436 30485 27437
rect 30419 27372 30420 27436
rect 30484 27372 30485 27436
rect 30419 27371 30485 27372
rect 28947 26212 29013 26213
rect 28947 26148 28948 26212
rect 29012 26148 29013 26212
rect 28947 26147 29013 26148
rect 28763 24308 28829 24309
rect 28763 24244 28764 24308
rect 28828 24244 28829 24308
rect 28763 24243 28829 24244
rect 27843 23628 27909 23629
rect 27843 23564 27844 23628
rect 27908 23564 27909 23628
rect 27843 23563 27909 23564
rect 26555 20636 26621 20637
rect 26555 20572 26556 20636
rect 26620 20572 26621 20636
rect 26555 20571 26621 20572
rect 27107 19820 27173 19821
rect 27107 19756 27108 19820
rect 27172 19756 27173 19820
rect 27107 19755 27173 19756
rect 26923 16420 26989 16421
rect 26923 16356 26924 16420
rect 26988 16356 26989 16420
rect 26923 16355 26989 16356
rect 26371 15196 26437 15197
rect 26371 15132 26372 15196
rect 26436 15132 26437 15196
rect 26371 15131 26437 15132
rect 26371 14380 26437 14381
rect 26371 14316 26372 14380
rect 26436 14316 26437 14380
rect 26371 14315 26437 14316
rect 26187 13972 26253 13973
rect 26187 13908 26188 13972
rect 26252 13908 26253 13972
rect 26187 13907 26253 13908
rect 26190 9485 26250 13907
rect 26374 10165 26434 14315
rect 26926 14109 26986 16355
rect 26923 14108 26989 14109
rect 26923 14044 26924 14108
rect 26988 14044 26989 14108
rect 26923 14043 26989 14044
rect 26739 13700 26805 13701
rect 26739 13636 26740 13700
rect 26804 13636 26805 13700
rect 26739 13635 26805 13636
rect 26371 10164 26437 10165
rect 26371 10100 26372 10164
rect 26436 10100 26437 10164
rect 26371 10099 26437 10100
rect 26742 9621 26802 13635
rect 27110 12341 27170 19755
rect 27846 15333 27906 23563
rect 28766 23493 28826 24243
rect 28950 23901 29010 26147
rect 31526 25941 31586 29003
rect 31523 25940 31589 25941
rect 31523 25876 31524 25940
rect 31588 25876 31589 25940
rect 31523 25875 31589 25876
rect 29315 24988 29381 24989
rect 29315 24924 29316 24988
rect 29380 24924 29381 24988
rect 29315 24923 29381 24924
rect 28947 23900 29013 23901
rect 28947 23836 28948 23900
rect 29012 23836 29013 23900
rect 28947 23835 29013 23836
rect 28763 23492 28829 23493
rect 28763 23428 28764 23492
rect 28828 23428 28829 23492
rect 28763 23427 28829 23428
rect 29131 23492 29197 23493
rect 29131 23428 29132 23492
rect 29196 23428 29197 23492
rect 29131 23427 29197 23428
rect 28579 21452 28645 21453
rect 28579 21388 28580 21452
rect 28644 21388 28645 21452
rect 28579 21387 28645 21388
rect 28211 19412 28277 19413
rect 28211 19348 28212 19412
rect 28276 19348 28277 19412
rect 28211 19347 28277 19348
rect 27291 15332 27357 15333
rect 27291 15268 27292 15332
rect 27356 15268 27357 15332
rect 27291 15267 27357 15268
rect 27843 15332 27909 15333
rect 27843 15268 27844 15332
rect 27908 15268 27909 15332
rect 27843 15267 27909 15268
rect 27107 12340 27173 12341
rect 27107 12276 27108 12340
rect 27172 12276 27173 12340
rect 27107 12275 27173 12276
rect 27294 11661 27354 15267
rect 27843 12884 27909 12885
rect 27843 12820 27844 12884
rect 27908 12820 27909 12884
rect 27843 12819 27909 12820
rect 27291 11660 27357 11661
rect 27291 11596 27292 11660
rect 27356 11596 27357 11660
rect 27291 11595 27357 11596
rect 27846 10029 27906 12819
rect 28027 12748 28093 12749
rect 28027 12684 28028 12748
rect 28092 12684 28093 12748
rect 28027 12683 28093 12684
rect 28030 10301 28090 12683
rect 28214 11389 28274 19347
rect 28395 16148 28461 16149
rect 28395 16084 28396 16148
rect 28460 16084 28461 16148
rect 28395 16083 28461 16084
rect 28211 11388 28277 11389
rect 28211 11324 28212 11388
rect 28276 11324 28277 11388
rect 28211 11323 28277 11324
rect 28027 10300 28093 10301
rect 28027 10236 28028 10300
rect 28092 10236 28093 10300
rect 28027 10235 28093 10236
rect 27843 10028 27909 10029
rect 27843 9964 27844 10028
rect 27908 9964 27909 10028
rect 27843 9963 27909 9964
rect 26739 9620 26805 9621
rect 26739 9556 26740 9620
rect 26804 9556 26805 9620
rect 26739 9555 26805 9556
rect 26187 9484 26253 9485
rect 26187 9420 26188 9484
rect 26252 9420 26253 9484
rect 26187 9419 26253 9420
rect 26190 9077 26250 9419
rect 28398 9213 28458 16083
rect 28582 15061 28642 21387
rect 28763 18868 28829 18869
rect 28763 18804 28764 18868
rect 28828 18804 28829 18868
rect 28763 18803 28829 18804
rect 28766 16557 28826 18803
rect 28763 16556 28829 16557
rect 28763 16492 28764 16556
rect 28828 16492 28829 16556
rect 28763 16491 28829 16492
rect 28579 15060 28645 15061
rect 28579 14996 28580 15060
rect 28644 14996 28645 15060
rect 28579 14995 28645 14996
rect 28395 9212 28461 9213
rect 28395 9148 28396 9212
rect 28460 9148 28461 9212
rect 28395 9147 28461 9148
rect 26187 9076 26253 9077
rect 26187 9012 26188 9076
rect 26252 9012 26253 9076
rect 26187 9011 26253 9012
rect 28582 8397 28642 14995
rect 28766 10029 28826 16491
rect 29134 11661 29194 23427
rect 29318 15197 29378 24923
rect 31526 24853 31586 25875
rect 31339 24852 31405 24853
rect 31339 24788 31340 24852
rect 31404 24788 31405 24852
rect 31339 24787 31405 24788
rect 31523 24852 31589 24853
rect 31523 24788 31524 24852
rect 31588 24788 31589 24852
rect 31523 24787 31589 24788
rect 31342 23357 31402 24787
rect 31339 23356 31405 23357
rect 31339 23292 31340 23356
rect 31404 23292 31405 23356
rect 31339 23291 31405 23292
rect 29499 22676 29565 22677
rect 29499 22612 29500 22676
rect 29564 22612 29565 22676
rect 29499 22611 29565 22612
rect 29315 15196 29381 15197
rect 29315 15132 29316 15196
rect 29380 15132 29381 15196
rect 29315 15131 29381 15132
rect 29502 11661 29562 22611
rect 29867 21860 29933 21861
rect 29867 21796 29868 21860
rect 29932 21796 29933 21860
rect 29867 21795 29933 21796
rect 29131 11660 29197 11661
rect 29131 11596 29132 11660
rect 29196 11596 29197 11660
rect 29131 11595 29197 11596
rect 29499 11660 29565 11661
rect 29499 11596 29500 11660
rect 29564 11596 29565 11660
rect 29499 11595 29565 11596
rect 28763 10028 28829 10029
rect 28763 9964 28764 10028
rect 28828 9964 28829 10028
rect 28763 9963 28829 9964
rect 28579 8396 28645 8397
rect 28579 8332 28580 8396
rect 28644 8332 28645 8396
rect 28579 8331 28645 8332
rect 28766 7581 28826 9963
rect 29502 8261 29562 11595
rect 29499 8260 29565 8261
rect 29499 8196 29500 8260
rect 29564 8196 29565 8260
rect 29499 8195 29565 8196
rect 28763 7580 28829 7581
rect 28763 7516 28764 7580
rect 28828 7516 28829 7580
rect 28763 7515 28829 7516
rect 29870 7037 29930 21795
rect 31894 21045 31954 30091
rect 32075 28388 32141 28389
rect 32075 28324 32076 28388
rect 32140 28324 32141 28388
rect 32075 28323 32141 28324
rect 32078 28117 32138 28323
rect 32075 28116 32141 28117
rect 32075 28052 32076 28116
rect 32140 28052 32141 28116
rect 32075 28051 32141 28052
rect 32262 25941 32322 30091
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 32443 29748 32509 29749
rect 32443 29684 32444 29748
rect 32508 29684 32509 29748
rect 32443 29683 32509 29684
rect 32446 29069 32506 29683
rect 32443 29068 32509 29069
rect 32443 29004 32444 29068
rect 32508 29004 32509 29068
rect 32443 29003 32509 29004
rect 34928 28864 35248 29888
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35387 29612 35453 29613
rect 35387 29548 35388 29612
rect 35452 29548 35453 29612
rect 35387 29547 35453 29548
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 33363 28388 33429 28389
rect 33363 28324 33364 28388
rect 33428 28324 33429 28388
rect 33363 28323 33429 28324
rect 32259 25940 32325 25941
rect 32259 25876 32260 25940
rect 32324 25876 32325 25940
rect 32259 25875 32325 25876
rect 32075 24444 32141 24445
rect 32075 24380 32076 24444
rect 32140 24380 32141 24444
rect 32075 24379 32141 24380
rect 31891 21044 31957 21045
rect 31891 20980 31892 21044
rect 31956 20980 31957 21044
rect 31891 20979 31957 20980
rect 31891 20908 31957 20909
rect 31891 20844 31892 20908
rect 31956 20844 31957 20908
rect 31891 20843 31957 20844
rect 31523 20772 31589 20773
rect 31523 20708 31524 20772
rect 31588 20708 31589 20772
rect 31523 20707 31589 20708
rect 30419 19412 30485 19413
rect 30419 19348 30420 19412
rect 30484 19348 30485 19412
rect 30419 19347 30485 19348
rect 30422 10981 30482 19347
rect 31155 15332 31221 15333
rect 31155 15268 31156 15332
rect 31220 15268 31221 15332
rect 31155 15267 31221 15268
rect 30419 10980 30485 10981
rect 30419 10916 30420 10980
rect 30484 10916 30485 10980
rect 30419 10915 30485 10916
rect 29867 7036 29933 7037
rect 29867 6972 29868 7036
rect 29932 6972 29933 7036
rect 29867 6971 29933 6972
rect 31158 6901 31218 15267
rect 31526 8805 31586 20707
rect 31894 20229 31954 20843
rect 31891 20228 31957 20229
rect 31891 20164 31892 20228
rect 31956 20164 31957 20228
rect 31891 20163 31957 20164
rect 31894 12341 31954 20163
rect 32078 12477 32138 24379
rect 32443 22676 32509 22677
rect 32443 22612 32444 22676
rect 32508 22612 32509 22676
rect 32443 22611 32509 22612
rect 32259 19412 32325 19413
rect 32259 19348 32260 19412
rect 32324 19348 32325 19412
rect 32259 19347 32325 19348
rect 32075 12476 32141 12477
rect 32075 12412 32076 12476
rect 32140 12412 32141 12476
rect 32075 12411 32141 12412
rect 31891 12340 31957 12341
rect 31891 12276 31892 12340
rect 31956 12276 31957 12340
rect 31891 12275 31957 12276
rect 31523 8804 31589 8805
rect 31523 8740 31524 8804
rect 31588 8740 31589 8804
rect 31523 8739 31589 8740
rect 31155 6900 31221 6901
rect 31155 6836 31156 6900
rect 31220 6836 31221 6900
rect 31155 6835 31221 6836
rect 32262 6629 32322 19347
rect 32446 7309 32506 22611
rect 33366 19821 33426 28323
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 35390 25533 35450 29547
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35387 25532 35453 25533
rect 35387 25468 35388 25532
rect 35452 25468 35453 25532
rect 35387 25467 35453 25468
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34099 23492 34165 23493
rect 34099 23428 34100 23492
rect 34164 23428 34165 23492
rect 34099 23427 34165 23428
rect 33731 22540 33797 22541
rect 33731 22476 33732 22540
rect 33796 22476 33797 22540
rect 33731 22475 33797 22476
rect 33363 19820 33429 19821
rect 33363 19756 33364 19820
rect 33428 19756 33429 19820
rect 33363 19755 33429 19756
rect 33366 11797 33426 19755
rect 33734 15469 33794 22475
rect 33731 15468 33797 15469
rect 33731 15404 33732 15468
rect 33796 15404 33797 15468
rect 33731 15403 33797 15404
rect 33363 11796 33429 11797
rect 33363 11732 33364 11796
rect 33428 11732 33429 11796
rect 33363 11731 33429 11732
rect 34102 11117 34162 23427
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34651 20772 34717 20773
rect 34651 20708 34652 20772
rect 34716 20708 34717 20772
rect 34651 20707 34717 20708
rect 34654 12069 34714 20707
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34651 12068 34717 12069
rect 34651 12004 34652 12068
rect 34716 12004 34717 12068
rect 34651 12003 34717 12004
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34099 11116 34165 11117
rect 34099 11052 34100 11116
rect 34164 11052 34165 11116
rect 34099 11051 34165 11052
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 32443 7308 32509 7309
rect 32443 7244 32444 7308
rect 32508 7244 32509 7308
rect 32443 7243 32509 7244
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 32259 6628 32325 6629
rect 32259 6564 32260 6628
rect 32324 6564 32325 6628
rect 32259 6563 32325 6564
rect 25819 6356 25885 6357
rect 25819 6292 25820 6356
rect 25884 6292 25885 6356
rect 25819 6291 25885 6292
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 22139 5812 22205 5813
rect 22139 5748 22140 5812
rect 22204 5748 22205 5812
rect 22139 5747 22205 5748
rect 25451 5812 25517 5813
rect 25451 5748 25452 5812
rect 25516 5748 25517 5812
rect 25451 5747 25517 5748
rect 17907 5404 17973 5405
rect 17907 5340 17908 5404
rect 17972 5340 17973 5404
rect 17907 5339 17973 5340
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 37043 20500 37109 20501
rect 37043 20436 37044 20500
rect 37108 20436 37109 20500
rect 37043 20435 37109 20436
rect 37046 19957 37106 20435
rect 37043 19956 37109 19957
rect 37043 19892 37044 19956
rect 37108 19892 37109 19956
rect 37043 19891 37109 19892
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__clkinv_4  _1351_
timestamp 18001
transform -1 0 22540 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 18001
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1353_
timestamp 18001
transform 1 0 25484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 18001
transform -1 0 25392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 18001
transform -1 0 8740 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 18001
transform 1 0 25668 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 18001
transform 1 0 25944 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 18001
transform 1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 18001
transform 1 0 27692 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 18001
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1361_
timestamp 18001
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 18001
transform -1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1363_
timestamp 18001
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 18001
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1365_
timestamp 18001
transform -1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 18001
transform -1 0 34500 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_2  _1367_
timestamp 18001
transform -1 0 31740 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_1  _1368_
timestamp 18001
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1369_
timestamp 18001
transform 1 0 26956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1370_
timestamp 18001
transform -1 0 26864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1371_
timestamp 18001
transform -1 0 25668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_4  _1372_
timestamp 18001
transform -1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__and2b_1  _1373_
timestamp 18001
transform -1 0 29348 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _1374_
timestamp 18001
transform 1 0 26956 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _1375_
timestamp 18001
transform -1 0 25944 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_2  _1376_
timestamp 18001
transform 1 0 33028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_4  _1377_
timestamp 18001
transform -1 0 27508 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1378_
timestamp 18001
transform -1 0 27232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1379_
timestamp 18001
transform 1 0 21528 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1380_
timestamp 18001
transform -1 0 26220 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_2  _1381_
timestamp 18001
transform -1 0 29716 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1382_
timestamp 18001
transform -1 0 27232 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1383_
timestamp 18001
transform -1 0 30544 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1384_
timestamp 18001
transform -1 0 29716 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1385_
timestamp 18001
transform -1 0 28336 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1386_
timestamp 18001
transform 1 0 23644 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1387_
timestamp 18001
transform -1 0 29440 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _1388_
timestamp 18001
transform -1 0 27600 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_4  _1389_
timestamp 18001
transform 1 0 29624 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nand4b_2  _1390_
timestamp 18001
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1391_
timestamp 18001
transform -1 0 27876 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1392_
timestamp 18001
transform -1 0 24196 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1393_
timestamp 18001
transform -1 0 25576 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1394_
timestamp 18001
transform 1 0 24380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1395_
timestamp 18001
transform -1 0 21436 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 18001
transform 1 0 25300 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _1397_
timestamp 18001
transform -1 0 26680 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _1398_
timestamp 18001
transform -1 0 26772 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1399_
timestamp 18001
transform 1 0 26956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _1400_
timestamp 18001
transform -1 0 34224 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_4  _1401_
timestamp 18001
transform -1 0 26864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _1402_
timestamp 18001
transform -1 0 27416 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor4b_4  _1403_
timestamp 18001
transform -1 0 32752 0 1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__or4b_4  _1404_
timestamp 18001
transform 1 0 26312 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 18001
transform -1 0 27416 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1406_
timestamp 18001
transform -1 0 21528 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _1407_
timestamp 18001
transform -1 0 31740 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or4bb_4  _1408_
timestamp 18001
transform -1 0 26864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1409_
timestamp 18001
transform -1 0 26128 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1410_
timestamp 18001
transform -1 0 21528 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1411_
timestamp 18001
transform 1 0 21068 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1412_
timestamp 18001
transform 1 0 24196 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o41ai_2  _1413_
timestamp 18001
transform -1 0 22264 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__or4b_4  _1414_
timestamp 18001
transform -1 0 29072 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and2_1  _1415_
timestamp 18001
transform -1 0 30084 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1416_
timestamp 18001
transform -1 0 26864 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1417_
timestamp 18001
transform 1 0 27416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1418_
timestamp 18001
transform -1 0 26680 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_2  _1419_
timestamp 18001
transform -1 0 30452 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _1420_
timestamp 18001
transform -1 0 26864 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1421_
timestamp 18001
transform 1 0 25300 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _1422_
timestamp 18001
transform 1 0 25116 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1423_
timestamp 18001
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _1424_
timestamp 18001
transform 1 0 23276 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__clkinv_4  _1425_
timestamp 18001
transform 1 0 25116 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1426_
timestamp 18001
transform -1 0 26128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1427_
timestamp 18001
transform 1 0 24840 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1428_
timestamp 18001
transform -1 0 24840 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1429_
timestamp 18001
transform 1 0 24472 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _1430_
timestamp 18001
transform -1 0 30820 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1431_
timestamp 18001
transform 1 0 27508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1432_
timestamp 18001
transform -1 0 27232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1433_
timestamp 18001
transform -1 0 33672 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_4  _1434_
timestamp 18001
transform 1 0 30820 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_2  _1435_
timestamp 18001
transform -1 0 27876 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o41a_1  _1436_
timestamp 18001
transform 1 0 25944 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _1437_
timestamp 18001
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_4  _1438_
timestamp 18001
transform 1 0 25760 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__or4b_1  _1439_
timestamp 18001
transform -1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1440_
timestamp 18001
transform 1 0 26036 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1441_
timestamp 18001
transform 1 0 25300 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1442_
timestamp 18001
transform 1 0 25852 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1443_
timestamp 18001
transform 1 0 25024 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 18001
transform 1 0 25300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_2  _1445_
timestamp 18001
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__o2111a_1  _1446_
timestamp 18001
transform 1 0 25852 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1447_
timestamp 18001
transform -1 0 25484 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1448_
timestamp 18001
transform -1 0 16560 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 18001
transform 1 0 16652 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1450_
timestamp 18001
transform -1 0 24288 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1451_
timestamp 18001
transform 1 0 24472 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1452_
timestamp 18001
transform 1 0 19780 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1453_
timestamp 18001
transform -1 0 20884 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1454_
timestamp 18001
transform -1 0 31372 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1455_
timestamp 18001
transform -1 0 21528 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 18001
transform -1 0 27784 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1457_
timestamp 18001
transform -1 0 21436 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1458_
timestamp 18001
transform 1 0 21528 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1459_
timestamp 18001
transform -1 0 28796 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1460_
timestamp 18001
transform 1 0 26220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1461_
timestamp 18001
transform -1 0 24104 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1462_
timestamp 18001
transform 1 0 27876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1463_
timestamp 18001
transform -1 0 29164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1464_
timestamp 18001
transform -1 0 22448 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1465_
timestamp 18001
transform -1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1466_
timestamp 18001
transform -1 0 27324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1467_
timestamp 18001
transform 1 0 26772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1468_
timestamp 18001
transform -1 0 22264 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1469_
timestamp 18001
transform 1 0 28428 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1470_
timestamp 18001
transform 1 0 20884 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1471_
timestamp 18001
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1472_
timestamp 18001
transform -1 0 26772 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1473_
timestamp 18001
transform -1 0 25576 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1474_
timestamp 18001
transform 1 0 28980 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1475_
timestamp 18001
transform 1 0 26128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1476_
timestamp 18001
transform 1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1477_
timestamp 18001
transform -1 0 26680 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1478_
timestamp 18001
transform 1 0 20516 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1479_
timestamp 18001
transform -1 0 25300 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1480_
timestamp 18001
transform -1 0 23644 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1481_
timestamp 18001
transform -1 0 25944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1482_
timestamp 18001
transform -1 0 24932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1483_
timestamp 18001
transform 1 0 27692 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1484_
timestamp 18001
transform 1 0 25208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1485_
timestamp 18001
transform -1 0 28612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1486_
timestamp 18001
transform -1 0 25392 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1487_
timestamp 18001
transform -1 0 18768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1488_
timestamp 18001
transform -1 0 26956 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1489_
timestamp 18001
transform 1 0 18492 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1490_
timestamp 18001
transform -1 0 27784 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 18001
transform 1 0 27324 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1492_
timestamp 18001
transform -1 0 27416 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1493_
timestamp 18001
transform 1 0 26496 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1494_
timestamp 18001
transform 1 0 22632 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1495_
timestamp 18001
transform -1 0 27416 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1496_
timestamp 18001
transform -1 0 27324 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1497_
timestamp 18001
transform -1 0 21620 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1498_
timestamp 18001
transform -1 0 21712 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1499_
timestamp 18001
transform -1 0 29532 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1500_
timestamp 18001
transform -1 0 28336 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1501_
timestamp 18001
transform 1 0 25024 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1502_
timestamp 18001
transform 1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1503_
timestamp 18001
transform -1 0 28888 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1504_
timestamp 18001
transform 1 0 23736 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _1505_
timestamp 18001
transform -1 0 27508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1506_
timestamp 18001
transform -1 0 21712 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1507_
timestamp 18001
transform -1 0 24840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1508_
timestamp 18001
transform -1 0 25484 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1509_
timestamp 18001
transform -1 0 24656 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1510_
timestamp 18001
transform 1 0 24380 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1511_
timestamp 18001
transform -1 0 24656 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1512_
timestamp 18001
transform -1 0 23920 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1513_
timestamp 18001
transform -1 0 22632 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1514_
timestamp 18001
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1515_
timestamp 18001
transform -1 0 21896 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1516_
timestamp 18001
transform 1 0 22172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1517_
timestamp 18001
transform 1 0 18952 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1518_
timestamp 18001
transform -1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _1519_
timestamp 18001
transform 1 0 27324 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 18001
transform 1 0 27784 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1521_
timestamp 18001
transform 1 0 25852 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1522_
timestamp 18001
transform -1 0 23736 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1523_
timestamp 18001
transform 1 0 22264 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1524_
timestamp 18001
transform 1 0 18492 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _1525_
timestamp 18001
transform -1 0 26956 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1526_
timestamp 18001
transform -1 0 19780 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a32oi_4  _1527_
timestamp 18001
transform 1 0 19688 0 -1 27200
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_2  _1528_
timestamp 18001
transform -1 0 26496 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1529_
timestamp 18001
transform 1 0 26312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1530_
timestamp 18001
transform -1 0 26772 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1531_
timestamp 18001
transform 1 0 25852 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1532_
timestamp 18001
transform 1 0 25852 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1533_
timestamp 18001
transform -1 0 21896 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 18001
transform -1 0 22264 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1535_
timestamp 18001
transform 1 0 21344 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1536_
timestamp 18001
transform -1 0 25300 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_4  _1537_
timestamp 18001
transform 1 0 24380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 18001
transform -1 0 20976 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1539_
timestamp 18001
transform 1 0 23000 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1540_
timestamp 18001
transform -1 0 33488 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1541_
timestamp 18001
transform 1 0 27692 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1542_
timestamp 18001
transform -1 0 27784 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1543_
timestamp 18001
transform 1 0 26956 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 18001
transform 1 0 24104 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 18001
transform 1 0 24656 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1546_
timestamp 18001
transform 1 0 20884 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 18001
transform 1 0 21712 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1548_
timestamp 18001
transform 1 0 20148 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1549_
timestamp 18001
transform -1 0 25024 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1550_
timestamp 18001
transform -1 0 35512 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1551_
timestamp 18001
transform 1 0 35052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1552_
timestamp 18001
transform -1 0 35328 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1553_
timestamp 18001
transform -1 0 35052 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1554_
timestamp 18001
transform -1 0 30452 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1555_
timestamp 18001
transform -1 0 33304 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1556_
timestamp 18001
transform 1 0 35052 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1557_
timestamp 18001
transform -1 0 30912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1558_
timestamp 18001
transform -1 0 34960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1559_
timestamp 18001
transform -1 0 34868 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1560_
timestamp 18001
transform 1 0 35512 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1561_
timestamp 18001
transform 1 0 34868 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1562_
timestamp 18001
transform 1 0 34960 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1563_
timestamp 18001
transform 1 0 33120 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1564_
timestamp 18001
transform 1 0 33580 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1565_
timestamp 18001
transform -1 0 35328 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1566_
timestamp 18001
transform -1 0 33488 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1567_
timestamp 18001
transform 1 0 33396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1568_
timestamp 18001
transform -1 0 32200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1569_
timestamp 18001
transform 1 0 34684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1570_
timestamp 18001
transform -1 0 31556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1571_
timestamp 18001
transform 1 0 28428 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1572_
timestamp 18001
transform -1 0 32016 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1573_
timestamp 18001
transform -1 0 33396 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1574_
timestamp 18001
transform 1 0 32108 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1575_
timestamp 18001
transform -1 0 32844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 18001
transform 1 0 32752 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1577_
timestamp 18001
transform -1 0 28704 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1578_
timestamp 18001
transform -1 0 29808 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1579_
timestamp 18001
transform 1 0 30452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1580_
timestamp 18001
transform -1 0 28612 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1581_
timestamp 18001
transform -1 0 30636 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1582_
timestamp 18001
transform 1 0 28888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1583_
timestamp 18001
transform -1 0 27784 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 18001
transform 1 0 27784 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1585_
timestamp 18001
transform 1 0 33396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1586_
timestamp 18001
transform 1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1587_
timestamp 18001
transform 1 0 30728 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1588_
timestamp 18001
transform -1 0 34592 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1589_
timestamp 18001
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1590_
timestamp 18001
transform -1 0 34868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1591_
timestamp 18001
transform 1 0 33488 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1592_
timestamp 18001
transform 1 0 32660 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 18001
transform 1 0 32752 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1594_
timestamp 18001
transform 1 0 27232 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1595_
timestamp 18001
transform 1 0 27876 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1596_
timestamp 18001
transform -1 0 31280 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1597_
timestamp 18001
transform 1 0 28980 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1598_
timestamp 18001
transform -1 0 29992 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1599_
timestamp 18001
transform 1 0 30360 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1600_
timestamp 18001
transform 1 0 31096 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1601_
timestamp 18001
transform 1 0 33488 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1602_
timestamp 18001
transform 1 0 30176 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1603_
timestamp 18001
transform -1 0 28888 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1604_
timestamp 18001
transform 1 0 33488 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1605_
timestamp 18001
transform 1 0 31924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _1606_
timestamp 18001
transform -1 0 31924 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 18001
transform 1 0 32108 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 18001
transform -1 0 32936 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 18001
transform 1 0 28796 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1610_
timestamp 18001
transform 1 0 27416 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1611_
timestamp 18001
transform 1 0 27968 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1612_
timestamp 18001
transform -1 0 30176 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1613_
timestamp 18001
transform 1 0 29716 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1614_
timestamp 18001
transform 1 0 31004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1615_
timestamp 18001
transform 1 0 29808 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1616_
timestamp 18001
transform 1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1617_
timestamp 18001
transform -1 0 31096 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1618_
timestamp 18001
transform -1 0 30636 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1619_
timestamp 18001
transform 1 0 30820 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1620_
timestamp 18001
transform 1 0 30636 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1621_
timestamp 18001
transform -1 0 31648 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _1622_
timestamp 18001
transform -1 0 30360 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1623_
timestamp 18001
transform -1 0 34040 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1624_
timestamp 18001
transform 1 0 34500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1625_
timestamp 18001
transform -1 0 33120 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1626_
timestamp 18001
transform 1 0 27968 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1627_
timestamp 18001
transform -1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1628_
timestamp 18001
transform 1 0 31096 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 18001
transform 1 0 29532 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 18001
transform 1 0 34776 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1631_
timestamp 18001
transform 1 0 35512 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1632_
timestamp 18001
transform 1 0 32200 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1633_
timestamp 18001
transform -1 0 28428 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1634_
timestamp 18001
transform 1 0 27968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 18001
transform -1 0 28244 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1636_
timestamp 18001
transform -1 0 33212 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1637_
timestamp 18001
transform -1 0 32016 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1638_
timestamp 18001
transform -1 0 30912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1639_
timestamp 18001
transform -1 0 29808 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 18001
transform 1 0 27600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1641_
timestamp 18001
transform 1 0 31096 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1642_
timestamp 18001
transform -1 0 34040 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1643_
timestamp 18001
transform -1 0 32752 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _1644_
timestamp 18001
transform 1 0 31648 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1645_
timestamp 18001
transform 1 0 32844 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1646_
timestamp 18001
transform 1 0 27600 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1647_
timestamp 18001
transform 1 0 33212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 18001
transform -1 0 28336 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1649_
timestamp 18001
transform 1 0 28796 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1650_
timestamp 18001
transform -1 0 29716 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1651_
timestamp 18001
transform 1 0 27968 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1652_
timestamp 18001
transform -1 0 33856 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1653_
timestamp 18001
transform 1 0 29440 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1654_
timestamp 18001
transform 1 0 35052 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1655_
timestamp 18001
transform 1 0 31004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1656_
timestamp 18001
transform 1 0 29624 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1657_
timestamp 18001
transform 1 0 29716 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1658_
timestamp 18001
transform -1 0 28704 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1659_
timestamp 18001
transform 1 0 33672 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1660_
timestamp 18001
transform 1 0 32568 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1661_
timestamp 18001
transform -1 0 33304 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1662_
timestamp 18001
transform 1 0 33304 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1663_
timestamp 18001
transform 1 0 33028 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1664_
timestamp 18001
transform 1 0 35144 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1665_
timestamp 18001
transform 1 0 34868 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1666_
timestamp 18001
transform -1 0 30268 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1667_
timestamp 18001
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1668_
timestamp 18001
transform 1 0 32844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1669_
timestamp 18001
transform 1 0 33212 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1670_
timestamp 18001
transform -1 0 34040 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1671_
timestamp 18001
transform -1 0 34500 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1672_
timestamp 18001
transform -1 0 33120 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1673_
timestamp 18001
transform 1 0 33304 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1674_
timestamp 18001
transform -1 0 33396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1675_
timestamp 18001
transform 1 0 31648 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1676_
timestamp 18001
transform 1 0 30912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 18001
transform 1 0 28888 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1678_
timestamp 18001
transform -1 0 28980 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1679_
timestamp 18001
transform 1 0 28520 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1680_
timestamp 18001
transform -1 0 30084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1681_
timestamp 18001
transform 1 0 30636 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1682_
timestamp 18001
transform 1 0 27784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1683_
timestamp 18001
transform 1 0 30452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1684_
timestamp 18001
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1685_
timestamp 18001
transform 1 0 29256 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1686_
timestamp 18001
transform -1 0 32660 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1687_
timestamp 18001
transform -1 0 33764 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1688_
timestamp 18001
transform -1 0 32752 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1689_
timestamp 18001
transform 1 0 32292 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1690_
timestamp 18001
transform -1 0 28612 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1691_
timestamp 18001
transform 1 0 33948 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1692_
timestamp 18001
transform -1 0 33212 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1693_
timestamp 18001
transform -1 0 32844 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1694_
timestamp 18001
transform 1 0 28796 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1695_
timestamp 18001
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1696_
timestamp 18001
transform 1 0 32292 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1697_
timestamp 18001
transform -1 0 32752 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1698_
timestamp 18001
transform -1 0 33580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1699_
timestamp 18001
transform -1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1700_
timestamp 18001
transform 1 0 30544 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1701_
timestamp 18001
transform -1 0 29992 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1702_
timestamp 18001
transform 1 0 28152 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1703_
timestamp 18001
transform -1 0 31832 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1704_
timestamp 18001
transform -1 0 31740 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1705_
timestamp 18001
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1706_
timestamp 18001
transform 1 0 27968 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1707_
timestamp 18001
transform 1 0 28244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1708_
timestamp 18001
transform 1 0 30176 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1709_
timestamp 18001
transform 1 0 28612 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1710_
timestamp 18001
transform 1 0 28152 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1711_
timestamp 18001
transform -1 0 29072 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1712_
timestamp 18001
transform 1 0 29072 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1713_
timestamp 18001
transform -1 0 29348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1714_
timestamp 18001
transform -1 0 29440 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1715_
timestamp 18001
transform -1 0 34592 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1716_
timestamp 18001
transform 1 0 34132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1717_
timestamp 18001
transform -1 0 33304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1718_
timestamp 18001
transform 1 0 28060 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1719_
timestamp 18001
transform -1 0 34592 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1720_
timestamp 18001
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1721_
timestamp 18001
transform -1 0 35512 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1722_
timestamp 18001
transform 1 0 34960 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1723_
timestamp 18001
transform -1 0 30360 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1724_
timestamp 18001
transform 1 0 34224 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1725_
timestamp 18001
transform 1 0 31280 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1726_
timestamp 18001
transform -1 0 34132 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1727_
timestamp 18001
transform -1 0 33856 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1728_
timestamp 18001
transform 1 0 34316 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1729_
timestamp 18001
transform -1 0 36064 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1730_
timestamp 18001
transform -1 0 35512 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1731_
timestamp 18001
transform -1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1732_
timestamp 18001
transform 1 0 33856 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1733_
timestamp 18001
transform -1 0 31004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1734_
timestamp 18001
transform -1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1735_
timestamp 18001
transform 1 0 31096 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1736_
timestamp 18001
transform -1 0 35420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1737_
timestamp 18001
transform 1 0 34868 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1738_
timestamp 18001
transform 1 0 31372 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1739_
timestamp 18001
transform 1 0 31648 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1740_
timestamp 18001
transform 1 0 32200 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1741_
timestamp 18001
transform 1 0 30636 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1742_
timestamp 18001
transform -1 0 29716 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1743_
timestamp 18001
transform -1 0 30728 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1744_
timestamp 18001
transform -1 0 31004 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1745_
timestamp 18001
transform 1 0 32108 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1746_
timestamp 18001
transform 1 0 29716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1747_
timestamp 18001
transform -1 0 30912 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1748_
timestamp 18001
transform 1 0 30636 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1749_
timestamp 18001
transform -1 0 33672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1750_
timestamp 18001
transform 1 0 29716 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1751_
timestamp 18001
transform -1 0 31832 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1752_
timestamp 18001
transform 1 0 29440 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1753_
timestamp 18001
transform 1 0 33304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1754_
timestamp 18001
transform 1 0 29256 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1755_
timestamp 18001
transform -1 0 31280 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1756_
timestamp 18001
transform -1 0 30912 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1757_
timestamp 18001
transform -1 0 35696 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1758_
timestamp 18001
transform 1 0 30728 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1759_
timestamp 18001
transform 1 0 31924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1760_
timestamp 18001
transform 1 0 32200 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1761_
timestamp 18001
transform 1 0 32476 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1762_
timestamp 18001
transform -1 0 32936 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1763_
timestamp 18001
transform 1 0 25116 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _1764_
timestamp 18001
transform 1 0 24656 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1765_
timestamp 18001
transform -1 0 16192 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1766_
timestamp 18001
transform -1 0 27600 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _1767_
timestamp 18001
transform -1 0 26588 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1768_
timestamp 18001
transform 1 0 15548 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _1769_
timestamp 18001
transform -1 0 26772 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1770_
timestamp 18001
transform -1 0 20516 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1771_
timestamp 18001
transform 1 0 15732 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1772_
timestamp 18001
transform -1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1773_
timestamp 18001
transform 1 0 15180 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1774_
timestamp 18001
transform -1 0 25208 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1775_
timestamp 18001
transform 1 0 15088 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1776_
timestamp 18001
transform 1 0 25116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1777_
timestamp 18001
transform -1 0 20516 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1778_
timestamp 18001
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1779_
timestamp 18001
transform -1 0 19320 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1780_
timestamp 18001
transform -1 0 15548 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1781_
timestamp 18001
transform -1 0 16284 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1782_
timestamp 18001
transform -1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1783_
timestamp 18001
transform -1 0 20516 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1784_
timestamp 18001
transform -1 0 17112 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1785_
timestamp 18001
transform 1 0 14444 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1786_
timestamp 18001
transform -1 0 17572 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1787_
timestamp 18001
transform -1 0 19320 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1788_
timestamp 18001
transform 1 0 17296 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1789_
timestamp 18001
transform -1 0 19136 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1790_
timestamp 18001
transform 1 0 14996 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1791_
timestamp 18001
transform -1 0 15456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1792_
timestamp 18001
transform 1 0 15824 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1793_
timestamp 18001
transform -1 0 17112 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1794_
timestamp 18001
transform 1 0 19320 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1795_
timestamp 18001
transform 1 0 20424 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1796_
timestamp 18001
transform 1 0 21344 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1797_
timestamp 18001
transform -1 0 20240 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1798_
timestamp 18001
transform 1 0 16008 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1799_
timestamp 18001
transform -1 0 17848 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1800_
timestamp 18001
transform 1 0 16744 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1801_
timestamp 18001
transform -1 0 18952 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1802_
timestamp 18001
transform -1 0 17664 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1803_
timestamp 18001
transform 1 0 17388 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1804_
timestamp 18001
transform 1 0 23092 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1805_
timestamp 18001
transform 1 0 24196 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1806_
timestamp 18001
transform -1 0 23092 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1807_
timestamp 18001
transform -1 0 22724 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1808_
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1809_
timestamp 18001
transform 1 0 19504 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1810_
timestamp 18001
transform -1 0 20332 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1811_
timestamp 18001
transform 1 0 19504 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1812_
timestamp 18001
transform -1 0 14352 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1813_
timestamp 18001
transform -1 0 19136 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1814_
timestamp 18001
transform 1 0 19228 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1815_
timestamp 18001
transform 1 0 17388 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1816_
timestamp 18001
transform -1 0 13340 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1817_
timestamp 18001
transform -1 0 11408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1818_
timestamp 18001
transform -1 0 18032 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1819_
timestamp 18001
transform 1 0 17204 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1820_
timestamp 18001
transform -1 0 21252 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1821_
timestamp 18001
transform 1 0 21712 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1822_
timestamp 18001
transform -1 0 20884 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1823_
timestamp 18001
transform -1 0 20884 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1824_
timestamp 18001
transform 1 0 20884 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1825_
timestamp 18001
transform 1 0 18952 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1826_
timestamp 18001
transform -1 0 15272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1827_
timestamp 18001
transform -1 0 14628 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1828_
timestamp 18001
transform -1 0 19136 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1829_
timestamp 18001
transform 1 0 16836 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1830_
timestamp 18001
transform 1 0 16100 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1831_
timestamp 18001
transform 1 0 16836 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1832_
timestamp 18001
transform -1 0 17756 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1833_
timestamp 18001
transform 1 0 18400 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1834_
timestamp 18001
transform -1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1835_
timestamp 18001
transform 1 0 18032 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1836_
timestamp 18001
transform -1 0 19044 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1837_
timestamp 18001
transform 1 0 20884 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1838_
timestamp 18001
transform 1 0 22172 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1839_
timestamp 18001
transform -1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1840_
timestamp 18001
transform -1 0 21436 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1841_
timestamp 18001
transform 1 0 19320 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1842_
timestamp 18001
transform -1 0 18492 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1843_
timestamp 18001
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1844_
timestamp 18001
transform 1 0 19412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1845_
timestamp 18001
transform -1 0 19872 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1846_
timestamp 18001
transform -1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a2111oi_1  _1847_
timestamp 18001
transform -1 0 16652 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1848_
timestamp 18001
transform -1 0 16560 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1849_
timestamp 18001
transform 1 0 16468 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1850_
timestamp 18001
transform -1 0 16008 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1851_
timestamp 18001
transform -1 0 16192 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1852_
timestamp 18001
transform -1 0 15916 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_4  _1853_
timestamp 18001
transform -1 0 16468 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_4  _1854_
timestamp 18001
transform -1 0 16284 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3b_4  _1855_
timestamp 18001
transform -1 0 16468 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__a221o_1  _1856_
timestamp 18001
transform 1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _1857_
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1858_
timestamp 18001
transform -1 0 16192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1859_
timestamp 18001
transform -1 0 14720 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1860_
timestamp 18001
transform 1 0 13064 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1861_
timestamp 18001
transform -1 0 26312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1862_
timestamp 18001
transform 1 0 20056 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1863_
timestamp 18001
transform -1 0 19136 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1864_
timestamp 18001
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1865_
timestamp 18001
transform -1 0 23092 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1866_
timestamp 18001
transform 1 0 17112 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1867_
timestamp 18001
transform -1 0 17020 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1868_
timestamp 18001
transform 1 0 17296 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1869_
timestamp 18001
transform 1 0 16008 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1870_
timestamp 18001
transform 1 0 17480 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1871_
timestamp 18001
transform -1 0 18400 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1872_
timestamp 18001
transform -1 0 17204 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1873_
timestamp 18001
transform 1 0 17296 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _1874_
timestamp 18001
transform -1 0 18308 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1875_
timestamp 18001
transform 1 0 12144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1876_
timestamp 18001
transform -1 0 16376 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1877_
timestamp 18001
transform 1 0 14352 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1878_
timestamp 18001
transform 1 0 14444 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1879_
timestamp 18001
transform 1 0 12512 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1880_
timestamp 18001
transform -1 0 13248 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1881_
timestamp 18001
transform -1 0 12512 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1882_
timestamp 18001
transform -1 0 12788 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1883_
timestamp 18001
transform -1 0 15640 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1884_
timestamp 18001
transform -1 0 14352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1885_
timestamp 18001
transform 1 0 17296 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1886_
timestamp 18001
transform 1 0 20148 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1887_
timestamp 18001
transform -1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1888_
timestamp 18001
transform -1 0 12696 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1889_
timestamp 18001
transform 1 0 11684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1890_
timestamp 18001
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1891_
timestamp 18001
transform 1 0 26128 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1892_
timestamp 18001
transform -1 0 21068 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1893_
timestamp 18001
transform -1 0 27140 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1894_
timestamp 18001
transform 1 0 25944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1895_
timestamp 18001
transform 1 0 26496 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1896_
timestamp 18001
transform 1 0 25852 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1897_
timestamp 18001
transform 1 0 25116 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1898_
timestamp 18001
transform -1 0 21528 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1899_
timestamp 18001
transform 1 0 19780 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _1900_
timestamp 18001
transform -1 0 14996 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1901_
timestamp 18001
transform -1 0 14904 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__o211a_1  _1902_
timestamp 18001
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1903_
timestamp 18001
transform -1 0 19136 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _1904_
timestamp 18001
transform 1 0 19228 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1905_
timestamp 18001
transform 1 0 18308 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1906_
timestamp 18001
transform 1 0 18124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1907_
timestamp 18001
transform -1 0 20240 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1908_
timestamp 18001
transform 1 0 18400 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1909_
timestamp 18001
transform -1 0 19780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1910_
timestamp 18001
transform 1 0 18676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1911_
timestamp 18001
transform 1 0 18216 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1912_
timestamp 18001
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1913_
timestamp 18001
transform 1 0 18124 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1914_
timestamp 18001
transform 1 0 19596 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1915_
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1916_
timestamp 18001
transform -1 0 10304 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1917_
timestamp 18001
transform -1 0 20516 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1918_
timestamp 18001
transform 1 0 23736 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1919_
timestamp 18001
transform 1 0 23460 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1920_
timestamp 18001
transform 1 0 23828 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1921_
timestamp 18001
transform 1 0 9660 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1922_
timestamp 18001
transform -1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1923_
timestamp 18001
transform 1 0 19688 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1924_
timestamp 18001
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1925_
timestamp 18001
transform -1 0 26312 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1926_
timestamp 18001
transform -1 0 28244 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1927_
timestamp 18001
transform -1 0 26864 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1928_
timestamp 18001
transform -1 0 27692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1929_
timestamp 18001
transform -1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1930_
timestamp 18001
transform 1 0 14076 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_4  _1931_
timestamp 18001
transform -1 0 10488 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1932_
timestamp 18001
transform -1 0 9016 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1933_
timestamp 18001
transform 1 0 8004 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1934_
timestamp 18001
transform -1 0 6532 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1935_
timestamp 18001
transform -1 0 14168 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1936_
timestamp 18001
transform -1 0 7360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1937_
timestamp 18001
transform -1 0 6900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1938_
timestamp 18001
transform -1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _1939_
timestamp 18001
transform -1 0 8740 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1940_
timestamp 18001
transform 1 0 3772 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_2  _1941_
timestamp 18001
transform 1 0 8924 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_4  _1942_
timestamp 18001
transform -1 0 9292 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__a221o_1  _1943_
timestamp 18001
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1944_
timestamp 18001
transform -1 0 5152 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1945_
timestamp 18001
transform 1 0 5336 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1946_
timestamp 18001
transform -1 0 21712 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _1947_
timestamp 18001
transform 1 0 22172 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _1948_
timestamp 18001
transform 1 0 21804 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1949_
timestamp 18001
transform 1 0 22356 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1950_
timestamp 18001
transform 1 0 22264 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1951_
timestamp 18001
transform -1 0 23368 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1952_
timestamp 18001
transform 1 0 22724 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1953_
timestamp 18001
transform 1 0 22448 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1954_
timestamp 18001
transform 1 0 21712 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _1955_
timestamp 18001
transform -1 0 21344 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1956_
timestamp 18001
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1957_
timestamp 18001
transform -1 0 23736 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1958_
timestamp 18001
transform -1 0 22080 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1959_
timestamp 18001
transform -1 0 23644 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1960_
timestamp 18001
transform -1 0 23184 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1961_
timestamp 18001
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1962_
timestamp 18001
transform -1 0 22816 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1963_
timestamp 18001
transform -1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1964_
timestamp 18001
transform 1 0 22080 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1965_
timestamp 18001
transform -1 0 26772 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _1966_
timestamp 18001
transform 1 0 23552 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1967_
timestamp 18001
transform -1 0 23644 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1968_
timestamp 18001
transform 1 0 23368 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1969_
timestamp 18001
transform 1 0 24288 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1970_
timestamp 18001
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1971_
timestamp 18001
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1972_
timestamp 18001
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1973_
timestamp 18001
transform 1 0 23644 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1974_
timestamp 18001
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1975_
timestamp 18001
transform 1 0 22172 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1976_
timestamp 18001
transform -1 0 20792 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1977_
timestamp 18001
transform 1 0 20056 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1978_
timestamp 18001
transform 1 0 19872 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1979_
timestamp 18001
transform 1 0 20056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1980_
timestamp 18001
transform -1 0 21712 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _1981_
timestamp 18001
transform 1 0 20700 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1982_
timestamp 18001
transform -1 0 12604 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _1983_
timestamp 18001
transform -1 0 22540 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 18001
transform -1 0 12328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1985_
timestamp 18001
transform -1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1986_
timestamp 18001
transform 1 0 17296 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1987_
timestamp 18001
transform -1 0 17296 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1988_
timestamp 18001
transform -1 0 18032 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _1989_
timestamp 18001
transform -1 0 17572 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1990_
timestamp 18001
transform -1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1991_
timestamp 18001
transform -1 0 10304 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1992_
timestamp 18001
transform 1 0 9384 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1993_
timestamp 18001
transform -1 0 10488 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1994_
timestamp 18001
transform 1 0 12052 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1995_
timestamp 18001
transform -1 0 21620 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1996_
timestamp 18001
transform -1 0 19780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1997_
timestamp 18001
transform -1 0 16652 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1998_
timestamp 18001
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1999_
timestamp 18001
transform -1 0 18400 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2000_
timestamp 18001
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2001_
timestamp 18001
transform 1 0 15088 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2002_
timestamp 18001
transform -1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_2  _2003_
timestamp 18001
transform 1 0 14904 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2004_
timestamp 18001
transform -1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2005_
timestamp 18001
transform -1 0 17664 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2006_
timestamp 18001
transform 1 0 16100 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _2007_
timestamp 18001
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2008_
timestamp 18001
transform 1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2009_
timestamp 18001
transform 1 0 14996 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2010_
timestamp 18001
transform 1 0 13064 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2011_
timestamp 18001
transform -1 0 13800 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2012_
timestamp 18001
transform 1 0 12512 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_2  _2013_
timestamp 18001
transform -1 0 18860 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _2014_
timestamp 18001
transform 1 0 20608 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2015_
timestamp 18001
transform 1 0 20516 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _2016_
timestamp 18001
transform 1 0 19688 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _2017_
timestamp 18001
transform 1 0 24656 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2018_
timestamp 18001
transform 1 0 24656 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _2019_
timestamp 18001
transform -1 0 24288 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2020_
timestamp 18001
transform 1 0 19596 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2021_
timestamp 18001
transform -1 0 19504 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2022_
timestamp 18001
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2023_
timestamp 18001
transform 1 0 19412 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2024_
timestamp 18001
transform -1 0 19504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2025_
timestamp 18001
transform 1 0 23828 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_4  _2026_
timestamp 18001
transform -1 0 26312 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__a31oi_4  _2027_
timestamp 18001
transform -1 0 24104 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__a31o_1  _2028_
timestamp 18001
transform 1 0 22540 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2029_
timestamp 18001
transform -1 0 19044 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _2030_
timestamp 18001
transform -1 0 18584 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _2031_
timestamp 18001
transform -1 0 18676 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2032_
timestamp 18001
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _2033_
timestamp 18001
transform 1 0 17848 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2034_
timestamp 18001
transform -1 0 18400 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2035_
timestamp 18001
transform 1 0 18400 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2036_
timestamp 18001
transform -1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2037_
timestamp 18001
transform -1 0 9384 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _2038_
timestamp 18001
transform -1 0 19136 0 1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _2039_
timestamp 18001
transform -1 0 9936 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2040_
timestamp 18001
transform -1 0 9384 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2041_
timestamp 18001
transform 1 0 9660 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2042_
timestamp 18001
transform 1 0 11960 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2043_
timestamp 18001
transform 1 0 11316 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2044_
timestamp 18001
transform -1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2045_
timestamp 18001
transform 1 0 12420 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2046_
timestamp 18001
transform -1 0 14720 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2047_
timestamp 18001
transform 1 0 12880 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2048_
timestamp 18001
transform -1 0 12512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2049_
timestamp 18001
transform -1 0 11776 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2050_
timestamp 18001
transform -1 0 6256 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2051_
timestamp 18001
transform 1 0 5152 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2052_
timestamp 18001
transform -1 0 6624 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2053_
timestamp 18001
transform 1 0 6624 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2054_
timestamp 18001
transform 1 0 17204 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2055_
timestamp 18001
transform -1 0 13156 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2oi_1  _2056_
timestamp 18001
transform 1 0 9568 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2057_
timestamp 18001
transform -1 0 9660 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2058_
timestamp 18001
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _2059_
timestamp 18001
transform 1 0 10764 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2060_
timestamp 18001
transform -1 0 8832 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2061_
timestamp 18001
transform -1 0 8832 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2062_
timestamp 18001
transform -1 0 8740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2063_
timestamp 18001
transform 1 0 11132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2064_
timestamp 18001
transform 1 0 11500 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2065_
timestamp 18001
transform 1 0 9936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2066_
timestamp 18001
transform -1 0 12144 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2067_
timestamp 18001
transform -1 0 11040 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2068_
timestamp 18001
transform -1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2069_
timestamp 18001
transform 1 0 10304 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2070_
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2071_
timestamp 18001
transform -1 0 10488 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2072_
timestamp 18001
transform -1 0 6900 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2073_
timestamp 18001
transform 1 0 4600 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2074_
timestamp 18001
transform -1 0 5152 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2075_
timestamp 18001
transform 1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2076_
timestamp 18001
transform -1 0 13432 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _2077_
timestamp 18001
transform 1 0 10028 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2078_
timestamp 18001
transform 1 0 13432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2079_
timestamp 18001
transform 1 0 14168 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2080_
timestamp 18001
transform 1 0 14904 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2081_
timestamp 18001
transform -1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2082_
timestamp 18001
transform 1 0 9200 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2083_
timestamp 18001
transform 1 0 7912 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2084_
timestamp 18001
transform 1 0 10488 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2085_
timestamp 18001
transform -1 0 13984 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2086_
timestamp 18001
transform -1 0 8740 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _2087_
timestamp 18001
transform 1 0 7360 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2088_
timestamp 18001
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2089_
timestamp 18001
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2090_
timestamp 18001
transform 1 0 9200 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2091_
timestamp 18001
transform -1 0 8464 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2092_
timestamp 18001
transform 1 0 9108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _2093_
timestamp 18001
transform 1 0 8464 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2094_
timestamp 18001
transform 1 0 4600 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2095_
timestamp 18001
transform -1 0 5336 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2096_
timestamp 18001
transform 1 0 4140 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2097_
timestamp 18001
transform 1 0 4784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2098_
timestamp 18001
transform -1 0 13156 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _2099_
timestamp 18001
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2100_
timestamp 18001
transform 1 0 16008 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2101_
timestamp 18001
transform -1 0 13892 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2102_
timestamp 18001
transform -1 0 18308 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2103_
timestamp 18001
transform 1 0 17388 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2104_
timestamp 18001
transform -1 0 17204 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2105_
timestamp 18001
transform 1 0 12420 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2106_
timestamp 18001
transform -1 0 11408 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2107_
timestamp 18001
transform 1 0 9844 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2108_
timestamp 18001
transform -1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2109_
timestamp 18001
transform -1 0 12144 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2110_
timestamp 18001
transform 1 0 10304 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2111_
timestamp 18001
transform -1 0 9568 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2112_
timestamp 18001
transform -1 0 9660 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2113_
timestamp 18001
transform -1 0 8648 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2114_
timestamp 18001
transform 1 0 8188 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2115_
timestamp 18001
transform 1 0 8556 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2116_
timestamp 18001
transform 1 0 9292 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2117_
timestamp 18001
transform -1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2118_
timestamp 18001
transform 1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2119_
timestamp 18001
transform 1 0 7544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2120_
timestamp 18001
transform 1 0 4416 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2121_
timestamp 18001
transform 1 0 4508 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2122_
timestamp 18001
transform -1 0 5336 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2123_
timestamp 18001
transform 1 0 5612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2124_
timestamp 18001
transform -1 0 15640 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2125_
timestamp 18001
transform 1 0 10212 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2126_
timestamp 18001
transform -1 0 16928 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2127_
timestamp 18001
transform 1 0 14076 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2128_
timestamp 18001
transform 1 0 14812 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2129_
timestamp 18001
transform 1 0 14720 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2130_
timestamp 18001
transform 1 0 11132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2131_
timestamp 18001
transform 1 0 9292 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2132_
timestamp 18001
transform -1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2133_
timestamp 18001
transform 1 0 10580 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2134_
timestamp 18001
transform -1 0 16560 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2135_
timestamp 18001
transform 1 0 7636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _2136_
timestamp 18001
transform 1 0 7820 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2137_
timestamp 18001
transform -1 0 8188 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2138_
timestamp 18001
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2139_
timestamp 18001
transform 1 0 8372 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2140_
timestamp 18001
transform -1 0 8188 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2141_
timestamp 18001
transform -1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2142_
timestamp 18001
transform 1 0 7452 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _2143_
timestamp 18001
transform 1 0 6900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _2144_
timestamp 18001
transform -1 0 7636 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a31oi_1  _2145_
timestamp 18001
transform 1 0 7544 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2146_
timestamp 18001
transform -1 0 7544 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _2147_
timestamp 18001
transform 1 0 10948 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2148_
timestamp 18001
transform 1 0 17020 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2149_
timestamp 18001
transform 1 0 11592 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2150_
timestamp 18001
transform -1 0 17388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _2151_
timestamp 18001
transform 1 0 11868 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _2152_
timestamp 18001
transform 1 0 10120 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2153_
timestamp 18001
transform -1 0 9936 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2154_
timestamp 18001
transform -1 0 12052 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2155_
timestamp 18001
transform 1 0 11132 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2156_
timestamp 18001
transform 1 0 7176 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2157_
timestamp 18001
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2158_
timestamp 18001
transform -1 0 17940 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2159_
timestamp 18001
transform -1 0 18492 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2160_
timestamp 18001
transform 1 0 10488 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2161_
timestamp 18001
transform 1 0 10120 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2162_
timestamp 18001
transform -1 0 17020 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2163_
timestamp 18001
transform 1 0 12696 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2164_
timestamp 18001
transform -1 0 14168 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2165_
timestamp 18001
transform 1 0 12880 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2166_
timestamp 18001
transform 1 0 7728 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _2167_
timestamp 18001
transform 1 0 7636 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _2168_
timestamp 18001
transform 1 0 8924 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2169_
timestamp 18001
transform -1 0 8004 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2170_
timestamp 18001
transform -1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2171_
timestamp 18001
transform -1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_2  _2172_
timestamp 18001
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2173_
timestamp 18001
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2174_
timestamp 18001
transform 1 0 17664 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2175_
timestamp 18001
transform -1 0 8556 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2176_
timestamp 18001
transform 1 0 18308 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _2177_
timestamp 18001
transform 1 0 17388 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2178_
timestamp 18001
transform -1 0 11224 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2179_
timestamp 18001
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2180_
timestamp 18001
transform 1 0 12144 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2181_
timestamp 18001
transform -1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _2182_
timestamp 18001
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2183_
timestamp 18001
transform -1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2184_
timestamp 18001
transform 1 0 10212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2185_
timestamp 18001
transform 1 0 15088 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2186_
timestamp 18001
transform -1 0 16836 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2187_
timestamp 18001
transform 1 0 15180 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2188_
timestamp 18001
transform -1 0 12604 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2189_
timestamp 18001
transform 1 0 5336 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2190_
timestamp 18001
transform -1 0 6072 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2191_
timestamp 18001
transform 1 0 5152 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o41ai_2  _2192_
timestamp 18001
transform -1 0 6256 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ba_1  _2193_
timestamp 18001
transform 1 0 16560 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2194_
timestamp 18001
transform -1 0 16376 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_2  _2195_
timestamp 18001
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _2196_
timestamp 18001
transform 1 0 12144 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _2197_
timestamp 18001
transform 1 0 11040 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__o2bb2a_1  _2198_
timestamp 18001
transform -1 0 13248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2199_
timestamp 18001
transform -1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2200_
timestamp 18001
transform -1 0 13248 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _2201_
timestamp 18001
transform -1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _2202_
timestamp 18001
transform -1 0 17848 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _2203_
timestamp 18001
transform -1 0 17848 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2204_
timestamp 18001
transform -1 0 17940 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _2205_
timestamp 18001
transform 1 0 16836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2206_
timestamp 18001
transform -1 0 13064 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2207_
timestamp 18001
transform -1 0 12512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _2208_
timestamp 18001
transform 1 0 12236 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_4  _2209_
timestamp 18001
transform 1 0 12052 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__a21bo_1  _2210_
timestamp 18001
transform -1 0 19504 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2211_
timestamp 18001
transform -1 0 18400 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2212_
timestamp 18001
transform 1 0 17572 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2213_
timestamp 18001
transform 1 0 19964 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _2214_
timestamp 18001
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2215_
timestamp 18001
transform -1 0 20332 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2216_
timestamp 18001
transform -1 0 18492 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2217_
timestamp 18001
transform -1 0 19136 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2218_
timestamp 18001
transform -1 0 13892 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2219_
timestamp 18001
transform -1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2220_
timestamp 18001
transform -1 0 13156 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_2  _2221_
timestamp 18001
transform 1 0 11868 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _2222_
timestamp 18001
transform 1 0 10580 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2223_
timestamp 18001
transform 1 0 10488 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2224_
timestamp 18001
transform 1 0 9752 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2225_
timestamp 18001
transform -1 0 10120 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2226_
timestamp 18001
transform -1 0 8832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2227_
timestamp 18001
transform 1 0 8280 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _2228_
timestamp 18001
transform -1 0 8648 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2229_
timestamp 18001
transform 1 0 7728 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2230_
timestamp 18001
transform 1 0 7084 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2231_
timestamp 18001
transform -1 0 6256 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2232_
timestamp 18001
transform -1 0 6624 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2233_
timestamp 18001
transform -1 0 8648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2234_
timestamp 18001
transform -1 0 10672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2235_
timestamp 18001
transform -1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _2236_
timestamp 18001
transform -1 0 15824 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2237_
timestamp 18001
transform 1 0 15272 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2238_
timestamp 18001
transform -1 0 14628 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2239_
timestamp 18001
transform 1 0 15548 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2240_
timestamp 18001
transform -1 0 16100 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _2241_
timestamp 18001
transform -1 0 15640 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _2242_
timestamp 18001
transform -1 0 16008 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _2243_
timestamp 18001
transform 1 0 12328 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2244_
timestamp 18001
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2245_
timestamp 18001
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _2246_
timestamp 18001
transform -1 0 14444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2247_
timestamp 18001
transform 1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2248_
timestamp 18001
transform -1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2249_
timestamp 18001
transform 1 0 12788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2250_
timestamp 18001
transform 1 0 12512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _2251_
timestamp 18001
transform 1 0 13248 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2252_
timestamp 18001
transform 1 0 19228 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2253_
timestamp 18001
transform -1 0 13064 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2254_
timestamp 18001
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _2255_
timestamp 18001
transform 1 0 10580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2256_
timestamp 18001
transform -1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2257_
timestamp 18001
transform -1 0 7820 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2258_
timestamp 18001
transform -1 0 10120 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2259_
timestamp 18001
transform -1 0 11684 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2260_
timestamp 18001
transform -1 0 6624 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2261_
timestamp 18001
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2262_
timestamp 18001
transform -1 0 7728 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2263_
timestamp 18001
transform -1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2264_
timestamp 18001
transform -1 0 8280 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2265_
timestamp 18001
transform -1 0 10212 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2266_
timestamp 18001
transform -1 0 11224 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2267_
timestamp 18001
transform -1 0 9016 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _2268_
timestamp 18001
transform -1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2269_
timestamp 18001
transform -1 0 7360 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2270_
timestamp 18001
transform 1 0 8188 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2271_
timestamp 18001
transform 1 0 10488 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2272_
timestamp 18001
transform 1 0 9936 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2273_
timestamp 18001
transform -1 0 10580 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2274_
timestamp 18001
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2275_
timestamp 18001
transform 1 0 19688 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2276_
timestamp 18001
transform -1 0 17020 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2277_
timestamp 18001
transform -1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2278_
timestamp 18001
transform 1 0 16192 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2279_
timestamp 18001
transform 1 0 15364 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2280_
timestamp 18001
transform 1 0 14628 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2281_
timestamp 18001
transform -1 0 18400 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2282_
timestamp 18001
transform -1 0 16100 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2283_
timestamp 18001
transform 1 0 17848 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _2284_
timestamp 18001
transform 1 0 17020 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _2285_
timestamp 18001
transform -1 0 13892 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2286_
timestamp 18001
transform -1 0 13248 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2287_
timestamp 18001
transform 1 0 11132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _2288_
timestamp 18001
transform 1 0 11500 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2289_
timestamp 18001
transform 1 0 11960 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2290_
timestamp 18001
transform 1 0 19228 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2291_
timestamp 18001
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2292_
timestamp 18001
transform 1 0 15548 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2293_
timestamp 18001
transform -1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2294_
timestamp 18001
transform 1 0 14168 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2295_
timestamp 18001
transform 1 0 14628 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2296_
timestamp 18001
transform 1 0 11592 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2297_
timestamp 18001
transform 1 0 14720 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2298_
timestamp 18001
transform 1 0 14168 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2299_
timestamp 18001
transform -1 0 12144 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2300_
timestamp 18001
transform 1 0 13432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _2301_
timestamp 18001
transform -1 0 13708 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2302_
timestamp 18001
transform 1 0 13340 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2303_
timestamp 18001
transform -1 0 24196 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2304_
timestamp 18001
transform -1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2305_
timestamp 18001
transform -1 0 14996 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _2306_
timestamp 18001
transform -1 0 14720 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2307_
timestamp 18001
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2308_
timestamp 18001
transform -1 0 20332 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2309_
timestamp 18001
transform -1 0 17296 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2310_
timestamp 18001
transform 1 0 14720 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2311_
timestamp 18001
transform 1 0 25668 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2312_
timestamp 18001
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _2313_
timestamp 18001
transform 1 0 17020 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2314_
timestamp 18001
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _2315_
timestamp 18001
transform 1 0 18032 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2316_
timestamp 18001
transform -1 0 17848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2317_
timestamp 18001
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2318_
timestamp 18001
transform -1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _2319_
timestamp 18001
transform -1 0 20148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2320_
timestamp 18001
transform -1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2321_
timestamp 18001
transform 1 0 19136 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2322_
timestamp 18001
transform -1 0 17388 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _2323_
timestamp 18001
transform -1 0 16744 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2324_
timestamp 18001
transform 1 0 14812 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2325_
timestamp 18001
transform 1 0 11776 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2326_
timestamp 18001
transform 1 0 15640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2327_
timestamp 18001
transform 1 0 11868 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2328_
timestamp 18001
transform 1 0 10580 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2329_
timestamp 18001
transform 1 0 11960 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2330_
timestamp 18001
transform 1 0 14536 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2331_
timestamp 18001
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _2332_
timestamp 18001
transform 1 0 22908 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2333_
timestamp 18001
transform 1 0 23828 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2334_
timestamp 18001
transform 1 0 24564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2335_
timestamp 18001
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2336_
timestamp 18001
transform 1 0 25024 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2337_
timestamp 18001
transform 1 0 23736 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2338_
timestamp 18001
transform -1 0 23184 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2339_
timestamp 18001
transform -1 0 22540 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _2340_
timestamp 18001
transform 1 0 20608 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2341_
timestamp 18001
transform 1 0 22816 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _2342_
timestamp 18001
transform -1 0 23828 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2343_
timestamp 18001
transform -1 0 24288 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2344_
timestamp 18001
transform -1 0 25392 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2345_
timestamp 18001
transform -1 0 24932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2346_
timestamp 18001
transform 1 0 17480 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2347_
timestamp 18001
transform 1 0 17572 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2348_
timestamp 18001
transform 1 0 16836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2349_
timestamp 18001
transform 1 0 16744 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2350_
timestamp 18001
transform 1 0 14444 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2351_
timestamp 18001
transform -1 0 14628 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2352_
timestamp 18001
transform 1 0 14628 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2353_
timestamp 18001
transform 1 0 14996 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2354_
timestamp 18001
transform -1 0 15824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2355_
timestamp 18001
transform -1 0 15916 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2356_
timestamp 18001
transform -1 0 17296 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2357_
timestamp 18001
transform 1 0 17756 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2358_
timestamp 18001
transform -1 0 17388 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2359_
timestamp 18001
transform 1 0 18492 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2360_
timestamp 18001
transform -1 0 19780 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2361_
timestamp 18001
transform 1 0 20240 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2362_
timestamp 18001
transform -1 0 20240 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2363_
timestamp 18001
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2364_
timestamp 18001
transform 1 0 24288 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2365_
timestamp 18001
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2366_
timestamp 18001
transform -1 0 25392 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2367_
timestamp 18001
transform 1 0 25392 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2368_
timestamp 18001
transform -1 0 23276 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2369_
timestamp 18001
transform -1 0 24288 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2370_
timestamp 18001
transform -1 0 22540 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2371_
timestamp 18001
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2372_
timestamp 18001
transform 1 0 18400 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2373_
timestamp 18001
transform 1 0 16284 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2374_
timestamp 18001
transform 1 0 14904 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2375_
timestamp 18001
transform -1 0 15456 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2376_
timestamp 18001
transform 1 0 18952 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _2377_
timestamp 18001
transform 1 0 20608 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2378_
timestamp 18001
transform 1 0 23184 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _2379_
timestamp 18001
transform 1 0 22816 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_2  _2380_
timestamp 18001
transform -1 0 23920 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_1  _2381_
timestamp 18001
transform 1 0 24104 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _2382_
timestamp 18001
transform 1 0 24196 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2383_
timestamp 18001
transform -1 0 22080 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2384_
timestamp 18001
transform -1 0 21712 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _2385_
timestamp 18001
transform 1 0 18216 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _2386_
timestamp 18001
transform 1 0 21804 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2387_
timestamp 18001
transform 1 0 25024 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2388_
timestamp 18001
transform -1 0 14536 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2389_
timestamp 18001
transform 1 0 10488 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2390_
timestamp 18001
transform 1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2391_
timestamp 18001
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _2392_
timestamp 18001
transform 1 0 11500 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2393_
timestamp 18001
transform 1 0 11960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2394_
timestamp 18001
transform 1 0 23460 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2395_
timestamp 18001
transform 1 0 24380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2396_
timestamp 18001
transform -1 0 23000 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2397_
timestamp 18001
transform -1 0 12144 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2398_
timestamp 18001
transform -1 0 9292 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2399_
timestamp 18001
transform -1 0 10120 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2400_
timestamp 18001
transform 1 0 10764 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2401_
timestamp 18001
transform 1 0 11500 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2402_
timestamp 18001
transform -1 0 21528 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2403_
timestamp 18001
transform -1 0 20332 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2404_
timestamp 18001
transform -1 0 8004 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2405_
timestamp 18001
transform 1 0 10580 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2406_
timestamp 18001
transform 1 0 11224 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2407_
timestamp 18001
transform 1 0 10764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _2408_
timestamp 18001
transform -1 0 8740 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _2409_
timestamp 18001
transform 1 0 8924 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2410_
timestamp 18001
transform -1 0 11408 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2411_
timestamp 18001
transform 1 0 11500 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2412_
timestamp 18001
transform -1 0 12144 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2413_
timestamp 18001
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _2414_
timestamp 18001
transform 1 0 18400 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _2415_
timestamp 18001
transform -1 0 19228 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2416_
timestamp 18001
transform 1 0 19412 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2417_
timestamp 18001
transform 1 0 19596 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _2418_
timestamp 18001
transform 1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2419_
timestamp 18001
transform -1 0 12144 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2420_
timestamp 18001
transform 1 0 11500 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2421_
timestamp 18001
transform 1 0 11132 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2422_
timestamp 18001
transform 1 0 20148 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2423_
timestamp 18001
transform 1 0 19964 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2424_
timestamp 18001
transform -1 0 17388 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2425_
timestamp 18001
transform 1 0 16928 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2426_
timestamp 18001
transform -1 0 19964 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2427_
timestamp 18001
transform 1 0 19228 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2428_
timestamp 18001
transform -1 0 18400 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2429_
timestamp 18001
transform -1 0 11224 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2430_
timestamp 18001
transform 1 0 10580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2431_
timestamp 18001
transform 1 0 10028 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2432_
timestamp 18001
transform 1 0 12328 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2433_
timestamp 18001
transform 1 0 10856 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2434_
timestamp 18001
transform 1 0 12696 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2435_
timestamp 18001
transform -1 0 13248 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2436_
timestamp 18001
transform -1 0 14720 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2437_
timestamp 18001
transform 1 0 14444 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2438_
timestamp 18001
transform -1 0 14628 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2439_
timestamp 18001
transform 1 0 16468 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2440_
timestamp 18001
transform 1 0 17480 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2441_
timestamp 18001
transform -1 0 17664 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2442_
timestamp 18001
transform -1 0 16284 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2443_
timestamp 18001
transform 1 0 10488 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2444_
timestamp 18001
transform 1 0 9936 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _2445_
timestamp 18001
transform -1 0 10212 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2446_
timestamp 18001
transform 1 0 13248 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2447_
timestamp 18001
transform 1 0 13064 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2448_
timestamp 18001
transform -1 0 15824 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2449_
timestamp 18001
transform -1 0 23552 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2450_
timestamp 18001
transform 1 0 22080 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2451_
timestamp 18001
transform 1 0 22908 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _2452_
timestamp 18001
transform 1 0 17848 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _2453_
timestamp 18001
transform -1 0 17480 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2454_
timestamp 18001
transform -1 0 18216 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2455_
timestamp 18001
transform 1 0 21068 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _2456_
timestamp 18001
transform 1 0 10488 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2457_
timestamp 18001
transform 1 0 9936 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2458_
timestamp 18001
transform -1 0 12696 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _2459_
timestamp 18001
transform 1 0 12420 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2460_
timestamp 18001
transform 1 0 12788 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2461_
timestamp 18001
transform -1 0 13340 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2462_
timestamp 18001
transform -1 0 13892 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2463_
timestamp 18001
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2464_
timestamp 18001
transform 1 0 22540 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2465_
timestamp 18001
transform 1 0 24380 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2466_
timestamp 18001
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2467_
timestamp 18001
transform 1 0 24748 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2468_
timestamp 18001
transform -1 0 24196 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _2469_
timestamp 18001
transform 1 0 9752 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2470_
timestamp 18001
transform 1 0 9660 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _2471_
timestamp 18001
transform 1 0 9384 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _2472_
timestamp 18001
transform -1 0 10212 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2473_
timestamp 18001
transform 1 0 9660 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2474_
timestamp 18001
transform 1 0 21712 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2475_
timestamp 18001
transform 1 0 22540 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2476_
timestamp 18001
transform 1 0 26128 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2477_
timestamp 18001
transform 1 0 26312 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2478_
timestamp 18001
transform 1 0 26036 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2479_
timestamp 18001
transform -1 0 24748 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2480_
timestamp 18001
transform 1 0 25668 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2481_
timestamp 18001
transform -1 0 25300 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2482_
timestamp 18001
transform 1 0 25024 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2483_
timestamp 18001
transform -1 0 10764 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2484_
timestamp 18001
transform -1 0 10488 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2485_
timestamp 18001
transform 1 0 10120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2486_
timestamp 18001
transform -1 0 10028 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2487_
timestamp 18001
transform -1 0 10304 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2488_
timestamp 18001
transform -1 0 9476 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2489_
timestamp 18001
transform 1 0 9016 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2490_
timestamp 18001
transform 1 0 25300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2491_
timestamp 18001
transform 1 0 25116 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2492_
timestamp 18001
transform 1 0 26220 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2493_
timestamp 18001
transform -1 0 26772 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2494_
timestamp 18001
transform -1 0 27140 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2495_
timestamp 18001
transform 1 0 25852 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2496_
timestamp 18001
transform 1 0 9476 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _2497_
timestamp 18001
transform -1 0 8832 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2498_
timestamp 18001
transform 1 0 8740 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2499_
timestamp 18001
transform 1 0 8096 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2500_
timestamp 18001
transform -1 0 22724 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _2501_
timestamp 18001
transform -1 0 26220 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _2502_
timestamp 18001
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2503_
timestamp 18001
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 18001
transform 1 0 4692 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2505_
timestamp 18001
transform 1 0 7268 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2507_
timestamp 18001
transform 1 0 4232 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2508_
timestamp 18001
transform 1 0 6348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2509_
timestamp 18001
transform -1 0 6900 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 18001
transform 1 0 4784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2511_
timestamp 18001
transform 1 0 5428 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _2512_
timestamp 18001
transform 1 0 26220 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2513_
timestamp 18001
transform 1 0 25576 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2514_
timestamp 18001
transform 1 0 14076 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2515_
timestamp 18001
transform 1 0 2484 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2516_
timestamp 18001
transform 1 0 7084 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 18001
transform 1 0 6624 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 18001
transform 1 0 2484 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2519_
timestamp 18001
transform 1 0 3772 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2520_
timestamp 18001
transform 1 0 1932 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2521_
timestamp 18001
transform 1 0 3772 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2522_
timestamp 18001
transform 1 0 3404 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2523_
timestamp 18001
transform 1 0 19504 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2524_
timestamp 18001
transform 1 0 24380 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _2525_
timestamp 18001
transform -1 0 22172 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _2526_
timestamp 18001
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2527_
timestamp 18001
transform -1 0 21528 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2528_
timestamp 18001
transform -1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_1  _2529_
timestamp 18001
transform 1 0 21160 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2530_
timestamp 18001
transform -1 0 22540 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2531_
timestamp 18001
transform 1 0 22356 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2532_
timestamp 18001
transform 1 0 22172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2533_
timestamp 18001
transform 1 0 25760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _2534_
timestamp 18001
transform 1 0 24932 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2535_
timestamp 18001
transform -1 0 22632 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _2536_
timestamp 18001
transform 1 0 22264 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2537_
timestamp 18001
transform 1 0 10580 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 18001
transform 1 0 6992 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2539_
timestamp 18001
transform 1 0 12144 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 18001
transform 1 0 7452 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2541_
timestamp 18001
transform 1 0 9568 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 18001
transform 1 0 8924 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2543_
timestamp 18001
transform 1 0 6348 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2544_
timestamp 18001
transform 1 0 6348 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2545_
timestamp 18001
transform 1 0 24656 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2546_
timestamp 18001
transform 1 0 24748 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2547_
timestamp 18001
transform 1 0 22448 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2548_
timestamp 18001
transform 1 0 22540 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2549_
timestamp 18001
transform 1 0 22540 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2550_
timestamp 18001
transform 1 0 22448 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2551_
timestamp 18001
transform -1 0 23736 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2552_
timestamp 18001
transform -1 0 21068 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2553_
timestamp 18001
transform -1 0 22724 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2554_
timestamp 18001
transform -1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2555_
timestamp 18001
transform -1 0 21344 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2556_
timestamp 18001
transform 1 0 20608 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2557_
timestamp 18001
transform 1 0 20792 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2558_
timestamp 18001
transform 1 0 20516 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2559_
timestamp 18001
transform -1 0 10028 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2560_
timestamp 18001
transform -1 0 9660 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2561_
timestamp 18001
transform 1 0 8740 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2562_
timestamp 18001
transform -1 0 19504 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2563_
timestamp 18001
transform -1 0 19044 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2564_
timestamp 18001
transform 1 0 17848 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _2565_
timestamp 18001
transform -1 0 9476 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2566_
timestamp 18001
transform 1 0 9568 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2567_
timestamp 18001
transform 1 0 9016 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _2568_
timestamp 18001
transform -1 0 18400 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _2569_
timestamp 18001
transform -1 0 17480 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2570_
timestamp 18001
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2571_
timestamp 18001
transform 1 0 9660 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2572_
timestamp 18001
transform 1 0 10120 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2573_
timestamp 18001
transform -1 0 16192 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2574_
timestamp 18001
transform 1 0 15640 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2575_
timestamp 18001
transform 1 0 13064 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2576_
timestamp 18001
transform 1 0 14168 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2577_
timestamp 18001
transform 1 0 10120 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2578_
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2579_
timestamp 18001
transform -1 0 11224 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2580_
timestamp 18001
transform -1 0 15640 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2581_
timestamp 18001
transform 1 0 15456 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2582_
timestamp 18001
transform -1 0 15180 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2583_
timestamp 18001
transform 1 0 12604 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2584_
timestamp 18001
transform -1 0 15916 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2585_
timestamp 18001
transform -1 0 15640 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2586_
timestamp 18001
transform -1 0 14628 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2587_
timestamp 18001
transform -1 0 12052 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2588_
timestamp 18001
transform 1 0 11960 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2589_
timestamp 18001
transform 1 0 14628 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2590_
timestamp 18001
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2591_
timestamp 18001
transform 1 0 19688 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _2592_
timestamp 18001
transform -1 0 15640 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2593_
timestamp 18001
transform 1 0 3220 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2594_
timestamp 18001
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2595_
timestamp 18001
transform 1 0 6256 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2596_
timestamp 18001
transform 1 0 2392 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2597_
timestamp 18001
transform 1 0 2208 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2598_
timestamp 18001
transform 1 0 2208 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2599_
timestamp 18001
transform 1 0 3864 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2600_
timestamp 18001
transform 1 0 2392 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _2601_
timestamp 18001
transform 1 0 21068 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _2602_
timestamp 18001
transform 1 0 20240 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2603_
timestamp 18001
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2604_
timestamp 18001
transform -1 0 22264 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2605_
timestamp 18001
transform 1 0 20884 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2606_
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_4  _2607_
timestamp 18001
transform -1 0 21712 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__a21bo_1  _2608_
timestamp 18001
transform 1 0 12788 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2609_
timestamp 18001
transform 1 0 8464 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2610_
timestamp 18001
transform 1 0 8740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2611_
timestamp 18001
transform 1 0 18124 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2612_
timestamp 18001
transform 1 0 7084 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2613_
timestamp 18001
transform -1 0 5704 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2614_
timestamp 18001
transform 1 0 6348 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2615_
timestamp 18001
transform 1 0 6992 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2616_
timestamp 18001
transform 1 0 4692 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2617_
timestamp 18001
transform 1 0 12972 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _2618_
timestamp 18001
transform -1 0 15272 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2619_
timestamp 18001
transform 1 0 13340 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_4  _2620_
timestamp 18001
transform -1 0 14996 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__or3b_2  _2621_
timestamp 18001
transform 1 0 13340 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2622_
timestamp 18001
transform 1 0 12328 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2623_
timestamp 18001
transform -1 0 13064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2624_
timestamp 18001
transform -1 0 13524 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2625_
timestamp 18001
transform -1 0 13616 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _2626_
timestamp 18001
transform 1 0 11776 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2627_
timestamp 18001
transform -1 0 13984 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2628_
timestamp 18001
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2629_
timestamp 18001
transform -1 0 13064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2630_
timestamp 18001
transform 1 0 12052 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2631_
timestamp 18001
transform 1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _2632_
timestamp 18001
transform -1 0 5796 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2633_
timestamp 18001
transform 1 0 4048 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2634_
timestamp 18001
transform 1 0 4784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2635_
timestamp 18001
transform -1 0 11040 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2636_
timestamp 18001
transform 1 0 10304 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2637_
timestamp 18001
transform -1 0 11040 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2638_
timestamp 18001
transform -1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2639_
timestamp 18001
transform -1 0 4784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2640_
timestamp 18001
transform -1 0 13156 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2641_
timestamp 18001
transform -1 0 5796 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2642_
timestamp 18001
transform -1 0 5520 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2643_
timestamp 18001
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2644_
timestamp 18001
transform 1 0 5428 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2645_
timestamp 18001
transform 1 0 8648 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2646_
timestamp 18001
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _2647_
timestamp 18001
transform 1 0 9016 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _2648_
timestamp 18001
transform -1 0 8280 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2649_
timestamp 18001
transform -1 0 7176 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2650_
timestamp 18001
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2651_
timestamp 18001
transform -1 0 8740 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2652_
timestamp 18001
transform 1 0 8924 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2653_
timestamp 18001
transform 1 0 7820 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2654_
timestamp 18001
transform 1 0 7360 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2655_
timestamp 18001
transform 1 0 6624 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2656_
timestamp 18001
transform 1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _2657_
timestamp 18001
transform 1 0 4784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2658_
timestamp 18001
transform 1 0 4416 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2659_
timestamp 18001
transform -1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2660_
timestamp 18001
transform 1 0 4876 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _2661_
timestamp 18001
transform -1 0 5060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2662_
timestamp 18001
transform 1 0 5796 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2663_
timestamp 18001
transform -1 0 8832 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2664_
timestamp 18001
transform -1 0 9108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2665_
timestamp 18001
transform -1 0 5796 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2666_
timestamp 18001
transform -1 0 4876 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2667_
timestamp 18001
transform -1 0 9936 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2668_
timestamp 18001
transform -1 0 7268 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2669_
timestamp 18001
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2670_
timestamp 18001
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2671_
timestamp 18001
transform -1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2672_
timestamp 18001
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2673_
timestamp 18001
transform 1 0 9108 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2674_
timestamp 18001
transform 1 0 7912 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2675_
timestamp 18001
transform 1 0 7452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _2676_
timestamp 18001
transform -1 0 7268 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2677_
timestamp 18001
transform -1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2678_
timestamp 18001
transform 1 0 6348 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2679_
timestamp 18001
transform -1 0 7636 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2680_
timestamp 18001
transform 1 0 6440 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2681_
timestamp 18001
transform 1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2682_
timestamp 18001
transform -1 0 10580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _2683_
timestamp 18001
transform 1 0 9660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2684_
timestamp 18001
transform -1 0 11132 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2685_
timestamp 18001
transform 1 0 5704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2686_
timestamp 18001
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2687_
timestamp 18001
transform 1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2688_
timestamp 18001
transform -1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2689_
timestamp 18001
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2690_
timestamp 18001
transform 1 0 11500 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2691_
timestamp 18001
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _2692_
timestamp 18001
transform 1 0 12512 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2693_
timestamp 18001
transform -1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _2694_
timestamp 18001
transform 1 0 12144 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2695_
timestamp 18001
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2696_
timestamp 18001
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2697_
timestamp 18001
transform 1 0 25944 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2698_
timestamp 18001
transform -1 0 24012 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _2699_
timestamp 18001
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _2700_
timestamp 18001
transform 1 0 2760 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2701_
timestamp 18001
transform 1 0 7636 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2702_
timestamp 18001
transform 1 0 5428 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2703_
timestamp 18001
transform 1 0 3956 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2704_
timestamp 18001
transform 1 0 2300 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2705_
timestamp 18001
transform 1 0 2116 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2706_
timestamp 18001
transform 1 0 4324 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2707_
timestamp 18001
transform 1 0 3404 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _2708_
timestamp 18001
transform -1 0 13248 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2709_
timestamp 18001
transform -1 0 13984 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2710_
timestamp 18001
transform -1 0 29440 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2711_
timestamp 18001
transform -1 0 29900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2712_
timestamp 18001
transform -1 0 18952 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2713_
timestamp 18001
transform 1 0 17204 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2714_
timestamp 18001
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_1  _2715_
timestamp 18001
transform 1 0 32108 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2716_
timestamp 18001
transform 1 0 34132 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2717_
timestamp 18001
transform -1 0 32384 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2718_
timestamp 18001
transform -1 0 30636 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2719_
timestamp 18001
transform 1 0 32568 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 18001
transform -1 0 28704 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2721_
timestamp 18001
transform 1 0 34132 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2722_
timestamp 18001
transform 1 0 34132 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 18001
transform 1 0 32752 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 18001
transform 1 0 29532 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 18001
transform 1 0 26956 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 18001
transform 1 0 26956 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2727_
timestamp 18001
transform -1 0 30360 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _2728_
timestamp 18001
transform -1 0 27784 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2729_
timestamp 18001
transform 1 0 19596 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2730_
timestamp 18001
transform 1 0 23276 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2731_
timestamp 18001
transform 1 0 24840 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2732_
timestamp 18001
transform 1 0 25024 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2733_
timestamp 18001
transform 1 0 21804 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2734_
timestamp 18001
transform 1 0 22080 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2735_
timestamp 18001
transform 1 0 13984 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2736_
timestamp 18001
transform 1 0 32108 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2737_
timestamp 18001
transform 1 0 32108 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2738_
timestamp 18001
transform 1 0 33580 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2739_
timestamp 18001
transform 1 0 32200 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2740_
timestamp 18001
transform -1 0 31372 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2741_
timestamp 18001
transform 1 0 28428 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2742_
timestamp 18001
transform 1 0 15180 0 1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2743_
timestamp 18001
transform 1 0 11684 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2744_
timestamp 18001
transform 1 0 15180 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2745_
timestamp 18001
transform 1 0 11408 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2746_
timestamp 18001
transform 1 0 13064 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2747_
timestamp 18001
transform 1 0 14076 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2748_
timestamp 18001
transform 1 0 25576 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2749_
timestamp 18001
transform 1 0 16192 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2750_
timestamp 18001
transform -1 0 14444 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2751_
timestamp 18001
transform 1 0 17296 0 -1 6528
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2752_
timestamp 18001
transform 1 0 17756 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2753_
timestamp 18001
transform 1 0 17756 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2754_
timestamp 18001
transform 1 0 18676 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2755_
timestamp 18001
transform 1 0 16836 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2756_
timestamp 18001
transform 1 0 16652 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2757_
timestamp 18001
transform 1 0 14720 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2758_
timestamp 18001
transform 1 0 14352 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2759_
timestamp 18001
transform 1 0 11224 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2760_
timestamp 18001
transform 1 0 15180 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2761_
timestamp 18001
transform 1 0 11408 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2762_
timestamp 18001
transform 1 0 9568 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2763_
timestamp 18001
transform 1 0 10120 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2764_
timestamp 18001
transform -1 0 14536 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2765_
timestamp 18001
transform 1 0 12880 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2766_
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2767_
timestamp 18001
transform 1 0 19596 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2768_
timestamp 18001
transform 1 0 13984 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2769_
timestamp 18001
transform 1 0 15088 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2770_
timestamp 18001
transform -1 0 23460 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2771_
timestamp 18001
transform 1 0 22816 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2772_
timestamp 18001
transform 1 0 24932 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2773_
timestamp 18001
transform 1 0 25760 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2774_
timestamp 18001
transform 1 0 4140 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2775_
timestamp 18001
transform 1 0 6440 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2776_
timestamp 18001
transform 1 0 5796 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2777_
timestamp 18001
transform 1 0 3588 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2778_
timestamp 18001
transform -1 0 7084 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2779_
timestamp 18001
transform 1 0 6348 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2780_
timestamp 18001
transform 1 0 3220 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 18001
transform -1 0 5612 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 18001
transform 1 0 1380 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 18001
transform 1 0 6348 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2784_
timestamp 18001
transform 1 0 4784 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2785_
timestamp 18001
transform 1 0 1380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2786_
timestamp 18001
transform 1 0 1472 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2787_
timestamp 18001
transform 1 0 1380 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2788_
timestamp 18001
transform 1 0 2760 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2789_
timestamp 18001
transform 1 0 1564 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2790_
timestamp 18001
transform -1 0 26036 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2791_
timestamp 18001
transform 1 0 10304 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2792_
timestamp 18001
transform 1 0 6348 0 -1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2793_
timestamp 18001
transform 1 0 11592 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2794_
timestamp 18001
transform 1 0 6440 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2795_
timestamp 18001
transform 1 0 8740 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2796_
timestamp 18001
transform 1 0 6624 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2797_
timestamp 18001
transform 1 0 4140 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2798_
timestamp 18001
transform 1 0 4876 0 1 34816
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2799_
timestamp 18001
transform -1 0 27692 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2800_
timestamp 18001
transform 1 0 23092 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2801_
timestamp 18001
transform 1 0 20148 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 18001
transform 1 0 18216 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 18001
transform -1 0 18492 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 18001
transform 1 0 13708 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2805_
timestamp 18001
transform 1 0 12052 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2806_
timestamp 18001
transform -1 0 17572 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2807_
timestamp 18001
transform 1 0 1380 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2808_
timestamp 18001
transform 1 0 8464 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2809_
timestamp 18001
transform 1 0 6348 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2810_
timestamp 18001
transform 1 0 1472 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2811_
timestamp 18001
transform 1 0 1380 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2812_
timestamp 18001
transform 1 0 1380 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2813_
timestamp 18001
transform 1 0 3220 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2814_
timestamp 18001
transform 1 0 1380 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2815_
timestamp 18001
transform -1 0 14352 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2816_
timestamp 18001
transform 1 0 6716 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2817_
timestamp 18001
transform 1 0 18584 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2818_
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2819_
timestamp 18001
transform -1 0 5796 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2820_
timestamp 18001
transform -1 0 7268 0 1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2821_
timestamp 18001
transform 1 0 6348 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2822_
timestamp 18001
transform -1 0 5888 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2823_
timestamp 18001
transform -1 0 6256 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2824_
timestamp 18001
transform 1 0 2944 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2825_
timestamp 18001
transform 1 0 5612 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2826_
timestamp 18001
transform 1 0 2576 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2827_
timestamp 18001
transform 1 0 2852 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2828_
timestamp 18001
transform 1 0 4416 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2829_
timestamp 18001
transform 1 0 4508 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2830_
timestamp 18001
transform 1 0 3772 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2831_
timestamp 18001
transform 1 0 24380 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2832_
timestamp 18001
transform -1 0 26220 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2833_
timestamp 18001
transform 1 0 1840 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2834_
timestamp 18001
transform 1 0 6992 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2835_
timestamp 18001
transform 1 0 5520 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2836_
timestamp 18001
transform 1 0 3404 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2837_
timestamp 18001
transform 1 0 1380 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2838_
timestamp 18001
transform 1 0 1380 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2839_
timestamp 18001
transform 1 0 3588 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2840_
timestamp 18001
transform 1 0 1840 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2841_
timestamp 18001
transform -1 0 13984 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2842_
timestamp 18001
transform 1 0 29532 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2843_
timestamp 18001
transform 1 0 13064 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _2844_
timestamp 18001
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 18001
transform 1 0 24932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 18001
transform 1 0 32660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 18001
transform -1 0 14720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 18001
transform 1 0 26036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 18001
transform 1 0 18124 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 18001
transform 1 0 18676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform 1 0 18768 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 18001
transform -1 0 7360 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 18001
transform -1 0 7636 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 18001
transform -1 0 12880 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 18001
transform -1 0 12512 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 18001
transform -1 0 6072 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 18001
transform -1 0 4784 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 18001
transform -1 0 7360 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 18001
transform 1 0 7820 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 18001
transform 1 0 23000 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 18001
transform -1 0 23460 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 18001
transform 1 0 27600 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 18001
transform -1 0 28152 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 18001
transform -1 0 24288 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 18001
transform -1 0 24288 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 18001
transform 1 0 29900 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 18001
transform 1 0 29532 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_6  clkload0
timestamp 18001
transform 1 0 6348 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload1
timestamp 18001
transform 1 0 6624 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload2
timestamp 18001
transform -1 0 11868 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload3
timestamp 18001
transform -1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload4
timestamp 18001
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload5
timestamp 18001
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload6
timestamp 18001
transform 1 0 8004 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_4  clkload7
timestamp 18001
transform -1 0 23000 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload8
timestamp 18001
transform 1 0 22448 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload9
timestamp 18001
transform -1 0 28336 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload10
timestamp 18001
transform 1 0 25944 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 18001
transform 1 0 23276 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload12
timestamp 18001
transform 1 0 23276 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload13
timestamp 18001
transform -1 0 32016 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload14
timestamp 18001
transform 1 0 28152 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 18001
transform -1 0 13984 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 18001
transform 1 0 17388 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 18001
transform -1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 18001
transform 1 0 21620 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 18001
transform -1 0 24288 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 18001
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 18001
transform -1 0 13800 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 18001
transform 1 0 28428 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 18001
transform -1 0 31740 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout28
timestamp 18001
transform -1 0 29808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 18001
transform -1 0 31372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 18001
transform 1 0 31280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 18001
transform -1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 18001
transform 1 0 31740 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 18001
transform -1 0 31740 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 18001
transform -1 0 32568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 18001
transform -1 0 32752 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout36
timestamp 18001
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 18001
transform -1 0 21252 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 18001
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 18001
transform 1 0 27600 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 18001
transform 1 0 29164 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout41
timestamp 18001
transform -1 0 17204 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 18001
transform 1 0 22448 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 18001
transform 1 0 25484 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 18001
transform -1 0 23552 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 18001
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 18001
transform -1 0 28152 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout47
timestamp 18001
transform 1 0 28428 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 18001
transform -1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 18001
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 18001
transform -1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 18001
transform -1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 18001
transform -1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 18001
transform -1 0 34408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout54
timestamp 18001
transform 1 0 28796 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 18001
transform -1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 18001
transform -1 0 22908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 18001
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 18001
transform 1 0 25208 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 18001
transform 1 0 30912 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 18001
transform -1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp 18001
transform -1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 18001
transform 1 0 27140 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 18001
transform -1 0 21804 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout64
timestamp 18001
transform -1 0 32384 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 18001
transform 1 0 33580 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 18001
transform -1 0 30912 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout67
timestamp 18001
transform 1 0 30084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 18001
transform -1 0 28980 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout69
timestamp 18001
transform 1 0 27140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 18001
transform -1 0 29072 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 18001
transform -1 0 29348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 18001
transform -1 0 28612 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 18001
transform -1 0 27140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 18001
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 18001
transform -1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout76
timestamp 18001
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout77
timestamp 18001
transform -1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 18001
transform -1 0 29164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 18001
transform 1 0 28428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout80
timestamp 18001
transform 1 0 30452 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 18001
transform 1 0 30268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout82
timestamp 18001
transform -1 0 27968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout83
timestamp 18001
transform -1 0 29808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout84
timestamp 18001
transform -1 0 34592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout85
timestamp 18001
transform -1 0 28336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 18001
transform -1 0 30268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 18001
transform -1 0 34868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 18001
transform -1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 18001
transform 1 0 32660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp 18001
transform -1 0 35236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 18001
transform 1 0 27876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 18001
transform 1 0 34132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 18001
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp 18001
transform -1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp 18001
transform -1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 18001
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 18001
transform -1 0 25668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 18001
transform 1 0 24012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp 18001
transform -1 0 25944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout100
timestamp 18001
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout101
timestamp 18001
transform -1 0 25576 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout102
timestamp 18001
transform 1 0 23460 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout103
timestamp 18001
transform 1 0 24748 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout104
timestamp 18001
transform -1 0 24012 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp 18001
transform -1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout106
timestamp 18001
transform 1 0 19964 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout107
timestamp 18001
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 18001
transform -1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 18001
transform -1 0 26588 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 18001
transform 1 0 26772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout111
timestamp 18001
transform -1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout112
timestamp 18001
transform 1 0 26956 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout113
timestamp 18001
transform -1 0 26864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 18001
transform -1 0 17204 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 18001
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 18001
transform -1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout117
timestamp 18001
transform 1 0 9660 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout118
timestamp 18001
transform -1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout119
timestamp 18001
transform -1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout120
timestamp 18001
transform -1 0 27508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout121
timestamp 18001
transform -1 0 35144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout122
timestamp 18001
transform -1 0 8464 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout123
timestamp 18001
transform -1 0 7084 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout124
timestamp 18001
transform -1 0 7820 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout125
timestamp 18001
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout126
timestamp 18001
transform 1 0 17572 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout127
timestamp 18001
transform -1 0 15548 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout128
timestamp 18001
transform -1 0 27508 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout129
timestamp 18001
transform 1 0 35696 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout130
timestamp 18001
transform -1 0 35696 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout131
timestamp 18001
transform -1 0 36156 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout132
timestamp 18001
transform -1 0 33120 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout133
timestamp 18001
transform 1 0 35420 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636986456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 18001
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 18001
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp 18001
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_126
timestamp 18001
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp 18001
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 18001
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 18001
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_161
timestamp 18001
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_205
timestamp 1636986456
transform 1 0 19964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 18001
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 18001
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636986456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 18001
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_253
timestamp 18001
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_259
timestamp 18001
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_266
timestamp 1636986456
transform 1 0 25576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 18001
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636986456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636986456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 18001
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636986456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636986456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 18001
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636986456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 18001
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_381
timestamp 18001
transform 1 0 36156 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp 18001
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_89
timestamp 18001
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 18001
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 18001
transform 1 0 12696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 18001
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_211
timestamp 1636986456
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_237
timestamp 18001
transform 1 0 22908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_251
timestamp 18001
transform 1 0 24196 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_373
timestamp 18001
transform 1 0 35420 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_381
timestamp 18001
transform 1 0 36156 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_97
timestamp 18001
transform 1 0 10028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 18001
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_204
timestamp 1636986456
transform 1 0 19872 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_216
timestamp 1636986456
transform 1 0 20976 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_228
timestamp 1636986456
transform 1 0 22080 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_240
timestamp 1636986456
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_287
timestamp 1636986456
transform 1 0 27508 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 18001
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_377
timestamp 18001
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 18001
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_11
timestamp 1636986456
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1636986456
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1636986456
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 18001
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 18001
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_101
timestamp 18001
transform 1 0 10396 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 18001
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 18001
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_155
timestamp 18001
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_211
timestamp 1636986456
transform 1 0 20516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_237
timestamp 18001
transform 1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_267
timestamp 18001
transform 1 0 25668 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_286
timestamp 1636986456
transform 1 0 27416 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_298
timestamp 1636986456
transform 1 0 28520 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_310
timestamp 1636986456
transform 1 0 29624 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_322
timestamp 1636986456
transform 1 0 30728 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 18001
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_373
timestamp 18001
transform 1 0 35420 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_381
timestamp 18001
transform 1 0 36156 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_109
timestamp 18001
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 18001
transform 1 0 13064 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp 18001
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_184
timestamp 18001
transform 1 0 18032 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 18001
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_216
timestamp 1636986456
transform 1 0 20976 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 18001
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 18001
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_259
timestamp 18001
transform 1 0 24932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_280
timestamp 1636986456
transform 1 0 26864 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_292
timestamp 1636986456
transform 1 0 27968 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 18001
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 18001
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_381
timestamp 18001
transform 1 0 36156 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 18001
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 18001
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 18001
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 18001
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_248
timestamp 18001
transform 1 0 23920 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_257
timestamp 18001
transform 1 0 24748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636986456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636986456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636986456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 18001
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_373
timestamp 18001
transform 1 0 35420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_381
timestamp 18001
transform 1 0 36156 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636986456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636986456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 18001
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 18001
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636986456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 18001
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 18001
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 18001
transform 1 0 14904 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_174
timestamp 18001
transform 1 0 17112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_180
timestamp 18001
transform 1 0 17664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 18001
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_201
timestamp 18001
transform 1 0 19596 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_222
timestamp 18001
transform 1 0 21528 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_235
timestamp 18001
transform 1 0 22724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_249
timestamp 18001
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 18001
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_267
timestamp 1636986456
transform 1 0 25668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_279
timestamp 1636986456
transform 1 0 26772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_291
timestamp 1636986456
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 18001
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 18001
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_329
timestamp 18001
transform 1 0 31372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 18001
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 18001
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 18001
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_381
timestamp 18001
transform 1 0 36156 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636986456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 18001
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636986456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636986456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636986456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636986456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 18001
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 18001
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 18001
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 18001
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 18001
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_175
timestamp 18001
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_212
timestamp 1636986456
transform 1 0 20608 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636986456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636986456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636986456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_261
timestamp 18001
transform 1 0 25116 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_270
timestamp 18001
transform 1 0 25944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_296
timestamp 18001
transform 1 0 28336 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636986456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 18001
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 18001
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_357
timestamp 1636986456
transform 1 0 33948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_369
timestamp 1636986456
transform 1 0 35052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_381
timestamp 18001
transform 1 0 36156 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636986456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636986456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636986456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 18001
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636986456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636986456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_109
timestamp 18001
transform 1 0 11132 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_132
timestamp 18001
transform 1 0 13248 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636986456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_176
timestamp 18001
transform 1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_182
timestamp 1636986456
transform 1 0 17848 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 18001
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1636986456
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_216
timestamp 18001
transform 1 0 20976 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_223
timestamp 18001
transform 1 0 21620 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 18001
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 18001
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_259
timestamp 18001
transform 1 0 24932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_290
timestamp 18001
transform 1 0 27784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_309
timestamp 18001
transform 1 0 29532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_320
timestamp 18001
transform 1 0 30544 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_329
timestamp 18001
transform 1 0 31372 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_337
timestamp 18001
transform 1 0 32108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_358
timestamp 18001
transform 1 0 34040 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636986456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_377
timestamp 18001
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_381
timestamp 18001
transform 1 0 36156 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636986456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 18001
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 18001
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636986456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636986456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636986456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636986456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 18001
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 18001
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1636986456
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_177
timestamp 1636986456
transform 1 0 17388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_189
timestamp 18001
transform 1 0 18492 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp 18001
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_214
timestamp 18001
transform 1 0 20792 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 18001
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_232
timestamp 18001
transform 1 0 22448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_236
timestamp 18001
transform 1 0 22816 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_241
timestamp 18001
transform 1 0 23276 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 18001
transform 1 0 24012 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_295
timestamp 18001
transform 1 0 28244 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_311
timestamp 18001
transform 1 0 29716 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636986456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_349
timestamp 18001
transform 1 0 33212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_373
timestamp 18001
transform 1 0 35420 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_381
timestamp 18001
transform 1 0 36156 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636986456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_53
timestamp 18001
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_71
timestamp 18001
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 18001
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 18001
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_89
timestamp 18001
transform 1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 18001
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 18001
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_141
timestamp 18001
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 18001
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_175
timestamp 18001
transform 1 0 17204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_181
timestamp 18001
transform 1 0 17756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 18001
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_205
timestamp 18001
transform 1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_213
timestamp 18001
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_225
timestamp 1636986456
transform 1 0 21804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_237
timestamp 1636986456
transform 1 0 22908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 18001
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_253
timestamp 18001
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_257
timestamp 18001
transform 1 0 24748 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_262
timestamp 1636986456
transform 1 0 25208 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_289
timestamp 18001
transform 1 0 27692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_299
timestamp 18001
transform 1 0 28612 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_344
timestamp 18001
transform 1 0 32752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_365
timestamp 18001
transform 1 0 34684 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_370
timestamp 1636986456
transform 1 0 35144 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636986456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_39
timestamp 18001
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 18001
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 18001
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 18001
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_67
timestamp 18001
transform 1 0 7268 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_95
timestamp 18001
transform 1 0 9844 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 18001
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_124
timestamp 18001
transform 1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_151
timestamp 18001
transform 1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_159
timestamp 18001
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 18001
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 18001
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 18001
transform 1 0 18768 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 18001
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_237
timestamp 18001
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_245
timestamp 18001
transform 1 0 23644 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_259
timestamp 18001
transform 1 0 24932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_267
timestamp 18001
transform 1 0 25668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_309
timestamp 18001
transform 1 0 29532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_321
timestamp 18001
transform 1 0 30636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 18001
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_337
timestamp 18001
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_371
timestamp 18001
transform 1 0 35236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_379
timestamp 18001
transform 1 0 35972 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 18001
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 18001
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 18001
transform 1 0 6716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_71
timestamp 18001
transform 1 0 7636 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 18001
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 18001
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 18001
transform 1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_128
timestamp 1636986456
transform 1 0 12880 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_165
timestamp 18001
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 18001
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_182
timestamp 18001
transform 1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636986456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_209
timestamp 18001
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_215
timestamp 18001
transform 1 0 20884 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_227
timestamp 18001
transform 1 0 21988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_233
timestamp 18001
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_239
timestamp 1636986456
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 18001
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_266
timestamp 18001
transform 1 0 25576 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_273
timestamp 18001
transform 1 0 26220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_287
timestamp 18001
transform 1 0 27508 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_296
timestamp 18001
transform 1 0 28336 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_305
timestamp 18001
transform 1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_321
timestamp 18001
transform 1 0 30636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_337
timestamp 18001
transform 1 0 32108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_343
timestamp 18001
transform 1 0 32660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_354
timestamp 18001
transform 1 0 33672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 18001
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1636986456
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_377
timestamp 18001
transform 1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_381
timestamp 18001
transform 1 0 36156 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 18001
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_35
timestamp 18001
transform 1 0 4324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 18001
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_67
timestamp 1636986456
transform 1 0 7268 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_79
timestamp 1636986456
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_91
timestamp 18001
transform 1 0 9476 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_97
timestamp 18001
transform 1 0 10028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 18001
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 18001
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_120
timestamp 1636986456
transform 1 0 12144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 18001
transform 1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_150
timestamp 18001
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 18001
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636986456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 18001
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_194
timestamp 18001
transform 1 0 18952 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_211
timestamp 1636986456
transform 1 0 20516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 18001
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_238
timestamp 18001
transform 1 0 23000 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 18001
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_249
timestamp 18001
transform 1 0 24012 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_256
timestamp 18001
transform 1 0 24656 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_264
timestamp 18001
transform 1 0 25392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_272
timestamp 18001
transform 1 0 26128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 18001
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 18001
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_294
timestamp 18001
transform 1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_312
timestamp 18001
transform 1 0 29808 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_319
timestamp 1636986456
transform 1 0 30452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 18001
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 18001
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_337
timestamp 18001
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_357
timestamp 18001
transform 1 0 33948 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_368
timestamp 1636986456
transform 1 0 34960 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_380
timestamp 18001
transform 1 0 36064 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 18001
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_62
timestamp 18001
transform 1 0 6808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 18001
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_99
timestamp 18001
transform 1 0 10212 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_126
timestamp 18001
transform 1 0 12696 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 18001
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 18001
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 18001
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_151
timestamp 18001
transform 1 0 14996 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_159
timestamp 18001
transform 1 0 15732 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_173
timestamp 18001
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_181
timestamp 18001
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 18001
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_222
timestamp 18001
transform 1 0 21528 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_234
timestamp 1636986456
transform 1 0 22632 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_246
timestamp 18001
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 18001
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 18001
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_268
timestamp 18001
transform 1 0 25760 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 18001
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_292
timestamp 18001
transform 1 0 27968 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 18001
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_309
timestamp 18001
transform 1 0 29532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_324
timestamp 18001
transform 1 0 30912 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1636986456
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1636986456
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 18001
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 18001
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1636986456
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 18001
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_381
timestamp 18001
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636986456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 18001
transform 1 0 5796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_68
timestamp 18001
transform 1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_82
timestamp 18001
transform 1 0 8648 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_90
timestamp 18001
transform 1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 18001
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 18001
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_142
timestamp 18001
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 18001
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 18001
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_175
timestamp 1636986456
transform 1 0 17204 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_187
timestamp 1636986456
transform 1 0 18308 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_199
timestamp 18001
transform 1 0 19412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_209
timestamp 18001
transform 1 0 20332 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 18001
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636986456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_237
timestamp 18001
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_241
timestamp 18001
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_248
timestamp 18001
transform 1 0 23920 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_256
timestamp 18001
transform 1 0 24656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 18001
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_311
timestamp 1636986456
transform 1 0 29716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_323
timestamp 1636986456
transform 1 0 30820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 18001
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_343
timestamp 1636986456
transform 1 0 32660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_355
timestamp 18001
transform 1 0 33764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_366
timestamp 18001
transform 1 0 34776 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_376
timestamp 18001
transform 1 0 35696 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 18001
transform 1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_46
timestamp 18001
transform 1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_50
timestamp 18001
transform 1 0 5704 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_56
timestamp 18001
transform 1 0 6256 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_64
timestamp 18001
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 18001
transform 1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 18001
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636986456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636986456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636986456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_121
timestamp 18001
transform 1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_130
timestamp 18001
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 18001
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636986456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_153
timestamp 18001
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_161
timestamp 18001
transform 1 0 15916 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 18001
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_179
timestamp 18001
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 18001
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 18001
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_265
timestamp 18001
transform 1 0 25484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 18001
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_317
timestamp 18001
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_324
timestamp 1636986456
transform 1 0 30912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_336
timestamp 18001
transform 1 0 32016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_344
timestamp 18001
transform 1 0 32752 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 18001
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1636986456
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 18001
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_381
timestamp 18001
transform 1 0 36156 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636986456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 18001
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_43
timestamp 18001
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_94
timestamp 18001
transform 1 0 9752 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 18001
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 18001
transform 1 0 11868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 18001
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_125
timestamp 18001
transform 1 0 12604 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_136
timestamp 1636986456
transform 1 0 13616 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_148
timestamp 18001
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_154
timestamp 18001
transform 1 0 15272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 18001
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636986456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 18001
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_194
timestamp 1636986456
transform 1 0 18952 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 18001
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_210
timestamp 18001
transform 1 0 20424 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 18001
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 18001
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_253
timestamp 18001
transform 1 0 24380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_266
timestamp 18001
transform 1 0 25576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 18001
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_309
timestamp 1636986456
transform 1 0 29532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_321
timestamp 18001
transform 1 0 30636 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 18001
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 18001
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_345
timestamp 18001
transform 1 0 32844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_361
timestamp 18001
transform 1 0 34316 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_373
timestamp 18001
transform 1 0 35420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_381
timestamp 18001
transform 1 0 36156 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 18001
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_50
timestamp 18001
transform 1 0 5704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 18001
transform 1 0 7636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 18001
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 18001
transform 1 0 12604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 18001
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 18001
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 18001
transform 1 0 17388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 18001
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_190
timestamp 18001
transform 1 0 18584 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_204
timestamp 18001
transform 1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_211
timestamp 18001
transform 1 0 20516 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 18001
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 18001
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_259
timestamp 1636986456
transform 1 0 24932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_271
timestamp 18001
transform 1 0 26036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_286
timestamp 18001
transform 1 0 27416 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 18001
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636986456
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1636986456
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_333
timestamp 18001
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_337
timestamp 18001
transform 1 0 32108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_350
timestamp 1636986456
transform 1 0 33304 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 18001
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1636986456
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_377
timestamp 18001
transform 1 0 35788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_381
timestamp 18001
transform 1 0 36156 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636986456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636986456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_39
timestamp 18001
transform 1 0 4692 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_45
timestamp 18001
transform 1 0 5244 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 18001
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 18001
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_67
timestamp 18001
transform 1 0 7268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_92
timestamp 18001
transform 1 0 9568 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_96
timestamp 18001
transform 1 0 9936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 18001
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_116
timestamp 1636986456
transform 1 0 11776 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_128
timestamp 1636986456
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_140
timestamp 18001
transform 1 0 13984 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_148
timestamp 18001
transform 1 0 14720 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 18001
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 18001
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_189
timestamp 1636986456
transform 1 0 18492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 18001
transform 1 0 19596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 18001
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 18001
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_225
timestamp 18001
transform 1 0 21804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_231
timestamp 18001
transform 1 0 22356 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_258
timestamp 18001
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_271
timestamp 18001
transform 1 0 26036 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_304
timestamp 1636986456
transform 1 0 29072 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_316
timestamp 18001
transform 1 0 30176 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 18001
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1636986456
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1636986456
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1636986456
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_373
timestamp 18001
transform 1 0 35420 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_381
timestamp 18001
transform 1 0 36156 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636986456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636986456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 18001
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_29
timestamp 18001
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_39
timestamp 18001
transform 1 0 4692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_43
timestamp 18001
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 18001
transform 1 0 5520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 18001
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_60
timestamp 1636986456
transform 1 0 6624 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_72
timestamp 1636986456
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 18001
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_92
timestamp 18001
transform 1 0 9568 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 18001
transform 1 0 10304 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_108
timestamp 1636986456
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_120
timestamp 18001
transform 1 0 12144 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_124
timestamp 18001
transform 1 0 12512 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 18001
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 18001
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636986456
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636986456
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 18001
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 18001
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_204
timestamp 18001
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_216
timestamp 18001
transform 1 0 20976 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_230
timestamp 1636986456
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 18001
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 18001
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_253
timestamp 18001
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_261
timestamp 18001
transform 1 0 25116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_270
timestamp 18001
transform 1 0 25944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_276
timestamp 18001
transform 1 0 26496 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_282
timestamp 1636986456
transform 1 0 27048 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_294
timestamp 1636986456
transform 1 0 28152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 18001
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636986456
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_321
timestamp 18001
transform 1 0 30636 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_329
timestamp 18001
transform 1 0 31372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_338
timestamp 18001
transform 1 0 32200 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_346
timestamp 18001
transform 1 0 32936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_354
timestamp 18001
transform 1 0 33672 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_358
timestamp 18001
transform 1 0 34040 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_365
timestamp 18001
transform 1 0 34684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_374
timestamp 18001
transform 1 0 35512 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 18001
transform 1 0 2484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_42
timestamp 18001
transform 1 0 4968 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 18001
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 18001
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_71
timestamp 18001
transform 1 0 7636 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 18001
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 18001
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 18001
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 18001
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 18001
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 18001
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 18001
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_180
timestamp 1636986456
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_192
timestamp 18001
transform 1 0 18768 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 18001
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_207
timestamp 1636986456
transform 1 0 20148 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 18001
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 18001
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636986456
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636986456
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_249
timestamp 18001
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_257
timestamp 18001
transform 1 0 24748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_266
timestamp 18001
transform 1 0 25576 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_274
timestamp 18001
transform 1 0 26312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 18001
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_284
timestamp 18001
transform 1 0 27232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_290
timestamp 18001
transform 1 0 27784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 18001
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_320
timestamp 18001
transform 1 0 30544 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_324
timestamp 1636986456
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_343
timestamp 1636986456
transform 1 0 32660 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_355
timestamp 1636986456
transform 1 0 33764 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_367
timestamp 1636986456
transform 1 0 34868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_379
timestamp 18001
transform 1 0 35972 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636986456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636986456
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 18001
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 18001
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_54
timestamp 18001
transform 1 0 6072 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 18001
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_98
timestamp 18001
transform 1 0 10120 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 18001
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_131
timestamp 18001
transform 1 0 13156 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 18001
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 18001
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 18001
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 18001
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_209
timestamp 18001
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_230
timestamp 18001
transform 1 0 22264 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_239
timestamp 1636986456
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 18001
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_253
timestamp 18001
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_289
timestamp 18001
transform 1 0 27692 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_297
timestamp 18001
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 18001
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_312
timestamp 18001
transform 1 0 29808 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_318
timestamp 18001
transform 1 0 30360 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_327
timestamp 1636986456
transform 1 0 31188 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_339
timestamp 1636986456
transform 1 0 32292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_351
timestamp 1636986456
transform 1 0 33396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 18001
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1636986456
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_377
timestamp 18001
transform 1 0 35788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_381
timestamp 18001
transform 1 0 36156 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 18001
transform 1 0 2484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 18001
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_40
timestamp 18001
transform 1 0 4784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 18001
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 18001
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 18001
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 18001
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 18001
transform 1 0 8188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 18001
transform 1 0 8556 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_89
timestamp 18001
transform 1 0 9292 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_97
timestamp 18001
transform 1 0 10028 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 18001
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_113
timestamp 18001
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_140
timestamp 18001
transform 1 0 13984 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 18001
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 18001
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_169
timestamp 18001
transform 1 0 16652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 18001
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_211
timestamp 18001
transform 1 0 20516 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_217
timestamp 18001
transform 1 0 21068 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_242
timestamp 18001
transform 1 0 23368 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_259
timestamp 1636986456
transform 1 0 24932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_271
timestamp 18001
transform 1 0 26036 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 18001
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_291
timestamp 18001
transform 1 0 27876 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_297
timestamp 18001
transform 1 0 28428 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_315
timestamp 18001
transform 1 0 30084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_323
timestamp 18001
transform 1 0 30820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 18001
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_337
timestamp 18001
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_345
timestamp 1636986456
transform 1 0 32844 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_357
timestamp 18001
transform 1 0 33948 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_365
timestamp 18001
transform 1 0 34684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_374
timestamp 18001
transform 1 0 35512 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636986456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_37
timestamp 1636986456
transform 1 0 4508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_49
timestamp 18001
transform 1 0 5612 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_53
timestamp 18001
transform 1 0 5980 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_63
timestamp 18001
transform 1 0 6900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_71
timestamp 18001
transform 1 0 7636 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 18001
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 18001
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_92
timestamp 18001
transform 1 0 9568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_101
timestamp 18001
transform 1 0 10396 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_107
timestamp 1636986456
transform 1 0 10948 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 18001
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 18001
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 18001
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 18001
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_166
timestamp 1636986456
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_184
timestamp 1636986456
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 18001
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_211
timestamp 1636986456
transform 1 0 20516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 18001
transform 1 0 21620 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_237
timestamp 1636986456
transform 1 0 22908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp 18001
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636986456
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 18001
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_269
timestamp 18001
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_285
timestamp 18001
transform 1 0 27324 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_293
timestamp 18001
transform 1 0 28060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 18001
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 18001
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1636986456
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_321
timestamp 18001
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_327
timestamp 18001
transform 1 0 31188 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_334
timestamp 1636986456
transform 1 0 31832 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_346
timestamp 18001
transform 1 0 32936 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_355
timestamp 18001
transform 1 0 33764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 18001
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1636986456
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 18001
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_381
timestamp 18001
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 18001
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 18001
transform 1 0 4232 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_74
timestamp 18001
transform 1 0 7912 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_80
timestamp 1636986456
transform 1 0 8464 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_92
timestamp 18001
transform 1 0 9568 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_100
timestamp 18001
transform 1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 18001
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 18001
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_117
timestamp 18001
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_130
timestamp 18001
transform 1 0 13064 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_135
timestamp 18001
transform 1 0 13524 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_145
timestamp 18001
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_151
timestamp 18001
transform 1 0 14996 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 18001
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 18001
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 18001
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_182
timestamp 18001
transform 1 0 17848 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_190
timestamp 18001
transform 1 0 18584 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 18001
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 18001
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_231
timestamp 1636986456
transform 1 0 22356 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_248
timestamp 18001
transform 1 0 23920 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_263
timestamp 18001
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 18001
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 18001
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_295
timestamp 18001
transform 1 0 28244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_301
timestamp 18001
transform 1 0 28796 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_309
timestamp 1636986456
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 18001
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1636986456
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1636986456
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1636986456
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_373
timestamp 18001
transform 1 0 35420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_381
timestamp 18001
transform 1 0 36156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 18001
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 18001
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 18001
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_44
timestamp 18001
transform 1 0 5152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_48
timestamp 18001
transform 1 0 5520 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_69
timestamp 18001
transform 1 0 7452 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 18001
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_91
timestamp 18001
transform 1 0 9476 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 18001
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 18001
transform 1 0 11960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_150
timestamp 18001
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_164
timestamp 18001
transform 1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 18001
transform 1 0 16744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 18001
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_205
timestamp 18001
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_212
timestamp 18001
transform 1 0 20608 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_220
timestamp 1636986456
transform 1 0 21344 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_232
timestamp 18001
transform 1 0 22448 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_240
timestamp 18001
transform 1 0 23184 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 18001
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 18001
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_285
timestamp 18001
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_296
timestamp 1636986456
transform 1 0 28336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 18001
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_317
timestamp 1636986456
transform 1 0 30268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_329
timestamp 18001
transform 1 0 31372 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 18001
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_344
timestamp 18001
transform 1 0 32752 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_350
timestamp 18001
transform 1 0 33304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_356
timestamp 18001
transform 1 0 33856 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_365
timestamp 18001
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_375
timestamp 18001
transform 1 0 35604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 18001
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 18001
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 18001
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_22
timestamp 18001
transform 1 0 3128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_26
timestamp 18001
transform 1 0 3496 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 18001
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 18001
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_68
timestamp 18001
transform 1 0 7360 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_100
timestamp 18001
transform 1 0 10304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 18001
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 18001
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 18001
transform 1 0 13248 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_158
timestamp 18001
transform 1 0 15640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 18001
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_184
timestamp 18001
transform 1 0 18032 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_192
timestamp 18001
transform 1 0 18768 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 18001
transform 1 0 20240 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 18001
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 18001
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_229
timestamp 18001
transform 1 0 22172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_237
timestamp 18001
transform 1 0 22908 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_257
timestamp 18001
transform 1 0 24748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_270
timestamp 18001
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 18001
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_284
timestamp 1636986456
transform 1 0 27232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_296
timestamp 18001
transform 1 0 28336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_304
timestamp 18001
transform 1 0 29072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_311
timestamp 1636986456
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_323
timestamp 1636986456
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 18001
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_349
timestamp 18001
transform 1 0 33212 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_365
timestamp 1636986456
transform 1 0 34684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_377
timestamp 18001
transform 1 0 35788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_381
timestamp 18001
transform 1 0 36156 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 18001
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_37
timestamp 18001
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_45
timestamp 18001
transform 1 0 5244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_68
timestamp 18001
transform 1 0 7360 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 18001
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_93
timestamp 1636986456
transform 1 0 9660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_105
timestamp 18001
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_110
timestamp 18001
transform 1 0 11224 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_118
timestamp 18001
transform 1 0 11960 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_124
timestamp 18001
transform 1 0 12512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_133
timestamp 18001
transform 1 0 13340 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 18001
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 18001
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_156
timestamp 18001
transform 1 0 15456 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_168
timestamp 18001
transform 1 0 16560 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_172
timestamp 18001
transform 1 0 16928 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 18001
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 18001
transform 1 0 19596 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 18001
transform 1 0 20056 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_214
timestamp 18001
transform 1 0 20792 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_225
timestamp 18001
transform 1 0 21804 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_236
timestamp 18001
transform 1 0 22816 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_242
timestamp 18001
transform 1 0 23368 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 18001
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_259
timestamp 18001
transform 1 0 24932 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636986456
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1636986456
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 18001
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 18001
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1636986456
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1636986456
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1636986456
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1636986456
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 18001
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 18001
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1636986456
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_377
timestamp 18001
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_381
timestamp 18001
transform 1 0 36156 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 18001
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_45
timestamp 18001
transform 1 0 5244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_57
timestamp 18001
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_63
timestamp 18001
transform 1 0 6900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_84
timestamp 18001
transform 1 0 8832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_88
timestamp 18001
transform 1 0 9200 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 18001
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 18001
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_121
timestamp 18001
transform 1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_138
timestamp 18001
transform 1 0 13800 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 18001
transform 1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_157
timestamp 18001
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 18001
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636986456
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_181
timestamp 18001
transform 1 0 17756 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_185
timestamp 18001
transform 1 0 18124 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_194
timestamp 18001
transform 1 0 18952 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 18001
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 18001
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 18001
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_249
timestamp 18001
transform 1 0 24012 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_254
timestamp 18001
transform 1 0 24472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_262
timestamp 18001
transform 1 0 25208 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_268
timestamp 18001
transform 1 0 25760 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 18001
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 18001
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_289
timestamp 18001
transform 1 0 27692 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_303
timestamp 1636986456
transform 1 0 28980 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_315
timestamp 18001
transform 1 0 30084 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_321
timestamp 18001
transform 1 0 30636 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 18001
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1636986456
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1636986456
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1636986456
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_373
timestamp 18001
transform 1 0 35420 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_381
timestamp 18001
transform 1 0 36156 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 18001
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 18001
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 18001
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 18001
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_94
timestamp 18001
transform 1 0 9752 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_127
timestamp 1636986456
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 18001
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 18001
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_183
timestamp 18001
transform 1 0 17940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 18001
transform 1 0 20240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_225
timestamp 18001
transform 1 0 21804 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_237
timestamp 1636986456
transform 1 0 22908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 18001
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 18001
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_259
timestamp 18001
transform 1 0 24932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_265
timestamp 18001
transform 1 0 25484 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_284
timestamp 1636986456
transform 1 0 27232 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_296
timestamp 1636986456
transform 1 0 28336 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1636986456
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1636986456
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_333
timestamp 18001
transform 1 0 31740 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_346
timestamp 18001
transform 1 0 32936 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 18001
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 18001
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_365
timestamp 18001
transform 1 0 34684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_379
timestamp 18001
transform 1 0 35972 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_15
timestamp 18001
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_35
timestamp 18001
transform 1 0 4324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_39
timestamp 18001
transform 1 0 4692 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp 18001
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636986456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_69
timestamp 18001
transform 1 0 7452 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_77
timestamp 18001
transform 1 0 8188 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 18001
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1636986456
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_142
timestamp 1636986456
transform 1 0 14168 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_154
timestamp 1636986456
transform 1 0 15272 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 18001
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_174
timestamp 18001
transform 1 0 17112 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_199
timestamp 18001
transform 1 0 19412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_207
timestamp 18001
transform 1 0 20148 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636986456
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_237
timestamp 18001
transform 1 0 22908 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_245
timestamp 18001
transform 1 0 23644 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_266
timestamp 18001
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_270
timestamp 18001
transform 1 0 25944 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 18001
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_289
timestamp 18001
transform 1 0 27692 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 18001
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_307
timestamp 18001
transform 1 0 29348 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_324
timestamp 1636986456
transform 1 0 30912 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1636986456
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1636986456
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1636986456
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_373
timestamp 18001
transform 1 0 35420 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_381
timestamp 18001
transform 1 0 36156 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 18001
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_49
timestamp 18001
transform 1 0 5612 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 18001
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_59
timestamp 18001
transform 1 0 6532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_63
timestamp 18001
transform 1 0 6900 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_68
timestamp 18001
transform 1 0 7360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 18001
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 18001
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_99
timestamp 18001
transform 1 0 10212 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_107
timestamp 18001
transform 1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_114
timestamp 18001
transform 1 0 11592 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_151
timestamp 18001
transform 1 0 14996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_157
timestamp 18001
transform 1 0 15548 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 18001
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_172
timestamp 18001
transform 1 0 16928 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_176
timestamp 1636986456
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 18001
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 18001
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_204
timestamp 18001
transform 1 0 19872 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_211
timestamp 1636986456
transform 1 0 20516 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_223
timestamp 1636986456
transform 1 0 21620 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_235
timestamp 18001
transform 1 0 22724 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_243
timestamp 18001
transform 1 0 23460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 18001
transform 1 0 25484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_273
timestamp 18001
transform 1 0 26220 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_281
timestamp 18001
transform 1 0 26956 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_287
timestamp 18001
transform 1 0 27508 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_296
timestamp 1636986456
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636986456
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_321
timestamp 18001
transform 1 0 30636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_327
timestamp 18001
transform 1 0 31188 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_332
timestamp 1636986456
transform 1 0 31648 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_344
timestamp 1636986456
transform 1 0 32752 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 18001
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1636986456
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 18001
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_381
timestamp 18001
transform 1 0 36156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 18001
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_34
timestamp 18001
transform 1 0 4232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 18001
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 18001
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_86
timestamp 1636986456
transform 1 0 9016 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_98
timestamp 1636986456
transform 1 0 10120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 18001
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_116
timestamp 18001
transform 1 0 11776 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 18001
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_174
timestamp 18001
transform 1 0 17112 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_184
timestamp 18001
transform 1 0 18032 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 18001
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 18001
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_233
timestamp 18001
transform 1 0 22540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 18001
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_249
timestamp 18001
transform 1 0 24012 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_253
timestamp 18001
transform 1 0 24380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 18001
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_290
timestamp 18001
transform 1 0 27784 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_295
timestamp 1636986456
transform 1 0 28244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_307
timestamp 18001
transform 1 0 29348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_316
timestamp 18001
transform 1 0 30176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_320
timestamp 18001
transform 1 0 30544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 18001
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 18001
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_346
timestamp 18001
transform 1 0 32936 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_357
timestamp 18001
transform 1 0 33948 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_363
timestamp 18001
transform 1 0 34500 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_367
timestamp 1636986456
transform 1 0 34868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_379
timestamp 18001
transform 1 0 35972 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636986456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 18001
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_44
timestamp 18001
transform 1 0 5152 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_52
timestamp 18001
transform 1 0 5888 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_60
timestamp 18001
transform 1 0 6624 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_100
timestamp 18001
transform 1 0 10304 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_126
timestamp 18001
transform 1 0 12696 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_132
timestamp 18001
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 18001
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 18001
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_169
timestamp 18001
transform 1 0 16652 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 18001
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_212
timestamp 18001
transform 1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_220
timestamp 18001
transform 1 0 21344 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 18001
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 18001
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636986456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636986456
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1636986456
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_289
timestamp 18001
transform 1 0 27692 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_300
timestamp 18001
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_325
timestamp 18001
transform 1 0 31004 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_335
timestamp 18001
transform 1 0 31924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_356
timestamp 18001
transform 1 0 33856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_380
timestamp 18001
transform 1 0 36064 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_24
timestamp 18001
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_28
timestamp 18001
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 18001
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 18001
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636986456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 18001
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_73
timestamp 18001
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_123
timestamp 1636986456
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_135
timestamp 18001
transform 1 0 13524 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 18001
transform 1 0 14904 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_158
timestamp 18001
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 18001
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 18001
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_204
timestamp 18001
transform 1 0 19872 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 18001
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 18001
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_230
timestamp 18001
transform 1 0 22264 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_236
timestamp 18001
transform 1 0 22816 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_244
timestamp 18001
transform 1 0 23552 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_256
timestamp 18001
transform 1 0 24656 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_263
timestamp 1636986456
transform 1 0 25300 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 18001
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 18001
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_286
timestamp 18001
transform 1 0 27416 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_302
timestamp 1636986456
transform 1 0 28888 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_314
timestamp 1636986456
transform 1 0 29992 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_326
timestamp 18001
transform 1 0 31096 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 18001
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1636986456
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1636986456
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1636986456
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_373
timestamp 18001
transform 1 0 35420 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_381
timestamp 18001
transform 1 0 36156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 18001
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 18001
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_67
timestamp 18001
transform 1 0 7268 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 18001
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_99
timestamp 18001
transform 1 0 10212 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_105
timestamp 18001
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_112
timestamp 18001
transform 1 0 11408 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_121
timestamp 18001
transform 1 0 12236 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_127
timestamp 18001
transform 1 0 12788 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 18001
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_146
timestamp 18001
transform 1 0 14536 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 18001
transform 1 0 15272 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_164
timestamp 1636986456
transform 1 0 16192 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_176
timestamp 18001
transform 1 0 17296 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 18001
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_201
timestamp 1636986456
transform 1 0 19596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_213
timestamp 1636986456
transform 1 0 20700 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_225
timestamp 1636986456
transform 1 0 21804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 18001
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_241
timestamp 18001
transform 1 0 23276 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 18001
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_290
timestamp 1636986456
transform 1 0 27784 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 18001
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 18001
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_316
timestamp 18001
transform 1 0 30176 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_320
timestamp 18001
transform 1 0 30544 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1636986456
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_338
timestamp 1636986456
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_350
timestamp 1636986456
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 18001
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1636986456
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_377
timestamp 18001
transform 1 0 35788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_381
timestamp 18001
transform 1 0 36156 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1636986456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_32
timestamp 18001
transform 1 0 4048 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1636986456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_69
timestamp 18001
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_77
timestamp 1636986456
transform 1 0 8188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_89
timestamp 18001
transform 1 0 9292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_99
timestamp 18001
transform 1 0 10212 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 18001
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_132
timestamp 18001
transform 1 0 13248 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_148
timestamp 18001
transform 1 0 14720 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 18001
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_175
timestamp 18001
transform 1 0 17204 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_184
timestamp 1636986456
transform 1 0 18032 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_210
timestamp 18001
transform 1 0 20424 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_37_221
timestamp 18001
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_242
timestamp 18001
transform 1 0 23368 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_258
timestamp 18001
transform 1 0 24840 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_264
timestamp 1636986456
transform 1 0 25392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 18001
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_289
timestamp 18001
transform 1 0 27692 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_300
timestamp 18001
transform 1 0 28704 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 18001
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_352
timestamp 18001
transform 1 0 33488 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_356
timestamp 18001
transform 1 0 33856 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_364
timestamp 18001
transform 1 0 34592 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 18001
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_46
timestamp 1636986456
transform 1 0 5336 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_58
timestamp 18001
transform 1 0 6440 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_64
timestamp 18001
transform 1 0 6992 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 18001
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 18001
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_105
timestamp 18001
transform 1 0 10764 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_116
timestamp 18001
transform 1 0 11776 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_120
timestamp 18001
transform 1 0 12144 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_132
timestamp 18001
transform 1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_144
timestamp 18001
transform 1 0 14352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_175
timestamp 18001
transform 1 0 17204 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_182
timestamp 18001
transform 1 0 17848 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_190
timestamp 18001
transform 1 0 18584 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_204
timestamp 18001
transform 1 0 19872 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_213
timestamp 18001
transform 1 0 20700 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_221
timestamp 18001
transform 1 0 21436 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_237
timestamp 18001
transform 1 0 22908 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 18001
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 18001
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 18001
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_257
timestamp 18001
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_264
timestamp 18001
transform 1 0 25392 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_274
timestamp 18001
transform 1 0 26312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_288
timestamp 18001
transform 1 0 27600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 18001
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_309
timestamp 18001
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_324
timestamp 18001
transform 1 0 30912 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_340
timestamp 1636986456
transform 1 0 32384 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_352
timestamp 1636986456
transform 1 0 33488 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_365
timestamp 18001
transform 1 0 34684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_374
timestamp 18001
transform 1 0 35512 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 18001
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_38
timestamp 18001
transform 1 0 4600 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 18001
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_91
timestamp 18001
transform 1 0 9476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_100
timestamp 18001
transform 1 0 10304 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_108
timestamp 18001
transform 1 0 11040 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 18001
transform 1 0 12788 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_142
timestamp 18001
transform 1 0 14168 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_150
timestamp 18001
transform 1 0 14904 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_208
timestamp 1636986456
transform 1 0 20240 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 18001
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_244
timestamp 18001
transform 1 0 23552 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_252
timestamp 18001
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 18001
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 18001
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_289
timestamp 18001
transform 1 0 27692 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_304
timestamp 1636986456
transform 1 0 29072 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_316
timestamp 18001
transform 1 0 30176 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_322
timestamp 18001
transform 1 0 30728 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_337
timestamp 18001
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_345
timestamp 18001
transform 1 0 32844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_359
timestamp 18001
transform 1 0 34132 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_367
timestamp 18001
transform 1 0 34868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_375
timestamp 18001
transform 1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1636986456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_15
timestamp 18001
transform 1 0 2484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 18001
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 18001
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_63
timestamp 18001
transform 1 0 6900 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_76
timestamp 18001
transform 1 0 8096 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 18001
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_103
timestamp 18001
transform 1 0 10580 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_125
timestamp 18001
transform 1 0 12604 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 18001
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_148
timestamp 18001
transform 1 0 14720 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_156
timestamp 18001
transform 1 0 15456 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_171
timestamp 1636986456
transform 1 0 16836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_183
timestamp 1636986456
transform 1 0 17940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 18001
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 18001
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_210
timestamp 1636986456
transform 1 0 20424 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 18001
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 18001
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 18001
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_266
timestamp 18001
transform 1 0 25576 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_275
timestamp 18001
transform 1 0 26404 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_283
timestamp 18001
transform 1 0 27140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_291
timestamp 18001
transform 1 0 27876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 18001
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1636986456
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 18001
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_329
timestamp 1636986456
transform 1 0 31372 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_358
timestamp 18001
transform 1 0 34040 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_32
timestamp 18001
transform 1 0 4048 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 18001
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_57
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_86
timestamp 18001
transform 1 0 9016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_90
timestamp 18001
transform 1 0 9384 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_99
timestamp 1636986456
transform 1 0 10212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 18001
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_127
timestamp 18001
transform 1 0 12788 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1636986456
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_149
timestamp 18001
transform 1 0 14812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 18001
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_169
timestamp 18001
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_200
timestamp 18001
transform 1 0 19504 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_209
timestamp 18001
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_217
timestamp 18001
transform 1 0 21068 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_232
timestamp 18001
transform 1 0 22448 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_250
timestamp 18001
transform 1 0 24104 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_263
timestamp 18001
transform 1 0 25300 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_269
timestamp 18001
transform 1 0 25852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 18001
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_290
timestamp 18001
transform 1 0 27784 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_296
timestamp 18001
transform 1 0 28336 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_303
timestamp 18001
transform 1 0 28980 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_311
timestamp 18001
transform 1 0 29716 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_319
timestamp 18001
transform 1 0 30452 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 18001
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_344
timestamp 18001
transform 1 0 32752 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_348
timestamp 18001
transform 1 0 33120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_3
timestamp 18001
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_11
timestamp 18001
transform 1 0 2116 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 18001
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp 18001
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_63
timestamp 18001
transform 1 0 6900 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 18001
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_90
timestamp 18001
transform 1 0 9384 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp 18001
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 18001
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 18001
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_148
timestamp 18001
transform 1 0 14720 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_159
timestamp 1636986456
transform 1 0 15732 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_200
timestamp 18001
transform 1 0 19504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_209
timestamp 18001
transform 1 0 20332 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_233
timestamp 18001
transform 1 0 22540 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_294
timestamp 1636986456
transform 1 0 28152 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 18001
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_314
timestamp 18001
transform 1 0 29992 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_320
timestamp 18001
transform 1 0 30544 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_358
timestamp 18001
transform 1 0 34040 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_365
timestamp 18001
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_372
timestamp 18001
transform 1 0 35328 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_381
timestamp 18001
transform 1 0 36156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_54
timestamp 18001
transform 1 0 6072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_84
timestamp 18001
transform 1 0 8832 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 18001
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_122
timestamp 18001
transform 1 0 12328 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_131
timestamp 1636986456
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_143
timestamp 1636986456
transform 1 0 14260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_155
timestamp 18001
transform 1 0 15364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_166
timestamp 18001
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_181
timestamp 18001
transform 1 0 17756 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_195
timestamp 18001
transform 1 0 19044 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_206
timestamp 1636986456
transform 1 0 20056 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_218
timestamp 18001
transform 1 0 21160 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636986456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_237
timestamp 18001
transform 1 0 22908 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_245
timestamp 18001
transform 1 0 23644 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_261
timestamp 18001
transform 1 0 25116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 18001
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_288
timestamp 18001
transform 1 0 27600 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_296
timestamp 18001
transform 1 0 28336 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_318
timestamp 18001
transform 1 0 30360 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_326
timestamp 18001
transform 1 0 31096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_337
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_351
timestamp 18001
transform 1 0 33396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_366
timestamp 18001
transform 1 0 34776 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_374
timestamp 18001
transform 1 0 35512 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1636986456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1636986456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_56
timestamp 18001
transform 1 0 6256 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_60
timestamp 18001
transform 1 0 6624 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_65
timestamp 18001
transform 1 0 7084 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 18001
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_92
timestamp 18001
transform 1 0 9568 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_99
timestamp 1636986456
transform 1 0 10212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_111
timestamp 18001
transform 1 0 11316 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_119
timestamp 18001
transform 1 0 12052 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_131
timestamp 18001
transform 1 0 13156 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 18001
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_156
timestamp 1636986456
transform 1 0 15456 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_182
timestamp 1636986456
transform 1 0 17848 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 18001
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1636986456
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_209
timestamp 18001
transform 1 0 20332 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_227
timestamp 18001
transform 1 0 21988 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_236
timestamp 1636986456
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 18001
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636986456
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_265
timestamp 18001
transform 1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_287
timestamp 18001
transform 1 0 27508 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 18001
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 18001
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_309
timestamp 18001
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_315
timestamp 18001
transform 1 0 30084 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_324
timestamp 1636986456
transform 1 0 30912 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_336
timestamp 18001
transform 1 0 32016 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 18001
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 18001
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_368
timestamp 18001
transform 1 0 34960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_375
timestamp 18001
transform 1 0 35604 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_3
timestamp 18001
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_11
timestamp 18001
transform 1 0 2116 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_21
timestamp 18001
transform 1 0 3036 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_43
timestamp 18001
transform 1 0 5060 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 18001
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_66
timestamp 18001
transform 1 0 7176 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_84
timestamp 18001
transform 1 0 8832 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_92
timestamp 18001
transform 1 0 9568 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_113
timestamp 18001
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_142
timestamp 1636986456
transform 1 0 14168 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_154
timestamp 1636986456
transform 1 0 15272 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 18001
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636986456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 18001
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_187
timestamp 1636986456
transform 1 0 18308 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_199
timestamp 18001
transform 1 0 19412 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_234
timestamp 18001
transform 1 0 22632 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_242
timestamp 18001
transform 1 0 23368 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_250
timestamp 18001
transform 1 0 24104 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_267
timestamp 18001
transform 1 0 25668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_291
timestamp 18001
transform 1 0 27876 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_295
timestamp 18001
transform 1 0 28244 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_299
timestamp 1636986456
transform 1 0 28612 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 18001
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 18001
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_337
timestamp 18001
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_343
timestamp 18001
transform 1 0 32660 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_357
timestamp 18001
transform 1 0 33948 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_380
timestamp 18001
transform 1 0 36064 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 18001
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_35
timestamp 18001
transform 1 0 4324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_73
timestamp 18001
transform 1 0 7820 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 18001
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 18001
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_110
timestamp 1636986456
transform 1 0 11224 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 18001
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 18001
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_156
timestamp 18001
transform 1 0 15456 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_187
timestamp 18001
transform 1 0 18308 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 18001
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_209
timestamp 18001
transform 1 0 20332 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_226
timestamp 1636986456
transform 1 0 21896 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_268
timestamp 18001
transform 1 0 25760 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_274
timestamp 18001
transform 1 0 26312 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_300
timestamp 18001
transform 1 0 28704 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_328
timestamp 18001
transform 1 0 31280 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_339
timestamp 1636986456
transform 1 0 32292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_351
timestamp 18001
transform 1 0 33396 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_375
timestamp 18001
transform 1 0 35604 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 18001
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_11
timestamp 18001
transform 1 0 2116 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_23
timestamp 18001
transform 1 0 3220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 18001
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 18001
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 18001
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_71
timestamp 18001
transform 1 0 7636 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_82
timestamp 1636986456
transform 1 0 8648 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_94
timestamp 18001
transform 1 0 9752 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_98
timestamp 18001
transform 1 0 10120 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_107
timestamp 18001
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 18001
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_113
timestamp 18001
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_121
timestamp 18001
transform 1 0 12236 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_129
timestamp 1636986456
transform 1 0 12972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_141
timestamp 1636986456
transform 1 0 14076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_153
timestamp 1636986456
transform 1 0 15180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 18001
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_177
timestamp 18001
transform 1 0 17388 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_197
timestamp 18001
transform 1 0 19228 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_205
timestamp 18001
transform 1 0 19964 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_213
timestamp 18001
transform 1 0 20700 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 18001
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 18001
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636986456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_237
timestamp 18001
transform 1 0 22908 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_247
timestamp 18001
transform 1 0 23828 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_252
timestamp 18001
transform 1 0 24288 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_257
timestamp 1636986456
transform 1 0 24748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 18001
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 18001
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 18001
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_285
timestamp 18001
transform 1 0 27324 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_305
timestamp 18001
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_319
timestamp 18001
transform 1 0 30452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_331
timestamp 18001
transform 1 0 31556 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_355
timestamp 18001
transform 1 0 33764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_361
timestamp 18001
transform 1 0 34316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_372
timestamp 18001
transform 1 0 35328 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 18001
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_49
timestamp 18001
transform 1 0 5612 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_79
timestamp 18001
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 18001
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_115
timestamp 18001
transform 1 0 11684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 18001
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636986456
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1636986456
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_165
timestamp 18001
transform 1 0 16284 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_178
timestamp 18001
transform 1 0 17480 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_187
timestamp 18001
transform 1 0 18308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 18001
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_203
timestamp 18001
transform 1 0 19780 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_209
timestamp 18001
transform 1 0 20332 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 18001
transform 1 0 21620 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_235
timestamp 18001
transform 1 0 22724 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 18001
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 18001
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_253
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_295
timestamp 18001
transform 1 0 28244 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 18001
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1636986456
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1636986456
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_333
timestamp 18001
transform 1 0 31740 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_348
timestamp 18001
transform 1 0 33120 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_357
timestamp 18001
transform 1 0 33948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_379
timestamp 18001
transform 1 0 35972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_3
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_24
timestamp 18001
transform 1 0 3312 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_96
timestamp 18001
transform 1 0 9936 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 18001
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 18001
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_137
timestamp 18001
transform 1 0 13708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_157
timestamp 18001
transform 1 0 15548 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_179
timestamp 18001
transform 1 0 17572 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_191
timestamp 18001
transform 1 0 18676 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_199
timestamp 18001
transform 1 0 19412 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 18001
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_225
timestamp 18001
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_239
timestamp 18001
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_247
timestamp 18001
transform 1 0 23828 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_259
timestamp 18001
transform 1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_268
timestamp 18001
transform 1 0 25760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_300
timestamp 18001
transform 1 0 28704 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_325
timestamp 18001
transform 1 0 31004 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 18001
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_350
timestamp 18001
transform 1 0 33304 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 18001
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_11
timestamp 18001
transform 1 0 2116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 18001
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_33
timestamp 18001
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_51
timestamp 18001
transform 1 0 5796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_55
timestamp 18001
transform 1 0 6164 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_82
timestamp 18001
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_90
timestamp 18001
transform 1 0 9384 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_110
timestamp 1636986456
transform 1 0 11224 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_122
timestamp 18001
transform 1 0 12328 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_132
timestamp 18001
transform 1 0 13248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_141
timestamp 18001
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_149
timestamp 18001
transform 1 0 14812 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_158
timestamp 18001
transform 1 0 15640 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_166
timestamp 18001
transform 1 0 16376 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_172
timestamp 18001
transform 1 0 16928 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_176
timestamp 18001
transform 1 0 17296 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 18001
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1636986456
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_239
timestamp 1636986456
transform 1 0 23092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 18001
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_260
timestamp 18001
transform 1 0 25024 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_268
timestamp 18001
transform 1 0 25760 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_333
timestamp 18001
transform 1 0 31740 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_347
timestamp 1636986456
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_359
timestamp 18001
transform 1 0 34132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_371
timestamp 18001
transform 1 0 35236 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636986456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_27
timestamp 18001
transform 1 0 3588 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 18001
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 18001
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_80
timestamp 18001
transform 1 0 8464 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_89
timestamp 18001
transform 1 0 9292 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_98
timestamp 1636986456
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 18001
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1636986456
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1636986456
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1636986456
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1636986456
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 18001
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 18001
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1636986456
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 18001
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_189
timestamp 18001
transform 1 0 18492 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_213
timestamp 18001
transform 1 0 20700 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_221
timestamp 18001
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_225
timestamp 18001
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_233
timestamp 18001
transform 1 0 22540 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_248
timestamp 18001
transform 1 0 23920 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_271
timestamp 18001
transform 1 0 26036 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 18001
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 18001
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1636986456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1636986456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1636986456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_41
timestamp 18001
transform 1 0 4876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 18001
transform 1 0 9476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_98
timestamp 18001
transform 1 0 10120 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_106
timestamp 18001
transform 1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_112
timestamp 1636986456
transform 1 0 11408 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_124
timestamp 1636986456
transform 1 0 12512 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 18001
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_141
timestamp 18001
transform 1 0 14076 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_147
timestamp 1636986456
transform 1 0 14628 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_159
timestamp 18001
transform 1 0 15732 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_167
timestamp 18001
transform 1 0 16468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_178
timestamp 18001
transform 1 0 17480 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_185
timestamp 18001
transform 1 0 18124 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_193
timestamp 18001
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1636986456
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_209
timestamp 18001
transform 1 0 20332 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_220
timestamp 1636986456
transform 1 0 21344 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_232
timestamp 18001
transform 1 0 22448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 18001
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 18001
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 18001
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 18001
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_287
timestamp 18001
transform 1 0 27508 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_328
timestamp 1636986456
transform 1 0 31280 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_340
timestamp 18001
transform 1 0 32384 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 18001
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1636986456
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 18001
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_381
timestamp 18001
transform 1 0 36156 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1636986456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1636986456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_39
timestamp 18001
transform 1 0 4692 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_50
timestamp 18001
transform 1 0 5704 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_68
timestamp 18001
transform 1 0 7360 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_97
timestamp 18001
transform 1 0 10028 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 18001
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_120
timestamp 18001
transform 1 0 12144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_128
timestamp 18001
transform 1 0 12880 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 18001
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_194
timestamp 18001
transform 1 0 18952 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_203
timestamp 18001
transform 1 0 19780 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 18001
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_235
timestamp 18001
transform 1 0 22724 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_248
timestamp 18001
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_259
timestamp 18001
transform 1 0 24932 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_272
timestamp 18001
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 18001
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_346
timestamp 18001
transform 1 0 32936 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_363
timestamp 1636986456
transform 1 0 34500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_375
timestamp 18001
transform 1 0 35604 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_381
timestamp 18001
transform 1 0 36156 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1636986456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_52
timestamp 18001
transform 1 0 5888 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_56
timestamp 18001
transform 1 0 6256 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_63
timestamp 18001
transform 1 0 6900 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 18001
transform 1 0 8188 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 18001
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_97
timestamp 18001
transform 1 0 10028 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 18001
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_149
timestamp 18001
transform 1 0 14812 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_156
timestamp 18001
transform 1 0 15456 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_176
timestamp 18001
transform 1 0 17296 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_181
timestamp 18001
transform 1 0 17756 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 18001
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_211
timestamp 18001
transform 1 0 20516 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_222
timestamp 18001
transform 1 0 21528 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_227
timestamp 18001
transform 1 0 21988 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_264
timestamp 1636986456
transform 1 0 25392 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_276
timestamp 18001
transform 1 0 26496 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_284
timestamp 18001
transform 1 0 27232 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_294
timestamp 18001
transform 1 0 28152 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_373
timestamp 18001
transform 1 0 35420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_381
timestamp 18001
transform 1 0 36156 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636986456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636986456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1636986456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 18001
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 18001
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_80
timestamp 18001
transform 1 0 8464 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_93
timestamp 18001
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 18001
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_132
timestamp 1636986456
transform 1 0 13248 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_144
timestamp 18001
transform 1 0 14352 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 18001
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_173
timestamp 18001
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_184
timestamp 18001
transform 1 0 18032 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_206
timestamp 18001
transform 1 0 20056 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_210
timestamp 18001
transform 1 0 20424 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 18001
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 18001
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_239
timestamp 18001
transform 1 0 23092 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 18001
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 18001
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 18001
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_366
timestamp 1636986456
transform 1 0 34776 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_378
timestamp 18001
transform 1 0 35880 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636986456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1636986456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1636986456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_53
timestamp 18001
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_61
timestamp 18001
transform 1 0 6716 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_73
timestamp 18001
transform 1 0 7820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_81
timestamp 18001
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1636986456
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_97
timestamp 18001
transform 1 0 10028 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_113
timestamp 1636986456
transform 1 0 11500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_125
timestamp 18001
transform 1 0 12604 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 18001
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 18001
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_159
timestamp 1636986456
transform 1 0 15732 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_171
timestamp 18001
transform 1 0 16836 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_179
timestamp 18001
transform 1 0 17572 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 18001
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_197
timestamp 18001
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_205
timestamp 18001
transform 1 0 19964 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_228
timestamp 18001
transform 1 0 22080 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_265
timestamp 18001
transform 1 0 25484 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_289
timestamp 18001
transform 1 0 27692 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_297
timestamp 18001
transform 1 0 28428 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 18001
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_330
timestamp 1636986456
transform 1 0 31464 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_342
timestamp 1636986456
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 18001
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 18001
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1636986456
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_377
timestamp 18001
transform 1 0 35788 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_381
timestamp 18001
transform 1 0 36156 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1636986456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1636986456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1636986456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1636986456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 18001
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 18001
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_86
timestamp 18001
transform 1 0 9016 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_57_99
timestamp 18001
transform 1 0 10212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_107
timestamp 18001
transform 1 0 10948 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_144
timestamp 18001
transform 1 0 14352 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_150
timestamp 18001
transform 1 0 14904 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 18001
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 18001
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_169
timestamp 18001
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_174
timestamp 1636986456
transform 1 0 17112 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_186
timestamp 1636986456
transform 1 0 18216 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_198
timestamp 1636986456
transform 1 0 19320 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_210
timestamp 18001
transform 1 0 20424 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_214
timestamp 18001
transform 1 0 20792 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_230
timestamp 18001
transform 1 0 22264 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_265
timestamp 1636986456
transform 1 0 25484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 18001
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1636986456
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1636986456
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1636986456
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1636986456
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 18001
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 18001
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1636986456
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1636986456
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1636986456
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_373
timestamp 18001
transform 1 0 35420 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_381
timestamp 18001
transform 1 0 36156 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636986456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1636986456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_53
timestamp 18001
transform 1 0 5980 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 18001
transform 1 0 9292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_101
timestamp 18001
transform 1 0 10396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_105
timestamp 18001
transform 1 0 10764 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_114
timestamp 18001
transform 1 0 11592 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_120
timestamp 1636986456
transform 1 0 12144 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 18001
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_141
timestamp 18001
transform 1 0 14076 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_184
timestamp 18001
transform 1 0 18032 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_220
timestamp 18001
transform 1 0 21344 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_228
timestamp 18001
transform 1 0 22080 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_232
timestamp 18001
transform 1 0 22448 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_240
timestamp 18001
transform 1 0 23184 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1636986456
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_265
timestamp 18001
transform 1 0 25484 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1636986456
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 18001
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 18001
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1636986456
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1636986456
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1636986456
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1636986456
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_377
timestamp 18001
transform 1 0 35788 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_381
timestamp 18001
transform 1 0 36156 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636986456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1636986456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1636986456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 18001
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 18001
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_66
timestamp 18001
transform 1 0 7176 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_74
timestamp 18001
transform 1 0 7912 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_100
timestamp 1636986456
transform 1 0 10304 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_130
timestamp 1636986456
transform 1 0 13064 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_142
timestamp 18001
transform 1 0 14168 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 18001
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 18001
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_169
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_173
timestamp 18001
transform 1 0 17020 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_177
timestamp 18001
transform 1 0 17388 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_185
timestamp 18001
transform 1 0 18124 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_198
timestamp 1636986456
transform 1 0 19320 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_210
timestamp 1636986456
transform 1 0 20424 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 18001
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_235
timestamp 18001
transform 1 0 22724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_239
timestamp 18001
transform 1 0 23092 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_246
timestamp 1636986456
transform 1 0 23736 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_258
timestamp 18001
transform 1 0 24840 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1636986456
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1636986456
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1636986456
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1636986456
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 18001
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 18001
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1636986456
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1636986456
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1636986456
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_373
timestamp 18001
transform 1 0 35420 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_381
timestamp 18001
transform 1 0 36156 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1636986456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1636986456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_73
timestamp 18001
transform 1 0 7820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_81
timestamp 18001
transform 1 0 8556 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_85
timestamp 18001
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_91
timestamp 18001
transform 1 0 9476 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_99
timestamp 18001
transform 1 0 10212 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_107
timestamp 18001
transform 1 0 10948 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_116
timestamp 18001
transform 1 0 11776 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_120
timestamp 18001
transform 1 0 12144 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 18001
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_147
timestamp 1636986456
transform 1 0 14628 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_159
timestamp 18001
transform 1 0 15732 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_174
timestamp 18001
transform 1 0 17112 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 18001
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 18001
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 18001
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_208
timestamp 1636986456
transform 1 0 20240 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_220
timestamp 18001
transform 1 0 21344 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_227
timestamp 18001
transform 1 0 21988 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_240
timestamp 1636986456
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_267
timestamp 18001
transform 1 0 25668 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_283
timestamp 1636986456
transform 1 0 27140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_295
timestamp 1636986456
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 18001
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1636986456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1636986456
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1636986456
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1636986456
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 18001
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_377
timestamp 18001
transform 1 0 35788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_381
timestamp 18001
transform 1 0 36156 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636986456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636986456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1636986456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1636986456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 18001
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 18001
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_80
timestamp 18001
transform 1 0 8464 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1636986456
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 18001
transform 1 0 11500 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_121
timestamp 18001
transform 1 0 12236 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_127
timestamp 18001
transform 1 0 12788 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_148
timestamp 18001
transform 1 0 14720 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 18001
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_178
timestamp 18001
transform 1 0 17480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_186
timestamp 18001
transform 1 0 18216 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_197
timestamp 18001
transform 1 0 19228 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_216
timestamp 18001
transform 1 0 20976 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 18001
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1636986456
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1636986456
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1636986456
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1636986456
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 18001
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 18001
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_373
timestamp 18001
transform 1 0 35420 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_381
timestamp 18001
transform 1 0 36156 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1636986456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1636986456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1636986456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_53
timestamp 18001
transform 1 0 5980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_57
timestamp 18001
transform 1 0 6348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_81
timestamp 18001
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_94
timestamp 18001
transform 1 0 9752 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_123
timestamp 18001
transform 1 0 12420 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_129
timestamp 18001
transform 1 0 12972 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_137
timestamp 18001
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 18001
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_173
timestamp 18001
transform 1 0 17020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_177
timestamp 18001
transform 1 0 17388 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_186
timestamp 18001
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 18001
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_214
timestamp 18001
transform 1 0 20792 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_243
timestamp 18001
transform 1 0 23460 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_62_258
timestamp 18001
transform 1 0 24840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_270
timestamp 18001
transform 1 0 25944 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1636986456
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1636986456
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 18001
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 18001
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1636986456
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1636986456
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1636986456
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1636986456
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 18001
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1636986456
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_377
timestamp 18001
transform 1 0 35788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_381
timestamp 18001
transform 1 0 36156 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_27
timestamp 18001
transform 1 0 3588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 18001
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_106
timestamp 18001
transform 1 0 10856 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_113
timestamp 18001
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_137
timestamp 18001
transform 1 0 13708 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 18001
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 18001
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 18001
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_180
timestamp 18001
transform 1 0 17664 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 18001
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_233
timestamp 18001
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1636986456
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1636986456
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1636986456
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1636986456
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 18001
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 18001
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1636986456
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1636986456
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1636986456
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_373
timestamp 18001
transform 1 0 35420 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_381
timestamp 18001
transform 1 0 36156 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1636986456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1636986456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1636986456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 18001
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_66
timestamp 18001
transform 1 0 7176 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_78
timestamp 18001
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_85
timestamp 18001
transform 1 0 8924 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_91
timestamp 18001
transform 1 0 9476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_101
timestamp 18001
transform 1 0 10396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_113
timestamp 18001
transform 1 0 11500 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_119
timestamp 18001
transform 1 0 12052 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_129
timestamp 18001
transform 1 0 12972 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 18001
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1636986456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1636986456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 18001
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_169
timestamp 18001
transform 1 0 16652 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_179
timestamp 1636986456
transform 1 0 17572 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_191
timestamp 18001
transform 1 0 18676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 18001
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1636986456
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1636986456
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 18001
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1636986456
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1636986456
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 18001
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1636986456
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1636986456
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 18001
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1636986456
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1636986456
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 18001
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1636986456
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1636986456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 18001
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_337
timestamp 1636986456
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_349
timestamp 1636986456
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 18001
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1636986456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_377
timestamp 18001
transform 1 0 35788 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_381
timestamp 18001
transform 1 0 36156 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform -1 0 19964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform -1 0 17756 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 35420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform -1 0 26588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform -1 0 26956 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform -1 0 13984 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 15364 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 18001
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 18001
transform -1 0 4324 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 18001
transform -1 0 11408 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 18001
transform -1 0 18860 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 18001
transform -1 0 18860 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 18001
transform -1 0 8924 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 18001
transform -1 0 12696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 18001
transform -1 0 16468 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 18001
transform -1 0 4692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 18001
transform -1 0 16652 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 18001
transform -1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 18001
transform 1 0 12144 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 18001
transform -1 0 8188 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 18001
transform -1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 18001
transform -1 0 13984 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 18001
transform -1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 18001
transform -1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 18001
transform -1 0 3496 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 18001
transform -1 0 4048 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 18001
transform 1 0 3772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 18001
transform 1 0 27416 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 18001
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 18001
transform -1 0 3680 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 18001
transform -1 0 6164 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 18001
transform -1 0 9660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 18001
transform -1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 18001
transform -1 0 7360 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 18001
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 18001
transform -1 0 9016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 18001
transform -1 0 18492 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 18001
transform -1 0 6256 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 18001
transform -1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 18001
transform -1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 18001
transform 1 0 5060 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 18001
transform -1 0 5796 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 18001
transform -1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 18001
transform -1 0 5888 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 18001
transform -1 0 29348 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 18001
transform -1 0 7820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 18001
transform -1 0 34776 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 18001
transform 1 0 19872 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 18001
transform -1 0 19964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 18001
transform 1 0 12512 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 18001
transform -1 0 5428 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 18001
transform -1 0 11040 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 18001
transform -1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 18001
transform -1 0 35696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 18001
transform -1 0 35788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 18001
transform -1 0 36248 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 18001
transform -1 0 36248 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 18001
transform -1 0 36248 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 18001
transform -1 0 36248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 18001
transform -1 0 36248 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 18001
transform -1 0 36248 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 18001
transform -1 0 36248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 18001
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 18001
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 18001
transform 1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 18001
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 18001
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 18001
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 18001
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 18001
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 18001
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 36524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 36524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 36524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 36524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 36524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 36524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 36524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 36524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 36524 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 36524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 36524 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 36524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 36524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 36524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 36524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 36524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 36524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 36524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 36524 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 36524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 36524 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 36524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 36524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 36524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 36524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 36524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 36524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 36524 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 36524 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 36524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 36524 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 36524 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 36524 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 36524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 36524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 36524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 36524 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 36524 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 36524 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 36524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 36524 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 36524 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 36524 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 36524 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 36524 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 36524 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 36524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 36524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 36524 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 36524 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 36524 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 36524 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 36524 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 36524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 36524 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 36524 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 36524 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 36524 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 36524 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 36524 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 36524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 36524 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_143
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_144
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_145
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_146
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_147
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_148
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_149
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_150
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_151
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_152
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_153
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_154
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_155
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_156
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_157
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_158
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_159
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_160
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_161
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_162
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_163
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_164
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_165
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_168
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_169
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_170
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_171
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_172
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_173
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_174
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_175
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_176
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_177
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_178
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_179
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_180
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_181
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_182
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_183
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_184
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_185
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_186
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_187
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_188
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_189
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_190
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_191
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_192
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_193
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_194
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_195
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_196
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_197
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_198
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_199
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_200
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_201
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_202
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_203
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_204
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_205
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_206
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_207
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_208
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_209
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_210
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_211
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_212
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_213
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_214
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_215
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_216
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_217
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_218
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_219
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_220
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_221
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_222
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_223
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_224
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_225
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_226
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_227
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_228
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_229
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_230
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_231
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_232
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_233
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_234
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_235
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_236
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_237
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_238
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_239
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_240
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_241
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_242
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_243
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_244
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_245
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_246
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_247
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_248
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_249
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_250
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_251
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_252
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_253
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_254
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_255
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_256
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_257
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_258
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_259
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_260
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_261
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_262
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_263
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_264
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_265
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_266
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_267
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_268
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_269
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_270
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_271
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_272
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_273
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_274
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_275
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_276
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_277
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_278
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_279
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_280
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_281
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_282
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_283
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_284
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_285
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_286
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_287
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_288
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_289
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_290
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_291
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_292
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_293
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_294
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_295
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_296
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_297
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_298
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_299
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_300
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_301
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_302
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_303
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_304
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_305
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_306
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_307
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_308
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_309
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_310
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_311
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_312
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_313
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_314
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_315
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_316
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_317
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_318
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_319
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_320
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_321
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_322
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_323
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_324
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_325
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_326
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_327
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_328
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_329
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_330
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_331
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_332
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_333
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_334
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_335
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_336
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_337
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_338
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_339
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_340
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_341
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_342
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_343
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_344
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_345
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_346
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_347
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_348
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_349
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_350
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_351
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_352
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_353
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_354
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_355
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_356
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_357
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_358
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_359
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_360
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_361
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_362
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_363
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_364
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_365
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_366
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_367
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_368
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_369
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_370
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_371
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_372
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_373
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_374
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_375
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_376
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_377
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_378
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_379
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_380
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_381
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_382
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_383
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_384
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_385
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_386
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_387
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_388
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_389
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_390
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_391
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_392
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_393
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_394
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_395
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_396
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_397
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_398
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_399
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_400
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_401
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_402
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_403
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_404
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_405
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_406
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_407
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_408
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_409
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_410
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_411
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_412
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_413
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_414
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_415
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_416
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_417
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_418
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_419
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_420
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_421
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_422
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_423
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_424
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_425
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_426
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_427
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_428
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_429
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_430
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_431
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_432
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_433
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_434
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_435
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_436
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_437
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_438
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_439
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_440
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_441
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_442
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_443
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_444
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_445
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_446
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_447
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_448
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_449
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_450
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_451
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_452
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_453
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_454
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_455
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_456
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_457
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_458
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_459
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_460
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_461
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_462
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_463
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_464
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_465
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_466
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_467
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_468
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_469
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_470
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_471
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_472
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_473
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_474
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_475
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_476
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_477
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_478
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_479
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_480
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_481
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_482
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_483
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_484
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_485
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_486
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_487
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_488
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_489
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_490
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_491
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_492
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_493
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_494
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_495
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_496
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_497
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_498
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_499
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_500
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_501
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_502
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_503
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_504
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_505
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_506
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_507
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_508
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_509
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_510
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_511
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_512
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_513
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_514
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_515
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_516
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_517
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_518
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_519
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_520
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_521
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_522
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_523
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_524
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_525
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_526
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_527
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_528
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_529
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_530
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_531
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_532
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_533
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_534
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_535
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_536
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_537
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_538
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_539
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_540
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_541
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_542
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_543
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_544
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_545
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_546
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_547
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_548
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_549
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_550
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_551
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_552
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_553
timestamp 18001
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_554
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_555
timestamp 18001
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_556
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_557
timestamp 18001
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_558
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_559
timestamp 18001
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_560
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_561
timestamp 18001
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_562
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_563
timestamp 18001
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_564
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 cs
port 3 nsew signal input
flabel metal3 s 36895 23808 37695 23928 0 FreeSans 480 0 0 0 dataBusIn[0]
port 4 nsew signal input
flabel metal3 s 36895 25168 37695 25288 0 FreeSans 480 0 0 0 dataBusIn[1]
port 5 nsew signal input
flabel metal3 s 36895 26528 37695 26648 0 FreeSans 480 0 0 0 dataBusIn[2]
port 6 nsew signal input
flabel metal3 s 36895 27208 37695 27328 0 FreeSans 480 0 0 0 dataBusIn[3]
port 7 nsew signal input
flabel metal3 s 36895 22448 37695 22568 0 FreeSans 480 0 0 0 dataBusIn[4]
port 8 nsew signal input
flabel metal3 s 36895 23128 37695 23248 0 FreeSans 480 0 0 0 dataBusIn[5]
port 9 nsew signal input
flabel metal3 s 36895 25848 37695 25968 0 FreeSans 480 0 0 0 dataBusIn[6]
port 10 nsew signal input
flabel metal3 s 36895 24488 37695 24608 0 FreeSans 480 0 0 0 dataBusIn[7]
port 11 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 dataBusOut[0]
port 12 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 dataBusOut[1]
port 13 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 dataBusOut[2]
port 14 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 dataBusOut[3]
port 15 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 dataBusOut[4]
port 16 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 dataBusOut[5]
port 17 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 dataBusOut[6]
port 18 nsew signal output
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 dataBusOut[7]
port 19 nsew signal output
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 dataBusSelect
port 20 nsew signal output
flabel metal2 s 12898 39039 12954 39839 0 FreeSans 224 90 0 0 gpio[0]
port 21 nsew signal bidirectional
flabel metal2 s 12254 39039 12310 39839 0 FreeSans 224 90 0 0 gpio[10]
port 22 nsew signal bidirectional
flabel metal2 s 8390 39039 8446 39839 0 FreeSans 224 90 0 0 gpio[11]
port 23 nsew signal bidirectional
flabel metal2 s 10966 39039 11022 39839 0 FreeSans 224 90 0 0 gpio[12]
port 24 nsew signal bidirectional
flabel metal2 s 9678 39039 9734 39839 0 FreeSans 224 90 0 0 gpio[13]
port 25 nsew signal bidirectional
flabel metal2 s 5814 39039 5870 39839 0 FreeSans 224 90 0 0 gpio[14]
port 26 nsew signal bidirectional
flabel metal2 s 6458 39039 6514 39839 0 FreeSans 224 90 0 0 gpio[15]
port 27 nsew signal bidirectional
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 gpio[16]
port 28 nsew signal bidirectional
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 gpio[17]
port 29 nsew signal bidirectional
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 gpio[18]
port 30 nsew signal bidirectional
flabel metal3 s 36895 21088 37695 21208 0 FreeSans 480 0 0 0 gpio[19]
port 31 nsew signal bidirectional
flabel metal2 s 9034 39039 9090 39839 0 FreeSans 224 90 0 0 gpio[1]
port 32 nsew signal bidirectional
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio[20]
port 33 nsew signal bidirectional
flabel metal3 s 36895 20408 37695 20528 0 FreeSans 480 0 0 0 gpio[21]
port 34 nsew signal bidirectional
flabel metal3 s 36895 21768 37695 21888 0 FreeSans 480 0 0 0 gpio[22]
port 35 nsew signal bidirectional
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpio[23]
port 36 nsew signal bidirectional
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpio[24]
port 37 nsew signal bidirectional
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio[25]
port 38 nsew signal bidirectional
flabel metal2 s 21270 39039 21326 39839 0 FreeSans 224 90 0 0 gpio[2]
port 39 nsew signal bidirectional
flabel metal2 s 10322 39039 10378 39839 0 FreeSans 224 90 0 0 gpio[3]
port 40 nsew signal bidirectional
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 gpio[4]
port 41 nsew signal bidirectional
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 gpio[5]
port 42 nsew signal bidirectional
flabel metal2 s 7746 39039 7802 39839 0 FreeSans 224 90 0 0 gpio[6]
port 43 nsew signal bidirectional
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 gpio[7]
port 44 nsew signal bidirectional
flabel metal2 s 11610 39039 11666 39839 0 FreeSans 224 90 0 0 gpio[8]
port 45 nsew signal bidirectional
flabel metal2 s 7102 39039 7158 39839 0 FreeSans 224 90 0 0 gpio[9]
port 46 nsew signal bidirectional
flabel metal3 s 36895 3408 37695 3528 0 FreeSans 480 0 0 0 nrst
port 47 nsew signal input
rlabel metal1 18814 36992 18814 36992 0 VGND
rlabel metal1 18814 37536 18814 37536 0 VPWR
rlabel metal1 32430 31450 32430 31450 0 _0000_
rlabel metal1 27646 29274 27646 29274 0 _0001_
rlabel metal1 27370 31994 27370 31994 0 _0002_
rlabel metal2 29394 29988 29394 29988 0 _0003_
rlabel metal1 34362 30158 34362 30158 0 _0004_
rlabel metal1 31740 31858 31740 31858 0 _0005_
rlabel metal1 29716 32334 29716 32334 0 _0006_
rlabel metal1 33028 30294 33028 30294 0 _0007_
rlabel metal1 28296 27642 28296 27642 0 _0008_
rlabel metal1 34592 24378 34592 24378 0 _0009_
rlabel metal1 34730 27642 34730 27642 0 _0010_
rlabel metal1 33258 31858 33258 31858 0 _0011_
rlabel metal1 30084 29818 30084 29818 0 _0012_
rlabel metal2 27370 25500 27370 25500 0 _0013_
rlabel metal2 20378 4964 20378 4964 0 _0014_
rlabel metal2 23598 4794 23598 4794 0 _0015_
rlabel metal1 24932 5134 24932 5134 0 _0016_
rlabel metal2 25346 5100 25346 5100 0 _0017_
rlabel metal2 22126 5338 22126 5338 0 _0018_
rlabel metal1 22356 4522 22356 4522 0 _0019_
rlabel metal2 32430 8330 32430 8330 0 _0020_
rlabel metal1 32614 6222 32614 6222 0 _0021_
rlabel metal1 33948 7446 33948 7446 0 _0022_
rlabel metal1 32561 6970 32561 6970 0 _0023_
rlabel metal3 31257 15300 31257 15300 0 _0024_
rlabel metal3 32361 19380 32361 19380 0 _0025_
rlabel metal2 14674 20196 14674 20196 0 _0026_
rlabel metal1 14582 18394 14582 18394 0 _0027_
rlabel metal2 25990 30940 25990 30940 0 _0028_
rlabel metal2 16514 4828 16514 4828 0 _0029_
rlabel metal2 14122 5406 14122 5406 0 _0030_
rlabel metal2 17618 6494 17618 6494 0 _0031_
rlabel metal1 18216 3910 18216 3910 0 _0032_
rlabel metal2 19918 4420 19918 4420 0 _0033_
rlabel metal2 14674 4760 14674 4760 0 _0034_
rlabel metal2 11546 4760 11546 4760 0 _0035_
rlabel metal1 15548 3434 15548 3434 0 _0036_
rlabel metal1 11822 3162 11822 3162 0 _0037_
rlabel metal2 9890 3230 9890 3230 0 _0038_
rlabel metal1 11217 5882 11217 5882 0 _0039_
rlabel metal1 14398 4046 14398 4046 0 _0040_
rlabel metal1 13340 3094 13340 3094 0 _0041_
rlabel via2 19366 33813 19366 33813 0 _0042_
rlabel metal2 20010 36516 20010 36516 0 _0043_
rlabel metal1 14444 35258 14444 35258 0 _0044_
rlabel metal1 15226 35802 15226 35802 0 _0045_
rlabel metal1 22816 35802 22816 35802 0 _0046_
rlabel metal2 23230 36244 23230 36244 0 _0047_
rlabel metal1 25208 36346 25208 36346 0 _0048_
rlabel metal2 26082 34204 26082 34204 0 _0049_
rlabel metal1 4692 24378 4692 24378 0 _0050_
rlabel metal2 7314 24548 7314 24548 0 _0051_
rlabel metal2 6118 28764 6118 28764 0 _0052_
rlabel metal1 4048 29206 4048 29206 0 _0053_
rlabel metal1 6440 27098 6440 27098 0 _0054_
rlabel metal1 6762 25466 6762 25466 0 _0055_
rlabel metal2 4830 26724 4830 26724 0 _0056_
rlabel metal2 5290 28798 5290 28798 0 _0057_
rlabel via1 1695 22202 1695 22202 0 _0058_
rlabel metal1 7130 23188 7130 23188 0 _0059_
rlabel metal1 6670 18836 6670 18836 0 _0060_
rlabel metal2 1702 20332 1702 20332 0 _0061_
rlabel metal1 1794 21624 1794 21624 0 _0062_
rlabel metal2 1702 23324 1702 23324 0 _0063_
rlabel metal1 3450 23290 3450 23290 0 _0064_
rlabel metal1 3450 20332 3450 20332 0 _0065_
rlabel metal2 24978 29988 24978 29988 0 _0066_
rlabel metal2 10626 36652 10626 36652 0 _0067_
rlabel metal2 7038 35428 7038 35428 0 _0068_
rlabel metal2 11914 36958 11914 36958 0 _0069_
rlabel metal2 7498 36652 7498 36652 0 _0070_
rlabel metal2 9062 36890 9062 36890 0 _0071_
rlabel metal1 7958 36346 7958 36346 0 _0072_
rlabel metal2 4462 36958 4462 36958 0 _0073_
rlabel metal1 5934 34714 5934 34714 0 _0074_
rlabel metal1 26358 32538 26358 32538 0 _0075_
rlabel metal1 23552 33558 23552 33558 0 _0076_
rlabel metal2 20562 32674 20562 32674 0 _0077_
rlabel metal1 18577 32198 18577 32198 0 _0078_
rlabel metal1 17940 32198 17940 32198 0 _0079_
rlabel metal2 14582 31076 14582 31076 0 _0080_
rlabel metal2 12558 32096 12558 32096 0 _0081_
rlabel metal1 15732 34034 15732 34034 0 _0082_
rlabel metal1 3266 24820 3266 24820 0 _0083_
rlabel metal1 8878 18938 8878 18938 0 _0084_
rlabel metal1 6486 29818 6486 29818 0 _0085_
rlabel metal2 1794 29342 1794 29342 0 _0086_
rlabel metal1 1978 27098 1978 27098 0 _0087_
rlabel metal2 2254 25636 2254 25636 0 _0088_
rlabel metal2 3910 25636 3910 25636 0 _0089_
rlabel metal1 2070 28186 2070 28186 0 _0090_
rlabel metal1 13754 33082 13754 33082 0 _0091_
rlabel metal1 7958 33626 7958 33626 0 _0092_
rlabel metal2 18814 30056 18814 30056 0 _0093_
rlabel metal2 7130 32164 7130 32164 0 _0094_
rlabel metal1 5520 30294 5520 30294 0 _0095_
rlabel metal1 6670 31926 6670 31926 0 _0096_
rlabel metal2 7038 33252 7038 33252 0 _0097_
rlabel metal2 5566 32028 5566 32028 0 _0098_
rlabel metal1 6026 15674 6026 15674 0 _0099_
rlabel metal1 3726 14586 3726 14586 0 _0100_
rlabel metal1 6348 16218 6348 16218 0 _0101_
rlabel metal1 3397 13702 3397 13702 0 _0102_
rlabel metal1 3174 11832 3174 11832 0 _0103_
rlabel metal1 5658 9486 5658 9486 0 _0104_
rlabel metal1 5198 8602 5198 8602 0 _0105_
rlabel metal1 8050 9928 8050 9928 0 _0106_
rlabel metal1 2162 18632 2162 18632 0 _0107_
rlabel metal1 7498 17850 7498 17850 0 _0108_
rlabel metal2 5842 17884 5842 17884 0 _0109_
rlabel metal2 3726 18462 3726 18462 0 _0110_
rlabel metal2 1702 16558 1702 16558 0 _0111_
rlabel metal1 1932 17850 1932 17850 0 _0112_
rlabel metal1 4508 16762 4508 16762 0 _0113_
rlabel metal2 2714 16694 2714 16694 0 _0114_
rlabel metal2 13662 20060 13662 20060 0 _0115_
rlabel metal1 29808 30906 29808 30906 0 _0116_
rlabel metal2 13386 8670 13386 8670 0 _0117_
rlabel metal1 14168 26350 14168 26350 0 _0118_
rlabel metal1 15088 26486 15088 26486 0 _0119_
rlabel via1 10626 26214 10626 26214 0 _0120_
rlabel metal2 11086 21692 11086 21692 0 _0121_
rlabel metal1 2392 23630 2392 23630 0 _0122_
rlabel metal2 8694 14926 8694 14926 0 _0123_
rlabel metal1 10994 16660 10994 16660 0 _0124_
rlabel metal1 8694 26384 8694 26384 0 _0125_
rlabel metal1 7912 26554 7912 26554 0 _0126_
rlabel metal2 6578 32164 6578 32164 0 _0127_
rlabel metal1 10902 32232 10902 32232 0 _0128_
rlabel metal1 10074 16762 10074 16762 0 _0129_
rlabel metal1 9154 12920 9154 12920 0 _0130_
rlabel metal1 8602 10608 8602 10608 0 _0131_
rlabel metal1 9430 12138 9430 12138 0 _0132_
rlabel metal1 8878 11526 8878 11526 0 _0133_
rlabel metal2 5244 27302 5244 27302 0 _0134_
rlabel metal1 4692 22202 4692 22202 0 _0135_
rlabel metal1 4830 22644 4830 22644 0 _0136_
rlabel metal1 7590 22440 7590 22440 0 _0137_
rlabel metal1 11730 27438 11730 27438 0 _0138_
rlabel metal1 10580 26826 10580 26826 0 _0139_
rlabel metal1 17250 27438 17250 27438 0 _0140_
rlabel metal1 13064 27642 13064 27642 0 _0141_
rlabel metal1 17848 23698 17848 23698 0 _0142_
rlabel metal1 17204 23834 17204 23834 0 _0143_
rlabel metal1 16514 27540 16514 27540 0 _0144_
rlabel via1 11362 21521 11362 21521 0 _0145_
rlabel metal1 11500 21454 11500 21454 0 _0146_
rlabel metal1 8464 16082 8464 16082 0 _0147_
rlabel metal1 8418 15470 8418 15470 0 _0148_
rlabel metal1 11040 18802 11040 18802 0 _0149_
rlabel metal1 10028 18394 10028 18394 0 _0150_
rlabel metal1 8694 26554 8694 26554 0 _0151_
rlabel metal2 8970 27846 8970 27846 0 _0152_
rlabel metal1 8464 31858 8464 31858 0 _0153_
rlabel metal1 8234 30124 8234 30124 0 _0154_
rlabel metal1 9660 18326 9660 18326 0 _0155_
rlabel metal2 8142 14671 8142 14671 0 _0156_
rlabel metal1 7820 12138 7820 12138 0 _0157_
rlabel metal1 8556 12886 8556 12886 0 _0158_
rlabel metal1 8142 12750 8142 12750 0 _0159_
rlabel metal1 4876 20434 4876 20434 0 _0160_
rlabel metal1 5152 20434 5152 20434 0 _0161_
rlabel metal1 5474 20570 5474 20570 0 _0162_
rlabel metal1 10580 20978 10580 20978 0 _0163_
rlabel metal1 11086 29716 11086 29716 0 _0164_
rlabel metal1 9982 28186 9982 28186 0 _0165_
rlabel metal1 15318 29172 15318 29172 0 _0166_
rlabel metal1 14950 29002 14950 29002 0 _0167_
rlabel metal2 15410 28322 15410 28322 0 _0168_
rlabel metal1 9844 28390 9844 28390 0 _0169_
rlabel metal2 11178 21420 11178 21420 0 _0170_
rlabel metal1 3266 20774 3266 20774 0 _0171_
rlabel metal2 9246 15708 9246 15708 0 _0172_
rlabel metal1 11132 20774 11132 20774 0 _0173_
rlabel metal2 15962 28832 15962 28832 0 _0174_
rlabel metal1 8372 28730 8372 28730 0 _0175_
rlabel metal1 8188 31790 8188 31790 0 _0176_
rlabel metal1 8832 17306 8832 17306 0 _0177_
rlabel metal1 9660 17034 9660 17034 0 _0178_
rlabel metal2 8602 16762 8602 16762 0 _0179_
rlabel metal2 7774 15980 7774 15980 0 _0180_
rlabel metal1 11362 29138 11362 29138 0 _0181_
rlabel metal2 7774 20502 7774 20502 0 _0182_
rlabel metal2 7222 20604 7222 20604 0 _0183_
rlabel metal1 7360 20978 7360 20978 0 _0184_
rlabel metal1 11454 21012 11454 21012 0 _0185_
rlabel metal1 7728 20774 7728 20774 0 _0186_
rlabel metal1 10718 28628 10718 28628 0 _0187_
rlabel metal1 17388 28050 17388 28050 0 _0188_
rlabel metal2 12190 28764 12190 28764 0 _0189_
rlabel metal2 12282 28356 12282 28356 0 _0190_
rlabel metal1 11638 20774 11638 20774 0 _0191_
rlabel metal1 9844 16558 9844 16558 0 _0192_
rlabel metal2 9982 15946 9982 15946 0 _0193_
rlabel metal2 15870 7123 15870 7123 0 _0194_
rlabel metal2 10902 18496 10902 18496 0 _0195_
rlabel viali 8596 29138 8596 29138 0 _0196_
rlabel metal1 17894 30260 17894 30260 0 _0197_
rlabel metal2 17710 28900 17710 28900 0 _0198_
rlabel metal1 17986 30328 17986 30328 0 _0199_
rlabel metal2 10166 16762 10166 16762 0 _0200_
rlabel metal1 9338 13906 9338 13906 0 _0201_
rlabel metal1 13110 23664 13110 23664 0 _0202_
rlabel metal2 13202 23868 13202 23868 0 _0203_
rlabel metal1 13432 23562 13432 23562 0 _0204_
rlabel metal1 11960 19822 11960 19822 0 _0205_
rlabel metal1 7682 20570 7682 20570 0 _0206_
rlabel metal2 7682 22236 7682 22236 0 _0207_
rlabel metal1 8372 23562 8372 23562 0 _0208_
rlabel metal2 7958 21760 7958 21760 0 _0209_
rlabel metal2 12006 24412 12006 24412 0 _0210_
rlabel metal2 11914 23868 11914 23868 0 _0211_
rlabel metal1 9016 18598 9016 18598 0 _0212_
rlabel metal1 11684 16558 11684 16558 0 _0213_
rlabel metal1 18354 28730 18354 28730 0 _0214_
rlabel metal2 18170 28611 18170 28611 0 _0215_
rlabel metal2 17986 29444 17986 29444 0 _0216_
rlabel metal2 11224 32980 11224 32980 0 _0217_
rlabel metal1 11178 16558 11178 16558 0 _0218_
rlabel metal2 11454 19618 11454 19618 0 _0219_
rlabel metal1 12282 7412 12282 7412 0 _0220_
rlabel metal2 12006 18428 12006 18428 0 _0221_
rlabel metal1 11500 16558 11500 16558 0 _0222_
rlabel metal1 10534 15504 10534 15504 0 _0223_
rlabel metal1 10718 13906 10718 13906 0 _0224_
rlabel metal1 15640 24786 15640 24786 0 _0225_
rlabel metal1 15870 24310 15870 24310 0 _0226_
rlabel metal2 12926 24378 12926 24378 0 _0227_
rlabel metal1 11362 25262 11362 25262 0 _0228_
rlabel metal1 5704 21862 5704 21862 0 _0229_
rlabel metal2 5658 23868 5658 23868 0 _0230_
rlabel metal1 5750 20026 5750 20026 0 _0231_
rlabel metal2 12558 22678 12558 22678 0 _0232_
rlabel metal2 16330 26044 16330 26044 0 _0233_
rlabel metal1 16330 25772 16330 25772 0 _0234_
rlabel metal2 12098 25755 12098 25755 0 _0235_
rlabel metal1 12052 24922 12052 24922 0 _0236_
rlabel metal1 12696 16082 12696 16082 0 _0237_
rlabel metal1 12696 17102 12696 17102 0 _0238_
rlabel metal1 12236 15946 12236 15946 0 _0239_
rlabel metal1 13110 16558 13110 16558 0 _0240_
rlabel metal2 16882 25143 16882 25143 0 _0241_
rlabel metal1 17388 25466 17388 25466 0 _0242_
rlabel metal1 17618 23290 17618 23290 0 _0243_
rlabel metal2 17434 25024 17434 25024 0 _0244_
rlabel metal1 13018 17680 13018 17680 0 _0245_
rlabel metal1 12788 16218 12788 16218 0 _0246_
rlabel metal2 12558 17034 12558 17034 0 _0247_
rlabel metal2 13018 15674 13018 15674 0 _0248_
rlabel metal2 12926 16116 12926 16116 0 _0249_
rlabel metal2 18768 17646 18768 17646 0 _0250_
rlabel metal1 18078 15130 18078 15130 0 _0251_
rlabel metal2 17986 17340 17986 17340 0 _0252_
rlabel metal1 19826 11186 19826 11186 0 _0253_
rlabel metal2 19274 11407 19274 11407 0 _0254_
rlabel metal2 18906 17697 18906 17697 0 _0255_
rlabel metal1 19090 17680 19090 17680 0 _0256_
rlabel metal2 13662 17119 13662 17119 0 _0257_
rlabel metal2 13478 16524 13478 16524 0 _0258_
rlabel metal1 13110 14314 13110 14314 0 _0259_
rlabel metal1 12604 14586 12604 14586 0 _0260_
rlabel metal2 11362 14246 11362 14246 0 _0261_
rlabel metal1 10765 14994 10765 14994 0 _0262_
rlabel metal2 10902 14858 10902 14858 0 _0263_
rlabel metal2 9798 14212 9798 14212 0 _0264_
rlabel metal1 8970 15028 8970 15028 0 _0265_
rlabel metal1 9108 14450 9108 14450 0 _0266_
rlabel metal1 7498 13872 7498 13872 0 _0267_
rlabel metal1 8188 15606 8188 15606 0 _0268_
rlabel metal1 8326 15334 8326 15334 0 _0269_
rlabel metal1 5750 12818 5750 12818 0 _0270_
rlabel metal1 5934 11628 5934 11628 0 _0271_
rlabel metal2 6578 11356 6578 11356 0 _0272_
rlabel metal1 10718 10064 10718 10064 0 _0273_
rlabel metal1 11500 9554 11500 9554 0 _0274_
rlabel metal2 11914 10846 11914 10846 0 _0275_
rlabel metal2 15686 14688 15686 14688 0 _0276_
rlabel metal1 15686 13736 15686 13736 0 _0277_
rlabel metal1 15502 13906 15502 13906 0 _0278_
rlabel metal2 15962 14178 15962 14178 0 _0279_
rlabel metal2 15594 17034 15594 17034 0 _0280_
rlabel metal2 15226 15742 15226 15742 0 _0281_
rlabel metal2 5934 11118 5934 11118 0 _0282_
rlabel metal1 8188 13906 8188 13906 0 _0283_
rlabel metal2 12098 12444 12098 12444 0 _0284_
rlabel metal2 11270 12036 11270 12036 0 _0285_
rlabel metal1 15364 8466 15364 8466 0 _0286_
rlabel metal1 16100 8806 16100 8806 0 _0287_
rlabel metal1 13478 10608 13478 10608 0 _0288_
rlabel metal2 13294 10370 13294 10370 0 _0289_
rlabel metal1 4876 13226 4876 13226 0 _0290_
rlabel metal2 13570 10200 13570 10200 0 _0291_
rlabel metal1 13110 13294 13110 13294 0 _0292_
rlabel metal1 9016 14790 9016 14790 0 _0293_
rlabel metal1 10488 12614 10488 12614 0 _0294_
rlabel metal1 10074 8500 10074 8500 0 _0295_
rlabel metal1 13202 10676 13202 10676 0 _0296_
rlabel metal1 6578 12852 6578 12852 0 _0297_
rlabel viali 7863 13928 7863 13928 0 _0298_
rlabel metal1 6578 13328 6578 13328 0 _0299_
rlabel metal1 6394 12784 6394 12784 0 _0300_
rlabel metal1 6118 12886 6118 12886 0 _0301_
rlabel metal2 6670 10948 6670 10948 0 _0302_
rlabel metal2 7774 11084 7774 11084 0 _0303_
rlabel metal2 8326 9452 8326 9452 0 _0304_
rlabel metal2 10902 8602 10902 8602 0 _0305_
rlabel metal2 10718 8058 10718 8058 0 _0306_
rlabel metal2 6946 8092 6946 8092 0 _0307_
rlabel metal1 6762 10608 6762 10608 0 _0308_
rlabel metal1 7360 10438 7360 10438 0 _0309_
rlabel metal1 9660 8058 9660 8058 0 _0310_
rlabel metal1 10396 8058 10396 8058 0 _0311_
rlabel metal1 10074 8058 10074 8058 0 _0312_
rlabel metal1 15042 18190 15042 18190 0 _0313_
rlabel metal2 16054 8092 16054 8092 0 _0314_
rlabel via1 15778 7514 15778 7514 0 _0315_
rlabel metal1 16744 8058 16744 8058 0 _0316_
rlabel metal2 14950 7038 14950 7038 0 _0317_
rlabel metal1 16330 7786 16330 7786 0 _0318_
rlabel metal1 14674 7922 14674 7922 0 _0319_
rlabel metal1 18262 11526 18262 11526 0 _0320_
rlabel metal1 15640 10642 15640 10642 0 _0321_
rlabel metal2 17526 9214 17526 9214 0 _0322_
rlabel metal1 13892 7378 13892 7378 0 _0323_
rlabel viali 12458 7378 12458 7378 0 _0324_
rlabel metal1 11960 7242 11960 7242 0 _0325_
rlabel metal2 11546 7582 11546 7582 0 _0326_
rlabel via2 12558 7395 12558 7395 0 _0327_
rlabel metal1 17434 4182 17434 4182 0 _0328_
rlabel metal1 16422 6290 16422 6290 0 _0329_
rlabel metal1 15226 7344 15226 7344 0 _0330_
rlabel metal1 14720 7310 14720 7310 0 _0331_
rlabel metal2 13294 6834 13294 6834 0 _0332_
rlabel metal2 14766 9724 14766 9724 0 _0333_
rlabel metal1 14099 9554 14099 9554 0 _0334_
rlabel metal1 12558 10098 12558 10098 0 _0335_
rlabel metal2 13478 9860 13478 9860 0 _0336_
rlabel metal2 13846 8364 13846 8364 0 _0337_
rlabel metal2 13294 20706 13294 20706 0 _0338_
rlabel metal1 14260 19822 14260 19822 0 _0339_
rlabel metal1 18400 24378 18400 24378 0 _0340_
rlabel metal1 15548 18190 15548 18190 0 _0341_
rlabel metal1 17434 5236 17434 5236 0 _0342_
rlabel metal3 15755 6868 15755 6868 0 _0343_
rlabel metal2 17710 3910 17710 3910 0 _0344_
rlabel metal1 19918 4080 19918 4080 0 _0345_
rlabel metal3 16928 19380 16928 19380 0 _0346_
rlabel metal1 16652 11186 16652 11186 0 _0347_
rlabel metal1 12558 5712 12558 5712 0 _0348_
rlabel metal1 23690 25466 23690 25466 0 _0349_
rlabel metal1 24656 25874 24656 25874 0 _0350_
rlabel metal2 23690 25500 23690 25500 0 _0351_
rlabel metal2 22218 23341 22218 23341 0 _0352_
rlabel metal1 24334 19278 24334 19278 0 _0353_
rlabel metal2 23782 21284 23782 21284 0 _0354_
rlabel metal1 23092 20570 23092 20570 0 _0355_
rlabel metal1 22172 20570 22172 20570 0 _0356_
rlabel metal2 20838 20808 20838 20808 0 _0357_
rlabel metal1 23460 21114 23460 21114 0 _0358_
rlabel metal1 23322 23222 23322 23222 0 _0359_
rlabel metal1 24978 31994 24978 31994 0 _0360_
rlabel metal1 25011 31654 25011 31654 0 _0361_
rlabel metal2 21666 32164 21666 32164 0 _0362_
rlabel metal1 18446 34544 18446 34544 0 _0363_
rlabel metal2 17986 34408 17986 34408 0 _0364_
rlabel metal1 16882 33626 16882 33626 0 _0365_
rlabel metal1 16330 34510 16330 34510 0 _0366_
rlabel metal1 14950 34476 14950 34476 0 _0367_
rlabel metal1 14674 32844 14674 32844 0 _0368_
rlabel metal1 15134 32844 15134 32844 0 _0369_
rlabel metal2 15410 32538 15410 32538 0 _0370_
rlabel metal1 15778 31450 15778 31450 0 _0371_
rlabel metal1 15824 31790 15824 31790 0 _0372_
rlabel metal2 16882 32164 16882 32164 0 _0373_
rlabel metal1 17342 32368 17342 32368 0 _0374_
rlabel metal1 18354 31824 18354 31824 0 _0375_
rlabel via1 18906 31875 18906 31875 0 _0376_
rlabel metal1 19780 31450 19780 31450 0 _0377_
rlabel metal1 19274 31892 19274 31892 0 _0378_
rlabel metal1 19596 31654 19596 31654 0 _0379_
rlabel metal1 22402 31280 22402 31280 0 _0380_
rlabel metal1 25622 32436 25622 32436 0 _0381_
rlabel metal2 23966 31926 23966 31926 0 _0382_
rlabel metal1 25208 31926 25208 31926 0 _0383_
rlabel metal1 24196 32198 24196 32198 0 _0384_
rlabel metal1 22770 31926 22770 31926 0 _0385_
rlabel metal1 22310 31824 22310 31824 0 _0386_
rlabel metal1 19596 31790 19596 31790 0 _0387_
rlabel metal1 18906 31994 18906 31994 0 _0388_
rlabel via2 16698 31875 16698 31875 0 _0389_
rlabel metal1 15962 32436 15962 32436 0 _0390_
rlabel metal1 15042 34612 15042 34612 0 _0391_
rlabel metal2 15410 33966 15410 33966 0 _0392_
rlabel metal1 19366 35802 19366 35802 0 _0393_
rlabel metal1 22126 21386 22126 21386 0 _0394_
rlabel metal1 23046 30124 23046 30124 0 _0395_
rlabel metal1 20838 35530 20838 35530 0 _0396_
rlabel metal1 21666 33320 21666 33320 0 _0397_
rlabel metal1 23782 16218 23782 16218 0 _0398_
rlabel metal1 24794 32402 24794 32402 0 _0399_
rlabel metal1 18354 32946 18354 32946 0 _0400_
rlabel metal1 21114 33320 21114 33320 0 _0401_
rlabel metal2 18446 34170 18446 34170 0 _0402_
rlabel viali 18908 33966 18908 33966 0 _0403_
rlabel metal2 20976 32402 20976 32402 0 _0404_
rlabel metal2 13938 23817 13938 23817 0 _0405_
rlabel metal2 11868 25806 11868 25806 0 _0406_
rlabel metal1 10856 25126 10856 25126 0 _0407_
rlabel metal1 12512 21862 12512 21862 0 _0408_
rlabel metal1 12190 33490 12190 33490 0 _0409_
rlabel metal1 10948 37094 10948 37094 0 _0410_
rlabel metal1 24150 32878 24150 32878 0 _0411_
rlabel metal1 23736 32742 23736 32742 0 _0412_
rlabel metal2 20838 31076 20838 31076 0 _0413_
rlabel metal1 10672 31654 10672 31654 0 _0414_
rlabel metal2 9246 30838 9246 30838 0 _0415_
rlabel metal1 10396 30838 10396 30838 0 _0416_
rlabel metal2 11638 32096 11638 32096 0 _0417_
rlabel metal2 11914 34476 11914 34476 0 _0418_
rlabel metal1 20562 31280 20562 31280 0 _0419_
rlabel metal1 10166 31790 10166 31790 0 _0420_
rlabel metal2 10166 32062 10166 32062 0 _0421_
rlabel metal1 11270 32844 11270 32844 0 _0422_
rlabel metal2 11270 33456 11270 33456 0 _0423_
rlabel metal2 11086 34000 11086 34000 0 _0424_
rlabel metal1 8694 31688 8694 31688 0 _0425_
rlabel metal2 9522 32776 9522 32776 0 _0426_
rlabel metal1 11638 33354 11638 33354 0 _0427_
rlabel metal1 12006 33626 12006 33626 0 _0428_
rlabel metal1 17802 33898 17802 33898 0 _0429_
rlabel metal1 19274 35666 19274 35666 0 _0430_
rlabel metal2 18354 35258 18354 35258 0 _0431_
rlabel metal2 19918 35292 19918 35292 0 _0432_
rlabel metal2 20102 35462 20102 35462 0 _0433_
rlabel metal2 11454 24548 11454 24548 0 _0434_
rlabel metal1 11696 33898 11696 33898 0 _0435_
rlabel metal2 11546 34918 11546 34918 0 _0436_
rlabel metal2 11730 34782 11730 34782 0 _0437_
rlabel metal1 20332 35802 20332 35802 0 _0438_
rlabel metal1 17388 36006 17388 36006 0 _0439_
rlabel metal2 18170 37026 18170 37026 0 _0440_
rlabel metal1 19550 36244 19550 36244 0 _0441_
rlabel metal1 17986 36244 17986 36244 0 _0442_
rlabel metal2 14674 36346 14674 36346 0 _0443_
rlabel metal1 10488 26350 10488 26350 0 _0444_
rlabel metal1 10166 29138 10166 29138 0 _0445_
rlabel metal1 9798 33456 9798 33456 0 _0446_
rlabel metal1 14030 35734 14030 35734 0 _0447_
rlabel metal1 12742 35020 12742 35020 0 _0448_
rlabel metal1 14122 35802 14122 35802 0 _0449_
rlabel metal1 13938 35122 13938 35122 0 _0450_
rlabel metal2 14214 35360 14214 35360 0 _0451_
rlabel metal2 14398 35530 14398 35530 0 _0452_
rlabel metal1 17664 35122 17664 35122 0 _0453_
rlabel metal1 17848 36346 17848 36346 0 _0454_
rlabel metal1 15410 35564 15410 35564 0 _0455_
rlabel metal1 15824 35666 15824 35666 0 _0456_
rlabel viali 10166 29611 10166 29611 0 _0457_
rlabel metal1 8970 37162 8970 37162 0 _0458_
rlabel metal1 9706 33626 9706 33626 0 _0459_
rlabel metal1 13386 35530 13386 35530 0 _0460_
rlabel metal1 15456 35666 15456 35666 0 _0461_
rlabel metal2 23138 35258 23138 35258 0 _0462_
rlabel metal1 22954 35020 22954 35020 0 _0463_
rlabel metal2 21482 35428 21482 35428 0 _0464_
rlabel metal2 17894 35360 17894 35360 0 _0465_
rlabel metal1 17802 35734 17802 35734 0 _0466_
rlabel metal1 21206 35632 21206 35632 0 _0467_
rlabel metal1 21873 35598 21873 35598 0 _0468_
rlabel metal1 10166 27472 10166 27472 0 _0469_
rlabel metal1 10212 27574 10212 27574 0 _0470_
rlabel metal1 10396 34374 10396 34374 0 _0471_
rlabel metal2 12834 35020 12834 35020 0 _0472_
rlabel metal1 13018 35088 13018 35088 0 _0473_
rlabel metal1 13662 35088 13662 35088 0 _0474_
rlabel metal1 17618 34986 17618 34986 0 _0475_
rlabel metal2 23966 35462 23966 35462 0 _0476_
rlabel metal1 24932 35666 24932 35666 0 _0477_
rlabel metal1 24748 35666 24748 35666 0 _0478_
rlabel metal1 24472 35598 24472 35598 0 _0479_
rlabel metal1 23598 35768 23598 35768 0 _0480_
rlabel metal1 9844 25466 9844 25466 0 _0481_
rlabel metal1 9798 26554 9798 26554 0 _0482_
rlabel metal2 10258 34816 10258 34816 0 _0483_
rlabel metal1 9936 35258 9936 35258 0 _0484_
rlabel metal1 20010 35156 20010 35156 0 _0485_
rlabel metal2 22586 35462 22586 35462 0 _0486_
rlabel metal1 26404 35802 26404 35802 0 _0487_
rlabel metal1 26082 36108 26082 36108 0 _0488_
rlabel metal1 26036 35462 26036 35462 0 _0489_
rlabel metal1 25308 35802 25308 35802 0 _0490_
rlabel metal1 25760 35530 25760 35530 0 _0491_
rlabel metal1 25162 35258 25162 35258 0 _0492_
rlabel metal2 25622 35292 25622 35292 0 _0493_
rlabel metal1 10442 23120 10442 23120 0 _0494_
rlabel metal3 10005 33252 10005 33252 0 _0495_
rlabel metal2 8326 36856 8326 36856 0 _0496_
rlabel metal1 9384 34714 9384 34714 0 _0497_
rlabel metal1 9246 34612 9246 34612 0 _0498_
rlabel metal2 9338 35428 9338 35428 0 _0499_
rlabel metal2 20746 35326 20746 35326 0 _0500_
rlabel metal2 25530 35700 25530 35700 0 _0501_
rlabel metal2 26818 34816 26818 34816 0 _0502_
rlabel metal1 26220 35258 26220 35258 0 _0503_
rlabel metal1 26466 34986 26466 34986 0 _0504_
rlabel metal1 26128 34578 26128 34578 0 _0505_
rlabel metal1 8372 24106 8372 24106 0 _0506_
rlabel via2 8326 34595 8326 34595 0 _0507_
rlabel metal1 8602 34510 8602 34510 0 _0508_
rlabel via2 8694 34459 8694 34459 0 _0509_
rlabel metal1 25898 34612 25898 34612 0 _0510_
rlabel metal2 19274 17748 19274 17748 0 _0511_
rlabel metal1 8004 18938 8004 18938 0 _0512_
rlabel metal1 25622 16116 25622 16116 0 _0513_
rlabel metal2 14674 16405 14674 16405 0 _0514_
rlabel metal1 7452 18802 7452 18802 0 _0515_
rlabel metal1 21804 27914 21804 27914 0 _0516_
rlabel metal1 22264 23698 22264 23698 0 _0517_
rlabel metal1 23322 21318 23322 21318 0 _0518_
rlabel metal2 21482 18972 21482 18972 0 _0519_
rlabel metal1 22494 18938 22494 18938 0 _0520_
rlabel metal1 21758 18632 21758 18632 0 _0521_
rlabel metal1 22456 21658 22456 21658 0 _0522_
rlabel metal2 22678 21658 22678 21658 0 _0523_
rlabel metal2 22862 26452 22862 26452 0 _0524_
rlabel metal1 25944 28594 25944 28594 0 _0525_
rlabel metal1 25024 28730 25024 28730 0 _0526_
rlabel metal2 22310 29308 22310 29308 0 _0527_
rlabel metal1 10764 37298 10764 37298 0 _0528_
rlabel metal2 24886 32538 24886 32538 0 _0529_
rlabel metal2 22494 33558 22494 33558 0 _0530_
rlabel metal1 23184 34170 23184 34170 0 _0531_
rlabel metal1 22632 32538 22632 32538 0 _0532_
rlabel metal1 23276 33626 23276 33626 0 _0533_
rlabel metal2 21298 30906 21298 30906 0 _0534_
rlabel metal1 22356 31382 22356 31382 0 _0535_
rlabel metal1 21712 32198 21712 32198 0 _0536_
rlabel metal1 21160 30906 21160 30906 0 _0537_
rlabel metal2 21022 31348 21022 31348 0 _0538_
rlabel metal2 20838 32198 20838 32198 0 _0539_
rlabel metal2 9614 32198 9614 32198 0 _0540_
rlabel metal1 9292 32334 9292 32334 0 _0541_
rlabel via2 9338 32283 9338 32283 0 _0542_
rlabel metal1 19182 33014 19182 33014 0 _0543_
rlabel via2 17894 32861 17894 32861 0 _0544_
rlabel metal1 9384 30906 9384 30906 0 _0545_
rlabel metal1 9200 31246 9200 31246 0 _0546_
rlabel via2 14582 30787 14582 30787 0 _0547_
rlabel metal1 17388 31994 17388 31994 0 _0548_
rlabel metal1 17250 30906 17250 30906 0 _0549_
rlabel metal1 9982 31178 9982 31178 0 _0550_
rlabel metal1 13294 31416 13294 31416 0 _0551_
rlabel metal2 16146 31994 16146 31994 0 _0552_
rlabel metal1 15042 30702 15042 30702 0 _0553_
rlabel metal2 14214 30906 14214 30906 0 _0554_
rlabel metal1 10672 31790 10672 31790 0 _0555_
rlabel metal2 12926 31756 12926 31756 0 _0556_
rlabel metal1 11270 31994 11270 31994 0 _0557_
rlabel metal1 14950 32504 14950 32504 0 _0558_
rlabel metal2 15134 32572 15134 32572 0 _0559_
rlabel metal1 13110 32300 13110 32300 0 _0560_
rlabel metal1 15410 33354 15410 33354 0 _0561_
rlabel metal2 15134 33796 15134 33796 0 _0562_
rlabel metal1 14444 33966 14444 33966 0 _0563_
rlabel metal2 12006 32164 12006 32164 0 _0564_
rlabel metal1 13662 32538 13662 32538 0 _0565_
rlabel metal1 20608 13158 20608 13158 0 _0566_
rlabel metal1 15318 10642 15318 10642 0 _0567_
rlabel metal1 14490 10744 14490 10744 0 _0568_
rlabel metal1 20930 19142 20930 19142 0 _0569_
rlabel metal1 20470 19278 20470 19278 0 _0570_
rlabel metal2 21298 20944 21298 20944 0 _0571_
rlabel metal1 21942 23630 21942 23630 0 _0572_
rlabel metal2 20930 29376 20930 29376 0 _0573_
rlabel metal1 21758 23834 21758 23834 0 _0574_
rlabel metal1 5290 32402 5290 32402 0 _0575_
rlabel metal1 8786 33456 8786 33456 0 _0576_
rlabel metal1 13846 13838 13846 13838 0 _0577_
rlabel metal1 14260 14518 14260 14518 0 _0578_
rlabel metal1 13018 14518 13018 14518 0 _0579_
rlabel metal1 13018 13736 13018 13736 0 _0580_
rlabel metal1 9545 13770 9545 13770 0 _0581_
rlabel metal2 12742 14586 12742 14586 0 _0582_
rlabel metal2 12098 14994 12098 14994 0 _0583_
rlabel metal1 9384 13294 9384 13294 0 _0584_
rlabel via2 8050 14909 8050 14909 0 _0585_
rlabel metal1 12666 14994 12666 14994 0 _0586_
rlabel metal2 13570 11662 13570 11662 0 _0587_
rlabel metal1 12604 15130 12604 15130 0 _0588_
rlabel metal1 12282 15436 12282 15436 0 _0589_
rlabel metal1 12098 15368 12098 15368 0 _0590_
rlabel metal1 5842 13872 5842 13872 0 _0591_
rlabel metal1 4738 13294 4738 13294 0 _0592_
rlabel metal2 4554 14008 4554 14008 0 _0593_
rlabel metal2 10810 14042 10810 14042 0 _0594_
rlabel metal1 11040 13294 11040 13294 0 _0595_
rlabel metal1 8602 13430 8602 13430 0 _0596_
rlabel metal1 4784 14382 4784 14382 0 _0597_
rlabel metal1 5796 13294 5796 13294 0 _0598_
rlabel metal1 5704 13974 5704 13974 0 _0599_
rlabel metal2 6118 13702 6118 13702 0 _0600_
rlabel metal1 5845 14042 5845 14042 0 _0601_
rlabel metal1 6394 14314 6394 14314 0 _0602_
rlabel metal2 8050 14382 8050 14382 0 _0603_
rlabel metal1 9476 13498 9476 13498 0 _0604_
rlabel metal1 8648 13974 8648 13974 0 _0605_
rlabel metal2 8234 14008 8234 14008 0 _0606_
rlabel metal2 7130 15334 7130 15334 0 _0607_
rlabel via2 9430 15555 9430 15555 0 _0608_
rlabel metal1 8050 14416 8050 14416 0 _0609_
rlabel metal2 7866 14756 7866 14756 0 _0610_
rlabel metal1 6854 15028 6854 15028 0 _0611_
rlabel metal2 5290 14586 5290 14586 0 _0612_
rlabel metal1 5244 14042 5244 14042 0 _0613_
rlabel metal2 4646 14076 4646 14076 0 _0614_
rlabel metal2 5382 11696 5382 11696 0 _0615_
rlabel metal1 4876 11730 4876 11730 0 _0616_
rlabel metal2 4738 12002 4738 12002 0 _0617_
rlabel metal1 5750 11764 5750 11764 0 _0618_
rlabel metal1 8924 12410 8924 12410 0 _0619_
rlabel metal1 5520 11526 5520 11526 0 _0620_
rlabel metal1 5244 11866 5244 11866 0 _0621_
rlabel metal2 8234 8330 8234 8330 0 _0622_
rlabel metal1 6900 9146 6900 9146 0 _0623_
rlabel via1 7129 9554 7129 9554 0 _0624_
rlabel metal2 7222 10234 7222 10234 0 _0625_
rlabel metal1 7682 10098 7682 10098 0 _0626_
rlabel metal2 8142 11594 8142 11594 0 _0627_
rlabel metal1 8234 11186 8234 11186 0 _0628_
rlabel metal1 7912 10234 7912 10234 0 _0629_
rlabel metal1 7360 9554 7360 9554 0 _0630_
rlabel metal1 8786 7990 8786 7990 0 _0631_
rlabel metal1 7130 7922 7130 7922 0 _0632_
rlabel metal2 7130 8262 7130 8262 0 _0633_
rlabel metal1 5934 8330 5934 8330 0 _0634_
rlabel metal1 10396 10234 10396 10234 0 _0635_
rlabel metal2 10902 11492 10902 11492 0 _0636_
rlabel metal1 11086 10676 11086 10676 0 _0637_
rlabel metal1 6394 10132 6394 10132 0 _0638_
rlabel metal1 5658 8398 5658 8398 0 _0639_
rlabel metal2 9062 8772 9062 8772 0 _0640_
rlabel metal1 8878 8058 8878 8058 0 _0641_
rlabel metal1 8464 8874 8464 8874 0 _0642_
rlabel metal2 12650 9724 12650 9724 0 _0643_
rlabel metal2 12742 11356 12742 11356 0 _0644_
rlabel metal1 12282 10574 12282 10574 0 _0645_
rlabel metal2 12374 10234 12374 10234 0 _0646_
rlabel metal1 9246 9996 9246 9996 0 _0647_
rlabel metal1 8651 9894 8651 9894 0 _0648_
rlabel metal1 25714 15674 25714 15674 0 _0649_
rlabel metal1 25254 16490 25254 16490 0 _0650_
rlabel metal1 2714 17748 2714 17748 0 _0651_
rlabel metal2 13662 20604 13662 20604 0 _0652_
rlabel metal1 29486 30770 29486 30770 0 _0653_
rlabel metal1 17756 9078 17756 9078 0 _0654_
rlabel metal1 16008 9010 16008 9010 0 _0655_
rlabel metal2 11454 21148 11454 21148 0 _0656_
rlabel metal2 21574 11050 21574 11050 0 _0657_
rlabel metal2 36662 17680 36662 17680 0 _0658_
rlabel metal1 24840 23698 24840 23698 0 _0659_
rlabel metal2 8602 19686 8602 19686 0 _0660_
rlabel metal1 24702 31790 24702 31790 0 _0661_
rlabel metal1 24702 32810 24702 32810 0 _0662_
rlabel metal2 8326 19346 8326 19346 0 _0663_
rlabel metal1 13892 20978 13892 20978 0 _0664_
rlabel metal1 17986 3570 17986 3570 0 _0665_
rlabel metal1 20194 4080 20194 4080 0 _0666_
rlabel metal2 33810 29342 33810 29342 0 _0667_
rlabel metal1 13432 5882 13432 5882 0 _0668_
rlabel metal1 30222 31790 30222 31790 0 _0669_
rlabel metal3 25001 19244 25001 19244 0 _0670_
rlabel metal1 30038 31926 30038 31926 0 _0671_
rlabel metal1 36524 17170 36524 17170 0 _0672_
rlabel via2 22034 8245 22034 8245 0 _0673_
rlabel metal2 27554 19482 27554 19482 0 _0674_
rlabel metal1 28428 8942 28428 8942 0 _0675_
rlabel metal1 26542 13294 26542 13294 0 _0676_
rlabel metal1 18745 19346 18745 19346 0 _0677_
rlabel metal2 33350 14047 33350 14047 0 _0678_
rlabel metal1 27186 13838 27186 13838 0 _0679_
rlabel via2 20194 16541 20194 16541 0 _0680_
rlabel metal1 15594 14824 15594 14824 0 _0681_
rlabel metal1 21336 10710 21336 10710 0 _0682_
rlabel metal1 29854 20808 29854 20808 0 _0683_
rlabel metal1 21758 19346 21758 19346 0 _0684_
rlabel metal1 34362 17272 34362 17272 0 _0685_
rlabel metal3 30153 19380 30153 19380 0 _0686_
rlabel metal1 15778 21080 15778 21080 0 _0687_
rlabel metal1 23322 18054 23322 18054 0 _0688_
rlabel metal2 32522 8908 32522 8908 0 _0689_
rlabel metal1 16882 7446 16882 7446 0 _0690_
rlabel via1 18546 20502 18546 20502 0 _0691_
rlabel metal1 27600 14994 27600 14994 0 _0692_
rlabel metal1 20838 19414 20838 19414 0 _0693_
rlabel metal1 24334 14994 24334 14994 0 _0694_
rlabel metal1 21436 22610 21436 22610 0 _0695_
rlabel metal2 24886 27744 24886 27744 0 _0696_
rlabel metal2 21022 22780 21022 22780 0 _0697_
rlabel metal1 24978 14926 24978 14926 0 _0698_
rlabel metal1 25208 10030 25208 10030 0 _0699_
rlabel metal2 32522 14790 32522 14790 0 _0700_
rlabel via1 32982 22678 32982 22678 0 _0701_
rlabel metal1 34178 17238 34178 17238 0 _0702_
rlabel metal1 26174 7514 26174 7514 0 _0703_
rlabel metal1 17158 14450 17158 14450 0 _0704_
rlabel metal2 19274 8211 19274 8211 0 _0705_
rlabel metal1 26542 10030 26542 10030 0 _0706_
rlabel metal2 25990 16252 25990 16252 0 _0707_
rlabel metal2 19458 10948 19458 10948 0 _0708_
rlabel metal2 31142 10693 31142 10693 0 _0709_
rlabel metal1 25668 9554 25668 9554 0 _0710_
rlabel via2 18078 13515 18078 13515 0 _0711_
rlabel metal1 17618 12852 17618 12852 0 _0712_
rlabel metal2 21206 11900 21206 11900 0 _0713_
rlabel metal2 24242 13804 24242 13804 0 _0714_
rlabel metal1 22908 13226 22908 13226 0 _0715_
rlabel metal1 28106 9554 28106 9554 0 _0716_
rlabel metal1 29486 18258 29486 18258 0 _0717_
rlabel metal1 27462 14450 27462 14450 0 _0718_
rlabel metal1 27278 14314 27278 14314 0 _0719_
rlabel via3 26381 15164 26381 15164 0 _0720_
rlabel via3 29509 8228 29509 8228 0 _0721_
rlabel metal1 16974 7208 16974 7208 0 _0722_
rlabel metal2 23598 12988 23598 12988 0 _0723_
rlabel metal1 25392 12206 25392 12206 0 _0724_
rlabel metal2 24426 12580 24426 12580 0 _0725_
rlabel metal1 24932 2414 24932 2414 0 _0726_
rlabel metal1 28750 23630 28750 23630 0 _0727_
rlabel metal1 24150 23290 24150 23290 0 _0728_
rlabel metal2 24794 21420 24794 21420 0 _0729_
rlabel metal1 17664 24786 17664 24786 0 _0730_
rlabel metal4 32108 18428 32108 18428 0 _0731_
rlabel metal2 34546 19992 34546 19992 0 _0732_
rlabel metal2 34546 18309 34546 18309 0 _0733_
rlabel metal1 32752 9146 32752 9146 0 _0734_
rlabel metal2 31372 19278 31372 19278 0 _0735_
rlabel metal1 25944 19346 25944 19346 0 _0736_
rlabel metal1 26082 10642 26082 10642 0 _0737_
rlabel metal1 26864 11730 26864 11730 0 _0738_
rlabel metal1 25944 11594 25944 11594 0 _0739_
rlabel metal2 26358 18972 26358 18972 0 _0740_
rlabel metal1 26266 18632 26266 18632 0 _0741_
rlabel metal2 25898 17476 25898 17476 0 _0742_
rlabel metal2 26266 18564 26266 18564 0 _0743_
rlabel metal1 25438 17748 25438 17748 0 _0744_
rlabel metal2 25714 17850 25714 17850 0 _0745_
rlabel metal2 24978 17952 24978 17952 0 _0746_
rlabel via1 25246 18666 25246 18666 0 _0747_
rlabel metal1 25024 19346 25024 19346 0 _0748_
rlabel metal1 23782 19856 23782 19856 0 _0749_
rlabel metal2 17066 20978 17066 20978 0 _0750_
rlabel metal1 24104 20026 24104 20026 0 _0751_
rlabel metal1 24472 19482 24472 19482 0 _0752_
rlabel metal1 19780 12954 19780 12954 0 _0753_
rlabel metal1 20792 8466 20792 8466 0 _0754_
rlabel metal3 32407 22644 32407 22644 0 _0755_
rlabel metal1 21528 9146 21528 9146 0 _0756_
rlabel metal2 26818 16592 26818 16592 0 _0757_
rlabel metal1 21390 8398 21390 8398 0 _0758_
rlabel metal1 21988 9146 21988 9146 0 _0759_
rlabel metal1 26450 16048 26450 16048 0 _0760_
rlabel metal1 26358 13498 26358 13498 0 _0761_
rlabel metal2 23046 11696 23046 11696 0 _0762_
rlabel metal1 28704 8058 28704 8058 0 _0763_
rlabel metal2 22034 22797 22034 22797 0 _0764_
rlabel metal1 19642 12172 19642 12172 0 _0765_
rlabel metal1 28152 12614 28152 12614 0 _0766_
rlabel metal1 27600 15674 27600 15674 0 _0767_
rlabel metal1 26772 13498 26772 13498 0 _0768_
rlabel metal1 21712 8262 21712 8262 0 _0769_
rlabel via2 29210 16099 29210 16099 0 _0770_
rlabel metal1 20976 21522 20976 21522 0 _0771_
rlabel metal1 21712 15470 21712 15470 0 _0772_
rlabel metal2 35098 14943 35098 14943 0 _0773_
rlabel metal1 17940 13294 17940 13294 0 _0774_
rlabel metal1 20102 9622 20102 9622 0 _0775_
rlabel metal1 24472 12614 24472 12614 0 _0776_
rlabel metal2 22770 17442 22770 17442 0 _0777_
rlabel metal1 14076 12206 14076 12206 0 _0778_
rlabel metal1 20930 11628 20930 11628 0 _0779_
rlabel metal1 22264 14994 22264 14994 0 _0780_
rlabel metal1 23046 6630 23046 6630 0 _0781_
rlabel metal1 14950 9996 14950 9996 0 _0782_
rlabel via1 24794 6902 24794 6902 0 _0783_
rlabel metal1 16008 12818 16008 12818 0 _0784_
rlabel metal1 23368 10506 23368 10506 0 _0785_
rlabel metal1 31326 10064 31326 10064 0 _0786_
rlabel metal1 19918 10608 19918 10608 0 _0787_
rlabel metal2 18722 9078 18722 9078 0 _0788_
rlabel via2 32890 20757 32890 20757 0 _0789_
rlabel metal1 17986 10098 17986 10098 0 _0790_
rlabel metal1 14950 13906 14950 13906 0 _0791_
rlabel metal1 17710 13498 17710 13498 0 _0792_
rlabel metal2 17618 14637 17618 14637 0 _0793_
rlabel metal1 26358 15674 26358 15674 0 _0794_
rlabel metal2 22126 15232 22126 15232 0 _0795_
rlabel metal1 25668 16694 25668 16694 0 _0796_
rlabel metal1 34270 22712 34270 22712 0 _0797_
rlabel metal1 18768 14382 18768 14382 0 _0798_
rlabel metal2 22494 11322 22494 11322 0 _0799_
rlabel metal1 28888 8602 28888 8602 0 _0800_
rlabel metal1 17250 8840 17250 8840 0 _0801_
rlabel metal1 24334 9520 24334 9520 0 _0802_
rlabel metal1 24748 8602 24748 8602 0 _0803_
rlabel metal1 28060 7242 28060 7242 0 _0804_
rlabel metal1 23184 8466 23184 8466 0 _0805_
rlabel metal1 27968 20298 27968 20298 0 _0806_
rlabel metal2 21482 14688 21482 14688 0 _0807_
rlabel metal1 24886 7412 24886 7412 0 _0808_
rlabel metal2 25438 8432 25438 8432 0 _0809_
rlabel metal2 24426 9996 24426 9996 0 _0810_
rlabel metal2 24426 9231 24426 9231 0 _0811_
rlabel metal1 23782 9350 23782 9350 0 _0812_
rlabel metal2 22218 10336 22218 10336 0 _0813_
rlabel metal1 22724 10234 22724 10234 0 _0814_
rlabel metal1 21712 14586 21712 14586 0 _0815_
rlabel metal2 22218 11866 22218 11866 0 _0816_
rlabel metal3 23851 18020 23851 18020 0 _0817_
rlabel metal1 18860 8874 18860 8874 0 _0818_
rlabel metal2 27646 30600 27646 30600 0 _0819_
rlabel metal1 28474 30294 28474 30294 0 _0820_
rlabel metal2 26266 27030 26266 27030 0 _0821_
rlabel via2 23322 17323 23322 17323 0 _0822_
rlabel metal1 21252 26962 21252 26962 0 _0823_
rlabel metal2 18906 26758 18906 26758 0 _0824_
rlabel metal1 20102 26962 20102 26962 0 _0825_
rlabel metal1 19780 27438 19780 27438 0 _0826_
rlabel metal1 20746 26418 20746 26418 0 _0827_
rlabel metal1 26956 28050 26956 28050 0 _0828_
rlabel metal1 25944 28662 25944 28662 0 _0829_
rlabel metal2 19918 29478 19918 29478 0 _0830_
rlabel metal2 25898 27098 25898 27098 0 _0831_
rlabel metal2 21942 24888 21942 24888 0 _0832_
rlabel metal2 21482 27200 21482 27200 0 _0833_
rlabel metal2 21758 26588 21758 26588 0 _0834_
rlabel metal1 27278 25806 27278 25806 0 _0835_
rlabel via2 17250 21539 17250 21539 0 _0836_
rlabel metal2 36478 17340 36478 17340 0 _0837_
rlabel metal1 31832 20910 31832 20910 0 _0838_
rlabel metal1 27876 19890 27876 19890 0 _0839_
rlabel metal1 27646 24650 27646 24650 0 _0840_
rlabel metal2 20562 6409 20562 6409 0 _0841_
rlabel metal2 19182 24752 19182 24752 0 _0842_
rlabel metal1 35098 25228 35098 25228 0 _0843_
rlabel metal1 35236 25466 35236 25466 0 _0844_
rlabel metal1 35052 27846 35052 27846 0 _0845_
rlabel metal1 34316 27438 34316 27438 0 _0846_
rlabel metal1 30498 27404 30498 27404 0 _0847_
rlabel metal1 32706 29206 32706 29206 0 _0848_
rlabel metal2 34362 26758 34362 26758 0 _0849_
rlabel metal1 30452 25670 30452 25670 0 _0850_
rlabel metal1 34040 26282 34040 26282 0 _0851_
rlabel metal1 34546 26962 34546 26962 0 _0852_
rlabel metal1 35696 27030 35696 27030 0 _0853_
rlabel metal1 35742 26758 35742 26758 0 _0854_
rlabel metal1 32292 17170 32292 17170 0 _0855_
rlabel metal2 35098 18360 35098 18360 0 _0856_
rlabel metal1 28497 31756 28497 31756 0 _0857_
rlabel metal1 31694 28050 31694 28050 0 _0858_
rlabel metal2 32062 27846 32062 27846 0 _0859_
rlabel metal1 33580 27846 33580 27846 0 _0860_
rlabel metal1 31372 27846 31372 27846 0 _0861_
rlabel metal1 31234 29546 31234 29546 0 _0862_
rlabel metal1 32430 27982 32430 27982 0 _0863_
rlabel metal2 32982 26486 32982 26486 0 _0864_
rlabel metal1 32384 27846 32384 27846 0 _0865_
rlabel metal2 32798 29750 32798 29750 0 _0866_
rlabel metal1 28014 31654 28014 31654 0 _0867_
rlabel metal1 30130 29104 30130 29104 0 _0868_
rlabel metal1 30636 29274 30636 29274 0 _0869_
rlabel metal1 28704 27098 28704 27098 0 _0870_
rlabel metal1 30820 29478 30820 29478 0 _0871_
rlabel metal1 27738 31280 27738 31280 0 _0872_
rlabel metal1 27830 31348 27830 31348 0 _0873_
rlabel metal2 34546 29444 34546 29444 0 _0874_
rlabel metal1 34408 29818 34408 29818 0 _0875_
rlabel metal1 31050 29206 31050 29206 0 _0876_
rlabel metal2 34822 20655 34822 20655 0 _0877_
rlabel via1 33061 9554 33061 9554 0 _0878_
rlabel metal2 34730 20026 34730 20026 0 _0879_
rlabel metal1 32752 29614 32752 29614 0 _0880_
rlabel metal1 32200 29818 32200 29818 0 _0881_
rlabel metal2 28014 14841 28014 14841 0 _0882_
rlabel metal2 28566 26894 28566 26894 0 _0883_
rlabel metal1 29348 15470 29348 15470 0 _0884_
rlabel metal1 29900 29138 29900 29138 0 _0885_
rlabel metal1 29348 27846 29348 27846 0 _0886_
rlabel metal1 31188 30226 31188 30226 0 _0887_
rlabel metal1 32200 28934 32200 28934 0 _0888_
rlabel metal1 30176 27642 30176 27642 0 _0889_
rlabel metal1 32522 30260 32522 30260 0 _0890_
rlabel metal1 30958 29716 30958 29716 0 _0891_
rlabel metal2 32706 30838 32706 30838 0 _0892_
rlabel metal1 29532 27302 29532 27302 0 _0893_
rlabel metal2 30176 20842 30176 20842 0 _0894_
rlabel metal2 30406 29359 30406 29359 0 _0895_
rlabel metal1 30176 28934 30176 28934 0 _0896_
rlabel metal1 33902 16014 33902 16014 0 _0897_
rlabel metal1 30360 26554 30360 26554 0 _0898_
rlabel metal1 31419 23664 31419 23664 0 _0899_
rlabel metal1 31096 22202 31096 22202 0 _0900_
rlabel metal1 31464 20910 31464 20910 0 _0901_
rlabel metal1 28221 21590 28221 21590 0 _0902_
rlabel via2 33718 25245 33718 25245 0 _0903_
rlabel metal1 32982 25874 32982 25874 0 _0904_
rlabel metal1 32430 26010 32430 26010 0 _0905_
rlabel metal2 28382 22950 28382 22950 0 _0906_
rlabel metal2 31142 21114 31142 21114 0 _0907_
rlabel metal1 32614 18836 32614 18836 0 _0908_
rlabel metal1 33350 18632 33350 18632 0 _0909_
rlabel metal1 35558 18632 35558 18632 0 _0910_
rlabel metal1 34224 18734 34224 18734 0 _0911_
rlabel metal2 35190 16218 35190 16218 0 _0912_
rlabel metal1 28014 20468 28014 20468 0 _0913_
rlabel metal1 33626 20502 33626 20502 0 _0914_
rlabel metal1 27646 16660 27646 16660 0 _0915_
rlabel metal1 32890 25296 32890 25296 0 _0916_
rlabel metal1 30958 25262 30958 25262 0 _0917_
rlabel metal2 31142 17408 31142 17408 0 _0918_
rlabel metal1 27922 18156 27922 18156 0 _0919_
rlabel metal1 32752 16558 32752 16558 0 _0920_
rlabel metal1 32522 24752 32522 24752 0 _0921_
rlabel metal1 32706 24208 32706 24208 0 _0922_
rlabel metal2 33074 23460 33074 23460 0 _0923_
rlabel metal1 32476 21318 32476 21318 0 _0924_
rlabel metal1 32890 22474 32890 22474 0 _0925_
rlabel metal2 32706 19244 32706 19244 0 _0926_
rlabel metal1 33948 18598 33948 18598 0 _0927_
rlabel metal1 29486 24752 29486 24752 0 _0928_
rlabel metal2 29210 24582 29210 24582 0 _0929_
rlabel metal1 31924 22406 31924 22406 0 _0930_
rlabel via2 28934 13787 28934 13787 0 _0931_
rlabel metal1 28934 16048 28934 16048 0 _0932_
rlabel metal3 34431 22508 34431 22508 0 _0933_
rlabel metal1 34914 20944 34914 20944 0 _0934_
rlabel metal2 31418 21284 31418 21284 0 _0935_
rlabel metal2 30222 22780 30222 22780 0 _0936_
rlabel metal1 29210 22508 29210 22508 0 _0937_
rlabel metal1 32476 20434 32476 20434 0 _0938_
rlabel metal1 32798 26384 32798 26384 0 _0939_
rlabel metal1 32752 20978 32752 20978 0 _0940_
rlabel metal1 33350 20808 33350 20808 0 _0941_
rlabel metal1 33028 13906 33028 13906 0 _0942_
rlabel viali 33625 15470 33625 15470 0 _0943_
rlabel metal2 35742 21114 35742 21114 0 _0944_
rlabel metal1 34822 16558 34822 16558 0 _0945_
rlabel metal2 33442 21250 33442 21250 0 _0946_
rlabel metal1 32292 23494 32292 23494 0 _0947_
rlabel metal2 33166 25398 33166 25398 0 _0948_
rlabel metal2 33994 26384 33994 26384 0 _0949_
rlabel metal1 33580 26010 33580 26010 0 _0950_
rlabel metal1 33258 25262 33258 25262 0 _0951_
rlabel viali 32798 25263 32798 25263 0 _0952_
rlabel metal2 33350 26112 33350 26112 0 _0953_
rlabel metal1 32154 25364 32154 25364 0 _0954_
rlabel metal1 31510 25296 31510 25296 0 _0955_
rlabel metal2 31786 13957 31786 13957 0 _0956_
rlabel metal1 29670 16218 29670 16218 0 _0957_
rlabel metal1 28566 14960 28566 14960 0 _0958_
rlabel metal1 30038 15062 30038 15062 0 _0959_
rlabel metal2 30682 14348 30682 14348 0 _0960_
rlabel metal2 31970 13566 31970 13566 0 _0961_
rlabel metal2 29486 14756 29486 14756 0 _0962_
rlabel metal2 32154 14110 32154 14110 0 _0963_
rlabel metal1 32798 14042 32798 14042 0 _0964_
rlabel metal1 32430 17204 32430 17204 0 _0965_
rlabel metal2 32614 16864 32614 16864 0 _0966_
rlabel metal1 32384 16218 32384 16218 0 _0967_
rlabel metal1 32338 24922 32338 24922 0 _0968_
rlabel metal1 32844 16966 32844 16966 0 _0969_
rlabel metal1 32982 17238 32982 17238 0 _0970_
rlabel metal1 33580 17170 33580 17170 0 _0971_
rlabel metal1 32614 12206 32614 12206 0 _0972_
rlabel metal1 32338 14790 32338 14790 0 _0973_
rlabel metal1 29992 11118 29992 11118 0 _0974_
rlabel metal1 31786 11832 31786 11832 0 _0975_
rlabel metal2 32706 11322 32706 11322 0 _0976_
rlabel metal2 33718 10404 33718 10404 0 _0977_
rlabel metal1 30636 18054 30636 18054 0 _0978_
rlabel metal2 32522 13124 32522 13124 0 _0979_
rlabel via1 28382 19346 28382 19346 0 _0980_
rlabel metal2 30682 10812 30682 10812 0 _0981_
rlabel metal1 31832 20230 31832 20230 0 _0982_
rlabel metal2 31050 10438 31050 10438 0 _0983_
rlabel metal1 32890 10778 32890 10778 0 _0984_
rlabel metal1 28152 19346 28152 19346 0 _0985_
rlabel metal2 30222 19890 30222 19890 0 _0986_
rlabel metal2 32154 17136 32154 17136 0 _0987_
rlabel metal1 29762 11730 29762 11730 0 _0988_
rlabel metal2 29210 11577 29210 11577 0 _0989_
rlabel metal1 29072 11730 29072 11730 0 _0990_
rlabel metal1 34638 11526 34638 11526 0 _0991_
rlabel via3 29325 24956 29325 24956 0 _0992_
rlabel metal1 32568 13498 32568 13498 0 _0993_
rlabel metal2 33902 16864 33902 16864 0 _0994_
rlabel metal1 34776 13294 34776 13294 0 _0995_
rlabel metal1 35834 14994 35834 14994 0 _0996_
rlabel metal1 34638 27438 34638 27438 0 _0997_
rlabel metal1 33534 20400 33534 20400 0 _0998_
rlabel metal1 34914 13498 34914 13498 0 _0999_
rlabel metal1 35282 13362 35282 13362 0 _1000_
rlabel metal1 34270 9588 34270 9588 0 _1001_
rlabel metal1 35098 10710 35098 10710 0 _1002_
rlabel metal1 33626 24684 33626 24684 0 _1003_
rlabel metal2 34362 10897 34362 10897 0 _1004_
rlabel metal2 33810 11424 33810 11424 0 _1005_
rlabel metal1 34684 10642 34684 10642 0 _1006_
rlabel metal1 35420 20842 35420 20842 0 _1007_
rlabel metal1 34408 11118 34408 11118 0 _1008_
rlabel metal1 33626 11322 33626 11322 0 _1009_
rlabel metal1 33764 20434 33764 20434 0 _1010_
rlabel metal1 33350 13226 33350 13226 0 _1011_
rlabel metal2 31878 14620 31878 14620 0 _1012_
rlabel via3 34707 20740 34707 20740 0 _1013_
rlabel metal1 35328 11866 35328 11866 0 _1014_
rlabel metal2 31694 12823 31694 12823 0 _1015_
rlabel metal1 32200 12206 32200 12206 0 _1016_
rlabel metal2 31510 17952 31510 17952 0 _1017_
rlabel metal1 30498 22508 30498 22508 0 _1018_
rlabel metal2 30314 23290 30314 23290 0 _1019_
rlabel metal1 32016 22678 32016 22678 0 _1020_
rlabel metal2 32338 19108 32338 19108 0 _1021_
rlabel metal2 30682 16150 30682 16150 0 _1022_
rlabel metal1 30544 16082 30544 16082 0 _1023_
rlabel metal2 31602 15674 31602 15674 0 _1024_
rlabel metal2 33166 14433 33166 14433 0 _1025_
rlabel metal1 30268 22202 30268 22202 0 _1026_
rlabel metal2 30774 18904 30774 18904 0 _1027_
rlabel metal1 33074 20366 33074 20366 0 _1028_
rlabel metal2 32246 16830 32246 16830 0 _1029_
rlabel metal1 30774 23086 30774 23086 0 _1030_
rlabel metal1 31096 21998 31096 21998 0 _1031_
rlabel metal1 32292 18802 32292 18802 0 _1032_
rlabel metal2 31234 18530 31234 18530 0 _1033_
rlabel metal1 32476 18938 32476 18938 0 _1034_
rlabel metal1 32614 16422 32614 16422 0 _1035_
rlabel metal2 32890 19686 32890 19686 0 _1036_
rlabel metal2 15180 12580 15180 12580 0 _1037_
rlabel metal1 15916 13498 15916 13498 0 _1038_
rlabel metal1 27140 23290 27140 23290 0 _1039_
rlabel metal1 20102 14348 20102 14348 0 _1040_
rlabel metal1 15824 11526 15824 11526 0 _1041_
rlabel metal1 16330 9554 16330 9554 0 _1042_
rlabel metal3 16790 9384 16790 9384 0 _1043_
rlabel metal1 15686 9554 15686 9554 0 _1044_
rlabel metal1 20010 12648 20010 12648 0 _1045_
rlabel metal1 15180 7786 15180 7786 0 _1046_
rlabel metal1 15456 19822 15456 19822 0 _1047_
rlabel metal1 15410 20026 15410 20026 0 _1048_
rlabel metal2 16146 12036 16146 12036 0 _1049_
rlabel metal1 19366 12376 19366 12376 0 _1050_
rlabel metal1 16008 12614 16008 12614 0 _1051_
rlabel metal1 16376 15674 16376 15674 0 _1052_
rlabel metal2 15502 14314 15502 14314 0 _1053_
rlabel metal2 15686 12988 15686 12988 0 _1054_
rlabel metal2 15318 15402 15318 15402 0 _1055_
rlabel metal1 16192 15470 16192 15470 0 _1056_
rlabel metal1 16790 21522 16790 21522 0 _1057_
rlabel metal2 15226 17204 15226 17204 0 _1058_
rlabel metal1 16836 18938 16836 18938 0 _1059_
rlabel metal1 19642 21352 19642 21352 0 _1060_
rlabel metal2 16330 15266 16330 15266 0 _1061_
rlabel metal1 16008 15538 16008 15538 0 _1062_
rlabel metal2 15042 16592 15042 16592 0 _1063_
rlabel metal1 14122 17000 14122 17000 0 _1064_
rlabel metal1 15916 20570 15916 20570 0 _1065_
rlabel metal2 16054 15130 16054 15130 0 _1066_
rlabel metal2 19734 16762 19734 16762 0 _1067_
rlabel metal2 21390 17952 21390 17952 0 _1068_
rlabel metal2 21758 17340 21758 17340 0 _1069_
rlabel metal1 16054 17272 16054 17272 0 _1070_
rlabel metal1 17388 16762 17388 16762 0 _1071_
rlabel metal1 17572 16558 17572 16558 0 _1072_
rlabel metal2 16422 14144 16422 14144 0 _1073_
rlabel metal1 17710 14552 17710 14552 0 _1074_
rlabel metal1 17940 14790 17940 14790 0 _1075_
rlabel metal1 17802 16422 17802 16422 0 _1076_
rlabel metal1 20102 27472 20102 27472 0 _1077_
rlabel metal1 21298 28424 21298 28424 0 _1078_
rlabel via1 22585 28526 22585 28526 0 _1079_
rlabel metal1 22540 24718 22540 24718 0 _1080_
rlabel viali 19734 23834 19734 23834 0 _1081_
rlabel metal2 19550 23562 19550 23562 0 _1082_
rlabel metal1 20240 23494 20240 23494 0 _1083_
rlabel metal3 14789 19244 14789 19244 0 _1084_
rlabel metal2 13938 16830 13938 16830 0 _1085_
rlabel metal1 17066 12784 17066 12784 0 _1086_
rlabel metal1 18768 12818 18768 12818 0 _1087_
rlabel metal1 13892 21998 13892 21998 0 _1088_
rlabel metal2 12466 22270 12466 22270 0 _1089_
rlabel metal1 12190 23596 12190 23596 0 _1090_
rlabel metal1 16790 20910 16790 20910 0 _1091_
rlabel metal1 18032 21114 18032 21114 0 _1092_
rlabel metal1 21114 28934 21114 28934 0 _1093_
rlabel metal2 20654 29308 20654 29308 0 _1094_
rlabel metal1 20654 29206 20654 29206 0 _1095_
rlabel metal1 21574 28560 21574 28560 0 _1096_
rlabel metal1 18952 22474 18952 22474 0 _1097_
rlabel metal2 17710 8092 17710 8092 0 _1098_
rlabel metal2 14674 12002 14674 12002 0 _1099_
rlabel metal1 15318 12342 15318 12342 0 _1100_
rlabel metal2 18722 16354 18722 16354 0 _1101_
rlabel metal1 16928 12614 16928 12614 0 _1102_
rlabel metal1 16882 12104 16882 12104 0 _1103_
rlabel metal1 17710 12682 17710 12682 0 _1104_
rlabel metal1 18676 9350 18676 9350 0 _1105_
rlabel metal2 18446 11968 18446 11968 0 _1106_
rlabel metal2 18078 12614 18078 12614 0 _1107_
rlabel metal1 18538 12954 18538 12954 0 _1108_
rlabel metal1 16974 29750 16974 29750 0 _1109_
rlabel metal1 21252 26486 21252 26486 0 _1110_
rlabel metal2 20930 22916 20930 22916 0 _1111_
rlabel metal1 20378 22644 20378 22644 0 _1112_
rlabel metal1 19734 22610 19734 22610 0 _1113_
rlabel metal1 15134 16014 15134 16014 0 _1114_
rlabel metal1 19780 18054 19780 18054 0 _1115_
rlabel metal2 19918 19278 19918 19278 0 _1116_
rlabel metal1 16698 23052 16698 23052 0 _1117_
rlabel metal1 20010 19958 20010 19958 0 _1118_
rlabel metal1 15640 21114 15640 21114 0 _1119_
rlabel metal1 16790 23154 16790 23154 0 _1120_
rlabel metal2 16422 24106 16422 24106 0 _1121_
rlabel metal1 15824 23698 15824 23698 0 _1122_
rlabel metal1 15364 25670 15364 25670 0 _1123_
rlabel metal1 15686 21964 15686 21964 0 _1124_
rlabel metal2 15502 22916 15502 22916 0 _1125_
rlabel via1 13940 26962 13940 26962 0 _1126_
rlabel metal1 12282 29104 12282 29104 0 _1127_
rlabel metal1 15318 25330 15318 25330 0 _1128_
rlabel metal1 13524 24786 13524 24786 0 _1129_
rlabel via1 16695 27438 16695 27438 0 _1130_
rlabel metal1 16974 27846 16974 27846 0 _1131_
rlabel metal2 14122 24582 14122 24582 0 _1132_
rlabel metal2 13018 23834 13018 23834 0 _1133_
rlabel metal1 22770 23256 22770 23256 0 _1134_
rlabel metal1 19458 23596 19458 23596 0 _1135_
rlabel metal1 18492 22950 18492 22950 0 _1136_
rlabel metal1 17342 15674 17342 15674 0 _1137_
rlabel metal1 20286 18224 20286 18224 0 _1138_
rlabel metal1 17572 19754 17572 19754 0 _1139_
rlabel metal1 16882 10676 16882 10676 0 _1140_
rlabel metal1 17296 14246 17296 14246 0 _1141_
rlabel metal1 16283 11118 16283 11118 0 _1142_
rlabel metal2 17434 9588 17434 9588 0 _1143_
rlabel metal1 17526 10710 17526 10710 0 _1144_
rlabel via2 17342 10013 17342 10013 0 _1145_
rlabel metal2 17986 21369 17986 21369 0 _1146_
rlabel metal1 12190 21454 12190 21454 0 _1147_
rlabel metal2 12650 22848 12650 22848 0 _1148_
rlabel metal1 15318 15606 15318 15606 0 _1149_
rlabel metal1 14444 17306 14444 17306 0 _1150_
rlabel metal1 12742 23052 12742 23052 0 _1151_
rlabel metal2 12558 23800 12558 23800 0 _1152_
rlabel metal1 12834 20910 12834 20910 0 _1153_
rlabel metal1 12006 22542 12006 22542 0 _1154_
rlabel metal2 10350 24004 10350 24004 0 _1155_
rlabel metal1 14996 21658 14996 21658 0 _1156_
rlabel metal2 14306 22576 14306 22576 0 _1157_
rlabel metal2 19412 21658 19412 21658 0 _1158_
rlabel metal1 14536 21998 14536 21998 0 _1159_
rlabel metal1 11914 22032 11914 22032 0 _1160_
rlabel metal2 12466 24956 12466 24956 0 _1161_
rlabel metal2 9890 22338 9890 22338 0 _1162_
rlabel metal2 27002 22916 27002 22916 0 _1163_
rlabel metal1 26542 22746 26542 22746 0 _1164_
rlabel metal1 20424 10234 20424 10234 0 _1165_
rlabel metal1 26496 23290 26496 23290 0 _1166_
rlabel via1 26013 24378 26013 24378 0 _1167_
rlabel metal1 26358 24378 26358 24378 0 _1168_
rlabel metal2 25622 23868 25622 23868 0 _1169_
rlabel via2 19366 23477 19366 23477 0 _1170_
rlabel metal1 20654 10098 20654 10098 0 _1171_
rlabel metal2 17802 10608 17802 10608 0 _1172_
rlabel metal1 14536 21522 14536 21522 0 _1173_
rlabel metal1 10534 21522 10534 21522 0 _1174_
rlabel metal1 19182 8058 19182 8058 0 _1175_
rlabel metal1 17940 9010 17940 9010 0 _1176_
rlabel metal1 18354 9588 18354 9588 0 _1177_
rlabel metal1 18492 20570 18492 20570 0 _1178_
rlabel metal2 19458 19210 19458 19210 0 _1179_
rlabel metal2 19550 18530 19550 18530 0 _1180_
rlabel metal1 18630 19142 18630 19142 0 _1181_
rlabel metal1 19274 18836 19274 18836 0 _1182_
rlabel metal2 19136 16218 19136 16218 0 _1183_
rlabel metal2 18906 18870 18906 18870 0 _1184_
rlabel metal1 19366 19278 19366 19278 0 _1185_
rlabel metal3 19159 20604 19159 20604 0 _1186_
rlabel metal2 19734 21148 19734 21148 0 _1187_
rlabel via2 19274 20995 19274 20995 0 _1188_
rlabel metal2 9614 20502 9614 20502 0 _1189_
rlabel metal2 16606 14144 16606 14144 0 _1190_
rlabel metal1 23506 16059 23506 16059 0 _1191_
rlabel metal1 24104 15946 24104 15946 0 _1192_
rlabel via2 23874 21437 23874 21437 0 _1193_
rlabel metal2 9430 21930 9430 21930 0 _1194_
rlabel metal1 18538 14382 18538 14382 0 _1195_
rlabel via1 20286 14042 20286 14042 0 _1196_
rlabel metal3 16307 23052 16307 23052 0 _1197_
rlabel metal1 27692 28526 27692 28526 0 _1198_
rlabel metal1 27876 28730 27876 28730 0 _1199_
rlabel metal1 27646 29172 27646 29172 0 _1200_
rlabel via2 19458 23069 19458 23069 0 _1201_
rlabel metal1 14582 22644 14582 22644 0 _1202_
rlabel metal2 14214 22304 14214 22304 0 _1203_
rlabel metal1 6394 22032 6394 22032 0 _1204_
rlabel metal1 8418 20332 8418 20332 0 _1205_
rlabel metal1 8142 20570 8142 20570 0 _1206_
rlabel metal1 4646 19890 4646 19890 0 _1207_
rlabel metal1 8878 19822 8878 19822 0 _1208_
rlabel metal2 7038 20468 7038 20468 0 _1209_
rlabel metal1 6210 22644 6210 22644 0 _1210_
rlabel metal1 9343 23664 9343 23664 0 _1211_
rlabel via1 8052 22610 8052 22610 0 _1212_
rlabel metal2 2530 24208 2530 24208 0 _1213_
rlabel metal1 7334 20400 7334 20400 0 _1214_
rlabel metal1 7958 21556 7958 21556 0 _1215_
rlabel metal2 4554 19873 4554 19873 0 _1216_
rlabel metal1 5244 20026 5244 20026 0 _1217_
rlabel metal3 8924 20876 8924 20876 0 _1218_
rlabel metal1 22310 8296 22310 8296 0 _1219_
rlabel metal2 22494 8908 22494 8908 0 _1220_
rlabel metal2 22678 7072 22678 7072 0 _1221_
rlabel metal1 22356 6970 22356 6970 0 _1222_
rlabel via2 22770 8619 22770 8619 0 _1223_
rlabel metal2 23414 22848 23414 22848 0 _1224_
rlabel metal2 22770 11186 22770 11186 0 _1225_
rlabel metal1 22356 14586 22356 14586 0 _1226_
rlabel metal1 21850 15674 21850 15674 0 _1227_
rlabel metal1 21206 17782 21206 17782 0 _1228_
rlabel metal1 23782 21998 23782 21998 0 _1229_
rlabel metal1 23322 22066 23322 22066 0 _1230_
rlabel metal1 22632 20774 22632 20774 0 _1231_
rlabel metal1 22770 18054 22770 18054 0 _1232_
rlabel metal1 22586 18326 22586 18326 0 _1233_
rlabel metal2 22586 17408 22586 17408 0 _1234_
rlabel metal2 22402 19380 22402 19380 0 _1235_
rlabel metal2 23046 18649 23046 18649 0 _1236_
rlabel metal1 22816 21114 22816 21114 0 _1237_
rlabel metal1 26128 20434 26128 20434 0 _1238_
rlabel metal1 23736 20230 23736 20230 0 _1239_
rlabel metal1 21298 25228 21298 25228 0 _1240_
rlabel metal1 23874 30158 23874 30158 0 _1241_
rlabel metal1 24288 29070 24288 29070 0 _1242_
rlabel metal2 24978 26554 24978 26554 0 _1243_
rlabel metal1 23782 24174 23782 24174 0 _1244_
rlabel metal1 23230 27030 23230 27030 0 _1245_
rlabel metal1 23782 27098 23782 27098 0 _1246_
rlabel metal1 23598 30668 23598 30668 0 _1247_
rlabel metal2 21482 25432 21482 25432 0 _1248_
rlabel metal2 20654 20383 20654 20383 0 _1249_
rlabel metal1 20746 20468 20746 20468 0 _1250_
rlabel metal1 20378 21590 20378 21590 0 _1251_
rlabel metal1 20654 21658 20654 21658 0 _1252_
rlabel metal1 21528 25262 21528 25262 0 _1253_
rlabel metal1 17802 25874 17802 25874 0 _1254_
rlabel metal1 12604 27098 12604 27098 0 _1255_
rlabel metal1 17480 29206 17480 29206 0 _1256_
rlabel metal1 13202 26894 13202 26894 0 _1257_
rlabel metal1 17158 16490 17158 16490 0 _1258_
rlabel metal1 17296 19482 17296 19482 0 _1259_
rlabel metal1 17204 20026 17204 20026 0 _1260_
rlabel metal1 16744 26350 16744 26350 0 _1261_
rlabel metal2 15594 29444 15594 29444 0 _1262_
rlabel metal4 12604 26928 12604 26928 0 _1263_
rlabel metal1 10212 23834 10212 23834 0 _1264_
rlabel metal2 3910 20026 3910 20026 0 _1265_
rlabel metal1 10213 12206 10213 12206 0 _1266_
rlabel metal1 13110 18156 13110 18156 0 _1267_
rlabel metal1 19550 28560 19550 28560 0 _1268_
rlabel metal1 15502 17136 15502 17136 0 _1269_
rlabel metal1 16054 14518 16054 14518 0 _1270_
rlabel metal1 18354 16456 18354 16456 0 _1271_
rlabel metal1 16192 16762 16192 16762 0 _1272_
rlabel metal2 20378 16830 20378 16830 0 _1273_
rlabel metal1 15870 16218 15870 16218 0 _1274_
rlabel metal1 15594 16762 15594 16762 0 _1275_
rlabel metal1 12834 17102 12834 17102 0 _1276_
rlabel metal1 11868 18734 11868 18734 0 _1277_
rlabel metal2 17066 17340 17066 17340 0 _1278_
rlabel metal2 17158 17374 17158 17374 0 _1279_
rlabel metal1 12834 17612 12834 17612 0 _1280_
rlabel metal2 12190 16898 12190 16898 0 _1281_
rlabel metal1 14076 12614 14076 12614 0 _1282_
rlabel metal1 13018 17850 13018 17850 0 _1283_
rlabel metal1 11132 18666 11132 18666 0 _1284_
rlabel metal2 12374 18496 12374 18496 0 _1285_
rlabel metal1 18814 21114 18814 21114 0 _1286_
rlabel metal2 20470 18428 20470 18428 0 _1287_
rlabel metal1 20378 18054 20378 18054 0 _1288_
rlabel metal1 19872 18394 19872 18394 0 _1289_
rlabel metal1 24426 24718 24426 24718 0 _1290_
rlabel metal1 25530 27642 25530 27642 0 _1291_
rlabel metal2 19826 25466 19826 25466 0 _1292_
rlabel metal1 19550 25466 19550 25466 0 _1293_
rlabel metal2 18538 25024 18538 25024 0 _1294_
rlabel via2 20010 25789 20010 25789 0 _1295_
rlabel metal1 19274 26010 19274 26010 0 _1296_
rlabel metal1 9338 25364 9338 25364 0 _1297_
rlabel metal1 24150 17850 24150 17850 0 _1298_
rlabel metal1 23828 23018 23828 23018 0 _1299_
rlabel metal1 19090 24786 19090 24786 0 _1300_
rlabel metal2 18170 24412 18170 24412 0 _1301_
rlabel metal2 9154 24956 9154 24956 0 _1302_
rlabel metal2 17986 26214 17986 26214 0 _1303_
rlabel metal1 8234 29070 8234 29070 0 _1304_
rlabel metal2 18722 25194 18722 25194 0 _1305_
rlabel metal2 18262 27098 18262 27098 0 _1306_
rlabel metal1 18308 27982 18308 27982 0 _1307_
rlabel metal1 18078 29648 18078 29648 0 _1308_
rlabel metal1 7958 29274 7958 29274 0 _1309_
rlabel metal1 8510 28458 8510 28458 0 _1310_
rlabel metal2 16468 29138 16468 29138 0 _1311_
rlabel metal2 9338 29444 9338 29444 0 _1312_
rlabel metal1 11454 32912 11454 32912 0 _1313_
rlabel metal2 4922 32198 4922 32198 0 _1314_
rlabel metal1 11776 12818 11776 12818 0 _1315_
rlabel metal1 10718 9554 10718 9554 0 _1316_
rlabel metal1 10718 9690 10718 9690 0 _1317_
rlabel metal2 13386 25466 13386 25466 0 _1318_
rlabel metal1 13800 25262 13800 25262 0 _1319_
rlabel metal1 12466 23120 12466 23120 0 _1320_
rlabel metal1 11776 23018 11776 23018 0 _1321_
rlabel metal1 9062 23120 9062 23120 0 _1322_
rlabel metal2 5198 23766 5198 23766 0 _1323_
rlabel metal1 5934 23494 5934 23494 0 _1324_
rlabel metal1 6624 21998 6624 21998 0 _1325_
rlabel metal1 9614 22610 9614 22610 0 _1326_
rlabel metal1 13386 26894 13386 26894 0 _1327_
rlabel metal1 10626 22542 10626 22542 0 _1328_
rlabel metal1 9706 22746 9706 22746 0 _1329_
rlabel metal1 3864 23018 3864 23018 0 _1330_
rlabel metal1 10212 12682 10212 12682 0 _1331_
rlabel metal2 13662 8806 13662 8806 0 _1332_
rlabel metal1 8096 26758 8096 26758 0 _1333_
rlabel metal2 8234 26724 8234 26724 0 _1334_
rlabel metal1 11270 31858 11270 31858 0 _1335_
rlabel metal1 10994 32402 10994 32402 0 _1336_
rlabel metal2 11914 18870 11914 18870 0 _1337_
rlabel metal2 12098 19142 12098 19142 0 _1338_
rlabel metal2 10994 14127 10994 14127 0 _1339_
rlabel metal2 10994 12517 10994 12517 0 _1340_
rlabel metal2 9982 10404 9982 10404 0 _1341_
rlabel metal1 10350 11866 10350 11866 0 _1342_
rlabel metal1 10166 9588 10166 9588 0 _1343_
rlabel metal1 9246 8806 9246 8806 0 _1344_
rlabel metal1 4646 23120 4646 23120 0 _1345_
rlabel metal2 4554 21801 4554 21801 0 _1346_
rlabel metal1 5152 21522 5152 21522 0 _1347_
rlabel metal1 9798 21522 9798 21522 0 _1348_
rlabel metal1 10718 25976 10718 25976 0 _1349_
rlabel metal1 9936 25738 9936 25738 0 _1350_
rlabel metal3 644 35722 644 35722 0 clk
rlabel via2 20102 20213 20102 20213 0 clknet_0_clk
rlabel metal1 4324 8942 4324 8942 0 clknet_4_0_0_clk
rlabel metal1 32706 6834 32706 6834 0 clknet_4_10_0_clk
rlabel metal1 27094 11118 27094 11118 0 clknet_4_11_0_clk
rlabel metal1 18262 32436 18262 32436 0 clknet_4_12_0_clk
rlabel metal1 20562 34068 20562 34068 0 clknet_4_13_0_clk
rlabel metal2 34178 26928 34178 26928 0 clknet_4_14_0_clk
rlabel metal1 32154 32436 32154 32436 0 clknet_4_15_0_clk
rlabel metal2 2622 14450 2622 14450 0 clknet_4_1_0_clk
rlabel metal1 13110 8534 13110 8534 0 clknet_4_2_0_clk
rlabel metal1 16100 2482 16100 2482 0 clknet_4_3_0_clk
rlabel metal1 2070 22066 2070 22066 0 clknet_4_4_0_clk
rlabel metal2 1426 27982 1426 27982 0 clknet_4_5_0_clk
rlabel metal1 5244 35122 5244 35122 0 clknet_4_6_0_clk
rlabel metal1 6394 32266 6394 32266 0 clknet_4_7_0_clk
rlabel metal1 18722 3094 18722 3094 0 clknet_4_8_0_clk
rlabel via2 14122 18717 14122 18717 0 clknet_4_9_0_clk
rlabel via2 35558 24123 35558 24123 0 dataBusIn[0]
rlabel via2 35742 25245 35742 25245 0 dataBusIn[1]
rlabel metal1 36248 27438 36248 27438 0 dataBusIn[2]
rlabel metal2 36202 27659 36202 27659 0 dataBusIn[3]
rlabel via2 36202 22525 36202 22525 0 dataBusIn[4]
rlabel metal2 36202 23443 36202 23443 0 dataBusIn[5]
rlabel metal2 36202 26129 36202 26129 0 dataBusIn[6]
rlabel metal2 36110 24361 36110 24361 0 dataBusIn[7]
rlabel metal2 16146 1520 16146 1520 0 dataBusOut[0]
rlabel metal2 12926 1520 12926 1520 0 dataBusOut[1]
rlabel metal2 17434 959 17434 959 0 dataBusOut[2]
rlabel metal2 13570 1520 13570 1520 0 dataBusOut[3]
rlabel metal2 12282 1520 12282 1520 0 dataBusOut[4]
rlabel metal2 11638 1520 11638 1520 0 dataBusOut[5]
rlabel metal2 14214 1520 14214 1520 0 dataBusOut[6]
rlabel metal2 15502 1520 15502 1520 0 dataBusOut[7]
rlabel metal2 25162 1520 25162 1520 0 dataBusSelect
rlabel metal2 12650 33966 12650 33966 0 gpio[0]
rlabel metal2 12282 38158 12282 38158 0 gpio[10]
rlabel metal1 8188 37230 8188 37230 0 gpio[11]
rlabel metal1 10902 36822 10902 36822 0 gpio[12]
rlabel metal1 9568 36142 9568 36142 0 gpio[13]
rlabel metal1 6026 36754 6026 36754 0 gpio[14]
rlabel metal1 6716 34714 6716 34714 0 gpio[15]
rlabel metal2 16790 1299 16790 1299 0 gpio[16]
rlabel metal2 18722 1299 18722 1299 0 gpio[17]
rlabel metal2 24518 1588 24518 1588 0 gpio[18]
rlabel metal1 25898 21590 25898 21590 0 gpio[19]
rlabel metal2 9016 37332 9016 37332 0 gpio[1]
rlabel metal1 14674 5542 14674 5542 0 gpio[20]
rlabel via2 25438 19907 25438 19907 0 gpio[21]
rlabel metal3 36156 21896 36156 21896 0 gpio[22]
rlabel metal3 820 4148 820 4148 0 gpio[23]
rlabel metal1 23828 2822 23828 2822 0 gpio[24]
rlabel metal2 21298 35413 21298 35413 0 gpio[2]
rlabel metal1 9384 32470 9384 32470 0 gpio[3]
rlabel metal2 3726 30736 3726 30736 0 gpio[4]
rlabel metal1 6716 31790 6716 31790 0 gpio[5]
rlabel metal2 7774 37483 7774 37483 0 gpio[6]
rlabel metal1 3266 31790 3266 31790 0 gpio[7]
rlabel metal1 11362 37230 11362 37230 0 gpio[8]
rlabel metal1 7314 35122 7314 35122 0 gpio[9]
rlabel metal1 17572 25874 17572 25874 0 net1
rlabel metal1 16192 4454 16192 4454 0 net10
rlabel metal1 25806 26826 25806 26826 0 net100
rlabel metal2 24426 17119 24426 17119 0 net101
rlabel metal1 23920 19822 23920 19822 0 net102
rlabel metal1 18722 27336 18722 27336 0 net103
rlabel metal1 19136 13226 19136 13226 0 net104
rlabel metal1 17756 12818 17756 12818 0 net105
rlabel metal1 18078 14416 18078 14416 0 net106
rlabel metal1 16100 15130 16100 15130 0 net107
rlabel metal1 17112 11118 17112 11118 0 net108
rlabel metal1 20930 16456 20930 16456 0 net109
rlabel metal1 12834 4046 12834 4046 0 net11
rlabel metal1 26542 29104 26542 29104 0 net110
rlabel metal1 22011 29614 22011 29614 0 net111
rlabel metal2 26634 21930 26634 21930 0 net112
rlabel metal1 19642 29138 19642 29138 0 net113
rlabel metal1 16751 5610 16751 5610 0 net114
rlabel metal1 18223 2346 18223 2346 0 net115
rlabel metal1 19228 5678 19228 5678 0 net116
rlabel metal1 10035 19414 10035 19414 0 net117
rlabel metal1 8793 18326 8793 18326 0 net118
rlabel metal3 15295 18020 15295 18020 0 net119
rlabel metal1 17342 4012 17342 4012 0 net12
rlabel metal2 19366 4182 19366 4182 0 net120
rlabel metal2 34362 7650 34362 7650 0 net121
rlabel metal2 2990 20094 2990 20094 0 net122
rlabel metal2 6762 26112 6762 26112 0 net123
rlabel metal1 5704 28458 5704 28458 0 net124
rlabel metal1 8425 36754 8425 36754 0 net125
rlabel metal1 12275 36822 12275 36822 0 net126
rlabel metal1 14253 20502 14253 20502 0 net127
rlabel metal2 20378 35360 20378 35360 0 net128
rlabel metal1 32837 32470 32837 32470 0 net129
rlabel metal1 13524 3570 13524 3570 0 net13
rlabel metal1 20877 32810 20877 32810 0 net130
rlabel metal3 15801 21556 15801 21556 0 net131
rlabel via1 14380 26350 14380 26350 0 net132
rlabel via2 16790 27421 16790 27421 0 net133
rlabel metal1 19136 2618 19136 2618 0 net134
rlabel metal1 17020 2482 17020 2482 0 net135
rlabel metal1 34316 31450 34316 31450 0 net136
rlabel metal1 25714 3978 25714 3978 0 net137
rlabel metal1 26082 3094 26082 3094 0 net138
rlabel metal2 12742 3264 12742 3264 0 net139
rlabel metal1 12374 2448 12374 2448 0 net14
rlabel metal1 14582 3434 14582 3434 0 net140
rlabel metal2 14950 4352 14950 4352 0 net141
rlabel metal1 3404 19346 3404 19346 0 net142
rlabel metal2 10994 3706 10994 3706 0 net143
rlabel metal1 18124 3502 18124 3502 0 net144
rlabel metal1 18124 4182 18124 4182 0 net145
rlabel metal1 7866 23086 7866 23086 0 net146
rlabel metal1 12098 4250 12098 4250 0 net147
rlabel metal1 15502 5202 15502 5202 0 net148
rlabel metal1 4370 23086 4370 23086 0 net149
rlabel metal1 11960 2414 11960 2414 0 net15
rlabel metal1 15548 18394 15548 18394 0 net150
rlabel metal1 16376 4182 16376 4182 0 net151
rlabel metal2 12834 5848 12834 5848 0 net152
rlabel metal1 7268 18666 7268 18666 0 net153
rlabel metal1 4508 18666 4508 18666 0 net154
rlabel metal1 13938 5746 13938 5746 0 net155
rlabel metal1 3358 20026 3358 20026 0 net156
rlabel metal2 3818 20672 3818 20672 0 net157
rlabel metal2 2346 23936 2346 23936 0 net158
rlabel metal1 3128 22610 3128 22610 0 net159
rlabel metal1 14076 2414 14076 2414 0 net16
rlabel metal2 4462 21760 4462 21760 0 net160
rlabel metal1 28290 28050 28290 28050 0 net161
rlabel metal2 3818 15878 3818 15878 0 net162
rlabel metal1 2645 17578 2645 17578 0 net163
rlabel metal1 5106 16558 5106 16558 0 net164
rlabel metal1 8510 17578 8510 17578 0 net165
rlabel metal1 28750 29138 28750 29138 0 net166
rlabel metal2 6670 17782 6670 17782 0 net167
rlabel metal2 2714 17408 2714 17408 0 net168
rlabel metal1 7866 24174 7866 24174 0 net169
rlabel metal1 15410 2414 15410 2414 0 net17
rlabel metal2 17526 5372 17526 5372 0 net170
rlabel metal1 5336 24106 5336 24106 0 net171
rlabel metal1 6762 25262 6762 25262 0 net172
rlabel metal1 28382 31246 28382 31246 0 net173
rlabel metal1 5796 29274 5796 29274 0 net174
rlabel metal1 4968 28186 4968 28186 0 net175
rlabel metal1 6946 27098 6946 27098 0 net176
rlabel metal2 5198 26520 5198 26520 0 net177
rlabel metal1 28428 32742 28428 32742 0 net178
rlabel metal1 6946 29274 6946 29274 0 net179
rlabel metal1 25254 2380 25254 2380 0 net18
rlabel metal1 33350 31382 33350 31382 0 net180
rlabel metal1 20608 5678 20608 5678 0 net181
rlabel metal2 19274 4862 19274 4862 0 net182
rlabel metal1 13294 20434 13294 20434 0 net183
rlabel metal1 4554 25126 4554 25126 0 net184
rlabel metal2 9430 19142 9430 19142 0 net185
rlabel metal2 6486 15674 6486 15674 0 net186
rlabel metal1 11132 29070 11132 29070 0 net19
rlabel metal1 35374 26418 35374 26418 0 net2
rlabel metal1 17204 35666 17204 35666 0 net20
rlabel metal1 9430 33932 9430 33932 0 net21
rlabel via1 19642 36227 19642 36227 0 net22
rlabel metal1 22908 32946 22908 32946 0 net23
rlabel metal1 17986 27438 17986 27438 0 net24
rlabel metal1 8142 16456 8142 16456 0 net25
rlabel metal1 34454 9622 34454 9622 0 net26
rlabel metal1 31418 8942 31418 8942 0 net27
rlabel metal2 28198 13702 28198 13702 0 net28
rlabel metal1 32338 14960 32338 14960 0 net29
rlabel metal1 16974 28016 16974 28016 0 net3
rlabel metal1 28382 18326 28382 18326 0 net30
rlabel metal1 35192 18734 35192 18734 0 net31
rlabel metal2 29026 21216 29026 21216 0 net32
rlabel metal2 31786 22372 31786 22372 0 net33
rlabel metal2 32338 25364 32338 25364 0 net34
rlabel metal1 28382 31858 28382 31858 0 net35
rlabel metal1 32660 31790 32660 31790 0 net36
rlabel metal1 21390 33524 21390 33524 0 net37
rlabel metal1 13110 32402 13110 32402 0 net38
rlabel metal2 32430 29308 32430 29308 0 net39
rlabel viali 16504 29138 16504 29138 0 net4
rlabel metal1 34546 20434 34546 20434 0 net40
rlabel metal1 14996 21522 14996 21522 0 net41
rlabel metal1 15870 21998 15870 21998 0 net42
rlabel metal2 32522 24497 32522 24497 0 net43
rlabel metal1 17112 5134 17112 5134 0 net44
rlabel metal2 31832 25874 31832 25874 0 net45
rlabel metal1 28152 25126 28152 25126 0 net46
rlabel metal2 33350 24106 33350 24106 0 net47
rlabel metal2 14950 21699 14950 21699 0 net48
rlabel metal1 14168 17238 14168 17238 0 net49
rlabel viali 31234 22613 31234 22613 0 net5
rlabel metal1 13386 11696 13386 11696 0 net50
rlabel metal1 14398 19278 14398 19278 0 net51
rlabel metal1 19504 21998 19504 21998 0 net52
rlabel metal1 32246 28492 32246 28492 0 net53
rlabel metal1 33166 29104 33166 29104 0 net54
rlabel metal1 20608 19686 20608 19686 0 net55
rlabel metal1 17250 17748 17250 17748 0 net56
rlabel metal1 25070 14994 25070 14994 0 net57
rlabel metal1 18216 21930 18216 21930 0 net58
rlabel metal1 17986 17714 17986 17714 0 net59
rlabel metal1 35282 23596 35282 23596 0 net6
rlabel metal1 16146 13396 16146 13396 0 net60
rlabel metal1 24196 27846 24196 27846 0 net61
rlabel metal1 18538 27438 18538 27438 0 net62
rlabel metal1 26496 19822 26496 19822 0 net63
rlabel metal1 32154 22984 32154 22984 0 net64
rlabel metal2 21022 8687 21022 8687 0 net65
rlabel metal1 20470 8330 20470 8330 0 net66
rlabel metal1 30222 9350 30222 9350 0 net67
rlabel metal1 21574 18190 21574 18190 0 net68
rlabel metal2 27416 14382 27416 14382 0 net69
rlabel metal1 14076 25194 14076 25194 0 net7
rlabel metal1 20378 7854 20378 7854 0 net70
rlabel metal1 26588 16082 26588 16082 0 net71
rlabel metal1 26128 18054 26128 18054 0 net72
rlabel metal1 19680 19686 19680 19686 0 net73
rlabel metal1 32476 8942 32476 8942 0 net74
rlabel metal1 20102 8500 20102 8500 0 net75
rlabel metal1 21052 6698 21052 6698 0 net76
rlabel metal1 20930 11322 20930 11322 0 net77
rlabel metal1 23046 7310 23046 7310 0 net78
rlabel metal2 27186 22100 27186 22100 0 net79
rlabel metal1 12742 29546 12742 29546 0 net8
rlabel metal1 27048 19346 27048 19346 0 net80
rlabel metal1 29440 7990 29440 7990 0 net81
rlabel metal1 26220 8398 26220 8398 0 net82
rlabel metal2 28566 8330 28566 8330 0 net83
rlabel metal1 30084 8534 30084 8534 0 net84
rlabel metal1 27600 6766 27600 6766 0 net85
rlabel metal1 29762 7888 29762 7888 0 net86
rlabel metal1 34362 8330 34362 8330 0 net87
rlabel metal1 21482 7378 21482 7378 0 net88
rlabel metal2 28842 7616 28842 7616 0 net89
rlabel metal1 20286 4522 20286 4522 0 net9
rlabel metal2 31786 7616 31786 7616 0 net90
rlabel metal1 26588 6766 26588 6766 0 net91
rlabel metal1 32062 7820 32062 7820 0 net92
rlabel via1 18336 19346 18336 19346 0 net93
rlabel metal2 17664 23086 17664 23086 0 net94
rlabel metal1 17296 12954 17296 12954 0 net95
rlabel metal1 18584 8466 18584 8466 0 net96
rlabel metal1 23138 10030 23138 10030 0 net97
rlabel metal1 24380 11526 24380 11526 0 net98
rlabel metal2 21206 14144 21206 14144 0 net99
rlabel via2 36110 3451 36110 3451 0 nrst
rlabel metal1 19642 11118 19642 11118 0 top8227.PSRCurrentValue\[0\]
rlabel metal3 13800 16524 13800 16524 0 top8227.PSRCurrentValue\[1\]
rlabel via2 17342 7395 17342 7395 0 top8227.PSRCurrentValue\[2\]
rlabel metal3 13961 18020 13961 18020 0 top8227.PSRCurrentValue\[3\]
rlabel metal2 14122 9537 14122 9537 0 top8227.PSRCurrentValue\[6\]
rlabel metal2 14858 8449 14858 8449 0 top8227.PSRCurrentValue\[7\]
rlabel metal2 12558 20196 12558 20196 0 top8227.branchBackward
rlabel metal2 15778 19992 15778 19992 0 top8227.branchForward
rlabel metal2 30682 32572 30682 32572 0 top8227.demux.isAddressing
rlabel metal3 17204 17204 17204 17204 0 top8227.demux.nmi
rlabel metal1 17802 29716 17802 29716 0 top8227.demux.reset
rlabel metal3 16652 21692 16652 21692 0 top8227.demux.setInterruptFlag
rlabel metal1 34293 32334 34293 32334 0 top8227.demux.state_machine.currentAddress\[0\]
rlabel metal1 30130 29716 30130 29716 0 top8227.demux.state_machine.currentAddress\[10\]
rlabel metal1 28888 31314 28888 31314 0 top8227.demux.state_machine.currentAddress\[11\]
rlabel metal1 20792 28458 20792 28458 0 top8227.demux.state_machine.currentAddress\[12\]
rlabel metal1 33718 30294 33718 30294 0 top8227.demux.state_machine.currentAddress\[1\]
rlabel metal1 31050 31994 31050 31994 0 top8227.demux.state_machine.currentAddress\[2\]
rlabel metal1 28566 32266 28566 32266 0 top8227.demux.state_machine.currentAddress\[3\]
rlabel metal2 26910 28832 26910 28832 0 top8227.demux.state_machine.currentAddress\[4\]
rlabel metal2 26910 27812 26910 27812 0 top8227.demux.state_machine.currentAddress\[5\]
rlabel metal1 23184 29138 23184 29138 0 top8227.demux.state_machine.currentAddress\[6\]
rlabel metal1 23506 29036 23506 29036 0 top8227.demux.state_machine.currentAddress\[7\]
rlabel metal1 34914 31858 34914 31858 0 top8227.demux.state_machine.currentAddress\[8\]
rlabel metal1 31510 31110 31510 31110 0 top8227.demux.state_machine.currentAddress\[9\]
rlabel metal2 34178 7174 34178 7174 0 top8227.demux.state_machine.currentInstruction\[0\]
rlabel metal1 34224 6426 34224 6426 0 top8227.demux.state_machine.currentInstruction\[1\]
rlabel metal1 35098 7514 35098 7514 0 top8227.demux.state_machine.currentInstruction\[2\]
rlabel metal1 34224 6970 34224 6970 0 top8227.demux.state_machine.currentInstruction\[3\]
rlabel metal1 29992 8942 29992 8942 0 top8227.demux.state_machine.currentInstruction\[4\]
rlabel metal2 30222 6715 30222 6715 0 top8227.demux.state_machine.currentInstruction\[5\]
rlabel metal1 26036 16694 26036 16694 0 top8227.demux.state_machine.timeState\[0\]
rlabel metal1 17526 16116 17526 16116 0 top8227.demux.state_machine.timeState\[1\]
rlabel metal1 24518 4046 24518 4046 0 top8227.demux.state_machine.timeState\[2\]
rlabel metal1 24656 22066 24656 22066 0 top8227.demux.state_machine.timeState\[3\]
rlabel metal1 26772 4794 26772 4794 0 top8227.demux.state_machine.timeState\[4\]
rlabel metal1 20838 7446 20838 7446 0 top8227.demux.state_machine.timeState\[5\]
rlabel metal1 23414 4794 23414 4794 0 top8227.demux.state_machine.timeState\[6\]
rlabel metal2 16606 18564 16606 18564 0 top8227.freeCarry
rlabel metal2 17158 3230 17158 3230 0 top8227.instructionLoader.interruptInjector.interruptRequest
rlabel metal1 19734 5678 19734 5678 0 top8227.instructionLoader.interruptInjector.irqGenerated
rlabel metal2 20470 4658 20470 4658 0 top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
rlabel metal1 19780 2482 19780 2482 0 top8227.instructionLoader.interruptInjector.irqSync.nextQ2
rlabel metal1 19136 4726 19136 4726 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
rlabel metal1 18584 3502 18584 3502 0 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
rlabel metal1 15548 2958 15548 2958 0 top8227.instructionLoader.interruptInjector.nmiSync.in
rlabel metal1 16652 2958 16652 2958 0 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2
rlabel metal2 24886 30192 24886 30192 0 top8227.instructionLoader.interruptInjector.resetDetected
rlabel metal2 6026 25092 6026 25092 0 top8227.internalDataflow.accRegToDB\[0\]
rlabel metal1 12650 24140 12650 24140 0 top8227.internalDataflow.accRegToDB\[1\]
rlabel metal2 8142 29784 8142 29784 0 top8227.internalDataflow.accRegToDB\[2\]
rlabel via2 14122 29155 14122 29155 0 top8227.internalDataflow.accRegToDB\[3\]
rlabel metal2 2714 27302 2714 27302 0 top8227.internalDataflow.accRegToDB\[4\]
rlabel via2 13570 26979 13570 26979 0 top8227.internalDataflow.accRegToDB\[5\]
rlabel metal2 6210 26180 6210 26180 0 top8227.internalDataflow.accRegToDB\[6\]
rlabel metal1 3818 28016 3818 28016 0 top8227.internalDataflow.accRegToDB\[7\]
rlabel metal2 20838 34068 20838 34068 0 top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
rlabel metal2 16882 35088 16882 35088 0 top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
rlabel viali 13109 28526 13109 28526 0 top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
rlabel metal1 16330 35054 16330 35054 0 top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
rlabel metal2 19090 34459 19090 34459 0 top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
rlabel metal1 15410 30566 15410 30566 0 top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
rlabel metal1 25438 36006 25438 36006 0 top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
rlabel metal1 25622 34510 25622 34510 0 top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
rlabel metal2 20194 27812 20194 27812 0 top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
rlabel metal1 20562 28696 20562 28696 0 top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
rlabel metal1 18722 30124 18722 30124 0 top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
rlabel metal1 19550 31246 19550 31246 0 top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
rlabel metal1 17894 32266 17894 32266 0 top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
rlabel metal1 14536 31790 14536 31790 0 top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
rlabel metal1 14766 32470 14766 32470 0 top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
rlabel metal1 13294 21114 13294 21114 0 top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
rlabel metal1 5290 15878 5290 15878 0 top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
rlabel metal1 5014 15130 5014 15130 0 top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
rlabel metal1 7360 20502 7360 20502 0 top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
rlabel metal1 4830 20978 4830 20978 0 top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
rlabel metal2 2438 17068 2438 17068 0 top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
rlabel via2 6210 9435 6210 9435 0 top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
rlabel via1 5932 10030 5932 10030 0 top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
rlabel metal1 6164 20502 6164 20502 0 top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
rlabel metal1 5842 25262 5842 25262 0 top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
rlabel metal1 9108 24718 9108 24718 0 top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
rlabel metal1 7590 29206 7590 29206 0 top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
rlabel metal1 5566 28050 5566 28050 0 top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
rlabel metal1 7774 27404 7774 27404 0 top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
rlabel metal1 7682 25670 7682 25670 0 top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
rlabel metal1 5842 26996 5842 26996 0 top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
rlabel metal1 5244 29614 5244 29614 0 top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
rlabel metal1 15400 6970 15400 6970 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
rlabel metal2 12006 7650 12006 7650 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
rlabel metal2 15502 5916 15502 5916 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
rlabel metal1 11684 6426 11684 6426 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
rlabel metal2 13386 6494 13386 6494 0 top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
rlabel metal1 3864 18938 3864 18938 0 top8227.internalDataflow.stackBusModule.busInputs\[32\]
rlabel metal2 8786 17884 8786 17884 0 top8227.internalDataflow.stackBusModule.busInputs\[33\]
rlabel metal1 7728 17714 7728 17714 0 top8227.internalDataflow.stackBusModule.busInputs\[34\]
rlabel metal1 5060 19346 5060 19346 0 top8227.internalDataflow.stackBusModule.busInputs\[35\]
rlabel metal1 4968 17646 4968 17646 0 top8227.internalDataflow.stackBusModule.busInputs\[36\]
rlabel metal1 3266 18394 3266 18394 0 top8227.internalDataflow.stackBusModule.busInputs\[37\]
rlabel metal1 6164 17170 6164 17170 0 top8227.internalDataflow.stackBusModule.busInputs\[38\]
rlabel metal1 4186 16422 4186 16422 0 top8227.internalDataflow.stackBusModule.busInputs\[39\]
rlabel metal2 4002 22372 4002 22372 0 top8227.internalDataflow.stackBusModule.busInputs\[40\]
rlabel metal1 8464 23630 8464 23630 0 top8227.internalDataflow.stackBusModule.busInputs\[41\]
rlabel metal1 6762 18938 6762 18938 0 top8227.internalDataflow.stackBusModule.busInputs\[42\]
rlabel metal1 4462 19958 4462 19958 0 top8227.internalDataflow.stackBusModule.busInputs\[43\]
rlabel metal1 3910 21556 3910 21556 0 top8227.internalDataflow.stackBusModule.busInputs\[44\]
rlabel metal1 3956 23222 3956 23222 0 top8227.internalDataflow.stackBusModule.busInputs\[45\]
rlabel metal2 4554 24004 4554 24004 0 top8227.internalDataflow.stackBusModule.busInputs\[46\]
rlabel via1 4370 20570 4370 20570 0 top8227.internalDataflow.stackBusModule.busInputs\[47\]
rlabel metal1 13248 5338 13248 5338 0 top8227.negEdgeDetector.q1
rlabel metal1 26404 4046 26404 4046 0 top8227.pulse_slower.currentEnableState\[0\]
rlabel metal1 25392 4114 25392 4114 0 top8227.pulse_slower.currentEnableState\[1\]
rlabel metal2 36754 12733 36754 12733 0 top8227.pulse_slower.nextEnableState\[0\]
rlabel metal1 26726 3570 26726 3570 0 top8227.pulse_slower.nextEnableState\[1\]
<< properties >>
string FIXED_BBOX 0 0 37695 39839
<< end >>
