* NGSPICE file created from sample_proj.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt sample_proj VGND VPWR clk done enable nrst out[0] out[10] out[11] out[12]
+ out[13] out[14] out[15] out[16] out[17] out[18] out[19] out[1] out[20] out[21] out[22]
+ out[23] out[24] out[25] out[26] out[27] out[28] out[29] out[2] out[30] out[31] out[32]
+ out[33] out[3] out[4] out[5] out[6] out[7] out[8] out[9] prescaler[0] prescaler[10]
+ prescaler[11] prescaler[12] prescaler[13] prescaler[1] prescaler[2] prescaler[3]
+ prescaler[4] prescaler[5] prescaler[6] prescaler[7] prescaler[8] prescaler[9] stop
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1270_ net66 _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nand2b_1
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0985_ clk_divider.count_out\[15\] _0358_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__nand2_1
XFILLER_41_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0770_ _0133_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__and2b_1
X_1322_ clknet_2_0__leaf_clk clk_divider.next_count\[9\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[9\] sky130_fd_sc_hd__dfrtp_1
X_1253_ _0572_ _0596_ VGND VGND VPWR VPWR clk_divider.next_flag sky130_fd_sc_hd__nor2_1
X_1184_ clk_divider.count_out\[22\] _0522_ clk_divider.count_out\[23\] VGND VGND VPWR
+ VPWR _0533_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0968_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__inv_2
X_0899_ _0273_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__nand2_1
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0822_ _0196_ _0197_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_31_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0684_ _0005_ net14 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__nand2_1
X_0753_ _0099_ _0128_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_24_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1305_ _0617_ _0618_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__nor2_1
X_1236_ _0303_ _0542_ _0577_ _0578_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o2111ai_1
X_1167_ net60 net56 _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or4_1
XFILLER_12_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1098_ net61 net57 net54 _0032_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ _0028_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__xnor2_1
X_0805_ _0173_ _0180_ _0179_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a21o_1
X_0667_ net74 clk_divider.rollover_flag _0044_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__and3_1
X_0736_ _0101_ _0111_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__nor2_1
X_1219_ _0559_ _0560_ _0561_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__or4_1
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1004_ net78 _0035_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nor2_1
X_0719_ _0010_ _0011_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput20 net20 VGND VGND VPWR VPWR out[10] sky130_fd_sc_hd__buf_2
Xoutput31 net31 VGND VGND VPWR VPWR out[20] sky130_fd_sc_hd__buf_2
Xoutput42 net42 VGND VGND VPWR VPWR out[30] sky130_fd_sc_hd__buf_2
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0984_ clk_divider.count_out\[15\] _0358_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
XFILLER_27_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1321_ clknet_2_0__leaf_clk clk_divider.next_count\[8\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[8\] sky130_fd_sc_hd__dfrtp_1
X_1252_ _0576_ _0583_ _0588_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or4_1
X_1183_ clk_divider.count_out\[23\] clk_divider.count_out\[22\] _0522_ VGND VGND VPWR
+ VPWR _0532_ sky130_fd_sc_hd__and3_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0967_ _0238_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__xnor2_2
X_0898_ _0250_ _0253_ _0272_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0821_ _0168_ _0194_ _0149_ _0167_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a211o_1
X_0752_ _0118_ _0126_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__xnor2_2
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ _0056_ _0058_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__nor2_1
X_1304_ _0600_ _0604_ _0620_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__and3_1
X_1235_ _0445_ _0448_ _0449_ net8 VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a211o_1
X_1166_ clk_divider.count_out\[19\] _0509_ clk_divider.count_out\[20\] VGND VGND VPWR
+ VPWR _0518_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1097_ _0461_ VGND VGND VPWR VPWR clk_divider.next_count\[7\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1020_ _0193_ _0395_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__nand2_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0804_ _0170_ _0178_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__xnor2_1
X_0735_ net87 _0109_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__xnor2_1
X_0666_ clk_divider.rollover_flag _0044_ net74 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1218_ _0012_ clk_divider.next_count\[5\] clk_divider.next_count\[6\] _0011_ VGND
+ VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a2bb2o_1
X_1149_ clk_divider.count_out\[17\] clk_divider.count_out\[16\] _0495_ VGND VGND VPWR
+ VPWR _0504_ sky130_fd_sc_hd__and3_1
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1003_ _0012_ clk_divider.count_out\[5\] clk_divider.count_out\[4\] _0013_ VGND VGND
+ VPWR VPWR _0379_ sky130_fd_sc_hd__o22a_1
X_0718_ _0091_ _0093_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0649_ clk_divider.count_out\[12\] VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput32 net32 VGND VGND VPWR VPWR out[21] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR out[11] sky130_fd_sc_hd__buf_2
Xoutput43 net43 VGND VGND VPWR VPWR out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0983_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__inv_2
XFILLER_42_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ clknet_2_0__leaf_clk clk_divider.next_count\[7\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[7\] sky130_fd_sc_hd__dfrtp_2
X_1182_ _0531_ VGND VGND VPWR VPWR clk_divider.next_count\[22\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1251_ _0590_ _0591_ _0592_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__or4_1
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0897_ _0250_ _0253_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a21o_1
X_0966_ _0235_ _0341_ _0233_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0751_ _0118_ _0126_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__nand2_1
X_0820_ _0130_ _0132_ _0148_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__nand3_2
X_1303_ net69 net72 net74 net67 VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__and4b_1
X_0682_ net79 _0057_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__xnor2_2
X_1165_ clk_divider.count_out\[20\] clk_divider.count_out\[19\] _0509_ VGND VGND VPWR
+ VPWR _0517_ sky130_fd_sc_hd__and3_1
X_1234_ net91 _0516_ _0519_ _0521_ _0326_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a311o_1
X_1096_ net88 _0456_ _0459_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_22_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0949_ _0019_ _0321_ _0322_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__nand3_1
XFILLER_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0665_ count\[5\] _0041_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__nand2_1
X_0803_ _0178_ _0170_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__and2b_1
X_0734_ net87 _0109_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__nand2_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1217_ _0391_ clk_divider.next_count\[13\] clk_divider.next_count\[11\] _0367_ VGND
+ VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a2bb2o_1
X_1079_ clk_divider.count_out\[5\] clk_divider.count_out\[4\] _0435_ VGND VGND VPWR
+ VPWR _0446_ sky130_fd_sc_hd__and3_1
X_1148_ _0335_ _0408_ net54 _0023_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a211o_1
XFILLER_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ clk_divider.count_out\[9\] _0373_ _0377_ clk_divider.count_out\[8\] VGND VGND
+ VPWR VPWR _0378_ sky130_fd_sc_hd__a22o_1
X_0717_ _0081_ _0083_ _0090_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__and3_1
X_0648_ clk_divider.count_out\[13\] VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__inv_2
XFILLER_40_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput33 net33 VGND VGND VPWR VPWR out[22] sky130_fd_sc_hd__buf_2
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput22 net22 VGND VGND VPWR VPWR out[12] sky130_fd_sc_hd__buf_2
Xoutput44 net44 VGND VGND VPWR VPWR out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0982_ _0195_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__xnor2_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1250_ _0374_ _0469_ _0470_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o31ai_1
X_1181_ _0527_ _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21o_1
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0896_ net16 _0267_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__xnor2_1
X_0965_ _0196_ _0197_ _0226_ _0241_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_2_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0681_ net87 net15 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__xor2_2
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
X_0750_ _0119_ _0125_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__xnor2_2
X_1302_ _0615_ _0618_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__nor2_1
X_1233_ net88 _0471_ _0474_ _0475_ _0371_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__a311o_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1164_ net61 net57 net54 _0020_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__a211o_1
X_1095_ _0033_ net75 net63 VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__a21o_1
X_0948_ _0321_ _0322_ _0019_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__a21oi_1
X_0879_ _0253_ _0254_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__nand2_1
XFILLER_34_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0802_ _0176_ _0177_ _0175_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__a21oi_1
X_0664_ net73 net71 _0042_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__and3_1
X_0733_ net12 net11 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__xor2_1
X_1216_ _0013_ clk_divider.next_count\[4\] clk_divider.next_count\[11\] _0367_ VGND
+ VGND VPWR VPWR _0560_ sky130_fd_sc_hd__o22ai_1
X_1078_ net62 net58 net53 _0035_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a211o_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1147_ _0024_ net77 _0500_ _0502_ net65 VGND VGND VPWR VPWR clk_divider.next_count\[16\]
+ sky130_fd_sc_hd__a221oi_2
XFILLER_20_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ _0189_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__nand2_1
X_0716_ _0091_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_0647_ clk_divider.count_out\[14\] VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput34 net34 VGND VGND VPWR VPWR out[23] sky130_fd_sc_hd__buf_2
Xoutput23 net23 VGND VGND VPWR VPWR out[13] sky130_fd_sc_hd__buf_2
XFILLER_48_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput45 net45 VGND VGND VPWR VPWR out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ _0149_ _0196_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__and2b_1
XFILLER_8_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1180_ _0018_ net76 net64 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__a21o_1
XFILLER_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0964_ _0314_ _0316_ _0319_ _0339_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__nand4_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0895_ _0269_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout80 net6 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout91 net1 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0680_ net80 _0055_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__nand2_1
X_1301_ _0614_ _0618_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__nor2_1
X_1232_ _0370_ clk_divider.next_count\[10\] _0573_ _0574_ _0575_ VGND VGND VPWR VPWR
+ _0576_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_47_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1094_ net59 net55 _0457_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or4_1
X_1163_ _0514_ _0515_ VGND VGND VPWR VPWR clk_divider.next_count\[19\] sky130_fd_sc_hd__nor2_1
X_0947_ _0321_ _0322_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__nand2_1
X_0878_ _0005_ _0252_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__nand2_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_3_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0801_ _0171_ _0174_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__xor2_1
XFILLER_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0663_ _0041_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
X_0732_ _0008_ _0009_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__nor2_1
X_1146_ net60 net55 _0501_ net90 VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__o31a_1
X_1215_ _0363_ _0494_ _0542_ _0303_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__a22o_1
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ net88 _0441_ _0443_ _0444_ VGND VGND VPWR VPWR clk_divider.next_count\[4\]
+ sky130_fd_sc_hd__a31oi_1
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ net11 net3 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__or2_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0715_ _0081_ _0083_ _0090_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a21oi_1
X_0646_ clk_divider.count_out\[15\] VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__inv_2
X_1129_ _0027_ net75 net63 VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__a21o_1
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput35 net35 VGND VGND VPWR VPWR out[24] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR out[14] sky130_fd_sc_hd__buf_2
Xoutput46 net46 VGND VGND VPWR VPWR out[3] sky130_fd_sc_hd__buf_2
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0629_ net12 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XFILLER_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ _0348_ _0352_ _0355_ _0353_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_32_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0894_ _0262_ _0263_ _0268_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a21o_1
X_0963_ _0324_ _0325_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_2_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout70 net72 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
Xfanout81 net6 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1300_ _0613_ _0618_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__nor2_1
XFILLER_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1231_ _0514_ _0515_ _0344_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__o21ai_1
X_1162_ _0021_ net77 net65 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_47_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1093_ clk_divider.count_out\[7\] _0451_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nor2_1
X_0877_ _0005_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__or2_1
X_0946_ _0092_ _0247_ _0258_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__nand3_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0800_ net78 _0013_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__nor2_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0731_ _0009_ net10 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__nand2_1
X_0662_ count\[4\] _0039_ count\[5\] VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__or3b_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1214_ _0554_ _0556_ _0557_ _0555_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or4b_1
X_1145_ clk_divider.count_out\[16\] _0495_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__xnor2_1
X_1076_ _0036_ net75 net63 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a21o_1
X_0929_ _0300_ _0301_ _0304_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__and3_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0714_ net14 _0088_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__xnor2_1
X_0645_ clk_divider.count_out\[16\] VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
X_1128_ net59 net56 _0486_ net89 VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__o31a_1
X_1059_ net63 _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__nor2_1
XFILLER_15_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput36 net36 VGND VGND VPWR VPWR out[25] sky130_fd_sc_hd__buf_2
Xoutput25 net25 VGND VGND VPWR VPWR out[15] sky130_fd_sc_hd__buf_2
Xoutput47 net47 VGND VGND VPWR VPWR out[4] sky130_fd_sc_hd__buf_2
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0628_ net13 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__inv_2
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0893_ _0262_ _0263_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__nand3_1
X_0962_ _0327_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__nor2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout82 net5 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xfanout60 _0336_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1092_ clk_divider.count_out\[7\] clk_divider.count_out\[6\] _0446_ VGND VGND VPWR
+ VPWR _0457_ sky130_fd_sc_hd__and3_1
X_1230_ _0377_ clk_divider.next_count\[8\] VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nand2_1
X_1161_ _0021_ _0419_ _0513_ _0410_ net90 VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__o221a_1
X_0876_ _0250_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nand2_1
X_0945_ _0092_ _0247_ _0258_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_44_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0661_ _0039_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0730_ _0010_ net9 _0105_ _0103_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__a31o_1
X_1213_ _0425_ _0428_ _0429_ clk_divider.next_count\[0\] _0424_ VGND VGND VPWR VPWR
+ _0557_ sky130_fd_sc_hd__a311o_1
XFILLER_37_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1075_ net59 net55 _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or3_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1144_ net61 _0408_ net54 _0024_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a211o_1
X_0928_ clk_divider.count_out\[24\] _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0859_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__inv_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0713_ net14 _0088_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__and2_1
X_0644_ clk_divider.count_out\[17\] VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__inv_2
X_1127_ clk_divider.count_out\[13\] _0482_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__xnor2_1
X_1058_ net89 net62 net58 _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__and4_1
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput26 net26 VGND VGND VPWR VPWR out[16] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR out[5] sky130_fd_sc_hd__buf_2
Xoutput37 net37 VGND VGND VPWR VPWR out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0627_ net14 VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
XFILLER_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ _0020_ _0326_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__and2_1
X_0892_ net87 _0267_ _0264_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_2_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout72 count\[1\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xfanout61 _0335_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
Xfanout83 net2 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1091_ net62 net58 net53 _0033_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a211o_1
X_1160_ clk_divider.count_out\[19\] _0509_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__xnor2_1
X_0944_ _0314_ _0316_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__and3_1
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0875_ net80 _0004_ _0074_ _0249_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_30_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1289_ _0050_ _0616_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__and2_1
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0660_ net67 net69 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__or2_2
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1212_ _0354_ clk_divider.next_count\[16\] VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__xor2_1
XFILLER_37_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1074_ clk_divider.count_out\[4\] _0435_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__xnor2_1
X_1143_ _0498_ _0499_ VGND VGND VPWR VPWR clk_divider.next_count\[15\] sky130_fd_sc_hd__nor2_1
X_0927_ _0288_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__nor2_1
X_0789_ net3 _0164_ _0163_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__a21boi_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0858_ _0231_ _0232_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0712_ _0084_ _0086_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__xnor2_1
X_0643_ clk_divider.count_out\[18\] VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
X_1126_ net62 net58 net53 _0027_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a211o_1
X_1057_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] clk_divider.count_out\[2\]
+ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__and3_1
Xoutput38 net38 VGND VGND VPWR VPWR out[27] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR out[17] sky130_fd_sc_hd__buf_2
Xoutput49 net49 VGND VGND VPWR VPWR out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0626_ net15 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1109_ net62 net58 net53 _0030_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0960_ _0294_ _0333_ _0334_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or3_1
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0891_ _0265_ _0266_ _0264_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__o21a_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout73 count\[0\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xfanout62 _0335_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xfanout84 net2 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
X_1090_ _0455_ VGND VGND VPWR VPWR clk_divider.next_count\[6\] sky130_fd_sc_hd__inv_2
X_0874_ net80 _0004_ _0074_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__or4_1
X_0943_ clk_divider.count_out\[22\] _0318_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1288_ _0000_ net70 _0049_ _0606_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__and4_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1142_ _0025_ net77 net63 VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__a21o_1
X_1211_ _0363_ _0494_ _0531_ _0318_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__o22a_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1073_ net62 net58 net53 _0036_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_23_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0926_ _0278_ _0282_ _0287_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__and3_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0857_ _0231_ _0232_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__nor2_1
X_0788_ _0161_ _0162_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0711_ _0086_ _0084_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__and2b_1
X_0642_ clk_divider.count_out\[19\] VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__inv_2
X_1125_ _0028_ net77 _0481_ _0484_ net65 VGND VGND VPWR VPWR clk_divider.next_count\[12\]
+ sky130_fd_sc_hd__a221oi_4
X_1056_ _0037_ _0411_ clk_divider.count_out\[2\] VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o21bai_1
Xoutput28 net28 VGND VGND VPWR VPWR out[18] sky130_fd_sc_hd__buf_2
Xoutput39 net39 VGND VGND VPWR VPWR out[28] sky130_fd_sc_hd__buf_2
X_0909_ _0003_ _0261_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__or2_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0625_ net87 VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
XFILLER_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1039_ _0375_ _0378_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or3_1
X_1108_ _0469_ _0470_ VGND VGND VPWR VPWR clk_divider.next_count\[9\] sky130_fd_sc_hd__nor2_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_27_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0890_ net82 _0260_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__and2b_1
XFILLER_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout74 count\[0\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout63 net65 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
Xfanout85 net86 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0873_ net79 _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__xnor2_1
X_0942_ _0308_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__and2_1
XFILLER_9_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1287_ net66 _0606_ _0608_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__and3_1
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1072_ _0042_ counter_to_35.next_count\[0\] counter_to_35.next_count\[1\] VGND VGND
+ VPWR VPWR counter_to_35.next_flag sky130_fd_sc_hd__and3_1
X_1210_ _0430_ _0433_ _0434_ _0425_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a22o_1
X_1141_ _0025_ _0419_ _0497_ _0410_ net89 VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o221a_1
X_0925_ _0290_ _0298_ _0015_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a21o_1
X_0787_ _0161_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__nand2b_1
X_0856_ net11 _0222_ _0221_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a21boi_2
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1339_ clknet_2_2__leaf_clk clk_divider.next_count\[26\] net86 VGND VGND VPWR VPWR
+ clk_divider.count_out\[26\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0710_ net80 _0085_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__xnor2_1
X_0641_ clk_divider.count_out\[20\] VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__inv_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1124_ net59 net55 _0482_ _0483_ net89 VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__o41a_1
X_1055_ _0425_ _0428_ _0429_ VGND VGND VPWR VPWR clk_divider.next_count\[1\] sky130_fd_sc_hd__and3_1
Xoutput29 net29 VGND VGND VPWR VPWR out[19] sky130_fd_sc_hd__buf_2
X_0908_ _0053_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__nand2_1
X_0839_ _0007_ _0008_ _0208_ _0207_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o31ai_4
Xoutput18 net18 VGND VGND VPWR VPWR done sky130_fd_sc_hd__buf_2
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0624_ net79 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ _0382_ _0385_ _0413_ _0379_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or4b_1
X_1107_ _0031_ net76 net64 VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a21o_1
XFILLER_21_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout75 net77 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
Xfanout53 _0418_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
Xfanout64 net65 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_4
Xfanout86 net2 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ _0247_ _0258_ _0275_ _0280_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o211ai_1
X_0872_ net80 net82 net4 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o21ba_1
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1286_ _0605_ _0617_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__nor2_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1071_ count\[4\] _0438_ _0440_ VGND VGND VPWR VPWR counter_to_35.next_count\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ _0495_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or2_1
X_0924_ clk_divider.count_out\[25\] _0289_ _0298_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__or3b_1
X_0855_ net12 _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__xnor2_1
X_0786_ _0095_ _0116_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__xnor2_1
X_1338_ clknet_2_2__leaf_clk clk_divider.next_count\[25\] net86 VGND VGND VPWR VPWR
+ clk_divider.count_out\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1269_ net70 net68 net73 VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_41_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0640_ clk_divider.count_out\[21\] VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__inv_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1123_ clk_divider.count_out\[12\] _0477_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nor2_1
X_1054_ _0037_ _0411_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__nand2_1
XFILLER_18_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0907_ net79 net81 net5 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__a21o_1
Xoutput19 net19 VGND VGND VPWR VPWR out[0] sky130_fd_sc_hd__buf_2
X_0838_ _0199_ _0212_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__xnor2_4
X_0769_ _0108_ _0144_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0623_ clk_divider.count_out\[27\] VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__inv_2
X_1106_ _0031_ _0419_ _0468_ _0410_ net90 VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__o221a_1
XFILLER_42_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1037_ _0013_ clk_divider.count_out\[4\] _0380_ _0412_ VGND VGND VPWR VPWR _0413_
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout76 net77 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_4
Xfanout65 _0426_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
Xfanout54 _0418_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_2
Xfanout87 net16 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_4
X_0940_ clk_divider.count_out\[23\] _0313_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_1
X_0871_ _0242_ _0245_ _0094_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a21o_1
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1285_ net74 net72 net69 net67 VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or4bb_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1070_ count\[4\] _0438_ net17 VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__a21oi_1
X_0923_ _0290_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__nand2_1
X_0854_ _0227_ _0228_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__xor2_1
X_0785_ _0011_ _0012_ _0160_ _0159_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__o31a_1
X_1268_ _0605_ _0607_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__nor2_1
X_1337_ clknet_2_2__leaf_clk clk_divider.next_count\[24\] net86 VGND VGND VPWR VPWR
+ clk_divider.count_out\[24\] sky130_fd_sc_hd__dfrtp_1
X_1199_ net61 net57 _0544_ _0545_ net76 VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__a41oi_1
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1122_ clk_divider.count_out\[12\] _0477_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__and2_1
X_1053_ _0037_ _0411_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or2_1
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0906_ _0276_ _0280_ _0281_ _0269_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__o211a_1
X_0837_ _0199_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2_1
X_0699_ _0004_ _0074_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__nand2_1
X_0768_ _0141_ _0142_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__xnor2_2
XFILLER_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0622_ clk_divider.count_out\[0\] VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__inv_2
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _0466_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__or2_1
X_1036_ clk_divider.count_out\[0\] clk_divider.count_out\[1\] clk_divider.count_out\[3\]
+ clk_divider.count_out\[2\] VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__or4_1
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ _0184_ _0192_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_14_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout66 count\[3\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_4
Xfanout77 _0038_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0870_ _0242_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__nand2_1
X_1284_ net68 net70 _0616_ net73 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__and4b_1
X_0999_ _0030_ _0371_ _0374_ _0031_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a22o_1
XFILLER_46_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0922_ net81 _0053_ _0286_ _0288_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a211o_1
X_0853_ _0227_ _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__nand2_1
X_0784_ _0157_ _0158_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__xnor2_1
X_1267_ net74 net67 net71 net69 VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or4b_1
X_1336_ clknet_2_2__leaf_clk clk_divider.next_count\[23\] net86 VGND VGND VPWR VPWR
+ clk_divider.count_out\[23\] sky130_fd_sc_hd__dfrtp_1
X_1198_ clk_divider.count_out\[25\] _0538_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__or2_1
Xinput1 enable VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1121_ net62 net58 net53 _0028_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a211o_1
X_1052_ clk_divider.count_out\[0\] net75 _0419_ _0427_ _0411_ VGND VGND VPWR VPWR
+ clk_divider.next_count\[0\] sky130_fd_sc_hd__o311a_1
XFILLER_33_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0905_ _0273_ _0270_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__nand2b_1
X_0836_ net10 _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__xnor2_4
X_0767_ _0141_ _0142_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__nand2_1
X_0698_ net82 net4 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__nor2_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1319_ clknet_2_0__leaf_clk clk_divider.next_count\[6\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0621_ net73 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__inv_2
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1035_ _0001_ net75 net59 net55 VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or4_1
X_1104_ clk_divider.count_out\[9\] _0463_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nor2_1
X_0819_ _0168_ _0194_ _0167_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__a21o_1
XFILLER_29_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ clk_divider.count_out\[13\] _0391_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout67 count\[3\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xfanout56 _0409_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xfanout78 net8 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1283_ net70 _0040_ _0049_ _0606_ _0610_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o311a_1
X_0998_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__inv_2
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0921_ _0014_ _0292_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__xnor2_2
X_0852_ _0054_ _0070_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__xor2_1
X_0783_ _0157_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nand2_1
X_1335_ clknet_2_2__leaf_clk clk_divider.next_count\[22\] net85 VGND VGND VPWR VPWR
+ clk_divider.count_out\[22\] sky130_fd_sc_hd__dfrtp_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1266_ _0602_ _0605_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__nor2_1
XFILLER_36_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1197_ clk_divider.count_out\[25\] _0538_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_1
Xinput2 nrst VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ net88 _0476_ _0479_ _0480_ VGND VGND VPWR VPWR clk_divider.next_count\[11\]
+ sky130_fd_sc_hd__a31oi_1
X_1051_ _0001_ net75 net63 VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0904_ _0257_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__or2_1
X_0697_ net4 net87 net82 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__o21ai_1
X_0766_ _0008_ net11 _0125_ _0124_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a31o_1
X_0835_ _0200_ _0209_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__xor2_4
X_1318_ clknet_2_0__leaf_clk clk_divider.next_count\[5\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[5\] sky130_fd_sc_hd__dfrtp_1
X_1249_ net88 _0441_ _0443_ _0444_ net3 VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__a311o_1
XFILLER_24_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1103_ clk_divider.count_out\[9\] _0463_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and2_1
X_1034_ _0335_ net57 VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_16_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0818_ _0183_ _0193_ _0169_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__a21oi_2
X_0749_ _0110_ _0123_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__xor2_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1017_ clk_divider.count_out\[13\] _0391_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__nand2_1
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout79 net7 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
Xfanout68 count\[2\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xfanout57 _0408_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1282_ _0605_ _0615_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__nor2_1
X_0997_ _0190_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__or2_1
XFILLER_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0920_ _0294_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__or2_1
X_0851_ _0135_ _0219_ _0218_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a21bo_1
X_0782_ _0104_ _0105_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__xnor2_1
X_1265_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__inv_2
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1334_ clknet_2_2__leaf_clk clk_divider.next_count\[21\] net85 VGND VGND VPWR VPWR
+ clk_divider.count_out\[21\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1196_ net61 net57 net54 _0015_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__a211o_1
Xinput3 prescaler[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1050_ net89 _0350_ _0423_ net17 VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__a31o_1
X_0903_ _0091_ _0256_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__nor2_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0834_ _0200_ _0209_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nand2_1
X_0696_ _0063_ _0065_ _0066_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__o21bai_1
X_0765_ _0134_ _0140_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__xnor2_2
X_1317_ clknet_2_0__leaf_clk clk_divider.next_count\[4\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[4\] sky130_fd_sc_hd__dfrtp_2
X_1248_ _0359_ _0498_ _0499_ _0396_ clk_divider.next_count\[12\] VGND VGND VPWR VPWR
+ _0592_ sky130_fd_sc_hd__o32ai_1
X_1179_ net60 net56 _0528_ net91 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__o31a_1
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1102_ _0032_ net76 _0462_ _0465_ net64 VGND VGND VPWR VPWR clk_divider.next_count\[8\]
+ sky130_fd_sc_hd__a221oi_2
X_1033_ _0306_ _0320_ _0339_ _0407_ _0331_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a41o_1
X_0817_ _0184_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0679_ net15 net14 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__xor2_2
X_0748_ _0110_ _0123_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__nor2_1
XFILLER_44_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1016_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__inv_2
XFILLER_25_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout69 count\[2\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout58 _0408_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1281_ net74 net69 net71 net67 VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__or4bb_1
X_0996_ _0188_ _0189_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_21_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0850_ _0214_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__nor2_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0781_ _0011_ net78 _0156_ _0154_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__a31o_1
X_1264_ _0600_ _0603_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or2_2
Xinput4 prescaler[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_4
X_1333_ clknet_2_3__leaf_clk clk_divider.next_count\[20\] net85 VGND VGND VPWR VPWR
+ clk_divider.count_out\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1195_ _0542_ VGND VGND VPWR VPWR clk_divider.next_count\[24\] sky130_fd_sc_hd__inv_2
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0979_ _0024_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0902_ _0242_ _0245_ _0276_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a211o_1
X_0833_ _0120_ _0208_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__xnor2_2
X_0695_ _0054_ _0070_ _0069_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a21bo_1
X_0764_ _0122_ _0138_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__xor2_2
X_1178_ clk_divider.count_out\[22\] _0522_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__xnor2_1
X_1247_ _0323_ _0525_ _0526_ _0531_ _0318_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a32o_1
X_1316_ clknet_2_1__leaf_clk clk_divider.next_count\[3\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1032_ _0306_ _0320_ _0339_ _0407_ _0331_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a41oi_4
X_1101_ net59 net55 _0463_ _0464_ net88 VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_16_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0816_ _0185_ _0191_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__nor2_1
X_0747_ net4 _0121_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__xnor2_2
XPHY_EDGE_ROW_48_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0678_ _0005_ _0006_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_39_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1015_ _0194_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_4_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
XFILLER_22_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1280_ _0605_ _0614_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__nor2_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ _0152_ _0153_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__xor2_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1263_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__inv_2
Xinput5 prescaler[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
X_1194_ net90 _0537_ _0540_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__a31o_1
X_1332_ clknet_2_2__leaf_clk clk_divider.next_count\[19\] net86 VGND VGND VPWR VPWR
+ clk_divider.count_out\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0978_ _0198_ _0214_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__xor2_4
XFILLER_42_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0901_ _0094_ _0258_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__or2_1
X_0763_ _0122_ _0138_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__nor2_1
X_0832_ _0201_ _0206_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__xnor2_2
X_0694_ _0062_ _0068_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__xor2_1
X_1315_ clknet_2_1__leaf_clk clk_divider.next_count\[2\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[2\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_22_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1177_ net61 net57 net54 _0018_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a211o_1
X_1246_ _0344_ _0514_ _0515_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__o31ai_1
XFILLER_21_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1100_ clk_divider.count_out\[7\] _0451_ clk_divider.count_out\[8\] VGND VGND VPWR
+ VPWR _0464_ sky130_fd_sc_hd__a21oi_1
X_1031_ _0356_ _0402_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_16_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0815_ _0186_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__nand2_1
X_0746_ net4 _0121_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__nand2_1
X_0677_ net79 net80 net82 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__nand3_1
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1229_ _0498_ _0499_ _0359_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1014_ _0169_ _0183_ _0193_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__and3_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0729_ _0097_ _0102_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_4_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0994_ _0191_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__nand2_2
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1331_ clknet_2_3__leaf_clk clk_divider.next_count\[18\] net85 VGND VGND VPWR VPWR
+ clk_divider.count_out\[18\] sky130_fd_sc_hd__dfrtp_1
X_1262_ count\[5\] _0041_ _0598_ _0000_ _0043_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a221o_1
Xinput6 prescaler[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_1193_ _0016_ net76 net64 VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21o_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0977_ clk_divider.count_out\[17\] _0350_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nand2_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0900_ _0271_ _0275_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0693_ _0062_ _0068_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__nand2_1
X_0762_ net82 _0136_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__xnor2_2
X_0831_ _0201_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nand2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ clknet_2_1__leaf_clk clk_divider.next_count\[1\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_1176_ _0525_ _0526_ VGND VGND VPWR VPWR clk_divider.next_count\[21\] sky130_fd_sc_hd__and2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1245_ _0485_ _0487_ _0488_ _0392_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a211o_1
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1030_ _0348_ _0405_ _0404_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__o21a_1
X_0814_ _0188_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0676_ net17 _0052_ VGND VGND VPWR VPWR counter_to_35.next_count\[5\] sky130_fd_sc_hd__nor2_1
X_0745_ net13 net12 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__xor2_2
X_1228_ _0558_ _0563_ _0567_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or4_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1159_ _0022_ net77 net65 _0512_ VGND VGND VPWR VPWR clk_divider.next_count\[18\]
+ sky130_fd_sc_hd__a211oi_2
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1013_ _0030_ _0371_ _0375_ _0388_ _0368_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0659_ net88 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
X_0728_ _0010_ net9 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0993_ _0186_ _0190_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__or2_1
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1261_ _0000_ net66 net68 net70 VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or4b_1
X_1330_ clknet_2_3__leaf_clk clk_divider.next_count\[17\] net85 VGND VGND VPWR VPWR
+ clk_divider.count_out\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput7 prescaler[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_1192_ net60 net56 _0538_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or4_1
X_0976_ clk_divider.count_out\[17\] _0350_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__nor2_1
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0830_ _0202_ _0205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__xnor2_2
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0692_ _0063_ _0067_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__xnor2_1
X_0761_ net82 _0136_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__nand2_1
X_1313_ clknet_2_1__leaf_clk clk_divider.next_count\[0\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_1244_ _0584_ _0585_ _0586_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or4_1
X_1175_ _0019_ net76 net64 VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a21oi_1
X_0959_ _0294_ _0333_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nor3_4
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0813_ net11 net3 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__nand2_1
Xinput10 prescaler[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_4
X_0675_ clk_divider.rollover_flag _0043_ _0051_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__a21bo_1
X_0744_ _0007_ _0008_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__nor2_1
X_1227_ _0345_ clk_divider.next_count\[18\] _0568_ _0569_ _0570_ VGND VGND VPWR VPWR
+ _0571_ sky130_fd_sc_hd__a2111o_1
X_1158_ _0022_ _0419_ _0511_ _0410_ net90 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__o221a_1
XFILLER_29_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1089_ _0450_ _0453_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a21o_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1012_ _0382_ _0387_ _0378_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__o21ba_1
XFILLER_19_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0727_ _0097_ _0102_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0658_ clk_divider.count_out\[1\] VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__inv_2
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0992_ clk_divider.count_out\[11\] _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__nand2_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1260_ net73 _0601_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__nor2_1
X_1191_ clk_divider.count_out\[24\] _0532_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__nor2_1
Xinput8 prescaler[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0975_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__inv_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0760_ net14 net13 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__xor2_2
X_0691_ _0065_ _0066_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__nor2_1
X_1174_ _0019_ _0419_ _0524_ _0410_ net91 VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__o221ai_2
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1243_ net10 _0461_ clk_divider.next_count\[25\] _0299_ VGND VGND VPWR VPWR _0587_
+ sky130_fd_sc_hd__a22o_1
X_1312_ clknet_2_3__leaf_clk clk_divider.next_flag net85 VGND VGND VPWR VPWR clk_divider.rollover_flag
+ sky130_fd_sc_hd__dfrtp_1
X_0889_ _0003_ net82 net4 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__and3_1
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0958_ clk_divider.count_out\[27\] _0291_ _0293_ clk_divider.count_out\[26\] VGND
+ VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o211a_1
XFILLER_23_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0812_ _0174_ _0187_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__nand2_1
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0743_ _0008_ net11 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__nand2_1
Xinput11 prescaler[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_26_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0674_ count\[4\] net66 clk_divider.rollover_flag _0050_ count\[5\] VGND VGND VPWR
+ VPWR _0051_ sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_10_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1226_ _0469_ _0470_ _0374_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__o21a_1
X_1157_ _0509_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__or2_1
XFILLER_32_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1088_ _0034_ net75 net63 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__a21o_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1011_ net10 _0033_ _0381_ _0385_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o221a_1
XFILLER_19_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0726_ net15 _0100_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_4_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0657_ clk_divider.count_out\[4\] VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1209_ clk_divider.count_out\[27\] net90 _0550_ _0553_ _0425_ VGND VGND VPWR VPWR
+ clk_divider.next_count\[27\] sky130_fd_sc_hd__o221a_1
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0709_ net87 _0074_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__nor2_1
XFILLER_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0991_ _0192_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or2_2
XFILLER_39_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1190_ clk_divider.count_out\[24\] _0532_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__and2_1
Xinput9 prescaler[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_4
X_0974_ _0225_ _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_40_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0690_ net79 _0057_ _0064_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__and3_1
X_1311_ _0000_ net71 _0042_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__and3_1
X_1173_ _0522_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__or2_1
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1242_ _0313_ _0535_ _0536_ _0351_ _0508_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__a32o_1
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0888_ _0259_ net79 net4 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__or3b_1
X_0957_ _0301_ _0332_ _0296_ _0297_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a211oi_2
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0673_ net73 net68 net70 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and3_1
X_0811_ _0172_ _0173_ _0008_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__o21ai_1
X_0742_ _0009_ net10 _0113_ _0112_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a31o_1
Xinput12 prescaler[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1087_ net59 net55 _0451_ _0452_ net88 VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__o41a_1
X_1225_ _0291_ clk_divider.next_count\[27\] VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_1
X_1156_ clk_divider.count_out\[18\] _0504_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_43_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ net9 _0034_ _0384_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__or3_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0656_ clk_divider.count_out\[5\] VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__inv_2
X_0725_ net15 _0100_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__nand2_1
X_1208_ net61 net57 _0551_ _0552_ net76 VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__a41o_1
X_1139_ clk_divider.count_out\[15\] _0490_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__nor2_1
XFILLER_25_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0708_ _0072_ _0073_ _0075_ _0078_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ clk_divider.count_out\[22\] VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0990_ _0185_ _0191_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__and2_1
XFILLER_39_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0973_ _0198_ _0214_ _0213_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__o21ai_2
X_1310_ _0000_ net71 _0041_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__nor3_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1241_ _0010_ clk_divider.next_count\[7\] clk_divider.next_count\[12\] _0396_ VGND
+ VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a22o_1
X_1172_ clk_divider.count_out\[21\] _0517_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nor2_1
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0956_ _0303_ _0016_ _0300_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or3b_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0887_ _0259_ _0260_ _0261_ net4 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__a31o_1
XFILLER_46_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0810_ _0176_ _0177_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__xor2_1
XFILLER_14_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 prescaler[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_4
X_0672_ net66 net68 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__and2_1
X_0741_ _0010_ _0011_ _0116_ _0115_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__o31ai_2
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1224_ net64 _0548_ _0549_ _0292_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__o31a_1
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1086_ clk_divider.count_out\[6\] _0446_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__nor2_1
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1155_ clk_divider.count_out\[18\] _0504_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__and2_1
X_0939_ clk_divider.count_out\[23\] _0311_ _0312_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_15_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_38_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0655_ clk_divider.count_out\[6\] VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
X_0724_ net11 net10 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__xor2_1
X_1207_ _0002_ _0014_ _0544_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__or3_1
X_1069_ net67 _0437_ _0439_ VGND VGND VPWR VPWR counter_to_35.next_count\[3\] sky130_fd_sc_hd__o21a_1
X_1138_ clk_divider.count_out\[15\] _0490_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__and2_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0707_ net13 _0082_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0638_ clk_divider.count_out\[23\] VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__inv_2
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0972_ clk_divider.count_out\[19\] _0343_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a21o_1
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1171_ clk_divider.count_out\[21\] _0517_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and2_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1240_ _0299_ clk_divider.next_count\[25\] clk_divider.next_count\[27\] _0291_ VGND
+ VGND VPWR VPWR _0584_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0886_ net4 _0259_ _0260_ _0261_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__nand4_2
X_0955_ _0296_ _0297_ _0305_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and4bb_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 prescaler[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_4
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0740_ _0106_ _0114_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__xnor2_1
X_0671_ net71 _0046_ _0048_ VGND VGND VPWR VPWR counter_to_35.next_count\[1\] sky130_fd_sc_hd__o21ba_1
X_1154_ _0508_ VGND VGND VPWR VPWR clk_divider.next_count\[17\] sky130_fd_sc_hd__inv_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1223_ _0345_ clk_divider.next_count\[18\] _0564_ _0565_ _0566_ VGND VGND VPWR VPWR
+ _0567_ sky130_fd_sc_hd__o2111ai_1
X_1085_ clk_divider.count_out\[6\] _0446_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__and2_1
XFILLER_20_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0938_ _0311_ _0312_ clk_divider.count_out\[23\] VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0869_ _0196_ _0197_ _0226_ _0239_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__a41oi_4
XTAP_TAPCELL_ROW_7_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0723_ _0009_ _0010_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__nor2_1
X_0654_ clk_divider.count_out\[7\] VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__inv_2
X_1137_ _0494_ VGND VGND VPWR VPWR clk_divider.next_count\[14\] sky130_fd_sc_hd__inv_2
X_1206_ clk_divider.count_out\[26\] clk_divider.count_out\[25\] _0538_ clk_divider.count_out\[27\]
+ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__a31o_1
X_1068_ net17 _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__nor2_1
XFILLER_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0706_ _0071_ _0080_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__xor2_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0637_ clk_divider.count_out\[24\] VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ clk_divider.count_out\[19\] _0343_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__o21ai_1
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1170_ _0520_ _0521_ VGND VGND VPWR VPWR clk_divider.next_count\[20\] sky130_fd_sc_hd__nor2_1
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0885_ net80 net82 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__nand2b_1
X_0954_ _0314_ _0319_ _0328_ _0329_ _0315_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__a311o_1
X_1299_ net66 _0050_ _0619_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__and3b_1
XFILLER_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0670_ net71 _0046_ net17 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__a21o_1
Xinput15 prescaler[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1084_ net62 net58 net53 _0034_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a211o_1
X_1153_ _0503_ _0506_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a21o_1
X_1222_ _0525_ _0526_ _0323_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0937_ _0309_ _0310_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__nand2_1
X_0799_ _0171_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__nor2_1
X_0868_ _0236_ _0237_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_7_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0722_ net11 net10 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__nor2_1
X_0653_ clk_divider.count_out\[8\] VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__inv_2
X_1067_ net67 _0437_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__and2_1
X_1136_ _0489_ _0492_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__a21o_1
X_1205_ net61 net57 net54 _0002_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_47_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0636_ clk_divider.count_out\[25\] VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__inv_2
X_0705_ _0071_ _0080_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1119_ _0029_ net75 net65 VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ _0022_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0884_ net79 net80 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
X_0953_ _0017_ _0309_ _0310_ _0318_ _0018_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__a311oi_1
X_1298_ _0611_ _0618_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__nor2_1
XFILLER_23_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 prescaler[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
X_1221_ _0350_ clk_divider.next_count\[17\] VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
XFILLER_37_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1083_ _0445_ _0448_ _0449_ VGND VGND VPWR VPWR clk_divider.next_count\[5\] sky130_fd_sc_hd__a21oi_1
X_1152_ _0023_ net77 net65 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21o_1
X_0936_ _0273_ _0308_ _0271_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a21bo_1
X_0798_ _0008_ _0172_ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_21_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0867_ _0231_ _0232_ _0236_ _0237_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__o22a_1
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0721_ net14 _0096_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__nand2_1
X_0652_ clk_divider.count_out\[9\] VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__inv_2
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1204_ net64 _0548_ _0549_ VGND VGND VPWR VPWR clk_divider.next_count\[26\] sky130_fd_sc_hd__nor3_1
X_1066_ net17 _0436_ _0437_ VGND VGND VPWR VPWR counter_to_35.next_count\[2\] sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_35_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1135_ _0026_ net77 net63 VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a21o_1
X_0919_ clk_divider.count_out\[27\] _0291_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0704_ _0078_ _0079_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nor2_1
X_0635_ clk_divider.count_out\[26\] VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1118_ net59 net55 _0477_ _0478_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__or4_1
X_1049_ net89 _0424_ net17 VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0952_ _0325_ _0327_ _0324_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21o_1
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0883_ net82 net80 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nand2b_1
X_1297_ _0609_ _0618_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__nor2_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 stop VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
X_1220_ _0520_ _0521_ _0326_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__o21ai_1
X_1151_ net60 net56 _0504_ _0505_ net90 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__o41a_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1082_ _0035_ net75 net63 VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a21o_1
X_0935_ _0271_ _0273_ _0308_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__nand3b_1
X_0866_ _0239_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__nand2_1
X_0797_ net78 net3 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__and2_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ net10 net9 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__xor2_1
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0651_ clk_divider.count_out\[10\] VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
X_1134_ net60 net56 _0490_ _0491_ net89 VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__o41a_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1203_ clk_divider.count_out\[26\] net90 VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__nor2_1
X_1065_ net68 net72 _0047_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0918_ clk_divider.count_out\[27\] _0291_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__and2_1
X_0849_ _0223_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_3_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0703_ net87 net15 _0077_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0634_ net3 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1117_ clk_divider.count_out\[10\] _0466_ clk_divider.count_out\[11\] VGND VGND VPWR
+ VPWR _0478_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1048_ _0350_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0882_ _0256_ _0257_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__or2_1
X_0951_ _0020_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nor2_1
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1296_ _0607_ _0618_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1150_ clk_divider.count_out\[16\] _0495_ clk_divider.count_out\[17\] VGND VGND VPWR
+ VPWR _0505_ sky130_fd_sc_hd__a21oi_1
XFILLER_37_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1081_ net59 net55 _0446_ _0447_ net88 VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__o41a_1
X_0934_ _0273_ _0308_ _0271_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a21o_1
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0865_ _0223_ _0224_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a21oi_1
X_0796_ net78 net3 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nor2_1
X_1279_ _0000_ net68 net70 net66 VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or4b_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0650_ clk_divider.count_out\[11\] VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__inv_2
X_1064_ net71 _0047_ net68 VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__a21oi_1
X_1133_ clk_divider.count_out\[13\] _0482_ clk_divider.count_out\[14\] VGND VGND VPWR
+ VPWR _0491_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1202_ _0014_ _0419_ _0547_ _0410_ net90 VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__o221a_1
X_0779_ _0011_ net78 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__nand2_1
X_0848_ net10 _0211_ _0210_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a21boi_4
X_0917_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_9_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0702_ net87 net15 _0077_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__and3_1
X_0633_ net78 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1116_ clk_divider.count_out\[11\] clk_divider.count_out\[10\] _0466_ VGND VGND VPWR
+ VPWR _0477_ sky130_fd_sc_hd__and3_1
X_1047_ _0354_ _0358_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_31_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0881_ _0087_ _0089_ _0255_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__nor3b_1
X_0950_ _0094_ _0246_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__xnor2_2
XFILLER_32_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1295_ _0602_ _0618_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1080_ clk_divider.count_out\[4\] _0435_ clk_divider.count_out\[5\] VGND VGND VPWR
+ VPWR _0447_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0933_ _0271_ _0273_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__nand3_1
X_0795_ net13 _0151_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__xnor2_1
X_0864_ _0199_ _0212_ _0223_ _0224_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__o22a_1
X_1347_ clknet_2_3__leaf_clk counter_to_35.next_count\[5\] net86 VGND VGND VPWR VPWR
+ count\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1278_ _0605_ _0613_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__nor2_1
XFILLER_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1201_ _0014_ _0544_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__xnor2_1
X_1063_ _0425_ _0434_ VGND VGND VPWR VPWR clk_divider.next_count\[3\] sky130_fd_sc_hd__and2_1
X_1132_ clk_divider.count_out\[14\] clk_divider.count_out\[13\] _0482_ VGND VGND VPWR
+ VPWR _0490_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_25_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0916_ net7 _0289_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__o21a_1
XFILLER_33_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0778_ _0152_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__nor2_1
X_0847_ net11 _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__xnor2_4
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0701_ _0072_ _0076_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__xnor2_1
X_0632_ net9 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1115_ net62 net58 net53 _0029_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__a211o_1
X_1046_ _0362_ _0391_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_23_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1029_ _0024_ _0352_ _0354_ _0353_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_12_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ _0087_ _0089_ _0255_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__o21ba_1
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1294_ _0000_ net72 _0040_ _0619_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_18_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0932_ _0247_ _0279_ _0275_ _0257_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a211o_1
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0794_ _0155_ _0156_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__xnor2_1
X_0863_ _0234_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__nor2_1
X_1346_ clknet_2_3__leaf_clk counter_to_35.next_count\[4\] net86 VGND VGND VPWR VPWR
+ count\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1277_ net74 net69 net71 net67 VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__or4b_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1200_ _0015_ net76 _0543_ _0546_ net64 VGND VGND VPWR VPWR clk_divider.next_count\[25\]
+ sky130_fd_sc_hd__a221oi_2
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1062_ clk_divider.count_out\[3\] _0431_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__and2_1
X_1131_ net62 net58 net53 _0026_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a211o_1
XFILLER_18_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0915_ net5 _0288_ net79 net81 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o211ai_4
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0777_ net14 _0096_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__xnor2_1
X_0846_ _0215_ _0220_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__xor2_4
X_1329_ clknet_2_1__leaf_clk clk_divider.next_count\[16\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_42_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0700_ _0073_ _0075_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__nand2_1
X_0631_ net10 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1114_ net88 _0471_ _0474_ _0475_ VGND VGND VPWR VPWR clk_divider.next_count\[10\]
+ sky130_fd_sc_hd__a31oi_1
X_1045_ _0367_ _0370_ _0396_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_23_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0829_ _0137_ _0203_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__xor2_2
XFILLER_21_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1028_ clk_divider.count_out\[19\] _0343_ _0403_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1293_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0931_ _0296_ _0297_ _0305_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__or3b_1
X_0862_ _0236_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0793_ net3 _0164_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__xnor2_1
X_1276_ net68 net70 VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__nor2_1
X_1345_ clknet_2_3__leaf_clk counter_to_35.next_count\[3\] net86 VGND VGND VPWR VPWR
+ count\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1130_ _0485_ _0487_ _0488_ VGND VGND VPWR VPWR clk_divider.next_count\[13\] sky130_fd_sc_hd__a21oi_1
X_1061_ clk_divider.count_out\[3\] _0432_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__xor2_1
X_0914_ _0265_ _0288_ net81 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o21ai_1
X_0845_ _0215_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__nand2_1
X_0776_ net13 _0151_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__nand2_1
X_1259_ count\[5\] _0039_ count\[4\] net72 VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or4b_1
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1328_ clknet_2_1__leaf_clk clk_divider.next_count\[15\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0630_ net11 VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1113_ _0030_ net75 net63 VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a21o_1
X_1044_ _0011_ _0098_ _0172_ _0373_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and4_1
XFILLER_9_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0828_ _0137_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nor2_1
X_0759_ _0006_ _0007_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__nor2_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1027_ clk_divider.count_out\[19\] _0343_ _0345_ clk_divider.count_out\[18\] VGND
+ VGND VPWR VPWR _0403_ sky130_fd_sc_hd__a22o_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1292_ _0600_ _0604_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_18_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0930_ _0296_ _0297_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__nor3b_1
X_0861_ net13 _0082_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0792_ _0165_ _0166_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__xor2_2
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1275_ net66 _0050_ _0606_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__and3b_1
X_1344_ clknet_2_3__leaf_clk counter_to_35.next_count\[2\] net85 VGND VGND VPWR VPWR
+ count\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _0430_ _0433_ VGND VGND VPWR VPWR clk_divider.next_count\[2\] sky130_fd_sc_hd__and2_1
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0913_ _0265_ _0288_ net81 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__o21a_1
X_0844_ _0135_ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__xor2_2
X_0775_ net9 net78 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__xor2_1
X_1258_ _0597_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__or2_1
X_1189_ net61 net57 net54 _0016_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a211o_1
X_1327_ clknet_2_1__leaf_clk clk_divider.next_count\[14\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1043_ net61 net57 net53 VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__a21o_4
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1112_ net59 net55 _0472_ _0473_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__or4_1
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0827_ net80 _0055_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__xnor2_2
X_0758_ _0007_ net12 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__nand2_1
X_0689_ net79 _0057_ _0064_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1026_ _0026_ _0360_ _0363_ _0401_ _0361_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o311a_1
XFILLER_14_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1009_ net9 _0034_ _0383_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a211o_1
XFILLER_41_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1291_ _0598_ _0612_ _0616_ net73 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__and4b_1
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0860_ net12 _0230_ _0229_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__a21boi_2
XFILLER_13_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0791_ _0165_ _0166_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__nor2_1
X_1343_ clknet_2_3__leaf_clk counter_to_35.next_count\[1\] net85 VGND VGND VPWR VPWR
+ count\[1\] sky130_fd_sc_hd__dfrtp_1
X_1274_ _0605_ _0611_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__nor2_1
XFILLER_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0989_ _0360_ _0364_ _0361_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or3b_1
XFILLER_47_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0912_ _0278_ _0282_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a21oi_2
X_0843_ _0216_ _0217_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__xor2_2
X_0774_ _0011_ _0012_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1326_ clknet_2_1__leaf_clk clk_divider.next_count\[13\] net84 VGND VGND VPWR VPWR
+ clk_divider.count_out\[13\] sky130_fd_sc_hd__dfrtp_2
X_1257_ net71 _0039_ count\[4\] VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__o21a_1
X_1188_ _0535_ _0536_ VGND VGND VPWR VPWR clk_divider.next_count\[23\] sky130_fd_sc_hd__and2_1
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1111_ clk_divider.count_out\[10\] _0466_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__nor2_1
X_1042_ _0307_ _0340_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nor3_1
X_0688_ net4 net87 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__xor2_1
X_0826_ _0006_ net13 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__nand2_1
X_0757_ _0009_ _0010_ _0128_ _0127_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__o31a_1
X_1309_ _0000_ count\[5\] _0597_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1025_ _0393_ _0399_ _0400_ _0365_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a31o_1
X_0809_ _0173_ _0180_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1008_ _0010_ clk_divider.count_out\[7\] VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nor2_1
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1290_ net73 _0598_ _0612_ _0616_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__and4bb_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0790_ net78 _0131_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__xnor2_2
X_1273_ _0610_ net73 net68 VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or3b_1
X_1342_ clknet_2_3__leaf_clk counter_to_35.next_count\[0\] net85 VGND VGND VPWR VPWR
+ count\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_36_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0988_ clk_divider.count_out\[14\] _0362_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0911_ _0262_ _0284_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__a21o_1
X_0842_ _0216_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__nand2_1
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0773_ _0130_ _0132_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a21oi_1
X_1256_ net73 _0598_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__and2_1
X_1325_ clknet_2_0__leaf_clk clk_divider.next_count\[12\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1187_ _0017_ net76 net64 VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1110_ clk_divider.count_out\[10\] clk_divider.count_out\[9\] _0463_ VGND VGND VPWR
+ VPWR _0472_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_48_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1041_ _0356_ _0365_ _0398_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or4_1
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0825_ _0007_ net12 _0140_ _0139_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__a31o_1
X_0687_ _0004_ net15 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__nand2_1
X_0756_ net78 _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__nand2_1
X_1308_ count\[4\] net67 _0050_ _0604_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_39_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1239_ _0293_ clk_divider.next_count\[26\] _0580_ _0581_ _0582_ VGND VGND VPWR VPWR
+ _0583_ sky130_fd_sc_hd__a2111o_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1024_ clk_divider.count_out\[12\] _0394_ _0396_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nand3_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0808_ _0181_ _0182_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__xor2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0739_ _0106_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__nand2_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1007_ _0010_ clk_divider.count_out\[7\] clk_divider.count_out\[6\] _0011_ VGND VGND
+ VPWR VPWR _0383_ sky130_fd_sc_hd__a22o_1
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput50 net50 VGND VGND VPWR VPWR out[7] sky130_fd_sc_hd__buf_2
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1272_ net66 net70 VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nand2b_1
X_1341_ clknet_2_3__leaf_clk counter_to_35.next_flag net85 VGND VGND VPWR VPWR net18
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0987_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__inv_2
XFILLER_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0910_ _0262_ _0285_ _0284_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__a21oi_1
X_0841_ _0060_ _0061_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_11_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0772_ net9 _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1255_ count\[5\] _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ _0017_ _0419_ _0534_ _0410_ net90 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__o221ai_4
X_1324_ clknet_2_0__leaf_clk clk_divider.next_count\[11\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[11\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ clk_divider.count_out\[11\] _0367_ _0370_ clk_divider.count_out\[10\] _0415_
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0755_ _0117_ _0129_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__xor2_2
X_0824_ _0008_ _0009_ _0144_ _0143_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__o31ai_4
X_0686_ _0005_ net14 _0061_ _0059_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__a31o_1
XFILLER_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1307_ _0000_ net70 _0049_ _0619_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_39_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1169_ _0020_ net76 net64 VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__a21o_1
X_1238_ clk_divider.next_count\[8\] _0377_ net9 _0455_ VGND VGND VPWR VPWR _0582_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1023_ _0389_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or2_1
X_0807_ _0181_ _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__nand2_1
X_0738_ _0107_ _0113_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0669_ net17 _0045_ _0047_ VGND VGND VPWR VPWR counter_to_35.next_count\[0\] sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1006_ clk_divider.count_out\[8\] _0377_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nor2_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput51 net51 VGND VGND VPWR VPWR out[8] sky130_fd_sc_hd__buf_2
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput40 net40 VGND VGND VPWR VPWR out[29] sky130_fd_sc_hd__buf_2
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1340_ clknet_2_2__leaf_clk clk_divider.next_count\[27\] net86 VGND VGND VPWR VPWR
+ clk_divider.count_out\[27\] sky130_fd_sc_hd__dfrtp_2
X_1271_ _0605_ _0609_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__nor2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ _0168_ _0194_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__xnor2_2
XFILLER_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0840_ _0006_ net13 _0205_ _0204_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a31o_1
X_0771_ _0133_ _0145_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__xnor2_2
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1323_ clknet_2_0__leaf_clk clk_divider.next_count\[10\] net83 VGND VGND VPWR VPWR
+ clk_divider.count_out\[10\] sky130_fd_sc_hd__dfrtp_2
X_1254_ count\[4\] net72 _0039_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nor3_1
X_1185_ _0532_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__or2_1
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0969_ _0235_ _0341_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__xnor2_2
XFILLER_23_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0685_ _0056_ _0058_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__xor2_2
X_0754_ _0117_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__nand2_1
X_0823_ net9 _0147_ _0146_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a21oi_4
X_1306_ net66 _0608_ _0619_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__and3_1
X_1168_ net91 _0516_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__and3_1
X_1099_ clk_divider.count_out\[8\] clk_divider.count_out\[7\] _0451_ VGND VGND VPWR
+ VPWR _0463_ sky130_fd_sc_hd__and3_1
X_1237_ _0535_ _0536_ _0313_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1022_ clk_divider.count_out\[11\] _0367_ _0393_ _0394_ _0397_ VGND VGND VPWR VPWR
+ _0398_ sky130_fd_sc_hd__o2111ai_1
X_0668_ _0043_ _0046_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__and2b_1
X_0806_ _0150_ _0160_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__xnor2_1
X_0737_ _0101_ _0111_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__xor2_1
XFILLER_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ _0379_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__nor2_1
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput52 net52 VGND VGND VPWR VPWR out[9] sky130_fd_sc_hd__buf_2
Xoutput41 net41 VGND VGND VPWR VPWR out[2] sky130_fd_sc_hd__buf_2
Xoutput30 net30 VGND VGND VPWR VPWR out[1] sky130_fd_sc_hd__buf_2
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

