* NGSPICE file created from calculator_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt calculator_top ColOut[0] ColOut[1] ColOut[2] ColOut[3] RowIn[0] RowIn[1] RowIn[2]
+ RowIn[3] VGND VPWR clk complete display_output[0] display_output[10] display_output[11]
+ display_output[12] display_output[13] display_output[14] display_output[15] display_output[1]
+ display_output[2] display_output[3] display_output[4] display_output[5] display_output[6]
+ display_output[7] display_output[8] display_output[9] input_state_FPGA[0] input_state_FPGA[1]
+ input_state_FPGA[2] key_pressed nRST
X_2106_ input_ctrl_inst.debounce_cnt\[14\] _1057_ _1146_ VGND VGND VPWR VPWR _1164_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2037_ gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1 _1074_ VGND VGND
+ VPWR VPWR _1111_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_20_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1270_ gencon_inst.operand1\[10\] _0605_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_42_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1606_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0827_ VGND VGND
+ VPWR VPWR _0828_ sky130_fd_sc_hd__nor2_1
X_2724_ clknet_leaf_20_clk _0278_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2655_ clknet_leaf_28_clk net336 net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout105 net108 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xfanout149 net150 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
Xfanout116 net117 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
X_1468_ net396 net89 _0705_ net101 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a22o_1
X_1537_ gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__and2_1
Xfanout138 net157 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_4
Xfanout127 net137 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
X_2586_ clknet_leaf_31_clk _0145_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1399_ gencon_inst.mult_calc.out\[8\] net404 net104 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
Xhold170 input_ctrl_inst.scan_timer\[10\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2 VGND VGND VPWR
+ VPWR net349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold181 gencon_inst.mult_calc.compCount.in2\[1\] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2440_ clknet_leaf_1_clk _0038_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1253_ gencon_inst.operand1\[6\] net35 _0595_ _0596_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__o22a_1
X_1322_ gencon_inst.operand2\[4\] _0644_ _0647_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__or3_1
X_2371_ input_ctrl_inst.col_index\[13\] _0515_ net420 VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2707_ clknet_leaf_19_clk _0261_ net155 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2569_ clknet_leaf_21_clk _0132_ net152 VGND VGND VPWR VPWR gencon_inst.operand2\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_2638_ clknet_leaf_26_clk _0197_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1871_ net162 _0954_ _0985_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21ai_1
X_1940_ gencon_inst.operand2\[12\] net64 net41 net340 VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__a22o_1
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2423_ input_ctrl_inst.col_index\[30\] _0550_ _0523_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_67_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1236_ _0580_ _0581_ _0573_ _0576_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__a211o_1
X_1305_ gencon_inst.operand2\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0638_ sky130_fd_sc_hd__and2_1
X_2285_ _0445_ _0470_ _0472_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__and3_1
X_2354_ net310 _0506_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_50_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2070_ _1136_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__inv_2
XFILLER_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1854_ gencon_inst.operand1\[11\] net267 net62 VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
X_1785_ gencon_inst.operand2\[0\] gencon_inst.operand1\[0\] net76 VGND VGND VPWR VPWR
+ _0961_ sky130_fd_sc_hd__mux2_1
X_1923_ gencon_inst.operand2\[14\] _1204_ net74 gencon_inst.ALU_out\[14\] VGND VGND
+ VPWR VPWR _1021_ sky130_fd_sc_hd__a22o_1
X_2406_ input_ctrl_inst.col_index\[25\] _0537_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__xor2_1
X_1219_ _0562_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nor2_1
X_2268_ input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[8\] _0459_ VGND
+ VGND VPWR VPWR _0462_ sky130_fd_sc_hd__and3_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2199_ input_ctrl_inst.col_index\[25\] input_ctrl_inst.col_index\[27\] input_ctrl_inst.col_index\[26\]
+ input_ctrl_inst.col_index\[29\] VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or4_1
X_2337_ net95 net262 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1
+ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a22o_1
XFILLER_71_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold63 gencon_inst.ALU_in2\[9\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 gencon_inst.ALU_in1\[0\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold41 gencon_inst.mult_calc.INn2\[15\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1 VGND VGND VPWR VPWR
+ net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 gencon_inst.mult_calc.INn2\[3\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold85 gencon_inst.mult_calc.INn1\[15\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _0068_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1570_ net107 gencon_inst.add_calc.main.in2\[10\] VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nand2_1
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2122_ input_ctrl_inst.debounce_cnt\[17\] _1173_ input_ctrl_inst.debounce_cnt\[18\]
+ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__a21oi_1
X_2053_ _1047_ _1048_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__nand2_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1837_ gencon_inst.operand2\[10\] net202 net62 VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
X_1768_ gencon_inst.ALU_in2\[12\] gencon_inst.ALU_in1\[12\] net69 VGND VGND VPWR VPWR
+ _0948_ sky130_fd_sc_hd__mux2_1
X_1906_ net66 _0970_ net57 gencon_inst.mult_calc.out\[8\] VGND VGND VPWR VPWR _1010_
+ sky130_fd_sc_hd__a22o_1
X_1699_ _0852_ _0906_ _0908_ net85 VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a31o_1
XFILLER_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput20 net20 VGND VGND VPWR VPWR display_output[3] sky130_fd_sc_hd__buf_2
Xoutput7 net7 VGND VGND VPWR VPWR ColOut[1] sky130_fd_sc_hd__buf_2
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1622_ _0793_ _0797_ _0842_ _0794_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__o31a_1
X_2740_ clknet_leaf_21_clk _0294_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2671_ clknet_leaf_27_clk _0230_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1553_ net441 _0775_ net113 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
X_1484_ gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nand2_1
X_2105_ input_ctrl_inst.debounce_cnt\[13\] input_ctrl_inst.debounce_cnt\[14\] _1157_
+ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__and3_1
X_2036_ gencon_inst.mult_calc.compCount.in2\[10\] _1105_ _1109_ gencon_inst.mult_calc.compCount.in2\[11\]
+ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__o22a_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2723_ clknet_leaf_20_clk _0277_ net155 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1605_ gencon_inst.add_calc.main.in2\[1\] net105 VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__xor2_1
X_1536_ gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__nor2_1
X_2585_ clknet_leaf_31_clk _0144_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2654_ clknet_leaf_28_clk _0213_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout106 net108 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
Xfanout128 net129 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
Xfanout117 _1031_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
X_1398_ gencon_inst.mult_calc.out\[7\] net296 net104 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
X_1467_ _0702_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__xnor2_1
Xfanout139 net157 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_4
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2019_ gencon_inst.mult_calc.compCount.in2\[3\] _1083_ _1092_ gencon_inst.mult_calc.compCount.in2\[4\]
+ _1091_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_19_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold182 gencon_inst.add_calc.main.in2\[13\] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 _0185_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _0173_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 gencon_inst.mult_calc.compCount.in2\[5\] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1252_ gencon_inst.ALU_out\[6\] net71 net51 gencon_inst.mult_calc.out\[6\] net43
+ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a221o_1
X_1321_ _0387_ _0651_ net47 VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2370_ net351 _0515_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__xor2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2706_ clknet_leaf_19_clk _0260_ net155 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ clknet_leaf_23_clk _0131_ net153 VGND VGND VPWR VPWR gencon_inst.operand2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2637_ clknet_leaf_25_clk _0196_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1519_ _0747_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2499_ clknet_leaf_28_clk net263 net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1870_ _0953_ _0984_ _0983_ _0388_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2422_ net434 net54 _0523_ _0551_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a22o_1
X_2353_ _0505_ _0506_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nor2_1
X_1235_ _0573_ _0576_ _0580_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__o211a_1
X_1304_ gencon_inst.operand2\[1\] _0637_ net47 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
X_2284_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__inv_2
XFILLER_52_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1999_ gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
+ _1072_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__and3_1
XFILLER_75_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ _1019_ _1020_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__or2_1
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1853_ gencon_inst.operand1\[10\] net233 net62 VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
X_1784_ net39 VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__inv_2
XFILLER_69_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2405_ input_ctrl_inst.col_index\[25\] net54 VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__and2_1
X_2336_ net95 net268 net80 net275 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__a22o_1
X_1218_ gencon_inst.operand1\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0567_ sky130_fd_sc_hd__xnor2_1
X_2267_ input_ctrl_inst.scan_timer\[7\] _0459_ input_ctrl_inst.scan_timer\[8\] VGND
+ VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a21o_1
XFILLER_25_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2198_ input_ctrl_inst.col_index\[24\] _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nor2_1
XFILLER_52_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold64 gencon_inst.ALU_in1\[2\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 gencon_inst.ALU_in1\[13\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 net16 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 _0190_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1 VGND VGND VPWR VPWR
+ net188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _0364_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 gencon_inst.mult_calc.INn2\[1\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold97 gencon_inst.mult_calc.countSave\[11\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2121_ _1175_ _1174_ net415 VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux2_1
X_2052_ _1058_ _1121_ _1122_ _1046_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__o22a_1
X_1905_ gencon_inst.ALU_out\[8\] net73 net45 net25 VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1698_ net31 _0906_ _0908_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a21oi_1
X_1767_ net384 _0947_ net112 VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
X_1836_ gencon_inst.operand2\[9\] net220 net61 VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2319_ net115 net284 _0484_ _0494_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__a22o_1
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR display_output[4] sky130_fd_sc_hd__buf_2
Xoutput10 net10 VGND VGND VPWR VPWR complete sky130_fd_sc_hd__buf_2
XFILLER_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput8 net8 VGND VGND VPWR VPWR ColOut[2] sky130_fd_sc_hd__buf_2
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1621_ _0797_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nor2_1
X_1552_ gencon_inst.add_calc.main.a0.in1 gencon_inst.add_calc.main.in2\[0\] VGND VGND
+ VPWR VPWR _0775_ sky130_fd_sc_hd__xor2_1
X_2670_ clknet_leaf_27_clk _0229_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2104_ _1026_ net36 _1157_ _1162_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a31o_1
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1483_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__inv_2
XFILLER_27_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2035_ _1073_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1819_ gencon_inst.latched_operator_input\[0\] net277 net59 VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__mux2_1
X_2799_ clknet_leaf_21_clk _0353_ net152 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
XFILLER_26_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2722_ clknet_leaf_19_clk _0276_ net155 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1604_ gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1 _0823_ _0824_ VGND
+ VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nand3_1
Xfanout107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
Xfanout129 net137 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_2
X_1535_ net102 _0761_ _0762_ net298 net91 VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a32o_1
Xfanout118 net120 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_4
X_2584_ clknet_leaf_31_clk _0143_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2653_ clknet_leaf_28_clk _0212_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1466_ _0697_ _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__or2_1
X_1397_ gencon_inst.mult_calc.out\[6\] net383 net103 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2018_ gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1 _1068_ VGND VGND
+ VPWR VPWR _1092_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold172 input_ctrl_inst.read_input_flag VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 gencon_inst.mult_calc.INn2\[0\] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 gencon_inst.mult_calc.INn2\[12\] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 gencon_inst.mult_calc.INn2\[11\] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 input_ctrl_inst.col_index\[13\] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1320_ _0644_ _0647_ gencon_inst.operand2\[4\] VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o21a_1
XFILLER_5_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1251_ _0556_ _0593_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__nor3_1
XFILLER_49_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2705_ clknet_leaf_17_clk _0259_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2636_ clknet_leaf_24_clk _0195_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2567_ clknet_leaf_24_clk _0130_ net151 VGND VGND VPWR VPWR gencon_inst.operand2\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_1518_ gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__nand2_1
XFILLER_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2498_ clknet_leaf_29_clk _0073_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1449_ net398 net302 net99 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_74_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1303_ net55 _0635_ _0636_ net49 gencon_inst.mult_calc.out\[1\] VGND VGND VPWR VPWR
+ _0637_ sky130_fd_sc_hd__a32o_1
X_2283_ input_ctrl_inst.scan_timer\[13\] input_ctrl_inst.scan_timer\[14\] _0468_ VGND
+ VGND VPWR VPWR _0471_ sky130_fd_sc_hd__and3_1
X_2421_ _0549_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__nor2_1
X_2352_ input_ctrl_inst.col_index\[5\] input_ctrl_inst.col_index\[4\] _0504_ VGND
+ VGND VPWR VPWR _0506_ sky130_fd_sc_hd__and3_1
X_1234_ gencon_inst.operand1\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0581_ sky130_fd_sc_hd__or2_1
XFILLER_49_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2619_ clknet_leaf_25_clk net290 net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1998_ gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1 _1071_ VGND VGND
+ VPWR VPWR _1072_ sky130_fd_sc_hd__and2_1
XFILLER_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1852_ gencon_inst.operand1\[9\] net239 net61 VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
X_1921_ gencon_inst.ALU_out\[13\] net73 net66 _0975_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1783_ net116 _0954_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_12_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2266_ net418 _0459_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__xor2_1
X_2404_ input_ctrl_inst.col_index\[24\] net53 _0538_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__a21bo_1
X_2335_ net95 net260 net80 net261 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__a22o_1
X_1217_ gencon_inst.operand1\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0566_ sky130_fd_sc_hd__and2_1
X_2197_ _0402_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__or2_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold54 gencon_inst.ALU_in2\[3\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0320_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 gencon_inst.ALU_in1\[10\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 input_ctrl_inst.input_control_state\[0\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 gencon_inst.mult_calc.INn1\[10\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1 VGND VGND VPWR VPWR
+ net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1 VGND VGND VPWR VPWR
+ net200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 gencon_inst.mult_calc.countSave\[9\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 gencon_inst.mult_calc.countSave\[1\] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2120_ net36 _1173_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and2_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2051_ _1044_ _1048_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__nor2_1
XFILLER_19_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1835_ gencon_inst.operand2\[8\] net214 net61 VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
X_1904_ _1007_ _1008_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__or2_1
X_1697_ _0846_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__xnor2_2
X_1766_ gencon_inst.ALU_in2\[11\] gencon_inst.ALU_in1\[11\] net69 VGND VGND VPWR VPWR
+ _0947_ sky130_fd_sc_hd__mux2_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2318_ gencon_inst.keypad_input\[2\] net82 _0491_ _0493_ VGND VGND VPWR VPWR _0494_
+ sky130_fd_sc_hd__a22o_1
X_2249_ _1052_ _0448_ _0449_ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_23_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput11 net11 VGND VGND VPWR VPWR display_output[0] sky130_fd_sc_hd__buf_2
Xoutput22 net22 VGND VGND VPWR VPWR display_output[5] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR ColOut[3] sky130_fd_sc_hd__buf_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1620_ _0801_ _0805_ _0839_ _0802_ _0798_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o311a_1
X_1551_ _0628_ _0773_ _0774_ net417 VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o22a_1
X_1482_ gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__or2_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2103_ net37 _1161_ input_ctrl_inst.debounce_cnt\[13\] VGND VGND VPWR VPWR _1162_
+ sky130_fd_sc_hd__o21a_1
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1 _1072_ gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1
+ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__a21oi_1
X_1818_ gencon_inst.latched_operator_input\[2\] net117 _0388_ gencon_inst.latched_operator_input\[1\]
+ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__or4b_4
X_2798_ clknet_leaf_21_clk _0352_ net152 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1749_ net366 _0938_ net109 VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
XFILLER_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2721_ clknet_leaf_18_clk _0275_ net155 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2652_ clknet_leaf_32_clk _0211_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1603_ _0823_ _0824_ gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1 VGND
+ VGND VPWR VPWR _0825_ sky130_fd_sc_hd__a21oi_1
Xfanout108 gencon_inst.add_calc.diffSign VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
X_1534_ _0758_ _0759_ _0760_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a21o_1
X_1465_ gencon_inst.mult_calc.main.a0.in2 gencon_inst.mult_calc.main.a0.in1 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2
+ gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1 VGND VGND VPWR VPWR _0703_
+ sky130_fd_sc_hd__a22oi_1
Xfanout119 net120 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
X_2583_ clknet_leaf_31_clk _0142_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1396_ gencon_inst.mult_calc.out\[5\] net285 net103 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
XFILLER_27_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2017_ gencon_inst.mult_calc.compCount.in2\[3\] _1083_ _1086_ _1090_ _1087_ VGND
+ VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a221o_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold140 gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1 VGND VGND VPWR
+ VPWR net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _0372_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2 VGND VGND VPWR
+ VPWR net308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold195 gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1 VGND VGND VPWR VPWR
+ net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 gencon_inst.ALU_out\[15\] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 gencon_inst.add_calc.main.in2\[6\] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1250_ _1039_ _0586_ gencon_inst.operand1\[6\] VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o21ba_1
XFILLER_49_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2704_ clknet_leaf_17_clk _0258_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2635_ clknet_leaf_24_clk _0194_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_74_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2566_ clknet_leaf_24_clk _0129_ net151 VGND VGND VPWR VPWR gencon_inst.operand2\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_1517_ gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
+ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__nor2_1
X_2497_ clknet_leaf_29_clk _0072_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1448_ net385 net362 net99 VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1379_ net86 _1103_ net90 net255 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2420_ input_ctrl_inst.col_index\[29\] _0427_ _0537_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and3_1
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
X_1233_ gencon_inst.operand1\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0580_ sky130_fd_sc_hd__nand2_1
X_1302_ gencon_inst.operand2\[0\] gencon_inst.latched_keypad_input\[0\] _0633_ _0634_
+ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__nand4_1
X_2282_ input_ctrl_inst.scan_timer\[13\] input_ctrl_inst.scan_timer\[12\] _0466_ input_ctrl_inst.scan_timer\[14\]
+ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a31o_1
X_2351_ input_ctrl_inst.col_index\[4\] _0504_ net425 VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1997_ gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
+ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__and3_1
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2549_ clknet_leaf_13_clk _0112_ net148 VGND VGND VPWR VPWR gencon_inst.operand1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2618_ clknet_leaf_32_clk net354 net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1851_ gencon_inst.operand1\[8\] net238 net61 VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__mux2_1
X_1920_ net15 net46 net58 gencon_inst.mult_calc.out\[13\] VGND VGND VPWR VPWR _1019_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1782_ net63 VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__inv_2
X_2403_ net53 _0501_ _0536_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or4_1
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1216_ gencon_inst.operand1\[0\] net34 _0564_ _0565_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__o22a_1
X_2265_ _0445_ _0458_ _0460_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and3_1
X_2334_ net95 net254 net80 net259 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__a22o_1
X_2196_ input_ctrl_inst.col_index\[0\] input_ctrl_inst.col_index\[1\] net114 input_ctrl_inst.col_index\[3\]
+ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o31a_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 gencon_inst.mult_calc.INn1\[4\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1 VGND VGND VPWR VPWR
+ net179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold55 gencon_inst.ALU_in2\[0\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 gencon_inst.ALU_in2\[6\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold77 net14 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1 VGND VGND VPWR VPWR
+ net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold88 gencon_inst.mult_calc.countSave\[3\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 _0069_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 input_ctrl_inst.scan_timer\[17\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ _1044_ net30 VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1765_ net381 _0946_ net112 VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
X_1834_ gencon_inst.operand2\[7\] net229 net61 VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
X_1903_ net66 _0969_ net57 gencon_inst.mult_calc.out\[7\] VGND VGND VPWR VPWR _1008_
+ sky130_fd_sc_hd__a22o_1
X_1696_ _0785_ _0786_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nand2b_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ gencon_inst.mult_calc.finish _1210_ _0392_ _1204_ net55 VGND VGND VPWR VPWR
+ _0393_ sky130_fd_sc_hd__a221o_1
X_2317_ input_ctrl_inst.decoded_key\[2\] _1199_ input_ctrl_inst.decoded_key\[3\] VGND
+ VGND VPWR VPWR _0493_ sky130_fd_sc_hd__a21o_1
X_2248_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[0\] input_ctrl_inst.scan_timer\[15\]
+ input_ctrl_inst.scan_timer\[14\] VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or4bb_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput23 net23 VGND VGND VPWR VPWR display_output[6] sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR display_output[10] sky130_fd_sc_hd__buf_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1550_ gencon_inst.operator_input\[0\] gencon_inst.key_read _1204_ _0381_ net47 VGND
+ VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a41o_1
X_1481_ net395 net89 _0716_ net102 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a22o_1
X_2102_ _1157_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nor2_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ _1101_ _1104_ _1106_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__a21o_1
XFILLER_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2797_ clknet_leaf_16_clk _0351_ net150 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
X_1748_ gencon_inst.ALU_in2\[2\] gencon_inst.ALU_in1\[2\] net67 VGND VGND VPWR VPWR
+ _0938_ sky130_fd_sc_hd__mux2_1
X_1817_ _0977_ net242 net39 VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _0797_ _0798_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__and2b_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1602_ net105 gencon_inst.add_calc.main.in2\[2\] VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__nand2_1
X_2720_ clknet_leaf_17_clk _0274_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2582_ clknet_leaf_35_clk _0141_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2651_ clknet_leaf_30_clk _0210_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout109 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
X_1533_ _0758_ _0759_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand3_1
X_1464_ _0700_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__and2b_1
X_1395_ gencon_inst.mult_calc.out\[4\] net395 net103 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
X_2016_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn gencon_inst.mult_calc.compCount.in2\[0\]
+ _1089_ _1088_ gencon_inst.mult_calc.compCount.in2\[1\] VGND VGND VPWR VPWR _1090_
+ sky130_fd_sc_hd__a32o_1
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
Xhold174 gencon_inst.add_calc.main.in2\[14\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _0182_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2 VGND VGND VPWR
+ VPWR net320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 gencon_inst.mult_calc.adderSave\[12\] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 gencon_inst.mult_calc.adderSave\[1\] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 _0184_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold196 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2 VGND VGND VPWR
+ VPWR net353 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_5_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
X_2703_ clknet_leaf_14_clk _0257_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2565_ clknet_leaf_24_clk _0128_ net151 VGND VGND VPWR VPWR gencon_inst.operand2\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_2634_ clknet_leaf_24_clk _0193_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1516_ net102 _0745_ _0746_ net305 net91 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a32o_1
X_2496_ clknet_leaf_29_clk _0071_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1378_ net86 _1099_ net88 net252 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__a2bb2o_1
X_1447_ net382 net361 net99 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
XFILLER_70_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout80 net81 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_4
Xfanout91 _0688_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
X_1232_ gencon_inst.operand1\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0579_ sky130_fd_sc_hd__and2_1
X_1301_ gencon_inst.operand2\[0\] gencon_inst.latched_keypad_input\[0\] _0633_ _0634_
+ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_2281_ net334 _0468_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__xor2_1
X_2350_ net433 _0504_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_50_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1996_ gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1 _1068_ VGND VGND VPWR
+ VPWR _1070_ sky130_fd_sc_hd__and4_1
X_2548_ clknet_leaf_13_clk _0111_ net148 VGND VGND VPWR VPWR gencon_inst.operand1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2617_ clknet_leaf_25_clk _0176_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2479_ clknet_leaf_4_clk _0054_ VGND VGND VPWR VPWR gencon_inst.operator_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_75_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1850_ gencon_inst.operand1\[7\] net248 net61 VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
X_1781_ _0388_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2402_ input_ctrl_inst.col_index\[24\] _0500_ _0508_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__and3_2
X_2333_ net95 net265 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
+ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__a22o_1
X_1215_ gencon_inst.ALU_out\[0\] net71 net51 gencon_inst.mult_calc.out\[0\] VGND VGND
+ VPWR VPWR _0565_ sky130_fd_sc_hd__a22o_1
XFILLER_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2264_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__inv_2
XFILLER_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2195_ _0398_ _0401_ _0405_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__nand3_1
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1979_ net92 _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__nor2_2
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold56 gencon_inst.ALU_in2\[2\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 gencon_inst.ALU_in2\[10\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 gencon_inst.prev_operator_input\[2\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold12 input_ctrl_inst.input_control_state\[1\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 _0476_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold67 gencon_inst.ALU_in1\[12\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold78 gencon_inst.mult_calc.out\[15\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold89 _0063_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ gencon_inst.ALU_out\[7\] net73 net45 net24 VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__a22o_1
XFILLER_34_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1764_ gencon_inst.ALU_in2\[10\] gencon_inst.ALU_in1\[10\] net69 VGND VGND VPWR VPWR
+ _0946_ sky130_fd_sc_hd__mux2_1
X_1833_ gencon_inst.operand2\[6\] net223 net61 VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_1
XFILLER_30_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1695_ _0897_ _0899_ _0904_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__or3_1
X_2316_ net115 net270 _0484_ _0492_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__a22o_1
XFILLER_72_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2178_ equal_input gencon_inst.read_input VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nand2b_1
XFILLER_38_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2247_ input_ctrl_inst.scan_timer\[3\] input_ctrl_inst.scan_timer\[2\] input_ctrl_inst.scan_timer\[5\]
+ input_ctrl_inst.scan_timer\[4\] VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_23_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput13 net13 VGND VGND VPWR VPWR display_output[11] sky130_fd_sc_hd__buf_2
Xoutput24 net24 VGND VGND VPWR VPWR display_output[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ _0713_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__xnor2_1
X_2101_ net36 _1146_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and2b_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2032_ gencon_inst.mult_calc.compCount.in2\[9\] _1103_ _1105_ gencon_inst.mult_calc.compCount.in2\[10\]
+ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__a22o_1
X_1678_ _0887_ _0889_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__or2_1
X_1747_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0937_ net109 VGND
+ VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
X_1816_ gencon_inst.operand2\[15\] gencon_inst.operand1\[15\] net76 VGND VGND VPWR
+ VPWR _0977_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ clknet_leaf_24_clk _0350_ net151 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1601_ net105 gencon_inst.add_calc.main.in2\[2\] VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_57_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1532_ _0753_ _0756_ _0754_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2581_ clknet_leaf_31_clk _0140_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2650_ clknet_leaf_31_clk net380 net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1394_ gencon_inst.mult_calc.out\[3\] net388 net103 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
X_1463_ gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__nand2_1
X_2015_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.compCount.in2\[1\]
+ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_75_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold120 gencon_inst.addOrSub VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dlygate4sd3_1
X_2779_ clknet_leaf_11_clk _0333_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold186 gencon_inst.mult_calc.INn2\[6\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 gencon_inst.mult_calc.INn2\[2\] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 gencon_inst.mult_calc.INn2\[13\] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _0181_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _0177_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 input_ctrl_inst.col_index\[6\] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold142 gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR
+ VPWR net299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2702_ clknet_leaf_14_clk _0256_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2564_ clknet_leaf_13_clk _0127_ net148 VGND VGND VPWR VPWR gencon_inst.operand2\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_2633_ clknet_leaf_24_clk _0192_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1515_ _0742_ _0743_ _0744_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a21o_1
X_2495_ clknet_leaf_28_clk _0070_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1377_ net86 _1096_ net88 net269 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a2bb2o_1
X_1446_ net379 gencon_inst.mult_calc.INn2\[7\] net97 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XFILLER_70_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout70 _0920_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
Xfanout92 input_ctrl_inst.input_control_state\[2\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
XFILLER_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout81 _1061_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1231_ gencon_inst.operand1\[2\] net34 _0577_ _0578_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__o22a_1
X_1300_ gencon_inst.operand2\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0634_ sky130_fd_sc_hd__or2_1
X_2280_ _0468_ _0469_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__nor2_1
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2616_ clknet_leaf_32_clk net356 net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1 _1068_ VGND VGND
+ VPWR VPWR _1069_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2547_ clknet_leaf_13_clk _0110_ net148 VGND VGND VPWR VPWR gencon_inst.operand1\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_2478_ clknet_leaf_4_clk _0053_ VGND VGND VPWR VPWR gencon_inst.operator_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1429_ net200 net182 net98 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1780_ gencon_inst.latched_operator_input\[1\] gencon_inst.latched_operator_input\[0\]
+ net117 gencon_inst.latched_operator_input\[2\] VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__or4b_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2401_ _0500_ _0508_ input_ctrl_inst.col_index\[24\] VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__a21oi_1
X_2332_ net95 net255 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1
+ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__a22o_1
XFILLER_65_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ gencon_inst.operand1\[0\] gencon_inst.latched_keypad_input\[0\] net43 _0563_
+ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__o22a_1
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2263_ input_ctrl_inst.scan_timer\[5\] input_ctrl_inst.scan_timer\[4\] input_ctrl_inst.scan_timer\[6\]
+ _0455_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and4_1
X_2194_ _0403_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1978_ input_ctrl_inst.input_control_state\[0\] input_ctrl_inst.input_control_state\[1\]
+ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2b_1
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold57 gencon_inst.ALU_in2\[8\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 gencon_inst.ALU_in1\[6\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 gencon_inst.prev_operator_input\[0\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1 VGND VGND VPWR
+ VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 gencon_inst.mult_calc.INn1\[11\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold79 input_ctrl_inst.scan_timer\[11\] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 gencon_inst.mult_calc.main.a0.in1 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1901_ _1005_ _1006_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__or2_1
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ gencon_inst.operand2\[5\] net204 net60 VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_1
XFILLER_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1694_ gencon_inst.ALU_out\[11\] _0905_ net113 VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
X_1763_ net414 _0945_ net111 VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
X_2315_ gencon_inst.keypad_input\[1\] net82 _0489_ _0491_ VGND VGND VPWR VPWR _0492_
+ sky130_fd_sc_hd__a22o_1
X_2246_ _0437_ _0446_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__or3b_1
XFILLER_53_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2177_ _1203_ _1206_ _0378_ _0391_ VGND VGND VPWR VPWR gencon_inst.next_state\[0\]
+ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_11_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput25 net25 VGND VGND VPWR VPWR display_output[8] sky130_fd_sc_hd__buf_2
Xoutput14 net14 VGND VGND VPWR VPWR display_output[12] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2100_ _1157_ _1159_ net427 net37 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2031_ gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1 _1072_ VGND VGND
+ VPWR VPWR _1105_ sky130_fd_sc_hd__xnor2_1
X_2795_ clknet_leaf_16_clk _0349_ net150 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_50_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ _0976_ net196 net41 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
XFILLER_30_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1677_ _0891_ _0890_ gencon_inst.ALU_out\[8\] net84 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a2bb2o_1
X_1746_ gencon_inst.ALU_in2\[1\] gencon_inst.ALU_in1\[1\] net67 VGND VGND VPWR VPWR
+ _0937_ sky130_fd_sc_hd__mux2_1
X_2229_ net283 net311 net266 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__o21ba_1
XFILLER_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1600_ gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1 _0819_ _0820_ VGND
+ VGND VPWR VPWR _0822_ sky130_fd_sc_hd__nand3_1
X_1531_ gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__nand2_1
X_1462_ gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nor2_1
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2580_ clknet_leaf_34_clk _0139_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1393_ gencon_inst.mult_calc.out\[2\] net396 net103 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2014_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__xnor2_1
Xhold110 gencon_inst.ALU_in1\[11\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ clknet_leaf_23_clk _0332_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold187 gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1 VGND VGND VPWR VPWR
+ net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1 VGND VGND VPWR VPWR
+ net333 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 gencon_inst.add_calc.sameSignVal VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 gencon_inst.add_calc.state\[0\] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ net345 _0928_ net111 VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
Xhold121 _0297_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2 VGND VGND VPWR
+ VPWR net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2 VGND VGND VPWR
+ VPWR net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2 VGND VGND VPWR
+ VPWR net355 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_56_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2701_ clknet_leaf_15_clk _0255_ net150 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2632_ clknet_leaf_33_clk _0191_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2563_ clknet_leaf_24_clk _0126_ net148 VGND VGND VPWR VPWR gencon_inst.operand2\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_1514_ _0742_ _0743_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__nand3_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2494_ clknet_leaf_30_clk net256 net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1445_ net369 net343 net98 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ net86 _1080_ net88 net273 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout60 _0978_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
Xfanout82 _1054_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_2
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout93 net96 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
XFILLER_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ gencon_inst.ALU_out\[2\] net71 net51 gencon_inst.mult_calc.out\[2\] net43
+ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a221o_1
XFILLER_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1994_ gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1 _1067_ VGND VGND
+ VPWR VPWR _1068_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_15_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload30 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__clkinv_4
X_2615_ clknet_leaf_33_clk net301 net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2546_ clknet_leaf_12_clk _0109_ net133 VGND VGND VPWR VPWR gencon_inst.operand1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2477_ clknet_leaf_5_clk _0052_ VGND VGND VPWR VPWR equal_input sky130_fd_sc_hd__dfxtp_1
X_1428_ net187 net168 net98 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1359_ gencon_inst.operand2\[12\] _0681_ net48 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_74_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ _1036_ net53 _0534_ _0535_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_12_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1213_ net75 _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__and2_1
X_2262_ input_ctrl_inst.scan_timer\[5\] input_ctrl_inst.scan_timer\[4\] _0455_ input_ctrl_inst.scan_timer\[6\]
+ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a31o_1
X_2331_ net93 net252 net80 gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2193_ input_ctrl_inst.col_index\[5\] input_ctrl_inst.col_index\[4\] input_ctrl_inst.col_index\[7\]
+ input_ctrl_inst.col_index\[6\] VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or4_1
X_1977_ gencon_inst.key_read net82 _1052_ _1050_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__o211ai_1
X_2529_ clknet_leaf_37_clk _0100_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold47 gencon_inst.ALU_in2\[5\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold69 _0324_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 gencon_inst.mult_calc.INn1\[5\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 gencon_inst.mult_calc.INn1\[1\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 gencon_inst.mult_calc.INn1\[0\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold58 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1 VGND VGND VPWR
+ VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1831_ gencon_inst.operand2\[4\] net197 net59 VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
X_1900_ net66 _0968_ net57 gencon_inst.mult_calc.out\[6\] VGND VGND VPWR VPWR _1006_
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1693_ _0902_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__xnor2_1
X_1762_ gencon_inst.ALU_in2\[9\] gencon_inst.ALU_in1\[9\] net68 VGND VGND VPWR VPWR
+ _0945_ sky130_fd_sc_hd__mux2_1
X_2176_ _0384_ net55 _0390_ _0388_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__or4b_1
X_2314_ net82 _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__nor2_1
X_2245_ input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[6\] input_ctrl_inst.scan_timer\[9\]
+ input_ctrl_inst.scan_timer\[8\] VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__and4b_1
XFILLER_65_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput26 net26 VGND VGND VPWR VPWR display_output[9] sky130_fd_sc_hd__buf_2
Xoutput15 net15 VGND VGND VPWR VPWR display_output[13] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ gencon_inst.mult_calc.compCount.in2\[8\] _1099_ _1103_ gencon_inst.mult_calc.compCount.in2\[9\]
+ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__o22a_1
XFILLER_35_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1745_ net410 _0936_ net109 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_1
X_2794_ clknet_leaf_13_clk _0348_ net148 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
X_1814_ gencon_inst.operand2\[14\] gencon_inst.operand1\[14\] net77 VGND VGND VPWR
+ VPWR _0976_ sky130_fd_sc_hd__mux2_1
XFILLER_30_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1676_ _0852_ _0887_ _0889_ net84 VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__a31o_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2228_ net266 net311 VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2_1
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2159_ gencon_inst.gencon_state\[1\] gencon_inst.gencon_state\[2\] VGND VGND VPWR
+ VPWR _1207_ sky130_fd_sc_hd__nor2_1
XFILLER_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_33_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1392_ gencon_inst.mult_calc.out\[1\] net342 net103 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
X_1530_ gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__or2_1
X_1461_ net101 _0698_ _0699_ net342 net89 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a32o_1
XFILLER_67_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2013_ _1067_ _1084_ gencon_inst.mult_calc.compCount.in2\[2\] VGND VGND VPWR VPWR
+ _1087_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_50_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1728_ gencon_inst.ALU_in1\[7\] gencon_inst.ALU_in2\[7\] net68 VGND VGND VPWR VPWR
+ _0928_ sky130_fd_sc_hd__mux2_1
X_2777_ clknet_leaf_20_clk _0331_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold122 gencon_inst.mult_calc.INn2\[14\] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _0178_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _0174_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold111 gencon_inst.mult_calc.countSave\[13\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold100 gencon_inst.mult_calc.countSave\[2\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ net32 _0873_ _0875_ net84 VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__a31o_1
Xhold166 gencon_inst.add_calc.main.in2\[2\] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 gencon_inst.add_calc.main.in2\[7\] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 gencon_inst.mult_calc.INn2\[5\] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 input_ctrl_inst.scan_timer\[13\] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _0175_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ clknet_leaf_15_clk _0254_ net150 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2562_ clknet_leaf_13_clk _0125_ net148 VGND VGND VPWR VPWR gencon_inst.operand2\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_2631_ clknet_leaf_33_clk net177 net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_4_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
X_1513_ _0736_ _0740_ _0737_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__o21ai_1
X_2493_ clknet_leaf_30_clk net253 net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1375_ net86 _1081_ net88 net274 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__a2bb2o_1
X_1444_ net328 net312 net98 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2829_ clknet_leaf_5_clk input_ctrl_inst.next_state\[2\] net128 VGND VGND VPWR VPWR
+ input_ctrl_inst.input_control_state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_73_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout61 _0978_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
Xfanout72 _0558_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xfanout50 _0627_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_1
Xfanout94 net96 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_2
XFILLER_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1993_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR _1067_
+ sky130_fd_sc_hd__and3_1
Xclkload31 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__inv_6
X_2545_ clknet_leaf_11_clk _0108_ net134 VGND VGND VPWR VPWR gencon_inst.operand1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload20 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_12
X_2614_ clknet_leaf_33_clk net350 net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2476_ clknet_leaf_5_clk _0017_ net129 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1358_ _0679_ _0680_ gencon_inst.mult_calc.out\[12\] net50 VGND VGND VPWR VPWR _0681_
+ sky130_fd_sc_hd__a2bb2o_1
X_1427_ gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1 net176 net98 VGND
+ VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1289_ _0623_ _0624_ _0555_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__and3b_1
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload3 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_11_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1212_ gencon_inst.operand1\[0\] gencon_inst.latched_keypad_input\[0\] VGND VGND
+ VPWR VPWR _0562_ sky130_fd_sc_hd__nand2_1
X_2261_ net364 _0457_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__xnor2_1
X_2330_ net93 net269 net78 net276 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a22o_1
X_2192_ input_ctrl_inst.col_index\[0\] input_ctrl_inst.col_index\[1\] net114 input_ctrl_inst.col_index\[3\]
+ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_63_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ net92 input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nand3b_1
X_2528_ clknet_leaf_37_clk _0099_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_2459_ clknet_leaf_7_clk _0018_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold48 gencon_inst.ALU_in1\[14\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 gencon_inst.mult_calc.INn1\[9\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 gencon_inst.mult_calc.INn1\[2\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1 VGND VGND VPWR
+ VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 input_ctrl_inst.col_index\[15\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1761_ net344 _0944_ net111 VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ gencon_inst.operand2\[3\] net211 net60 VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1692_ _0844_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__xnor2_1
X_2313_ input_ctrl_inst.decoded_key\[2\] _0479_ input_ctrl_inst.decoded_key\[3\] VGND
+ VGND VPWR VPWR _0490_ sky130_fd_sc_hd__o21a_1
XFILLER_65_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2175_ gencon_inst.ALU_finish _0389_ _0380_ gencon_inst.read_input VGND VGND VPWR
+ VPWR _0390_ sky130_fd_sc_hd__a2bb2o_1
X_2244_ input_ctrl_inst.scan_timer\[11\] input_ctrl_inst.scan_timer\[10\] input_ctrl_inst.scan_timer\[13\]
+ input_ctrl_inst.scan_timer\[12\] VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__or4_1
X_1959_ net105 VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput16 net16 VGND VGND VPWR VPWR display_output[14] sky130_fd_sc_hd__buf_2
Xoutput27 net27 VGND VGND VPWR VPWR input_state_FPGA[0] sky130_fd_sc_hd__buf_2
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2793_ clknet_leaf_10_clk _0347_ net150 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
X_1744_ gencon_inst.ALU_in2\[0\] gencon_inst.ALU_in1\[0\] net67 VGND VGND VPWR VPWR
+ _0936_ sky130_fd_sc_hd__mux2_1
X_1813_ _0975_ net249 net41 VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ net31 _0887_ _0889_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ input_ctrl_inst.debounce_cnt\[10\] _1148_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__nor2_1
X_2158_ gencon_inst.read_input equal_input net76 VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_36_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2227_ net114 _0434_ input_ctrl_inst.col_index\[0\] input_ctrl_inst.col_index\[1\]
+ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__or4bb_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ _0696_ _0697_ _0694_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_26_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ gencon_inst.mult_calc.out\[0\] net303 net103 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ gencon_inst.mult_calc.compCount.in2\[2\] _1067_ _1084_ VGND VGND VPWR VPWR
+ _1086_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_33_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold134 gencon_inst.add_calc.main.in2\[10\] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ net32 _0873_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__a21oi_1
Xhold167 gencon_inst.add_calc.main.in2\[4\] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ net341 _0927_ net111 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
X_2776_ clknet_leaf_20_clk _0330_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[12\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_44_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold145 gencon_inst.mult_calc.INn2\[10\] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _0366_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _0375_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold101 gencon_inst.mult_calc.countSave\[4\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 gencon_inst.mult_calc.countSave\[7\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
X_1589_ net108 gencon_inst.add_calc.main.in2\[5\] VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or2_1
Xhold189 gencon_inst.add_calc.main.in2\[1\] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold178 gencon_inst.mult_calc.compCount.in2\[12\] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2561_ clknet_leaf_13_clk _0124_ net133 VGND VGND VPWR VPWR gencon_inst.operand2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2630_ clknet_leaf_33_clk _0189_ net127 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1512_ gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nand2_1
X_2492_ clknet_leaf_30_clk _0067_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1374_ net86 _1092_ net88 net258 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a2bb2o_1
X_1443_ net386 net378 net98 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2828_ clknet_leaf_5_clk input_ctrl_inst.next_state\[1\] net128 VGND VGND VPWR VPWR
+ input_ctrl_inst.input_control_state\[1\] sky130_fd_sc_hd__dfrtp_2
X_2759_ clknet_leaf_19_clk _0313_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_73_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout62 _0978_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout51 _0559_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_4
Xfanout73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xfanout40 net42 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout84 _1033_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout95 net96 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
XFILLER_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload10 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_15_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1992_ _1028_ _1066_ net78 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a21oi_1
Xclkload32 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__inv_6
X_2544_ clknet_leaf_11_clk _0107_ net132 VGND VGND VPWR VPWR gencon_inst.operand1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2475_ clknet_leaf_6_clk _0016_ net129 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload21 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_2
X_2613_ clknet_leaf_33_clk _0172_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1288_ gencon_inst.operand1\[12\] gencon_inst.operand1\[13\] _0612_ gencon_inst.operand1\[14\]
+ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a31o_1
X_1357_ gencon_inst.operand2\[12\] _0675_ net56 VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__o21ai_1
X_1426_ net175 net172 net97 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_28_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload4 clknet_leaf_1_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_4
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1211_ _1208_ net51 _0378_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__a21o_1
X_2260_ net115 _0443_ _0455_ input_ctrl_inst.scan_timer\[4\] _0457_ VGND VGND VPWR
+ VPWR _0036_ sky130_fd_sc_hd__o221a_1
X_2191_ input_ctrl_inst.col_index\[0\] input_ctrl_inst.col_index\[1\] net114 input_ctrl_inst.col_index\[3\]
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_63_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1975_ net92 input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__and3b_2
X_2458_ clknet_leaf_5_clk _0008_ net128 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold27 gencon_inst.mult_calc.INn1\[7\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 gencon_inst.mult_calc.INn1\[6\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1 VGND VGND VPWR VPWR
+ net195 sky130_fd_sc_hd__dlygate4sd3_1
X_1409_ net94 gencon_inst.mult_calc.adderSave\[2\] net349 net79 VGND VGND VPWR VPWR
+ _0173_ sky130_fd_sc_hd__a22o_1
X_2527_ clknet_leaf_37_clk _0098_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold49 gencon_inst.ALU_in2\[11\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2389_ input_ctrl_inst.col_index\[20\] net53 VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__and2_1
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1691_ _0789_ _0790_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__and2b_1
X_1760_ gencon_inst.ALU_in2\[8\] gencon_inst.ALU_in1\[8\] net68 VGND VGND VPWR VPWR
+ _0944_ sky130_fd_sc_hd__mux2_1
X_2312_ _1199_ _0479_ _0485_ input_ctrl_inst.decoded_key\[3\] VGND VGND VPWR VPWR
+ _0489_ sky130_fd_sc_hd__a31o_1
XFILLER_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2174_ _1029_ _0385_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or2_1
X_2243_ net115 _0443_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__or2_1
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput17 net17 VGND VGND VPWR VPWR display_output[15] sky130_fd_sc_hd__buf_2
X_1889_ _0997_ _0998_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
Xoutput28 net28 VGND VGND VPWR VPWR input_state_FPGA[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1958_ input_ctrl_inst.col_index\[31\] VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__inv_2
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2792_ clknet_leaf_10_clk _0346_ net136 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
X_1674_ _0840_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__xnor2_1
X_1743_ net331 _0935_ net111 VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
X_1812_ gencon_inst.operand2\[13\] gencon_inst.operand1\[13\] net77 VGND VGND VPWR
+ VPWR _0975_ sky130_fd_sc_hd__mux2_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2226_ input_ctrl_inst.col_index\[0\] net114 _0434_ input_ctrl_inst.col_index\[1\]
+ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__or4b_1
X_2088_ input_ctrl_inst.debounce_cnt\[10\] _1057_ _1146_ VGND VGND VPWR VPWR _1150_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2157_ _1029_ gencon_inst.gencon_state\[3\] gencon_inst.gencon_state\[2\] gencon_inst.gencon_state\[0\]
+ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_36_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1390_ net227 _0692_ net97 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ _1067_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1657_ _0835_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__xnor2_1
X_1588_ gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1 _0807_ _0808_ VGND
+ VGND VPWR VPWR _0810_ sky130_fd_sc_hd__nand3_1
Xhold124 input_ctrl_inst.debounce_cnt\[3\] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 gencon_inst.add_calc.main.in2\[12\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dlygate4sd3_1
X_1726_ gencon_inst.ALU_in1\[6\] gencon_inst.ALU_in2\[6\] net70 VGND VGND VPWR VPWR
+ _0927_ sky130_fd_sc_hd__mux2_1
X_2775_ clknet_leaf_20_clk _0329_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[11\] sky130_fd_sc_hd__dfxtp_1
Xhold113 gencon_inst.keypad_input\[1\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2 VGND VGND VPWR
+ VPWR net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 gencon_inst.mult_calc.adderSave\[0\] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1 VGND VGND VPWR
+ VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _0214_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 gencon_inst.mult_calc.adderSave\[13\] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2209_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[20\] input_ctrl_inst.col_index\[23\]
+ input_ctrl_inst.col_index\[22\] VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__and4_1
XFILLER_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_32_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2560_ clknet_leaf_3_clk _0123_ net133 VGND VGND VPWR VPWR gencon_inst.operand2\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1511_ gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__or2_1
X_2491_ clknet_leaf_30_clk _0066_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1442_ net389 net209 net97 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1373_ net86 _1083_ net88 net245 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2758_ clknet_leaf_19_clk _0312_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[10\] sky130_fd_sc_hd__dfxtp_1
X_2827_ clknet_leaf_5_clk input_ctrl_inst.next_state\[0\] net128 VGND VGND VPWR VPWR
+ input_ctrl_inst.input_control_state\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2689_ clknet_leaf_17_clk _0243_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1709_ _0915_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout85 _1033_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_52_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout52 _0559_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
Xfanout74 _0558_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
Xfanout63 _0957_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
Xfanout41 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xfanout96 gencon_inst.mult_calc.state\[4\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload33 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__clkinv_8
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload22 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__clkinvlp_4
X_2612_ clknet_leaf_34_clk _0171_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.a0.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload11 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_6
X_1991_ _1062_ _1063_ _1065_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nor3_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2474_ clknet_leaf_7_clk _0015_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1425_ net179 net171 net97 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
X_2543_ clknet_leaf_0_clk net159 net122 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_66_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1287_ gencon_inst.operand1\[13\] gencon_inst.operand1\[14\] _0616_ VGND VGND VPWR
+ VPWR _0623_ sky130_fd_sc_hd__and3_1
X_1356_ gencon_inst.operand2\[12\] _0675_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__and2_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload5 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload5/X sky130_fd_sc_hd__clkbuf_8
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2190_ input_ctrl_inst.col_index\[12\] _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__nor2_1
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1974_ _1048_ net83 VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nand2_1
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold28 gencon_inst.keypad_input\[3\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 gencon_inst.mult_calc.INn1\[8\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
X_2457_ clknet_leaf_0_clk _0030_ net122 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[3\]
+ sky130_fd_sc_hd__dfstp_1
Xhold39 gencon_inst.mult_calc.INn1\[14\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ net94 net342 net399 net79 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__a22o_1
X_2526_ clknet_leaf_37_clk _0097_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_2388_ net408 net53 _0527_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__a21bo_1
XFILLER_71_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1339_ gencon_inst.operand2\[8\] _0663_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__xor2_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1690_ _0897_ _0899_ net31 VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__o21ai_1
XFILLER_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2311_ net115 net282 _0484_ _0488_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__a22o_1
X_2242_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__inv_2
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2173_ _1029_ _1201_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or2_1
X_1957_ input_ctrl_inst.col_index\[23\] VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__inv_2
Xoutput18 net18 VGND VGND VPWR VPWR display_output[1] sky130_fd_sc_hd__buf_2
X_1888_ net65 _0963_ net57 gencon_inst.mult_calc.out\[2\] VGND VGND VPWR VPWR _0998_
+ sky130_fd_sc_hd__a22o_1
Xoutput29 net29 VGND VGND VPWR VPWR input_state_FPGA[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2509_ clknet_leaf_38_clk _0080_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_6_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2791_ clknet_leaf_10_clk _0345_ net135 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1811_ _0974_ net163 net41 VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
X_1673_ _0801_ _0802_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nand2b_1
X_1742_ gencon_inst.ALU_in1\[14\] gencon_inst.ALU_in2\[14\] net68 VGND VGND VPWR VPWR
+ _0935_ sky130_fd_sc_hd__mux2_1
XFILLER_7_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2225_ input_ctrl_inst.col_index\[1\] net114 _0434_ input_ctrl_inst.col_index\[0\]
+ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
X_2087_ _1148_ _1149_ net439 net37 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a2bb2o_1
X_2156_ gencon_inst.gencon_state\[2\] gencon_inst.gencon_state\[0\] gencon_inst.gencon_state\[1\]
+ _1030_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__and4b_4
XTAP_TAPCELL_ROW_36_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2010_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR _1084_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_75_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1725_ net348 _0926_ net110 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
X_2774_ clknet_leaf_20_clk _0328_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[10\] sky130_fd_sc_hd__dfxtp_1
X_1656_ _0813_ _0814_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__and2b_1
X_1587_ _0807_ _0808_ gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1 VGND
+ VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a21oi_1
Xhold158 gencon_inst.add_calc.main.in2\[11\] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 gencon_inst.add_calc.main.in2\[9\] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold125 gencon_inst.keypad_input\[0\] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _0183_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 gencon_inst.mult_calc.countSave\[0\] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 gencon_inst.mult_calc.countSave\[12\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 gencon_inst.mult_calc.compCount.in2\[0\] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2139_ net82 _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__nor2_1
X_2208_ _0400_ _0414_ _0417_ _0408_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1510_ net404 net91 _0741_ net102 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
X_2490_ clknet_leaf_31_clk _0065_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1441_ net363 net332 net97 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__mux2_1
XFILLER_67_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1372_ net101 _1085_ net88 net257 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2688_ clknet_leaf_16_clk _0242_ net149 VGND VGND VPWR VPWR gencon_inst.ALU_out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1708_ _0849_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__xnor2_1
X_2757_ clknet_leaf_14_clk _0311_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[9\] sky130_fd_sc_hd__dfxtp_1
X_2826_ clknet_leaf_3_clk _0376_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_1639_ _0825_ _0826_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__nand2b_1
XFILLER_73_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xfanout75 _0555_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout64 _0957_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xfanout42 _0959_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XFILLER_10_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout53 _0451_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xfanout97 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_4
Xfanout86 _1032_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1990_ gencon_inst.mult_calc.INn2\[13\] gencon_inst.mult_calc.INn2\[12\] gencon_inst.mult_calc.INn2\[14\]
+ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or4_1
Xclkload34 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__inv_8
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload12 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_8
X_2611_ clknet_leaf_2_clk _0170_ net125 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2542_ clknet_leaf_0_clk net160 net122 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[2\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload23 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__clkinv_8
X_2473_ clknet_leaf_7_clk _0014_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1355_ gencon_inst.operand2\[11\] _0678_ net48 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
X_1424_ net203 net193 net97 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ gencon_inst.operand1\[13\] net35 _0621_ _0622_ VGND VGND VPWR VPWR _0120_
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload6 clknet_leaf_33_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2809_ clknet_leaf_4_clk gencon_inst.next_state\[2\] net132 VGND VGND VPWR VPWR gencon_inst.gencon_state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ net92 input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__nor3b_1
X_2525_ clknet_leaf_37_clk _0096_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold29 gencon_inst.prev_operator_input\[1\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
X_1338_ gencon_inst.operand2\[7\] _0665_ net47 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
Xhold18 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR
+ net175 sky130_fd_sc_hd__dlygate4sd3_1
X_2456_ clknet_leaf_0_clk _0029_ net123 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[2\]
+ sky130_fd_sc_hd__dfstp_2
X_1407_ net94 net303 net397 net79 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a22o_1
X_2387_ _0526_ net33 _0525_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__nand3b_1
XFILLER_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1269_ gencon_inst.operand1\[10\] _0605_ net75 VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2172_ gencon_inst.gencon_state\[1\] _0385_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__or2_1
X_2310_ gencon_inst.keypad_input\[0\] _1053_ _0486_ _0487_ VGND VGND VPWR VPWR _0488_
+ sky130_fd_sc_hd__o22a_1
X_2241_ input_ctrl_inst.scan_timer\[3\] _1052_ _0440_ _0442_ VGND VGND VPWR VPWR _0443_
+ sky130_fd_sc_hd__or4_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1887_ gencon_inst.ALU_out\[2\] net72 net45 net19 VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a22o_1
X_1956_ net329 VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput19 net19 VGND VGND VPWR VPWR display_output[2] sky130_fd_sc_hd__buf_2
X_2508_ clknet_leaf_38_clk _0079_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2439_ clknet_leaf_1_clk _0037_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1741_ net339 _0934_ net112 VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
X_2790_ clknet_leaf_12_clk _0344_ net133 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
X_1810_ gencon_inst.operand2\[12\] gencon_inst.operand1\[12\] net77 VGND VGND VPWR
+ VPWR _0974_ sky130_fd_sc_hd__mux2_1
X_1672_ _0873_ _0875_ _0880_ _0884_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__or4_1
XFILLER_7_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2155_ gencon_inst.mult_calc.finish _1202_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__and2_1
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2224_ _0408_ _0425_ _0431_ _0433_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__or4b_1
X_2086_ input_ctrl_inst.debounce_cnt\[9\] _1144_ _1147_ _1124_ VGND VGND VPWR VPWR
+ _1149_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_53_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1939_ gencon_inst.operand2\[11\] net64 net40 net318 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a22o_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold126 gencon_inst.add_calc.next_finish VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dlygate4sd3_1
X_1724_ gencon_inst.ALU_in1\[5\] gencon_inst.ALU_in2\[5\] net67 VGND VGND VPWR VPWR
+ _0926_ sky130_fd_sc_hd__mux2_1
X_2773_ clknet_leaf_23_clk net240 VGND VGND VPWR VPWR gencon_inst.ALU_in1\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold104 gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1 VGND VGND VPWR
+ VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _0202_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ _0868_ _0871_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__or2_1
X_1586_ net106 gencon_inst.add_calc.main.in2\[6\] VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__nand2_1
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold148 gencon_inst.mult_calc.adderSave\[9\] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2 VGND VGND VPWR
+ VPWR net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1 VGND VGND VPWR
+ VPWR net294 sky130_fd_sc_hd__dlygate4sd3_1
X_2069_ input_ctrl_inst.debounce_cnt\[4\] input_ctrl_inst.debounce_cnt\[5\] _1130_
+ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__and3_1
X_2138_ input_ctrl_inst.col_index\[2\] _1188_ _1187_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__mux2_1
X_2207_ _0405_ _0415_ _0416_ input_ctrl_inst.col_index\[14\] VGND VGND VPWR VPWR _0417_
+ sky130_fd_sc_hd__and4b_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1371_ net86 _1088_ net88 net244 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a2bb2o_1
X_1440_ net338 net199 net97 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2825_ clknet_leaf_25_clk net280 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2687_ clknet_leaf_16_clk _0241_ net149 VGND VGND VPWR VPWR gencon_inst.ALU_out\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_1638_ net32 _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__nand2_1
X_1707_ _0778_ _0850_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__nor2_1
X_2756_ clknet_leaf_14_clk _0310_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[8\] sky130_fd_sc_hd__dfxtp_1
X_1569_ net107 gencon_inst.add_calc.main.in2\[10\] VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__or2_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout32 _0852_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout76 _1205_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_4
Xfanout43 _0561_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
Xfanout65 _0952_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
Xfanout54 _0451_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout98 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
Xfanout87 _1032_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_9_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload35 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload35/X sky130_fd_sc_hd__clkbuf_4
X_2472_ clknet_leaf_6_clk _0013_ net128 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload13 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_8
X_2541_ clknet_leaf_0_clk net161 net121 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2610_ clknet_leaf_25_clk _0169_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload24 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_12
XFILLER_68_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1285_ gencon_inst.ALU_out\[13\] net73 net52 gencon_inst.mult_calc.out\[13\] net44
+ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__a221o_1
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1354_ net56 _0676_ _0677_ net50 gencon_inst.mult_calc.out\[11\] VGND VGND VPWR VPWR
+ _0678_ sky130_fd_sc_hd__a32o_1
X_1423_ net103 gencon_inst.mult_calc.finish _0693_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_70_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2808_ clknet_leaf_4_clk gencon_inst.next_state\[1\] net132 VGND VGND VPWR VPWR gencon_inst.gencon_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload7 clknet_leaf_35_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_12
X_2739_ clknet_leaf_21_clk _0293_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1972_ net92 net30 _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2455_ clknet_leaf_5_clk _0028_ net128 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2524_ clknet_leaf_37_clk _0095_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1268_ net444 net34 _0607_ _0608_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__o22a_1
X_1337_ net55 _0662_ _0664_ net49 gencon_inst.mult_calc.out\[7\] VGND VGND VPWR VPWR
+ _0665_ sky130_fd_sc_hd__a32o_1
Xhold19 gencon_inst.mult_calc.INn1\[3\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ net235 net227 net103 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
X_2386_ input_ctrl_inst.col_index\[17\] input_ctrl_inst.col_index\[19\] input_ctrl_inst.col_index\[18\]
+ _0518_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__and4_1
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2171_ gencon_inst.gencon_state\[1\] _0385_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nor2_1
X_2240_ input_ctrl_inst.scan_timer\[11\] _0437_ _0441_ input_ctrl_inst.scan_timer\[8\]
+ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__or4b_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1886_ _0995_ _0996_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or2_1
X_1955_ input_ctrl_inst.decoded_key\[3\] VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2438_ clknet_leaf_1_clk _0036_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_2507_ clknet_leaf_39_clk _0078_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_56_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2369_ _0514_ _0515_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__nor2_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ gencon_inst.ALU_out\[7\] _0886_ net113 VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_62_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1740_ gencon_inst.ALU_in1\[13\] gencon_inst.ALU_in2\[13\] net68 VGND VGND VPWR VPWR
+ _0934_ sky130_fd_sc_hd__mux2_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2085_ input_ctrl_inst.debounce_cnt\[9\] _1144_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__and2_1
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2154_ gencon_inst.gencon_state\[1\] _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_36_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ input_ctrl_inst.col_index\[4\] _0403_ _0432_ _0422_ VGND VGND VPWR VPWR _0433_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_44_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1869_ _1024_ _0381_ gencon_inst.prev_operator_input\[2\] gencon_inst.prev_operator_input\[0\]
+ gencon_inst.prev_operator_input\[1\] VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__a2111o_1
X_1938_ gencon_inst.operand2\[10\] net63 net40 net302 VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__a22o_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1654_ gencon_inst.ALU_out\[4\] _0872_ net113 VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
X_1723_ net324 _0925_ net110 VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
Xhold138 gencon_inst.latched_operator_input\[2\] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dlygate4sd3_1
X_2772_ clknet_leaf_14_clk _0326_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 gencon_inst.keypad_input\[2\] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2 VGND VGND VPWR
+ VPWR net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold116 gencon_inst.mult_calc.countSave\[6\] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 gencon_inst.mult_calc.countSave\[14\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
X_1585_ net106 gencon_inst.add_calc.main.in2\[6\] VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__or2_1
XFILLER_58_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2206_ input_ctrl_inst.col_index\[13\] input_ctrl_inst.col_index\[12\] input_ctrl_inst.col_index\[15\]
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__and3_1
X_2068_ input_ctrl_inst.debounce_cnt\[4\] _1130_ input_ctrl_inst.debounce_cnt\[5\]
+ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__a21o_1
X_2137_ input_ctrl_inst.RowSync\[2\] input_ctrl_inst.RowSync\[0\] input_ctrl_inst.col_index\[2\]
+ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1370_ gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn net86 net304 net88
+ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2824_ clknet_leaf_26_clk _0374_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2686_ clknet_leaf_16_clk _0240_ net149 VGND VGND VPWR VPWR gencon_inst.ALU_out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1637_ _0775_ _0854_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__nand2b_1
X_1706_ _0906_ _0908_ _0913_ _0852_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__o31a_1
X_2755_ clknet_leaf_14_clk _0309_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1 _0787_ _0788_ VGND
+ VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nand3_1
XFILLER_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1499_ gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nand2_1
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout44 _0561_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout55 _0386_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
Xfanout33 _0523_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_2
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout66 _0952_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xfanout77 _1205_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_2
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout88 net91 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xfanout99 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2471_ clknet_leaf_6_clk _0012_ net128 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload14 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinv_8
Xclkload36 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__bufinv_16
X_2540_ clknet_leaf_0_clk net158 net121 VGND VGND VPWR VPWR input_ctrl_inst.RowSync\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_9_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload25 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__inv_12
X_1422_ net86 net78 VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__nand2_1
XFILLER_68_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1284_ gencon_inst.operand1\[13\] _0616_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_50_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1353_ gencon_inst.operand2\[10\] _0668_ gencon_inst.operand2\[11\] VGND VGND VPWR
+ VPWR _0677_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2807_ clknet_leaf_4_clk gencon_inst.next_state\[0\] net132 VGND VGND VPWR VPWR gencon_inst.gencon_state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2738_ clknet_leaf_26_clk _0292_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[11\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkload8 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2669_ clknet_leaf_26_clk _0228_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1971_ input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__nor2_1
X_2454_ clknet_leaf_0_clk _0027_ net122 VGND VGND VPWR VPWR input_ctrl_inst.decoded_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1405_ gencon_inst.mult_calc.out\[14\] net375 net104 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
X_2385_ input_ctrl_inst.col_index\[17\] input_ctrl_inst.col_index\[18\] _0518_ input_ctrl_inst.col_index\[19\]
+ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a31o_1
X_2523_ clknet_leaf_38_clk _0094_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_1267_ gencon_inst.ALU_out\[9\] net74 net52 gencon_inst.mult_calc.out\[9\] net44
+ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a221o_1
X_1336_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__inv_2
XFILLER_28_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 RowIn[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_39_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ gencon_inst.gencon_state\[0\] _1030_ gencon_inst.gencon_state\[2\] VGND VGND
+ VPWR VPWR _0385_ sky130_fd_sc_hd__nand3_1
X_1954_ gencon_inst.add_calc.state\[1\] VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__inv_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1885_ net65 _0962_ net57 gencon_inst.mult_calc.out\[1\] VGND VGND VPWR VPWR _0996_
+ sky130_fd_sc_hd__a22o_1
X_2437_ clknet_leaf_1_clk _0035_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2506_ clknet_leaf_38_clk _0077_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2368_ input_ctrl_inst.col_index\[11\] input_ctrl_inst.col_index\[12\] _0513_ VGND
+ VGND VPWR VPWR _0515_ sky130_fd_sc_hd__and3_1
XFILLER_71_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1319_ gencon_inst.operand2\[3\] _0650_ net47 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
X_2299_ net128 _1053_ equal_input VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_39_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1670_ _0884_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__xnor2_1
X_2222_ input_ctrl_inst.col_index\[5\] input_ctrl_inst.col_index\[7\] input_ctrl_inst.col_index\[6\]
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__and3_1
X_2084_ input_ctrl_inst.debounce_cnt\[9\] _1057_ _1146_ VGND VGND VPWR VPWR _1147_
+ sky130_fd_sc_hd__o21bai_1
X_2153_ gencon_inst.gencon_state\[0\] gencon_inst.gencon_state\[3\] gencon_inst.gencon_state\[2\]
+ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__or3b_1
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1937_ gencon_inst.operand2\[9\] net63 net40 net362 VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1868_ _1202_ _1210_ net65 _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__or4_1
X_1799_ _0968_ net173 net40 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2771_ clknet_leaf_14_clk _0325_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1653_ _0869_ _0871_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__xnor2_1
X_1584_ gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1 _0803_ _0804_ VGND
+ VGND VPWR VPWR _0806_ sky130_fd_sc_hd__nand3_1
X_1722_ gencon_inst.ALU_in1\[4\] gencon_inst.ALU_in2\[4\] net70 VGND VGND VPWR VPWR
+ _0925_ sky130_fd_sc_hd__mux2_1
Xhold139 gencon_inst.mult_calc.adderSave\[7\] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 gencon_inst.mult_calc.adderSave\[5\] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold117 gencon_inst.mult_calc.countSave\[5\] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold106 _0074_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
X_2205_ input_ctrl_inst.col_index\[9\] input_ctrl_inst.col_index\[8\] input_ctrl_inst.col_index\[11\]
+ input_ctrl_inst.col_index\[10\] VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and4_1
X_2067_ net36 _1133_ _1134_ net38 input_ctrl_inst.debounce_cnt\[4\] VGND VGND VPWR
+ VPWR _0021_ sky130_fd_sc_hd__a32o_1
X_2136_ _1027_ input_ctrl_inst.RowSync\[1\] input_ctrl_inst.RowSync\[3\] VGND VGND
+ VPWR VPWR _1187_ sky130_fd_sc_hd__o21a_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1705_ net443 _0914_ net113 VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
X_2754_ clknet_leaf_14_clk _0308_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[6\] sky130_fd_sc_hd__dfxtp_1
X_2823_ clknet_leaf_26_clk _0373_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2685_ clknet_leaf_16_clk _0239_ net150 VGND VGND VPWR VPWR gencon_inst.ALU_out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1636_ net84 _0856_ _0857_ _0855_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__o31a_1
X_1567_ _0787_ _0788_ gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1 VGND
+ VGND VPWR VPWR _0789_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2119_ _1172_ _1174_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__and2_1
X_1498_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout67 net70 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout45 _0991_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_4
Xfanout34 _0560_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_4
Xfanout56 _0386_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout78 net81 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout89 net91 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload15 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__inv_8
Xclkload26 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__inv_12
X_2470_ clknet_leaf_6_clk _0011_ net129 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload37 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__inv_8
X_1421_ net96 gencon_inst.mult_calc.adderSave\[14\] net316 net81 VGND VGND VPWR VPWR
+ _0185_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1283_ gencon_inst.operand1\[13\] _0616_ net75 VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1352_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__inv_2
X_2806_ clknet_leaf_11_clk _0360_ net134 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_2737_ clknet_leaf_26_clk _0291_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2668_ clknet_leaf_25_clk _0227_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload9 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_6
X_1619_ _0801_ _0805_ _0839_ _0802_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__o31a_1
XFILLER_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2599_ clknet_leaf_33_clk _0158_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1970_ _1048_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2522_ clknet_leaf_37_clk _0093_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1335_ gencon_inst.operand2\[7\] _0659_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__and2_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2384_ input_ctrl_inst.col_index\[18\] net53 net33 _0524_ VGND VGND VPWR VPWR _0093_
+ sky130_fd_sc_hd__a22o_1
X_2453_ clknet_leaf_34_clk net166 VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_1404_ gencon_inst.mult_calc.out\[13\] net314 net104 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
X_1266_ gencon_inst.operand1\[9\] _0601_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__o21a_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 RowIn[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1884_ gencon_inst.ALU_out\[1\] net72 net45 net18 VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__a22o_1
X_1953_ net101 VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__inv_2
X_2505_ clknet_leaf_39_clk _0076_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1318_ net55 _0648_ _0649_ net49 gencon_inst.mult_calc.out\[3\] VGND VGND VPWR VPWR
+ _0650_ sky130_fd_sc_hd__a32o_1
X_2298_ input_ctrl_inst.decoded_key\[1\] _1198_ _1053_ net128 VGND VGND VPWR VPWR
+ _0480_ sky130_fd_sc_hd__o211ai_1
X_2436_ clknet_leaf_39_clk _0034_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2367_ input_ctrl_inst.col_index\[11\] _0513_ input_ctrl_inst.col_index\[12\] VGND
+ VGND VPWR VPWR _0514_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1249_ _0579_ _0582_ gencon_inst.operand1\[4\] gencon_inst.operand1\[5\] gencon_inst.operand1\[6\]
+ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_39_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2152_ net329 _1200_ _1182_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o21a_1
X_2221_ _0406_ _0429_ net6 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__a21boi_1
X_2083_ _1046_ _1122_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__nand2_1
XFILLER_61_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1867_ gencon_inst.key_read _0389_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1936_ gencon_inst.operand2\[8\] net63 net40 net361 VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__a22o_1
X_1798_ gencon_inst.operand2\[6\] gencon_inst.operand1\[6\] net77 VGND VGND VPWR VPWR
+ _0968_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2419_ _0427_ _0537_ input_ctrl_inst.col_index\[29\] VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a21oi_1
XFILLER_12_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ net347 _0924_ net110 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
X_2770_ clknet_leaf_14_clk net226 VGND VGND VPWR VPWR gencon_inst.ALU_in1\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _0834_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__xnor2_1
X_1583_ _0803_ _0804_ gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1 VGND
+ VGND VPWR VPWR _0805_ sky130_fd_sc_hd__a21oi_1
Xhold129 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2 VGND VGND VPWR
+ VPWR net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1 VGND VGND VPWR
+ VPWR net275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold107 input_ctrl_inst.scan_timer\[16\] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
X_2135_ _1182_ _1186_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__nand2_1
X_2204_ input_ctrl_inst.col_index\[12\] _0403_ _0404_ _0413_ VGND VGND VPWR VPWR _0414_
+ sky130_fd_sc_hd__o31a_1
X_2066_ input_ctrl_inst.debounce_cnt\[4\] _1130_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__nand2_1
X_1919_ _1018_ net234 net46 VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2684_ clknet_leaf_15_clk _0238_ net150 VGND VGND VPWR VPWR gencon_inst.ALU_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1704_ _0911_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__xnor2_1
X_2753_ clknet_leaf_14_clk _0307_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[5\] sky130_fd_sc_hd__dfxtp_1
X_2822_ clknet_leaf_26_clk net319 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1635_ _0775_ net32 _0854_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a21oi_1
X_1566_ net107 gencon_inst.add_calc.main.in2\[11\] VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__nand2_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1497_ gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2118_ net37 _1170_ input_ctrl_inst.debounce_cnt\[16\] VGND VGND VPWR VPWR _1174_
+ sky130_fd_sc_hd__or3b_1
X_2049_ _1047_ _1118_ _1120_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_1_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout68 net70 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_4
Xfanout35 _0560_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xfanout57 _0992_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
Xfanout46 _0991_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xfanout79 net81 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload16 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinv_8
Xclkload38 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__inv_8
XFILLER_9_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload27 clknet_leaf_31_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__inv_8
X_1351_ gencon_inst.operand2\[11\] gencon_inst.operand2\[10\] _0668_ VGND VGND VPWR
+ VPWR _0675_ sky130_fd_sc_hd__and3_1
X_1420_ net95 gencon_inst.mult_calc.adderSave\[13\] net286 net81 VGND VGND VPWR VPWR
+ _0184_ sky130_fd_sc_hd__a22o_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1282_ gencon_inst.operand1\[12\] net35 _0618_ _0619_ VGND VGND VPWR VPWR _0119_
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2805_ clknet_leaf_21_clk _0359_ net152 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1618_ _0805_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__nor2_1
X_2736_ clknet_leaf_25_clk _0290_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2667_ clknet_leaf_25_clk _0226_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1549_ net55 _0771_ _0772_ _1202_ gencon_inst.mult_calc.out\[15\] VGND VGND VPWR
+ VPWR _0773_ sky130_fd_sc_hd__a32o_1
X_2598_ clknet_leaf_33_clk _0157_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold290 gencon_inst.operand2\[15\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2521_ clknet_leaf_38_clk _0092_ net118 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1265_ _0556_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nor2_1
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1334_ gencon_inst.operand2\[7\] _0659_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or2_1
X_1403_ gencon_inst.mult_calc.out\[12\] net298 net104 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2383_ input_ctrl_inst.col_index\[18\] _0521_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__xnor2_1
X_2452_ clknet_leaf_34_clk _0050_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 RowIn[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2719_ clknet_leaf_16_clk _0273_ net151 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_38_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1883_ _0993_ _0994_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or2_1
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1952_ net125 VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__inv_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2435_ clknet_leaf_39_clk _0033_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2504_ clknet_leaf_39_clk _0075_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_1248_ gencon_inst.operand1\[5\] net34 _0591_ _0592_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__o22a_1
X_1317_ _0645_ _0646_ _0638_ _0640_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_39_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2297_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[1\] VGND VGND
+ VPWR VPWR _0479_ sky130_fd_sc_hd__or2_1
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2366_ net371 _0513_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__xor2_1
XFILLER_71_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2082_ _1125_ _1143_ _1145_ net38 net407 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__a32o_1
X_2151_ _1053_ _1198_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__and3_1
X_2220_ input_ctrl_inst.col_index\[24\] _0408_ _0411_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__or3_1
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1866_ net185 gencon_inst.latched_keypad_input\[3\] _0954_ VGND VGND VPWR VPWR _0341_
+ sky130_fd_sc_hd__mux2_1
X_1935_ gencon_inst.operand2\[7\] net63 net40 net394 VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__a22o_1
X_1797_ _0967_ net182 net42 VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
X_2418_ net416 net54 net33 _0548_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a22o_1
X_2349_ _0503_ _0504_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__nor2_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1651_ _0817_ _0818_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nand2b_1
X_1720_ gencon_inst.ALU_in1\[3\] gencon_inst.ALU_in2\[3\] net67 VGND VGND VPWR VPWR
+ _0924_ sky130_fd_sc_hd__mux2_1
XFILLER_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 gencon_inst.mult_calc.countSave\[10\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
X_1582_ net106 gencon_inst.add_calc.main.in2\[7\] VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold119 gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1 VGND VGND VPWR
+ VPWR net276 sky130_fd_sc_hd__dlygate4sd3_1
X_2065_ input_ctrl_inst.debounce_cnt\[4\] _1130_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ input_ctrl_inst.decoded_key\[1\] _1053_ _1185_ VGND VGND VPWR VPWR _1186_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_26_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2203_ input_ctrl_inst.col_index\[4\] input_ctrl_inst.col_index\[12\] _0402_ _0407_
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or4_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1849_ gencon_inst.operand1\[6\] net225 net61 VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
X_1918_ gencon_inst.operand1\[12\] _0990_ net58 gencon_inst.mult_calc.out\[12\] _1017_
+ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a221o_1
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2821_ clknet_leaf_26_clk _0371_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ _0775_ net32 _0854_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and3_1
X_2683_ clknet_leaf_10_clk _0237_ net134 VGND VGND VPWR VPWR gencon_inst.ALU_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1703_ _0847_ _0912_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__xnor2_1
X_2752_ clknet_leaf_15_clk _0306_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[4\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
X_1565_ net107 gencon_inst.add_calc.main.in2\[11\] VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__or2_1
X_1496_ net383 net89 _0729_ net101 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a22o_1
XFILLER_66_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2117_ input_ctrl_inst.debounce_cnt\[15\] input_ctrl_inst.debounce_cnt\[16\] _1163_
+ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__and3_1
X_2048_ _1044_ _1058_ _1118_ _1119_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_1_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout69 net70 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_2
Xfanout36 _1125_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
Xfanout58 _0992_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout47 _0629_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinv_4
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload28 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__clkinv_8
X_1281_ gencon_inst.ALU_out\[12\] net73 net52 gencon_inst.mult_calc.out\[12\] net44
+ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__a221o_1
X_1350_ gencon_inst.operand2\[10\] _0674_ net48 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_1
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
X_2804_ clknet_leaf_21_clk _0358_ net153 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1617_ _0809_ _0813_ _0836_ _0810_ _0806_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__o311a_1
X_2735_ clknet_leaf_24_clk _0289_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2597_ clknet_leaf_2_clk _0156_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2666_ clknet_leaf_25_clk _0225_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1548_ gencon_inst.operand2\[15\] _0685_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__nand2_1
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ _0706_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold280 input_ctrl_inst.debounce_cnt\[2\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1402_ gencon_inst.mult_calc.out\[11\] net377 net104 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2520_ clknet_leaf_38_clk _0091_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2451_ clknet_leaf_34_clk _0049_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_1264_ gencon_inst.operand1\[7\] gencon_inst.operand1\[8\] gencon_inst.operand1\[9\]
+ _0593_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__and4_1
X_1333_ gencon_inst.operand2\[6\] net48 _0661_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o21a_1
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 RowIn[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_2382_ input_ctrl_inst.col_index\[17\] net53 _0522_ net33 VGND VGND VPWR VPWR _0092_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2718_ clknet_leaf_14_clk _0272_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2649_ clknet_leaf_31_clk _0208_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ net65 _0961_ net57 gencon_inst.mult_calc.out\[0\] VGND VGND VPWR VPWR _0994_
+ sky130_fd_sc_hd__a22o_1
X_1951_ gencon_inst.gencon_state\[3\] VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__inv_2
X_2434_ clknet_leaf_0_clk _0032_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2503_ clknet_leaf_0_clk net4 net122 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_2365_ _0512_ _0513_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__nor2_1
XFILLER_71_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1247_ gencon_inst.ALU_out\[5\] net71 net51 gencon_inst.mult_calc.out\[5\] net43
+ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__a221o_1
X_1316_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2296_ net165 _0477_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2081_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__inv_2
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2150_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[1\] VGND VGND
+ VPWR VPWR _1199_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1934_ gencon_inst.operand2\[6\] net63 net39 net343 VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a22o_1
XFILLER_21_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1796_ gencon_inst.operand2\[5\] gencon_inst.operand1\[5\] net76 VGND VGND VPWR VPWR
+ _0967_ sky130_fd_sc_hd__mux2_1
X_1865_ net284 gencon_inst.latched_keypad_input\[2\] _0954_ VGND VGND VPWR VPWR _0340_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2417_ _0427_ _0537_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__a21oi_1
X_2348_ _1192_ _0452_ _0498_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and3_1
XFILLER_52_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2279_ net393 _0466_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nor2_1
XFILLER_75_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1650_ net32 _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_1
X_1581_ net106 gencon_inst.add_calc.main.in2\[7\] VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__or2_1
Xhold109 gencon_inst.add_calc.start VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2202_ _0406_ _0409_ _0411_ _0412_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__or4_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2064_ net36 _1131_ _1132_ net37 net281 VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_49_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ input_ctrl_inst.col_index\[1\] _1048_ net82 VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or3_1
X_1917_ gencon_inst.operand2\[12\] _1204_ net73 gencon_inst.ALU_out\[12\] VGND VGND
+ VPWR VPWR _1017_ sky130_fd_sc_hd__a22o_1
XFILLER_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1848_ gencon_inst.operand1\[5\] net230 net60 VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
X_1779_ net117 _0953_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nor2_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2751_ clknet_leaf_11_clk _0305_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[3\] sky130_fd_sc_hd__dfxtp_1
X_2820_ clknet_leaf_22_clk _0370_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2682_ clknet_leaf_10_clk _0236_ net134 VGND VGND VPWR VPWR gencon_inst.ALU_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1633_ net113 gencon_inst.ALU_out\[1\] VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__or2_1
XFILLER_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1702_ _0781_ _0782_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__and2b_1
X_1564_ gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1 _0783_ _0784_ VGND
+ VGND VPWR VPWR _0786_ sky130_fd_sc_hd__nand3_1
XFILLER_39_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1495_ _0726_ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2116_ input_ctrl_inst.debounce_cnt\[15\] net36 _1163_ input_ctrl_inst.debounce_cnt\[16\]
+ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__a31o_1
Xfanout37 _1123_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
X_2047_ _1025_ _1045_ _1057_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__or3_1
Xfanout59 _0978_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
Xfanout48 _0629_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload18 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_8
XFILLER_70_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload29 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_6
X_1280_ _0616_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2803_ clknet_leaf_21_clk _0357_ net152 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
X_2734_ clknet_leaf_24_clk _0288_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_1616_ _0809_ _0813_ _0836_ _0810_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__o31a_1
X_1547_ gencon_inst.operand2\[15\] _0685_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__or2_1
X_2665_ clknet_leaf_24_clk _0224_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2596_ clknet_leaf_34_clk _0155_ net125 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1478_ _0697_ _0700_ _0703_ _0707_ _0701_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_65_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold281 gencon_inst.ALU_out\[14\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold270 input_ctrl_inst.debounce_cnt\[12\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1401_ gencon_inst.mult_calc.out\[10\] net391 net104 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2381_ net53 _0501_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__nor2_1
X_2450_ clknet_leaf_39_clk _0048_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_1263_ gencon_inst.operand1\[8\] net34 _0603_ _0604_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__o22a_1
X_1332_ gencon_inst.mult_calc.out\[6\] net49 _0658_ _0660_ _0628_ VGND VGND VPWR VPWR
+ _0661_ sky130_fd_sc_hd__a221o_1
Xinput5 nRST VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2717_ clknet_leaf_15_clk _0271_ net149 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2579_ clknet_leaf_34_clk _0138_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2648_ clknet_leaf_31_clk _0207_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1950_ gencon_inst.gencon_state\[1\] VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__inv_2
X_1881_ gencon_inst.ALU_out\[0\] net72 net45 net11 VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a22o_1
X_2502_ clknet_leaf_0_clk net3 net121 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2433_ _1208_ net51 _0378_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a21oi_1
X_1315_ _0638_ _0640_ _0645_ _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__o211a_1
X_2364_ input_ctrl_inst.col_index\[9\] input_ctrl_inst.col_index\[10\] _0511_ VGND
+ VGND VPWR VPWR _0513_ sky130_fd_sc_hd__and3_1
X_1246_ _0556_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__nor2_1
X_2295_ _0477_ _0478_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2080_ input_ctrl_inst.debounce_cnt\[7\] input_ctrl_inst.debounce_cnt\[8\] _1139_
+ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__and3_1
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1933_ gencon_inst.operand2\[5\] net64 net39 net312 VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a22o_1
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1864_ net270 gencon_inst.latched_keypad_input\[1\] _0954_ VGND VGND VPWR VPWR _0339_
+ sky130_fd_sc_hd__mux2_1
X_1795_ _0966_ net168 net42 VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2278_ input_ctrl_inst.scan_timer\[12\] _0466_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__and2_1
X_2416_ input_ctrl_inst.col_index\[28\] _0545_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__nor2_1
X_2347_ net114 _0499_ input_ctrl_inst.col_index\[3\] VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1229_ _0576_ net75 _0575_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and3b_1
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1580_ gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1 _0799_ _0800_ VGND
+ VGND VPWR VPWR _0802_ sky130_fd_sc_hd__nand3_1
XFILLER_7_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2132_ _1181_ _1184_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__nor2_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2201_ input_ctrl_inst.col_index\[24\] _0408_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__and2_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2063_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[2\]
+ input_ctrl_inst.debounce_cnt\[3\] VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__a31o_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1847_ gencon_inst.operand1\[4\] net219 net59 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
X_1916_ _1015_ _1016_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__or2_1
X_1778_ gencon_inst.read_input net65 VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nand2_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2681_ clknet_leaf_10_clk _0235_ net134 VGND VGND VPWR VPWR gencon_inst.ALU_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1701_ _0906_ _0908_ _0852_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__o21ai_1
X_2750_ clknet_leaf_11_clk _0304_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[2\] sky130_fd_sc_hd__dfxtp_1
X_1632_ _0829_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__xnor2_1
X_1563_ _0783_ _0784_ gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1 VGND
+ VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a21oi_1
X_1494_ _0718_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__or2_1
XFILLER_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2115_ net37 _1170_ _1171_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o21a_1
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout38 _1123_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_52_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2046_ _1025_ _1048_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__xnor2_1
Xfanout49 _0627_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload19 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__inv_4
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2802_ clknet_leaf_20_clk _0356_ net156 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
X_2733_ clknet_leaf_24_clk _0287_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_2664_ clknet_leaf_25_clk _0223_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1615_ _0813_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nor2_1
X_1546_ net109 net105 _0691_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__o21a_1
X_2595_ clknet_leaf_2_clk _0154_ net125 VGND VGND VPWR VPWR gencon_inst.mult_calc.diffSign
+ sky130_fd_sc_hd__dfrtp_1
X_1477_ _0711_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_6_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _1072_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_17_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold271 gencon_inst.ALU_in1\[15\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 gencon_inst.operand2\[15\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 input_ctrl_inst.debounce_cnt\[9\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1331_ _0387_ _0659_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__nor2_1
X_1400_ gencon_inst.mult_calc.out\[9\] net305 net104 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
X_2380_ _0520_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and2_1
X_1262_ gencon_inst.ALU_out\[8\] net74 net52 gencon_inst.mult_calc.out\[8\] net43
+ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__a221o_1
XFILLER_36_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2716_ clknet_leaf_15_clk _0270_ net150 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2647_ clknet_leaf_31_clk _0206_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2578_ clknet_leaf_4_clk _0137_ net129 VGND VGND VPWR VPWR gencon_inst.read_input
+ sky130_fd_sc_hd__dfrtp_4
X_1529_ net377 net90 _0757_ net102 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__a22o_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1030_ _1208_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2501_ clknet_leaf_0_clk net2 net121 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_56_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2432_ net75 net71 VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ gencon_inst.operand2\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0646_ sky130_fd_sc_hd__or2_1
X_2294_ input_ctrl_inst.scan_timer\[18\] _0475_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__or2_1
X_2363_ input_ctrl_inst.col_index\[9\] _0511_ net424 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1245_ _1039_ _0586_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_25_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1932_ gencon_inst.operand2\[4\] net63 net39 net378 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a22o_1
X_1863_ net282 gencon_inst.latched_keypad_input\[0\] _0954_ VGND VGND VPWR VPWR _0338_
+ sky130_fd_sc_hd__mux2_1
X_1794_ gencon_inst.operand2\[4\] gencon_inst.operand1\[4\] net76 VGND VGND VPWR VPWR
+ _0966_ sky130_fd_sc_hd__mux2_1
X_2415_ net411 net54 _0546_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a21bo_1
X_1228_ _0566_ _0568_ _0572_ _0574_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__o211a_1
X_2277_ _0466_ net237 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__nor2_1
X_2346_ net114 _0499_ _0502_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_32_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2062_ _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ input_ctrl_inst.decoded_key\[0\] net82 _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a21oi_1
X_2200_ input_ctrl_inst.col_index\[28\] input_ctrl_inst.col_index\[31\] input_ctrl_inst.col_index\[30\]
+ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or4_1
XFILLER_74_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_1846_ gencon_inst.operand1\[3\] net228 net60 VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
X_1915_ net66 _0973_ net58 gencon_inst.mult_calc.out\[11\] VGND VGND VPWR VPWR _1016_
+ sky130_fd_sc_hd__a22o_1
X_1777_ net65 VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__inv_2
XFILLER_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2329_ net93 net273 net78 net294 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
XFILLER_68_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2680_ clknet_leaf_10_clk _0234_ net135 VGND VGND VPWR VPWR gencon_inst.ALU_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1700_ _0910_ _0909_ gencon_inst.ALU_out\[12\] net85 VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a2bb2o_1
X_1631_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0827_ VGND VGND
+ VPWR VPWR _0853_ sky130_fd_sc_hd__xor2_1
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1562_ net107 gencon_inst.add_calc.main.in2\[12\] VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_3_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_1493_ _0706_ _0711_ _0714_ _0719_ _0712_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__o311a_1
X_2045_ net266 net283 net113 VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a21o_1
X_2114_ net36 _1163_ input_ctrl_inst.debounce_cnt\[15\] VGND VGND VPWR VPWR _1171_
+ sky130_fd_sc_hd__a21o_1
Xfanout39 net42 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1829_ gencon_inst.operand2\[2\] net213 net60 VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2801_ clknet_leaf_21_clk _0355_ net152 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XFILLER_74_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1614_ _0817_ _0821_ _0833_ _0818_ _0814_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__o311a_1
X_2594_ clknet_leaf_9_clk _0153_ net135 VGND VGND VPWR VPWR gencon_inst.add_calc.sameSignVal
+ sky130_fd_sc_hd__dfrtp_1
X_2732_ clknet_leaf_24_clk _0286_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2663_ clknet_leaf_33_clk _0222_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1476_ gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__nand2_1
X_1545_ net375 net90 _0770_ net102 VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2028_ gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1 _1071_ VGND VGND
+ VPWR VPWR _1102_ sky130_fd_sc_hd__nor2_1
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold272 input_ctrl_inst.debounce_cnt\[5\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 input_ctrl_inst.debounce_cnt\[8\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 input_ctrl_inst.scan_timer\[7\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 input_ctrl_inst.col_index\[26\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1261_ gencon_inst.operand1\[8\] _0597_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o21a_1
X_1330_ _0644_ _0647_ gencon_inst.operand2\[6\] gencon_inst.operand2\[5\] gencon_inst.operand2\[4\]
+ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__o2111a_1
XFILLER_64_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2715_ clknet_leaf_15_clk _0269_ net150 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2577_ clknet_leaf_9_clk _0005_ net131 VGND VGND VPWR VPWR gencon_inst.add_calc.next_finish
+ sky130_fd_sc_hd__dfrtp_1
X_2646_ clknet_leaf_33_clk _0205_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1528_ _0755_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__xor2_1
X_1459_ _0694_ _0696_ _0697_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or3_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2431_ _1030_ _0379_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nor2_2
X_2500_ clknet_leaf_0_clk net1 net121 VGND VGND VPWR VPWR input_ctrl_inst.RowMid\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_56_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1244_ gencon_inst.operand1\[4\] net34 _0588_ _0589_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__o22a_1
XFILLER_49_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1313_ gencon_inst.operand2\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0645_ sky130_fd_sc_hd__nand2_1
X_2362_ net372 _0511_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__xor2_1
X_2293_ net430 _0475_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__nand2_1
XFILLER_52_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2629_ clknet_leaf_2_clk _0188_ net127 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1862_ net295 _0382_ _0383_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a21bo_1
X_1793_ _0965_ net176 net42 VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
X_1931_ gencon_inst.operand2\[3\] _0958_ _0960_ net209 VGND VGND VPWR VPWR _0364_
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2414_ _0544_ _0545_ _0523_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or3b_1
XFILLER_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1227_ _0572_ _0574_ _0566_ _0568_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__a211o_1
XFILLER_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2276_ input_ctrl_inst.scan_timer\[10\] _0464_ net236 VGND VGND VPWR VPWR _0467_
+ sky130_fd_sc_hd__a21oi_1
X_2345_ net114 _0499_ _0501_ _0452_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[3\]
+ input_ctrl_inst.debounce_cnt\[2\] VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_53_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2130_ input_ctrl_inst.col_index\[0\] net30 _1053_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__and3_1
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1914_ gencon_inst.ALU_out\[11\] net74 net46 net13 VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1845_ gencon_inst.operand1\[2\] net221 net60 VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
X_1776_ _1204_ _0380_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__or2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2328_ net93 net274 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
+ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__a22o_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2259_ input_ctrl_inst.scan_timer\[4\] _0455_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__nand2_1
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ _0778_ _0781_ _0848_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__o31a_1
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1561_ net107 gencon_inst.add_calc.main.in2\[12\] VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__or2_1
XFILLER_39_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1492_ _0724_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__and2b_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2113_ input_ctrl_inst.debounce_cnt\[15\] _1163_ _1160_ VGND VGND VPWR VPWR _1170_
+ sky130_fd_sc_hd__a21oi_1
X_2044_ net101 _1116_ _1117_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a21o_1
X_1759_ net370 _0943_ net111 VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_1
X_1828_ gencon_inst.operand2\[1\] net217 net59 VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2800_ clknet_leaf_21_clk _0354_ net152 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
X_2731_ clknet_leaf_33_clk _0285_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ _0817_ _0821_ _0833_ _0818_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__o31a_1
XFILLER_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1544_ _0768_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__xnor2_1
X_2662_ clknet_leaf_32_clk _0221_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2593_ clknet_leaf_28_clk _0152_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1475_ gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
+ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nor2_1
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2027_ _1095_ _1097_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a21o_1
XFILLER_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold284 gencon_inst.ALU_out\[0\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 gencon_inst.operand1\[15\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold240 gencon_inst.mult_calc.main.a0.in2 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 input_ctrl_inst.col_index\[19\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 input_ctrl_inst.scan_timer\[18\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1260_ _0556_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__nor2_1
XFILLER_64_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ clknet_leaf_15_clk _0268_ net134 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2576_ clknet_leaf_9_clk _0001_ net131 VGND VGND VPWR VPWR gencon_inst.add_calc.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_1527_ _0747_ _0751_ _0748_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o21a_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2645_ clknet_leaf_34_clk _0204_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1389_ gencon_inst.mult_calc.INn2\[15\] gencon_inst.mult_calc.INn1\[15\] VGND VGND
+ VPWR VPWR _0692_ sky130_fd_sc_hd__xor2_1
X_1458_ gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__nor2_1
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2430_ gencon_inst.gencon_state\[3\] _1207_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__and2_1
X_2361_ _0510_ _0511_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__nor2_1
X_1243_ gencon_inst.ALU_out\[4\] net71 net51 gencon_inst.mult_calc.out\[4\] VGND VGND
+ VPWR VPWR _0589_ sky130_fd_sc_hd__a22o_1
X_1312_ gencon_inst.operand2\[3\] gencon_inst.latched_keypad_input\[3\] VGND VGND
+ VPWR VPWR _0644_ sky130_fd_sc_hd__and2_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2292_ _0475_ net191 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__nor2_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2559_ clknet_leaf_3_clk _0122_ net133 VGND VGND VPWR VPWR gencon_inst.operand2\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_2628_ clknet_leaf_2_clk _0187_ net125 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.a0.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1930_ gencon_inst.operand2\[2\] net63 net39 net332 VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a22o_1
X_1861_ net247 _0383_ _0382_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a21bo_1
X_1792_ gencon_inst.operand1\[3\] net76 _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21o_1
XFILLER_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2413_ input_ctrl_inst.col_index\[27\] _0542_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__and2_1
X_2344_ net114 _0430_ _0498_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__and4bb_1
X_1226_ gencon_inst.operand1\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0574_ sky130_fd_sc_hd__or2_1
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2275_ input_ctrl_inst.scan_timer\[11\] input_ctrl_inst.scan_timer\[10\] _0464_ VGND
+ VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and3_1
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2060_ net36 _1128_ _1129_ net37 net437 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_57_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1913_ _1013_ _1014_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1775_ net283 gencon_inst.ALU_finish _0951_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
X_1844_ gencon_inst.operand1\[1\] net241 net59 VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
XFILLER_69_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2258_ _0455_ _0456_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and2b_1
X_2327_ net93 net258 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
+ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a22o_1
XFILLER_40_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ input_ctrl_inst.col_index\[13\] input_ctrl_inst.col_index\[15\] input_ctrl_inst.col_index\[14\]
+ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__or4_1
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1560_ gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1 _0779_ _0780_ VGND
+ VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nand3_1
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2112_ _1166_ _1167_ _1169_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__or3_1
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1491_ gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__nand2_1
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2043_ gencon_inst.mult_calc.start net104 _1066_ net98 VGND VGND VPWR VPWR _1117_
+ sky130_fd_sc_hd__a22o_1
X_1827_ gencon_inst.operand2\[0\] net212 net59 VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
X_1689_ _0901_ _0900_ gencon_inst.ALU_out\[10\] net85 VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a2bb2o_1
X_1758_ gencon_inst.ALU_in2\[7\] gencon_inst.ALU_in1\[7\] net68 VGND VGND VPWR VPWR
+ _0943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2730_ clknet_leaf_3_clk _0284_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_2661_ clknet_leaf_33_clk _0220_ net142 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1612_ _0821_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__nor2_1
X_1474_ net388 net89 _0710_ net101 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a22o_1
X_1543_ _0763_ _0765_ _0764_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__o21ba_1
XFILLER_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2592_ clknet_leaf_28_clk _0151_ net147 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2026_ gencon_inst.mult_calc.compCount.in2\[7\] _1096_ _1099_ gencon_inst.mult_calc.compCount.in2\[8\]
+ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__a22o_1
Xhold285 gencon_inst.ALU_out\[2\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 input_ctrl_inst.debounce_cnt\[6\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 net17 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold274 net10 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold263 input_ctrl_inst.col_index\[14\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 gencon_inst.mult_calc.compCount.in2\[10\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2713_ clknet_leaf_10_clk _0267_ net134 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2644_ clknet_leaf_34_clk _0203_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2575_ clknet_leaf_9_clk net109 net135 VGND VGND VPWR VPWR gencon_inst.add_calc.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1526_ _0753_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nand2b_1
X_1457_ gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__and2_1
X_1388_ net445 net322 _0691_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2009_ gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1 _1067_ VGND VGND
+ VPWR VPWR _1083_ sky130_fd_sc_hd__xnor2_1
XFILLER_73_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1311_ gencon_inst.operand2\[2\] _0643_ net47 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
X_2291_ input_ctrl_inst.scan_timer\[16\] _0473_ net190 VGND VGND VPWR VPWR _0476_
+ sky130_fd_sc_hd__a21oi_1
X_2360_ input_ctrl_inst.col_index\[8\] _0444_ _0508_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__and3_1
X_1242_ gencon_inst.operand1\[4\] _0579_ _0582_ _0587_ VGND VGND VPWR VPWR _0588_
+ sky130_fd_sc_hd__o31a_1
XFILLER_49_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2627_ clknet_leaf_34_clk _0186_ net125 VGND VGND VPWR VPWR gencon_inst.mult_calc.finish
+ sky130_fd_sc_hd__dfrtp_2
X_2558_ clknet_leaf_22_clk _0121_ net153 VGND VGND VPWR VPWR gencon_inst.operand1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1509_ _0738_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__xnor2_1
X_2489_ clknet_leaf_31_clk _0064_ net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ net373 gencon_inst.operator_input\[0\] _0384_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1791_ gencon_inst.operand2\[3\] _1204_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__and2_1
XFILLER_69_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2274_ net327 _0464_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__xor2_1
X_2412_ input_ctrl_inst.col_index\[27\] _0542_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nor2_1
X_2343_ _0418_ _0424_ _0433_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
X_1225_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1989_ gencon_inst.mult_calc.INn2\[9\] gencon_inst.mult_calc.INn2\[8\] gencon_inst.mult_calc.INn2\[11\]
+ gencon_inst.mult_calc.INn2\[10\] VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__or4_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1843_ gencon_inst.operand1\[0\] net231 net59 VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
X_1912_ net66 _0972_ net58 gencon_inst.mult_calc.out\[10\] VGND VGND VPWR VPWR _1014_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1774_ net109 net113 VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_2257_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[2\] _0435_ input_ctrl_inst.scan_timer\[3\]
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a31o_1
X_2326_ net93 net245 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1
+ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a22o_1
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2188_ input_ctrl_inst.col_index\[9\] input_ctrl_inst.col_index\[8\] input_ctrl_inst.col_index\[11\]
+ input_ctrl_inst.col_index\[10\] VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or4_1
XFILLER_48_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1490_ gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
+ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__nor2_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2111_ _1058_ _1168_ input_ctrl_inst.debounce_cnt\[14\] _1046_ VGND VGND VPWR VPWR
+ _1169_ sky130_fd_sc_hd__o211a_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 input_ctrl_inst.RowMid\[0\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
X_2042_ gencon_inst.mult_calc.compCount.in2\[14\] _1076_ _1114_ _1115_ VGND VGND VPWR
+ VPWR _1116_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1826_ net117 net266 net59 VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__a21bo_1
XFILLER_30_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1688_ net31 _0897_ _0899_ net85 VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__a31o_1
X_1757_ net333 _0942_ net111 VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2309_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[2\] _1053_ VGND
+ VGND VPWR VPWR _0487_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1611_ _0825_ _0828_ _0830_ _0826_ _0822_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__o311a_1
X_2660_ clknet_leaf_33_clk _0219_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1473_ _0708_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__xnor2_1
X_1542_ gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1
+ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__xor2_1
X_2591_ clknet_leaf_29_clk _0150_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2025_ _1071_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_59_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_68_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold253 gencon_inst.add_calc.main.a0.in1 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd3_1
X_2789_ clknet_leaf_12_clk _0343_ net132 VGND VGND VPWR VPWR gencon_inst.operand1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1809_ _0973_ net181 net41 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
Xhold220 gencon_inst.mult_calc.adderSave\[11\] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 gencon_inst.mult_calc.adderSave\[3\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2 VGND VGND VPWR
+ VPWR net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 gencon_inst.ALU_out\[13\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 gencon_inst.add_calc.main.in2\[0\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 gencon_inst.mult_calc.start VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2712_ clknet_leaf_10_clk _0266_ net135 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2574_ clknet_leaf_9_clk _0000_ net131 VGND VGND VPWR VPWR gencon_inst.add_calc.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2643_ clknet_leaf_34_clk net272 net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1387_ _0690_ net109 VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__nand2b_1
X_1525_ gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__nand2_1
X_1456_ net101 _0694_ _0695_ net303 net89 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a32o_1
X_2008_ gencon_inst.mult_calc.compCount.in2\[5\] _1081_ VGND VGND VPWR VPWR _1082_
+ sky130_fd_sc_hd__or2_1
XFILLER_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1241_ net75 _0586_ net43 VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a21o_1
X_1310_ gencon_inst.mult_calc.out\[2\] net49 _0642_ net55 VGND VGND VPWR VPWR _0643_
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2290_ input_ctrl_inst.scan_timer\[17\] input_ctrl_inst.scan_timer\[16\] _0473_ VGND
+ VGND VPWR VPWR _0475_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_22_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2557_ clknet_leaf_20_clk _0120_ net153 VGND VGND VPWR VPWR gencon_inst.operand1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2626_ clknet_leaf_25_clk net317 net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1508_ _0731_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__or2_1
X_2488_ clknet_leaf_35_clk net246 net138 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1439_ net271 gencon_inst.mult_calc.INn2\[0\] net97 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_62_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1790_ _0963_ net172 net42 VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
XFILLER_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2411_ net440 net54 net33 _0543_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__a22o_1
X_1224_ gencon_inst.operand1\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0572_ sky130_fd_sc_hd__nand2_1
X_2273_ _0464_ _0465_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__nor2_1
X_2342_ _0497_ _0499_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1988_ gencon_inst.mult_calc.INn2\[1\] gencon_inst.mult_calc.INn2\[0\] gencon_inst.mult_calc.INn2\[3\]
+ gencon_inst.mult_calc.INn2\[2\] VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__or4_1
X_2609_ clknet_leaf_27_clk _0168_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_43_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1773_ net297 _0950_ net111 VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
X_1842_ net447 net251 net59 VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
X_1911_ gencon_inst.ALU_out\[10\] net73 net46 net12 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a22o_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_40_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2256_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[3\] input_ctrl_inst.scan_timer\[2\]
+ _0435_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__and4_1
X_2187_ _0396_ _0397_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__nor2_1
X_2325_ net93 net257 net78 net299 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__a22o_1
XFILLER_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2110_ _1040_ net30 VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__nor2_1
Xhold2 input_ctrl_inst.RowMid\[3\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ gencon_inst.mult_calc.compCount.in2\[14\] _1076_ _1111_ gencon_inst.mult_calc.compCount.in2\[13\]
+ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__o22a_1
X_1756_ gencon_inst.ALU_in2\[6\] gencon_inst.ALU_in1\[6\] net70 VGND VGND VPWR VPWR
+ _0942_ sky130_fd_sc_hd__mux2_1
X_1825_ net180 _0981_ _0955_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XFILLER_30_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1687_ net31 _0897_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a21oi_1
X_2308_ input_ctrl_inst.decoded_key\[1\] input_ctrl_inst.decoded_key\[3\] _0485_ VGND
+ VGND VPWR VPWR _0486_ sky130_fd_sc_hd__nor3_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2239_ input_ctrl_inst.scan_timer\[10\] _0438_ input_ctrl_inst.scan_timer\[9\] VGND
+ VGND VPWR VPWR _0441_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1610_ _0825_ _0828_ _0830_ _0826_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__o31a_1
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2590_ clknet_leaf_29_clk _0149_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ _0700_ _0704_ _0701_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__o21ai_1
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1541_ net102 _0766_ _0767_ net314 net90 VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a32o_1
XFILLER_62_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2024_ gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1 _1070_ gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__a21oi_1
Xhold210 gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1 VGND VGND VPWR VPWR
+ net367 sky130_fd_sc_hd__dlygate4sd3_1
X_1739_ net325 _0933_ net112 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
X_1808_ gencon_inst.operand2\[11\] gencon_inst.operand1\[11\] net77 VGND VGND VPWR
+ VPWR _0973_ sky130_fd_sc_hd__mux2_1
Xhold287 gencon_inst.operand1\[9\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
X_2788_ clknet_leaf_4_clk _0342_ net132 VGND VGND VPWR VPWR gencon_inst.key_read sky130_fd_sc_hd__dfrtp_2
Xhold221 gencon_inst.mult_calc.INn2\[4\] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold243 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 VGND VGND VPWR
+ VPWR net400 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 input_ctrl_inst.col_index\[21\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold254 input_ctrl_inst.col_index\[27\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 input_ctrl_inst.col_index\[4\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 gencon_inst.mult_calc.compCount.in2\[3\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2711_ clknet_leaf_9_clk _0265_ net135 VGND VGND VPWR VPWR gencon_inst.add_calc.main.a0.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2573_ clknet_leaf_22_clk _0136_ net153 VGND VGND VPWR VPWR gencon_inst.operand2\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_1524_ gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__nor2_1
X_2642_ clknet_leaf_25_clk _0201_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1386_ gencon_inst.addOrSub _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__xnor2_1
X_1455_ gencon_inst.mult_calc.main.a0.in2 gencon_inst.mult_calc.main.a0.in1 VGND VGND
+ VPWR VPWR _0695_ sky130_fd_sc_hd__or2_1
XFILLER_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2007_ gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1 _1069_ VGND VGND
+ VPWR VPWR _1081_ sky130_fd_sc_hd__xor2_1
XFILLER_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1240_ _0579_ _0582_ gencon_inst.operand1\[4\] VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2556_ clknet_leaf_22_clk _0119_ net153 VGND VGND VPWR VPWR gencon_inst.operand1\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_1507_ _0718_ _0724_ _0727_ _0732_ _0725_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__o311a_1
X_2487_ clknet_leaf_34_clk _0062_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2625_ clknet_leaf_27_clk net287 net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1438_ net215 net196 net100 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_1369_ net100 net102 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__nor2_1
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2410_ _0541_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__nor2_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2341_ _0452_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__and2_1
X_1223_ gencon_inst.operand1\[1\] _0571_ net34 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2272_ net376 _0462_ _0445_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1987_ gencon_inst.mult_calc.INn2\[5\] gencon_inst.mult_calc.INn2\[4\] gencon_inst.mult_calc.INn2\[7\]
+ gencon_inst.mult_calc.INn2\[6\] VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__or4_1
X_2539_ clknet_leaf_5_clk _0031_ net128 VGND VGND VPWR VPWR input_ctrl_inst.read_input_flag
+ sky130_fd_sc_hd__dfrtp_1
X_2608_ clknet_leaf_26_clk _0167_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_73_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1910_ _1011_ _1012_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1772_ gencon_inst.ALU_in2\[14\] gencon_inst.ALU_in1\[14\] net68 VGND VGND VPWR VPWR
+ _0950_ sky130_fd_sc_hd__mux2_1
X_1841_ gencon_inst.operand2\[14\] net208 net62 VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2324_ net93 net244 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
+ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__a22o_1
X_2255_ net374 _0453_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2186_ input_ctrl_inst.col_index\[17\] input_ctrl_inst.col_index\[16\] input_ctrl_inst.col_index\[19\]
+ input_ctrl_inst.col_index\[18\] VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or4_1
XFILLER_43_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 input_ctrl_inst.RowMid\[2\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ gencon_inst.mult_calc.compCount.in2\[13\] _1111_ _1113_ _1078_ VGND VGND VPWR
+ VPWR _1114_ sky130_fd_sc_hd__a22o_1
XFILLER_30_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1686_ _0843_ _0898_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__xnor2_1
X_1755_ net365 _0941_ net110 VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
X_1824_ gencon_inst.read_input gencon_inst.operator_input\[2\] VGND VGND VPWR VPWR
+ _0981_ sky130_fd_sc_hd__and2b_1
X_2307_ input_ctrl_inst.decoded_key\[0\] input_ctrl_inst.decoded_key\[2\] VGND VGND
+ VPWR VPWR _0485_ sky130_fd_sc_hd__nand2_1
X_2238_ input_ctrl_inst.scan_timer\[1\] input_ctrl_inst.scan_timer\[0\] input_ctrl_inst.scan_timer\[2\]
+ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or4_1
X_2169_ _0382_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1540_ _0763_ _0764_ _0765_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1471_ _0706_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__nand2b_1
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2023_ gencon_inst.mult_calc.compCount.in2\[6\] _1080_ _1096_ gencon_inst.mult_calc.compCount.in2\[7\]
+ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__o22a_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1807_ _0972_ net178 net41 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
X_1669_ _0878_ _0880_ net31 VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__o21ai_1
Xhold211 gencon_inst.ALU_finish VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1 VGND VGND VPWR
+ VPWR net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 gencon_inst.ALU_in1\[15\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
X_1738_ gencon_inst.ALU_in1\[12\] gencon_inst.ALU_in2\[12\] net69 VGND VGND VPWR VPWR
+ _0933_ sky130_fd_sc_hd__mux2_1
Xhold266 input_ctrl_inst.debounce_cnt\[11\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 gencon_inst.operator_input\[2\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__dlygate4sd3_1
X_2787_ clknet_leaf_4_clk _0341_ net132 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[3\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold233 gencon_inst.mult_calc.compCount.in2\[13\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold277 input_ctrl_inst.col_index\[29\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 gencon_inst.mult_calc.compCount.in2\[7\] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 gencon_inst.mult_calc.compCount.in2\[14\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2710_ clknet_leaf_17_clk _0264_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2572_ clknet_leaf_22_clk _0135_ net153 VGND VGND VPWR VPWR gencon_inst.operand2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1523_ net391 net90 _0752_ net102 VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a22o_1
X_1454_ gencon_inst.mult_calc.main.a0.in2 gencon_inst.mult_calc.main.a0.in1 VGND VGND
+ VPWR VPWR _0694_ sky130_fd_sc_hd__nand2_1
X_2641_ clknet_leaf_27_clk net250 net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_67_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1385_ gencon_inst.ALU_in2\[15\] gencon_inst.ALU_in1\[15\] VGND VGND VPWR VPWR _0689_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2006_ _1070_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__nand2b_1
XFILLER_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2624_ clknet_leaf_27_clk net293 net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_2555_ clknet_leaf_20_clk _0118_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1506_ _0736_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__and2b_1
X_2486_ clknet_leaf_34_clk _0061_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_1437_ gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1 net249 net100 VGND
+ VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1368_ gencon_inst.read_input _1054_ _1200_ _1035_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a22o_1
X_1299_ gencon_inst.operand2\[1\] gencon_inst.latched_keypad_input\[1\] VGND VGND
+ VPWR VPWR _0633_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2271_ input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[9\] input_ctrl_inst.scan_timer\[8\]
+ _0459_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__and4_1
X_2340_ input_ctrl_inst.col_index\[0\] input_ctrl_inst.col_index\[1\] VGND VGND VPWR
+ VPWR _0498_ sky130_fd_sc_hd__and2_1
X_1222_ gencon_inst.ALU_out\[1\] net71 net51 gencon_inst.mult_calc.out\[1\] _0570_
+ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__a221o_1
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1986_ net93 net97 VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
X_2607_ clknet_leaf_26_clk _0166_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2469_ clknet_leaf_7_clk _0010_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2538_ clknet_leaf_0_clk net92 net122 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire83 _1051_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_24_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1840_ gencon_inst.operand2\[13\] net218 net61 VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1771_ net357 _0949_ net112 VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2254_ _0453_ _0454_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__and2_1
X_2323_ net93 net304 net78 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a22o_1
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2185_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[20\] input_ctrl_inst.col_index\[23\]
+ input_ctrl_inst.col_index\[22\] VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or4_1
X_1969_ input_ctrl_inst.RowSync\[2\] input_ctrl_inst.RowSync\[0\] input_ctrl_inst.RowSync\[1\]
+ input_ctrl_inst.RowSync\[3\] VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__and4_4
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 input_ctrl_inst.RowMid\[1\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
X_1823_ net186 _0980_ _0955_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1685_ _0793_ _0794_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nand2b_1
X_1754_ gencon_inst.ALU_in2\[5\] gencon_inst.ALU_in1\[5\] net67 VGND VGND VPWR VPWR
+ _0941_ sky130_fd_sc_hd__mux2_1
X_2306_ input_ctrl_inst.input_control_state\[2\] _1048_ _1049_ _1181_ net116 VGND
+ VGND VPWR VPWR _0484_ sky130_fd_sc_hd__a311oi_4
X_2237_ input_ctrl_inst.scan_timer\[5\] input_ctrl_inst.scan_timer\[7\] input_ctrl_inst.scan_timer\[6\]
+ input_ctrl_inst.scan_timer\[4\] VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or4bb_1
X_2099_ input_ctrl_inst.debounce_cnt\[12\] _1153_ _1158_ _1124_ VGND VGND VPWR VPWR
+ _1159_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2168_ gencon_inst.operator_input\[2\] _0380_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nand2_1
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2022_ gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1 _1070_ VGND VGND
+ VPWR VPWR _1096_ sky130_fd_sc_hd__xnor2_1
Xhold201 gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1 VGND VGND VPWR
+ VPWR net358 sky130_fd_sc_hd__dlygate4sd3_1
X_1806_ gencon_inst.operand2\[10\] gencon_inst.operand1\[10\] net77 VGND VGND VPWR
+ VPWR _0972_ sky130_fd_sc_hd__mux2_1
X_2786_ clknet_leaf_4_clk _0340_ net132 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_28_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1668_ _0838_ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__xnor2_1
X_1599_ _0819_ _0820_ gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1 VGND
+ VGND VPWR VPWR _0821_ sky130_fd_sc_hd__a21oi_1
X_1737_ net315 _0932_ net112 VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold256 gencon_inst.operator_input\[1\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 gencon_inst.operand2\[15\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_37_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold234 gencon_inst.mult_calc.adderSave\[10\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 input_ctrl_inst.scan_timer\[15\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 gencon_inst.mult_calc.compCount.in2\[6\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 input_ctrl_inst.col_index\[10\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _0209_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 input_ctrl_inst.col_index\[8\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2640_ clknet_leaf_26_clk net164 net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
X_2571_ clknet_leaf_22_clk _0134_ net153 VGND VGND VPWR VPWR gencon_inst.operand2\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_1522_ _0749_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__xnor2_1
X_1453_ net412 net279 net99 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
XFILLER_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2005_ gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1 gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
+ _1068_ gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1 VGND VGND VPWR
+ VPWR _1079_ sky130_fd_sc_hd__a31o_1
X_1384_ net87 _1076_ net90 net262 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2769_ clknet_leaf_14_clk _0323_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2554_ clknet_leaf_20_clk _0117_ net152 VGND VGND VPWR VPWR gencon_inst.operand1\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_2623_ clknet_leaf_26_clk net309 net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1367_ gencon_inst.operand2\[14\] _0687_ net48 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_1
X_1436_ gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1 net163 net99 VGND
+ VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_28_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1505_ gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__nand2_1
X_2485_ clknet_leaf_35_clk _0060_ net126 VGND VGND VPWR VPWR gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1298_ gencon_inst.operand2\[0\] net47 _0630_ _0632_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1221_ _0568_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__nor2_1
X_2270_ _0445_ _0461_ _0463_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1985_ input_ctrl_inst.input_control_state\[2\] _1049_ _1053_ gencon_inst.key_read
+ _1047_ VGND VGND VPWR VPWR input_ctrl_inst.next_state\[2\] sky130_fd_sc_hd__a221o_1
X_2537_ clknet_leaf_0_clk net169 net122 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
X_2606_ clknet_leaf_26_clk _0165_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2468_ clknet_leaf_7_clk _0009_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1419_ net95 gencon_inst.mult_calc.adderSave\[12\] net292 net80 VGND VGND VPWR VPWR
+ _0183_ sky130_fd_sc_hd__a22o_1
X_2399_ input_ctrl_inst.col_index\[22\] net33 _0530_ input_ctrl_inst.col_index\[23\]
+ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__a31o_1
XFILLER_73_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1770_ gencon_inst.ALU_in2\[13\] gencon_inst.ALU_in1\[13\] net68 VGND VGND VPWR VPWR
+ _0949_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2184_ gencon_inst.mult_calc.finish net368 _0389_ VGND VGND VPWR VPWR gencon_inst.next_state\[3\]
+ sky130_fd_sc_hd__o21ba_1
X_2322_ _0484_ _0495_ _0496_ net185 net115 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a32o_1
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2253_ input_ctrl_inst.scan_timer\[1\] _0435_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or2_1
XFILLER_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1899_ gencon_inst.ALU_out\[6\] _0558_ net45 net23 VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a22o_1
X_1968_ _1044_ _1046_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 gencon_inst.prev_read_input VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1753_ net367 _0940_ net110 VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
X_1822_ gencon_inst.read_input gencon_inst.operator_input\[1\] VGND VGND VPWR VPWR
+ _0980_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_17_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1684_ _0887_ _0889_ _0894_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__or3_1
XFILLER_72_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2167_ gencon_inst.operator_input\[1\] _0380_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nand2_1
X_2305_ net401 net115 _0482_ _0483_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__a22o_1
X_2236_ input_ctrl_inst.scan_timer\[13\] input_ctrl_inst.scan_timer\[12\] input_ctrl_inst.scan_timer\[15\]
+ input_ctrl_inst.scan_timer\[14\] VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__or4bb_1
XPHY_EDGE_ROW_13_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2098_ input_ctrl_inst.debounce_cnt\[12\] _1057_ _1146_ VGND VGND VPWR VPWR _1158_
+ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_51_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2021_ gencon_inst.mult_calc.compCount.in2\[6\] _1080_ _1082_ _1094_ VGND VGND VPWR
+ VPWR _1095_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold224 gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1 VGND VGND VPWR
+ VPWR net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1 VGND VGND VPWR VPWR
+ net370 sky130_fd_sc_hd__dlygate4sd3_1
X_1736_ gencon_inst.ALU_in1\[11\] gencon_inst.ALU_in2\[11\] net69 VGND VGND VPWR VPWR
+ _0932_ sky130_fd_sc_hd__mux2_1
X_2785_ clknet_leaf_1_clk _0339_ net125 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_1805_ _0971_ net183 net40 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
Xhold202 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2 VGND VGND VPWR
+ VPWR net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 input_ctrl_inst.col_index\[7\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__dlygate4sd3_1
X_1667_ _0805_ _0806_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and2b_1
X_1598_ net105 gencon_inst.add_calc.main.in2\[3\] VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__nand2_1
Xhold257 gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1 VGND VGND VPWR VPWR
+ net414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 gencon_inst.operand2\[5\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 input_ctrl_inst.col_index\[5\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 gencon_inst.mult_calc.compCount.in2\[11\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2219_ _0412_ _0427_ _0428_ _0426_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__a31o_1
XFILLER_41_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2570_ clknet_leaf_21_clk _0133_ net152 VGND VGND VPWR VPWR gencon_inst.operand2\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_10_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1521_ gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
+ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__o21bai_1
X_1383_ net87 _1111_ net90 net268 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a2bb2o_1
X_1452_ net390 net288 net99 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_55_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2004_ gencon_inst.mult_calc.compCount.in2\[12\] _1077_ VGND VGND VPWR VPWR _1078_
+ sky130_fd_sc_hd__or2_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2699_ clknet_leaf_11_clk _0253_ net134 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1719_ net323 _0923_ net109 VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
X_2768_ clknet_leaf_14_clk _0322_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2553_ clknet_leaf_23_clk _0116_ net153 VGND VGND VPWR VPWR gencon_inst.operand1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2622_ clknet_leaf_26_clk net321 net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1504_ gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
+ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__nor2_1
X_1366_ _0685_ _0686_ gencon_inst.mult_calc.out\[14\] net50 VGND VGND VPWR VPWR _0687_
+ sky130_fd_sc_hd__a2bb2o_1
X_2484_ clknet_leaf_4_clk _0059_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_1435_ net192 net181 net100 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1297_ gencon_inst.operand2\[0\] gencon_inst.latched_keypad_input\[0\] _0628_ _0631_
+ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ _0562_ _0567_ _0556_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_35_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1984_ net92 net169 _1060_ VGND VGND VPWR VPWR input_ctrl_inst.next_state\[1\] sky130_fd_sc_hd__a21oi_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2467_ clknet_leaf_7_clk _0026_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2605_ clknet_leaf_25_clk _0164_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2536_ clknet_leaf_0_clk net167 net122 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1349_ gencon_inst.mult_calc.out\[10\] net50 _0672_ _0673_ VGND VGND VPWR VPWR _0674_
+ sky130_fd_sc_hd__a22o_1
X_1418_ net95 gencon_inst.mult_calc.adderSave\[11\] net308 net80 VGND VGND VPWR VPWR
+ _0182_ sky130_fd_sc_hd__a22o_1
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2398_ input_ctrl_inst.col_index\[22\] net53 _0533_ _0534_ VGND VGND VPWR VPWR _0097_
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2321_ gencon_inst.keypad_input\[3\] _1053_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or2_1
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2183_ _1202_ _0394_ _0395_ VGND VGND VPWR VPWR gencon_inst.next_state\[2\] sky130_fd_sc_hd__or3_1
X_2252_ input_ctrl_inst.scan_timer\[1\] _0435_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__nand2_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1898_ _1003_ _1004_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or2_1
X_1967_ input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ net92 VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nand3b_2
XFILLER_68_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2519_ clknet_leaf_36_clk _0090_ net126 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 gencon_inst.mult_calc.INn1\[12\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_1683_ _0896_ _0895_ gencon_inst.ALU_out\[9\] net85 VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a2bb2o_1
X_1752_ gencon_inst.ALU_in2\[4\] gencon_inst.ALU_in1\[4\] net70 VGND VGND VPWR VPWR
+ _0940_ sky130_fd_sc_hd__mux2_1
X_1821_ net170 _0979_ _0955_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
X_2304_ _1034_ input_ctrl_inst.decoded_key\[2\] VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ input_ctrl_inst.debounce_cnt\[12\] _1153_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__and2_1
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2166_ gencon_inst.operator_input\[2\] gencon_inst.operator_input\[1\] VGND VGND
+ VPWR VPWR _0381_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ input_ctrl_inst.scan_timer\[17\] input_ctrl_inst.scan_timer\[16\] input_ctrl_inst.scan_timer\[19\]
+ input_ctrl_inst.scan_timer\[18\] VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_51_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2020_ gencon_inst.mult_calc.compCount.in2\[5\] _1081_ _1092_ gencon_inst.mult_calc.compCount.in2\[4\]
+ _1093_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1666_ _0882_ _0881_ gencon_inst.ALU_out\[6\] net84 VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a2bb2o_1
X_1735_ net291 _0931_ net112 VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
Xhold258 input_ctrl_inst.debounce_cnt\[17\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__dlygate4sd3_1
X_1804_ gencon_inst.operand2\[9\] gencon_inst.operand1\[9\] net77 VGND VGND VPWR VPWR
+ _0971_ sky130_fd_sc_hd__mux2_1
X_2784_ clknet_leaf_2_clk _0338_ net125 VGND VGND VPWR VPWR gencon_inst.latched_keypad_input\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold269 gencon_inst.mult_calc.start VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 gencon_inst.mult_calc.adderSave\[8\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 input_ctrl_inst.scan_timer\[12\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _0179_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 input_ctrl_inst.col_index\[11\] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 gencon_inst.mult_calc.compCount.in2\[8\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlygate4sd3_1
X_1597_ net105 gencon_inst.add_calc.main.in2\[3\] VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__or2_1
X_2149_ input_ctrl_inst.decoded_key\[0\] _1034_ input_ctrl_inst.decoded_key\[2\] VGND
+ VGND VPWR VPWR _1198_ sky130_fd_sc_hd__or3b_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2218_ input_ctrl_inst.col_index\[29\] input_ctrl_inst.col_index\[31\] input_ctrl_inst.col_index\[30\]
+ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and3_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1520_ _0731_ _0736_ _0739_ _0743_ _0737_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_10_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1382_ net87 _1077_ net90 net260 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__a2bb2o_1
X_1451_ net335 gencon_inst.mult_calc.INn2\[12\] net100 VGND VGND VPWR VPWR _0214_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2003_ gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1 _1073_ VGND VGND
+ VPWR VPWR _1077_ sky130_fd_sc_hd__xnor2_1
X_1649_ _0858_ _0861_ _0865_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__or3_1
X_2698_ clknet_leaf_11_clk _0252_ net134 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1718_ gencon_inst.ALU_in1\[2\] gencon_inst.ALU_in2\[2\] net67 VGND VGND VPWR VPWR
+ _0923_ sky130_fd_sc_hd__mux2_1
X_2767_ clknet_leaf_15_clk _0321_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2552_ clknet_leaf_23_clk _0115_ net148 VGND VGND VPWR VPWR gencon_inst.operand1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2483_ clknet_leaf_4_clk _0058_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1503_ net101 _0734_ _0735_ net296 net88 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a32o_1
X_2621_ clknet_leaf_25_clk _0180_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
X_1296_ gencon_inst.operand2\[0\] gencon_inst.latched_keypad_input\[0\] _0387_ VGND
+ VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a21oi_1
X_1365_ gencon_inst.operand2\[14\] _0682_ net56 VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__o21ai_1
X_1434_ net194 net178 net100 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2819_ clknet_leaf_23_clk _0369_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ gencon_inst.key_read net82 _1056_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__o211a_1
X_2604_ clknet_leaf_25_clk _0163_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2466_ clknet_leaf_8_clk _0025_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1417_ net95 gencon_inst.mult_calc.adderSave\[10\] net320 net80 VGND VGND VPWR VPWR
+ _0181_ sky130_fd_sc_hd__a22o_1
X_2535_ clknet_leaf_36_clk _0106_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_1279_ gencon_inst.operand1\[12\] _0612_ net75 VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__o21ai_1
X_1348_ gencon_inst.operand2\[10\] _0668_ net56 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__o21a_1
X_2397_ input_ctrl_inst.col_index\[22\] _0530_ net33 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__a21boi_1
XFILLER_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout151 net156 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__buf_2
Xfanout140 net142 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
XFILLER_15_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2320_ _1199_ _0479_ _0483_ _1054_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__a31o_1
X_2251_ _0435_ _0436_ _0445_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and3b_1
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2182_ gencon_inst.read_input equal_input _1204_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o21a_1
X_1966_ input_ctrl_inst.input_control_state\[1\] input_ctrl_inst.input_control_state\[0\]
+ net92 VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__and3b_1
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1897_ gencon_inst.ALU_out\[5\] net72 net65 _0967_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a22o_1
XFILLER_56_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2449_ clknet_leaf_1_clk _0047_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2518_ clknet_leaf_36_clk _0089_ net120 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_54_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 _0199_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_70_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1820_ gencon_inst.read_input _1024_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1682_ net31 _0892_ _0894_ net85 VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__a31o_1
X_1751_ net352 _0939_ net110 VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
X_2303_ net413 net115 _1034_ _0482_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__a22o_1
X_2234_ net122 _1048_ net83 input_ctrl_inst.scan_timer\[0\] VGND VGND VPWR VPWR _0436_
+ sky130_fd_sc_hd__a31o_1
X_2096_ net423 net37 _1156_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a21bo_1
X_2165_ gencon_inst.gencon_state\[3\] _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ net94 VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2783_ clknet_leaf_4_clk _0337_ net129 VGND VGND VPWR VPWR gencon_inst.latched_operator_input\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1803_ _0970_ net174 net40 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1665_ net31 _0878_ _0880_ net84 VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__a31o_1
X_1596_ gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1 _0815_ _0816_ VGND
+ VGND VPWR VPWR _0818_ sky130_fd_sc_hd__nand3_1
X_1734_ gencon_inst.ALU_in1\[10\] gencon_inst.ALU_in2\[10\] net69 VGND VGND VPWR VPWR
+ _0931_ sky130_fd_sc_hd__mux2_1
Xhold237 gencon_inst.mult_calc.INn2\[7\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 gencon_inst.mult_calc.INn2\[8\] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 gencon_inst.mult_calc.adderSave\[6\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 input_ctrl_inst.col_index\[28\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold248 input_ctrl_inst.col_index\[16\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 input_ctrl_inst.col_index\[9\] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ input_ctrl_inst.col_index\[25\] input_ctrl_inst.col_index\[27\] input_ctrl_inst.col_index\[26\]
+ input_ctrl_inst.col_index\[28\] VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_64_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2079_ input_ctrl_inst.debounce_cnt\[7\] _1139_ input_ctrl_inst.debounce_cnt\[8\]
+ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__a21o_1
XFILLER_34_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2148_ input_ctrl_inst.decoded_key\[3\] net82 _1181_ _1197_ VGND VGND VPWR VPWR _0030_
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_24_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ net403 net318 net99 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XFILLER_67_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1381_ net87 _1109_ net90 net254 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_61_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2002_ gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1 _1075_ VGND VGND
+ VPWR VPWR _1076_ sky130_fd_sc_hd__xor2_1
X_2766_ clknet_leaf_11_clk net222 VGND VGND VPWR VPWR gencon_inst.ALU_in1\[2\] sky130_fd_sc_hd__dfxtp_1
X_1648_ _0867_ _0866_ gencon_inst.ALU_out\[3\] net84 VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__a2bb2o_1
X_1579_ _0799_ _0800_ gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1 VGND
+ VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a21oi_1
X_2697_ clknet_leaf_9_clk _0251_ net135 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1717_ net346 _0922_ net109 VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2620_ clknet_leaf_25_clk net360 net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2551_ clknet_leaf_14_clk _0114_ net148 VGND VGND VPWR VPWR gencon_inst.operand1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2482_ clknet_leaf_1_clk _0057_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_1433_ net195 net183 net99 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
X_1502_ _0730_ _0732_ _0733_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__a21o_1
X_1295_ gencon_inst.mult_calc.out\[0\] net49 VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__and2_1
X_1364_ gencon_inst.operand2\[14\] _0682_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2749_ clknet_leaf_11_clk _0303_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[1\] sky130_fd_sc_hd__dfxtp_1
X_2818_ clknet_leaf_24_clk _0368_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1982_ net30 _1051_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nand2_1
X_2603_ clknet_leaf_24_clk _0162_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2534_ clknet_leaf_36_clk _0105_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_2465_ clknet_leaf_8_clk _0024_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1347_ gencon_inst.operand2\[10\] _0668_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__nand2_1
X_1416_ net96 net305 net400 net81 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__a22o_1
X_2396_ input_ctrl_inst.col_index\[22\] _0530_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or2_1
X_1278_ gencon_inst.operand1\[12\] _0612_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__and2_1
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout130 net137 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout152 net153 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout141 net142 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__inv_2
XFILLER_65_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2181_ _0384_ _0393_ _0394_ VGND VGND VPWR VPWR gencon_inst.next_state\[1\] sky130_fd_sc_hd__or3_1
X_1965_ input_ctrl_inst.debounce_cnt\[14\] _1043_ _1040_ VGND VGND VPWR VPWR _1044_
+ sky130_fd_sc_hd__o21a_1
X_1896_ net22 net45 net57 gencon_inst.mult_calc.out\[5\] VGND VGND VPWR VPWR _1003_
+ sky130_fd_sc_hd__a22o_1
X_2517_ clknet_leaf_36_clk _0088_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_75_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2448_ clknet_leaf_1_clk _0046_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2379_ input_ctrl_inst.col_index\[17\] _0518_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_54_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 input_ctrl_inst.scan_timer\[19\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1750_ gencon_inst.ALU_in2\[3\] gencon_inst.ALU_in1\[3\] net67 VGND VGND VPWR VPWR
+ _0939_ sky130_fd_sc_hd__mux2_1
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1681_ net31 _0892_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2164_ gencon_inst.gencon_state\[1\] gencon_inst.gencon_state\[0\] gencon_inst.gencon_state\[2\]
+ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__or3_2
X_2302_ gencon_inst.operator_input\[0\] net115 input_ctrl_inst.decoded_key\[2\] _0482_
+ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__a22o_1
X_2233_ input_ctrl_inst.scan_timer\[0\] net122 _1048_ net83 VGND VGND VPWR VPWR _0435_
+ sky130_fd_sc_hd__and4_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2095_ _1124_ _1154_ _1155_ _1153_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__a211o_1
XFILLER_53_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1879_ _0557_ net65 VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__nor2_1
X_1948_ input_ctrl_inst.RowSync\[2\] VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__inv_2
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1733_ net326 _0930_ net111 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
X_2782_ clknet_leaf_6_clk _0336_ net129 VGND VGND VPWR VPWR gencon_inst.latched_operator_input\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1802_ gencon_inst.operand2\[8\] gencon_inst.operand1\[8\] net76 VGND VGND VPWR VPWR
+ _0970_ sky130_fd_sc_hd__mux2_1
XFILLER_43_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664_ net31 _0878_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a21oi_1
Xhold227 gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1 VGND VGND VPWR
+ VPWR net384 sky130_fd_sc_hd__dlygate4sd3_1
X_1595_ _0815_ _0816_ gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1 VGND
+ VGND VPWR VPWR _0817_ sky130_fd_sc_hd__a21oi_1
Xhold216 gencon_inst.latched_operator_input\[0\] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 gencon_inst.mult_calc.INn2\[9\] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 gencon_inst.mult_calc.adderSave\[4\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold249 gencon_inst.mult_calc.state\[0\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__dlygate4sd3_1
X_2147_ input_ctrl_inst.RowSync\[3\] _1191_ _1192_ _1196_ _1053_ VGND VGND VPWR VPWR
+ _1197_ sky130_fd_sc_hd__o311a_1
XFILLER_26_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2216_ input_ctrl_inst.col_index\[24\] _0408_ _0411_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_64_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2078_ _1125_ _1141_ _1142_ net38 input_ctrl_inst.debounce_cnt\[7\] VGND VGND VPWR
+ VPWR _0024_ sky130_fd_sc_hd__a32o_1
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1380_ net87 _1105_ net90 net265 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2001_ gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1 _1074_ VGND VGND
+ VPWR VPWR _1075_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2696_ clknet_leaf_9_clk _0250_ net135 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1716_ gencon_inst.ALU_in1\[1\] gencon_inst.ALU_in2\[1\] net67 VGND VGND VPWR VPWR
+ _0922_ sky130_fd_sc_hd__mux2_1
X_2765_ clknet_leaf_11_clk _0319_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1647_ net32 _0863_ _0865_ net84 VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a31o_1
X_1578_ net106 gencon_inst.add_calc.main.in2\[8\] VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__nand2_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ clknet_leaf_14_clk _0113_ net148 VGND VGND VPWR VPWR gencon_inst.operand1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1363_ gencon_inst.operand2\[13\] _0684_ net48 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
X_2481_ clknet_leaf_1_clk _0056_ VGND VGND VPWR VPWR gencon_inst.keypad_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_1432_ net188 net174 net99 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
X_1501_ _0730_ _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nand3_1
X_1294_ _1203_ net55 _0557_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_43_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2748_ clknet_leaf_11_clk _0302_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2679_ clknet_leaf_3_clk _0233_ net132 VGND VGND VPWR VPWR gencon_inst.operand2\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_2817_ clknet_leaf_24_clk _0367_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1981_ _1044_ _1057_ _1055_ _1047_ VGND VGND VPWR VPWR input_ctrl_inst.next_state\[0\]
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_43_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2602_ clknet_leaf_32_clk _0161_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2533_ clknet_leaf_37_clk _0104_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2464_ clknet_leaf_8_clk _0023_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1346_ gencon_inst.operand2\[9\] _0671_ net48 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux2_1
X_1415_ net96 gencon_inst.mult_calc.adderSave\[8\] net359 net81 VGND VGND VPWR VPWR
+ _0179_ sky130_fd_sc_hd__a22o_1
X_2395_ net422 net53 _0532_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__a21o_1
X_1277_ gencon_inst.operand1\[11\] net35 _0614_ _0615_ VGND VGND VPWR VPWR _0118_
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_31_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
Xfanout131 net137 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xfanout120 net127 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout153 net156 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout142 net157 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_57_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2180_ gencon_inst.mult_calc.finish gencon_inst.ALU_finish _0389_ _0388_ VGND VGND
+ VPWR VPWR _0394_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_48_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1895_ _1001_ _1002_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
X_1964_ _1041_ _1042_ input_ctrl_inst.debounce_cnt\[13\] VGND VGND VPWR VPWR _1043_
+ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_2447_ clknet_leaf_34_clk _0045_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2516_ clknet_leaf_36_clk _0087_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1329_ gencon_inst.operand2\[5\] _0651_ gencon_inst.operand2\[6\] VGND VGND VPWR
+ VPWR _0658_ sky130_fd_sc_hd__a21o_1
X_2378_ input_ctrl_inst.col_index\[17\] _0518_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 _0051_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1680_ _0841_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__xnor2_1
X_2301_ net116 _1181_ _1199_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__nor3_1
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2163_ gencon_inst.mult_calc.finish _1209_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
X_2232_ net103 net406 net426 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__o21ba_1
XFILLER_65_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2094_ input_ctrl_inst.debounce_cnt\[10\] _1148_ input_ctrl_inst.debounce_cnt\[11\]
+ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1947_ input_ctrl_inst.debounce_cnt\[13\] VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__inv_2
X_1878_ _1204_ _0557_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nor2_1
XFILLER_9_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1663_ _0837_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__xnor2_1
X_1732_ gencon_inst.ALU_in1\[9\] gencon_inst.ALU_in2\[9\] net68 VGND VGND VPWR VPWR
+ _0930_ sky130_fd_sc_hd__mux2_1
X_2781_ clknet_leaf_4_clk _0335_ net129 VGND VGND VPWR VPWR gencon_inst.latched_operator_input\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1801_ _0969_ net184 net40 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
Xhold217 input_ctrl_inst.scan_timer\[2\] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold206 gencon_inst.mult_calc.compCount.in2\[2\] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__dlygate4sd3_1
X_1594_ net105 gencon_inst.add_calc.main.in2\[4\] VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nand2_1
Xhold239 gencon_inst.mult_calc.adderSave\[2\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold228 gencon_inst.mult_calc.compCount.in2\[9\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_64_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2077_ input_ctrl_inst.debounce_cnt\[7\] _1139_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nand2_1
XFILLER_53_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2146_ input_ctrl_inst.RowSync\[2\] _1193_ _1194_ _1195_ VGND VGND VPWR VPWR _1196_
+ sky130_fd_sc_hd__a31o_1
X_2215_ _0418_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nand2_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2000_ gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1 _1073_ VGND VGND
+ VPWR VPWR _1074_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1646_ net32 _0863_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a21oi_1
X_1715_ net432 _0921_ net109 VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
X_2695_ clknet_leaf_9_clk _0249_ net134 VGND VGND VPWR VPWR gencon_inst.ALU_out\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2764_ clknet_leaf_11_clk _0318_ VGND VGND VPWR VPWR gencon_inst.ALU_in1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1577_ net106 gencon_inst.add_calc.main.in2\[8\] VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__or2_1
X_2129_ _1044_ _1045_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__nand2_1
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2480_ clknet_leaf_4_clk _0055_ VGND VGND VPWR VPWR gencon_inst.operator_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1500_ _0724_ _0728_ _0725_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__o21ai_1
X_1293_ _1203_ net49 VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__and2b_1
X_1362_ _0682_ _0683_ gencon_inst.mult_calc.out\[13\] net50 VGND VGND VPWR VPWR _0684_
+ sky130_fd_sc_hd__a2bb2o_1
X_1431_ net201 net184 net99 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
XFILLER_63_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2816_ clknet_leaf_24_clk net313 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1629_ _1038_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nor2_1
X_2747_ clknet_leaf_7_clk _0301_ VGND VGND VPWR VPWR gencon_inst.add_calc.start sky130_fd_sc_hd__dfxtp_1
X_2678_ clknet_leaf_32_clk _0004_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1980_ net92 _1056_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2463_ clknet_leaf_8_clk _0022_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2601_ clknet_leaf_24_clk _0160_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2532_ clknet_leaf_36_clk _0103_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1276_ gencon_inst.ALU_out\[11\] net73 net52 gencon_inst.mult_calc.out\[11\] net44
+ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__a221o_1
X_1345_ net56 _0669_ _0670_ net50 gencon_inst.mult_calc.out\[9\] VGND VGND VPWR VPWR
+ _0671_ sky130_fd_sc_hd__a32o_1
X_1414_ net94 gencon_inst.mult_calc.adderSave\[7\] net289 net79 VGND VGND VPWR VPWR
+ _0178_ sky130_fd_sc_hd__a22o_1
X_2394_ _0530_ _0531_ net33 VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_34_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout110 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xfanout154 net156 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net136 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout143 net147 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net123 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1963_ input_ctrl_inst.debounce_cnt\[9\] input_ctrl_inst.debounce_cnt\[11\] input_ctrl_inst.debounce_cnt\[10\]
+ input_ctrl_inst.debounce_cnt\[12\] VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__or4_1
X_1894_ net65 _0966_ net57 gencon_inst.mult_calc.out\[4\] VGND VGND VPWR VPWR _1002_
+ sky130_fd_sc_hd__a22o_1
X_2446_ clknet_leaf_2_clk _0044_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_2515_ clknet_leaf_36_clk _0086_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1259_ gencon_inst.operand1\[7\] gencon_inst.operand1\[8\] _0593_ VGND VGND VPWR
+ VPWR _0601_ sky130_fd_sc_hd__and3_1
X_1328_ _0628_ _0655_ _0657_ _0656_ net436 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__o32a_1
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2377_ _0452_ _0518_ _0519_ net405 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2300_ net115 _1182_ _0480_ _0481_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__o211a_1
X_2231_ net421 net406 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and2_1
X_2093_ input_ctrl_inst.debounce_cnt\[11\] _1057_ _1146_ VGND VGND VPWR VPWR _1154_
+ sky130_fd_sc_hd__o21bai_1
X_2162_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__inv_2
XFILLER_38_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1877_ _1030_ net431 _0379_ _0557_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a31o_1
X_1946_ input_ctrl_inst.debounce_cnt\[0\] VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_59_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2429_ _1029_ gencon_inst.gencon_state\[0\] gencon_inst.gencon_state\[3\] gencon_inst.gencon_state\[2\]
+ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or4_4
XFILLER_71_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ gencon_inst.operand2\[7\] gencon_inst.operand1\[7\] net76 VGND VGND VPWR VPWR
+ _0969_ sky130_fd_sc_hd__mux2_1
X_1662_ _0809_ _0810_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__nand2b_1
X_1731_ net337 _0929_ net111 VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
X_2780_ clknet_leaf_4_clk _0334_ VGND VGND VPWR VPWR gencon_inst.prev_read_input sky130_fd_sc_hd__dfxtp_1
Xhold207 input_ctrl_inst.scan_timer\[5\] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 gencon_inst.mult_calc.adderSave\[14\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold229 gencon_inst.mult_calc.compCount.in2\[4\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__dlygate4sd3_1
X_1593_ net105 gencon_inst.add_calc.main.in2\[4\] VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__or2_1
X_2214_ _0421_ _0398_ _0423_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2076_ input_ctrl_inst.debounce_cnt\[7\] _1139_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__or2_1
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2145_ input_ctrl_inst.RowSync\[2\] input_ctrl_inst.col_index\[3\] input_ctrl_inst.RowSync\[3\]
+ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__o21ai_1
X_1929_ gencon_inst.operand2\[1\] _0958_ _0960_ net199 VGND VGND VPWR VPWR _0362_
+ sky130_fd_sc_hd__o22a_1
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 gencon_inst.latched_operator_input\[1\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2763_ clknet_leaf_9_clk _0317_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1645_ _0832_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__xor2_1
X_2694_ clknet_leaf_17_clk _0248_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1576_ gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1 _0795_ _0796_ VGND
+ VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nand3_1
X_1714_ gencon_inst.ALU_in1\[0\] gencon_inst.ALU_in2\[0\] net67 VGND VGND VPWR VPWR
+ _0921_ sky130_fd_sc_hd__mux2_1
XFILLER_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2059_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[2\]
+ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a21o_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2128_ _1044_ _1045_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__and2_2
XFILLER_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1430_ net189 net173 net98 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
X_1361_ gencon_inst.operand2\[13\] _0679_ net56 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__o21ai_1
X_1292_ net55 _0557_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__nor2_1
XFILLER_51_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2746_ clknet_leaf_6_clk _0300_ VGND VGND VPWR VPWR gencon_inst.prev_operator_input\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_2815_ clknet_leaf_24_clk _0365_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1559_ _0779_ _0780_ gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1 VGND
+ VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a21oi_1
X_1628_ gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1 _0776_ _0777_ VGND
+ VGND VPWR VPWR _0850_ sky130_fd_sc_hd__and3_1
X_2677_ clknet_leaf_34_clk _0003_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2600_ clknet_leaf_32_clk _0159_ net140 VGND VGND VPWR VPWR gencon_inst.mult_calc.out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2462_ clknet_leaf_8_clk _0021_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ net94 gencon_inst.mult_calc.adderSave\[6\] net353 net79 VGND VGND VPWR VPWR
+ _0177_ sky130_fd_sc_hd__a22o_1
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2531_ clknet_leaf_36_clk _0102_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_2393_ input_ctrl_inst.col_index\[20\] _0526_ input_ctrl_inst.col_index\[21\] VGND
+ VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a21o_1
XFILLER_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1275_ _0612_ _0613_ net75 VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__and3b_1
X_1344_ gencon_inst.operand2\[8\] gencon_inst.operand2\[7\] _0659_ gencon_inst.operand2\[9\]
+ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__a31o_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2729_ clknet_leaf_3_clk _0283_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout155 net156 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
Xfanout111 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout133 net136 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xfanout122 net123 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout100 gencon_inst.mult_calc.state\[3\] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_2
Xfanout144 net147 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1962_ input_ctrl_inst.debounce_cnt\[5\] input_ctrl_inst.debounce_cnt\[7\] input_ctrl_inst.debounce_cnt\[6\]
+ input_ctrl_inst.debounce_cnt\[8\] VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1893_ gencon_inst.ALU_out\[4\] net72 net45 net21 VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2445_ clknet_leaf_2_clk _0043_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_2376_ _0418_ _0433_ _0452_ _0508_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__and4_1
X_2514_ clknet_leaf_39_clk _0085_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1258_ gencon_inst.operand1\[7\] net34 _0599_ _0600_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__o22a_1
X_1327_ gencon_inst.operand2\[5\] _0651_ _0387_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_67_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ net87 _1116_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__nor2_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2092_ input_ctrl_inst.debounce_cnt\[11\] input_ctrl_inst.debounce_cnt\[10\] _1148_
+ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__and3_1
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2161_ gencon_inst.gencon_state\[3\] _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__or2_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1945_ gencon_inst.operator_input\[0\] VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1876_ net43 _0987_ _0988_ _0989_ net419 VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_8_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2428_ _1029_ gencon_inst.gencon_state\[0\] gencon_inst.gencon_state\[3\] gencon_inst.gencon_state\[2\]
+ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__nor4_2
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2359_ net435 _0509_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__nor2_1
XFILLER_71_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1661_ _0873_ _0875_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__or2_1
X_1592_ gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1 _0811_ _0812_ VGND
+ VGND VPWR VPWR _0814_ sky130_fd_sc_hd__nand3_1
Xhold208 gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1 VGND VGND VPWR VPWR
+ net365 sky130_fd_sc_hd__dlygate4sd3_1
X_1730_ gencon_inst.ALU_in1\[8\] gencon_inst.ALU_in2\[8\] net68 VGND VGND VPWR VPWR
+ _0929_ sky130_fd_sc_hd__mux2_1
Xhold219 input_ctrl_inst.scan_timer\[9\] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2144_ input_ctrl_inst.RowSync\[0\] input_ctrl_inst.col_index\[3\] input_ctrl_inst.RowSync\[1\]
+ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__or3b_1
X_2213_ _0401_ _0422_ _0408_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_64_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2075_ _1125_ _1138_ _1140_ net38 net387 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__a32o_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1859_ net162 gencon_inst.read_input _0955_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__mux2_1
X_1928_ gencon_inst.operand2\[0\] net63 net39 net307 VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a22o_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold91 gencon_inst.ALU_in1\[7\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 _0467_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
X_1713_ gencon_inst.ALU_in1\[15\] _0690_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nand2_1
X_2762_ clknet_leaf_20_clk _0316_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[14\] sky130_fd_sc_hd__dfxtp_1
X_2693_ clknet_leaf_18_clk _0247_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1575_ _0795_ _0796_ gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1 VGND
+ VGND VPWR VPWR _0797_ sky130_fd_sc_hd__a21oi_2
X_1644_ _0821_ _0822_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__nand2b_1
X_2127_ _1045_ _1180_ _1178_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__o21a_1
XFILLER_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2058_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] input_ctrl_inst.debounce_cnt\[2\]
+ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nand3_1
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1360_ gencon_inst.operand2\[13\] gencon_inst.operand2\[12\] _0675_ VGND VGND VPWR
+ VPWR _0682_ sky130_fd_sc_hd__and3_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1291_ gencon_inst.operand1\[14\] net35 _0625_ _0626_ VGND VGND VPWR VPWR _0121_
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2745_ clknet_leaf_4_clk _0299_ VGND VGND VPWR VPWR gencon_inst.prev_operator_input\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2814_ clknet_leaf_33_clk net210 VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2676_ clknet_leaf_32_clk _0007_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1627_ _0781_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__nor2_1
X_1558_ net106 gencon_inst.add_calc.main.in2\[13\] VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__nand2_1
X_1489_ net101 _0722_ _0723_ net285 net89 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a32o_1
XFILLER_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_34_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_43_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ clknet_leaf_37_clk _0101_ net119 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2461_ clknet_leaf_8_clk _0020_ net130 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1343_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__inv_2
X_1412_ net94 net285 net306 net79 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__a22o_1
X_2392_ input_ctrl_inst.col_index\[21\] input_ctrl_inst.col_index\[20\] _0526_ VGND
+ VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and3_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ gencon_inst.operand1\[10\] _0605_ gencon_inst.operand1\[11\] VGND VGND VPWR
+ VPWR _0613_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_24_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2728_ clknet_leaf_2_clk _0282_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_2659_ clknet_leaf_2_clk _0218_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout112 gencon_inst.add_calc.state\[2\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xfanout134 net136 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
Xfanout101 net102 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net147 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_4
Xfanout123 net127 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1961_ input_ctrl_inst.debounce_cnt\[15\] input_ctrl_inst.debounce_cnt\[17\] input_ctrl_inst.debounce_cnt\[16\]
+ input_ctrl_inst.debounce_cnt\[18\] VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and4_1
X_1892_ _0999_ _1000_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2513_ clknet_leaf_39_clk _0084_ net123 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
X_1326_ _0651_ _0655_ net47 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__o21a_1
X_2444_ clknet_leaf_2_clk _0042_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_2375_ input_ctrl_inst.col_index\[16\] _0418_ _0508_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and3_1
X_1257_ gencon_inst.ALU_out\[7\] net74 net51 gencon_inst.mult_calc.out\[7\] net43
+ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a221o_1
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2160_ gencon_inst.gencon_state\[0\] _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__nand2_1
X_2091_ _1151_ _1152_ input_ctrl_inst.debounce_cnt\[10\] net38 VGND VGND VPWR VPWR
+ _0009_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1875_ gencon_inst.operator_input\[0\] gencon_inst.key_read _0380_ _0381_ net34 VGND
+ VGND VPWR VPWR _0989_ sky130_fd_sc_hd__a41o_1
X_1944_ net116 net421 _0960_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_16_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2427_ _1037_ net54 _0552_ _0554_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__o31a_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1309_ _0640_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__nor2_1
X_2358_ _0507_ _0509_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__nor2_1
X_2289_ net264 _0473_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__xor2_1
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1660_ _0877_ _0876_ gencon_inst.ALU_out\[5\] net84 VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a2bb2o_1
X_1591_ _0811_ _0812_ gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1 VGND
+ VGND VPWR VPWR _0813_ sky130_fd_sc_hd__a21oi_1
Xhold209 gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1 VGND VGND VPWR VPWR
+ net366 sky130_fd_sc_hd__dlygate4sd3_1
X_2143_ _1191_ _1192_ input_ctrl_inst.RowSync\[1\] VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__o21bai_1
X_2212_ _0404_ _0407_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nor2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2074_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1927_ net65 _0977_ net45 net409 _1023_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a221o_1
X_1858_ net419 net428 net59 VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_1
X_1789_ gencon_inst.operand2\[2\] gencon_inst.operand1\[2\] net76 VGND VGND VPWR VPWR
+ _0963_ sky130_fd_sc_hd__mux2_1
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold81 gencon_inst.ALU_in1\[8\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 gencon_inst.mult_calc.diffSign VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 gencon_inst.mult_calc.INn1\[13\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2830_ clknet_leaf_2_clk _0377_ VGND VGND VPWR VPWR gencon_inst.mult_calc.start sky130_fd_sc_hd__dfxtp_1
XFILLER_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1643_ _0858_ _0861_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__or2_1
X_2692_ clknet_leaf_17_clk _0246_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_1712_ net113 net330 net32 _0919_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__o22a_1
X_2761_ clknet_leaf_20_clk _0315_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 _0560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ net106 gencon_inst.add_calc.main.in2\[9\] VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__nand2_1
XFILLER_66_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2057_ net36 _1126_ _1127_ net37 input_ctrl_inst.debounce_cnt\[1\] VGND VGND VPWR
+ VPWR _0018_ sky130_fd_sc_hd__a32o_1
X_2126_ _1057_ _1122_ _1177_ _1179_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_24_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1290_ gencon_inst.ALU_out\[14\] net74 net52 gencon_inst.mult_calc.out\[14\] net43
+ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__a221o_1
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2813_ clknet_leaf_3_clk _0363_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_1626_ _0785_ _0789_ _0845_ _0786_ _0782_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__o311a_1
X_2744_ clknet_leaf_4_clk _0298_ VGND VGND VPWR VPWR gencon_inst.prev_operator_input\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2675_ clknet_leaf_32_clk _0006_ net141 VGND VGND VPWR VPWR gencon_inst.mult_calc.next_finish
+ sky130_fd_sc_hd__dfrtp_1
X_1557_ net106 gencon_inst.add_calc.main.in2\[13\] VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__or2_1
X_1488_ _0720_ _0721_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nand2_1
X_2109_ _1040_ _1045_ net30 input_ctrl_inst.debounce_cnt\[14\] VGND VGND VPWR VPWR
+ _1167_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_37_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2460_ clknet_leaf_8_clk _0019_ net131 VGND VGND VPWR VPWR input_ctrl_inst.debounce_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1273_ gencon_inst.operand1\[10\] gencon_inst.operand1\[11\] _0605_ VGND VGND VPWR
+ VPWR _0612_ sky130_fd_sc_hd__and3_1
X_1342_ gencon_inst.operand2\[9\] gencon_inst.operand2\[8\] gencon_inst.operand2\[7\]
+ _0659_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__and4_1
X_2391_ net33 _0529_ _0528_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a21o_1
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1411_ net94 gencon_inst.mult_calc.adderSave\[4\] net355 net79 VGND VGND VPWR VPWR
+ _0175_ sky130_fd_sc_hd__a22o_1
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1609_ _0828_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__nor2_1
Xfanout113 gencon_inst.add_calc.state\[1\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
X_2727_ clknet_leaf_2_clk _0281_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_2658_ clknet_leaf_34_clk _0217_ net124 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2589_ clknet_leaf_29_clk _0148_ net143 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout102 gencon_inst.mult_calc.state\[2\] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xfanout157 net5 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
Xfanout124 net125 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_40_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1960_ gencon_inst.operand1\[5\] VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__inv_2
X_1891_ net20 net45 net57 gencon_inst.mult_calc.out\[3\] _0964_ VGND VGND VPWR VPWR
+ _1000_ sky130_fd_sc_hd__a221o_1
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2443_ clknet_leaf_2_clk _0041_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_2512_ clknet_leaf_1_clk _0083_ net123 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1256_ _0597_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__nor2_1
X_1325_ gencon_inst.mult_calc.out\[5\] net49 VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__and2_1
X_2374_ net216 _0517_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__xor2_1
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ input_ctrl_inst.debounce_cnt\[10\] _1148_ _1150_ _1124_ VGND VGND VPWR VPWR
+ _1152_ sky130_fd_sc_hd__a22o_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1874_ gencon_inst.gencon_state\[0\] gencon_inst.mult_calc.out\[15\] _1207_ net71
+ gencon_inst.ALU_out\[15\] VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__a32o_1
X_1943_ net446 net63 net39 net198 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2426_ input_ctrl_inst.col_index\[30\] _0523_ _0550_ input_ctrl_inst.col_index\[31\]
+ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_67_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1239_ gencon_inst.operand1\[3\] net34 _0584_ _0585_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__o22a_1
X_1308_ _0638_ _0639_ _0633_ _0636_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__o211a_1
X_2357_ _0444_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__and2_1
X_2288_ _0473_ _0474_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__nor2_1
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1590_ net108 gencon_inst.add_calc.main.in2\[5\] VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__nand2_1
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2073_ input_ctrl_inst.debounce_cnt\[4\] input_ctrl_inst.debounce_cnt\[5\] input_ctrl_inst.debounce_cnt\[6\]
+ _1130_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__and4_1
X_2142_ input_ctrl_inst.col_index\[2\] input_ctrl_inst.col_index\[3\] VGND VGND VPWR
+ VPWR _1192_ sky130_fd_sc_hd__and2_1
X_2211_ input_ctrl_inst.col_index\[18\] _0419_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1857_ gencon_inst.operand1\[14\] net205 net62 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
X_1926_ _1204_ _0557_ _0988_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__o21a_1
X_1788_ _0962_ net171 net39 VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2409_ input_ctrl_inst.col_index\[25\] input_ctrl_inst.col_index\[26\] _0537_ VGND
+ VGND VPWR VPWR _0542_ sky130_fd_sc_hd__and3_1
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold60 gencon_inst.ALU_in2\[1\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 gencon_inst.ALU_in1\[3\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 gencon_inst.ALU_in1\[9\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 _0200_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2691_ clknet_leaf_18_clk _0245_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1642_ net442 _0862_ net113 VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
X_1711_ _1038_ gencon_inst.add_calc.sameSignVal net84 VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a21o_1
X_2760_ clknet_leaf_20_clk _0314_ VGND VGND VPWR VPWR gencon_inst.ALU_in2\[12\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_2 _0952_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1573_ net106 gencon_inst.add_calc.main.in2\[9\] VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__or2_1
XFILLER_66_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2056_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] VGND VGND
+ VPWR VPWR _1127_ sky130_fd_sc_hd__nand2_1
X_2125_ _1058_ _1121_ input_ctrl_inst.debounce_cnt\[18\] VGND VGND VPWR VPWR _1179_
+ sky130_fd_sc_hd__o21a_1
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1909_ net66 _0971_ net57 gencon_inst.mult_calc.out\[9\] VGND VGND VPWR VPWR _1012_
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2743_ clknet_leaf_7_clk net278 VGND VGND VPWR VPWR gencon_inst.addOrSub sky130_fd_sc_hd__dfxtp_1
X_2812_ clknet_leaf_2_clk _0362_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1625_ _0785_ _0789_ _0845_ _0786_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__o31a_1
X_1556_ _0776_ _0777_ gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1 VGND
+ VGND VPWR VPWR _0778_ sky130_fd_sc_hd__a21oi_1
X_2674_ clknet_leaf_34_clk _0002_ net125 VGND VGND VPWR VPWR gencon_inst.mult_calc.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1487_ _0720_ _0721_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or2_1
X_2108_ _1124_ _1164_ _1165_ _1163_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_37_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ _1107_ _1110_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_20_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1410_ net94 gencon_inst.mult_calc.adderSave\[3\] net300 net79 VGND VGND VPWR VPWR
+ _0174_ sky130_fd_sc_hd__a22o_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1272_ gencon_inst.operand1\[10\] net35 _0610_ _0611_ VGND VGND VPWR VPWR _0117_
+ sky130_fd_sc_hd__o22a_1
X_1341_ gencon_inst.operand2\[8\] net47 _0667_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__o21a_1
X_2390_ input_ctrl_inst.col_index\[20\] _0526_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__xor2_1
X_2726_ clknet_leaf_9_clk _0280_ net135 VGND VGND VPWR VPWR gencon_inst.ALU_finish
+ sky130_fd_sc_hd__dfrtp_1
X_1608_ gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1 _0827_ _0829_ VGND
+ VGND VPWR VPWR _0830_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout136 net137 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
X_1539_ _0763_ _0764_ _0765_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__or3_1
Xfanout103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
X_2588_ clknet_leaf_30_clk _0147_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout147 net157 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
Xfanout114 input_ctrl_inst.col_index\[2\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
X_2657_ clknet_leaf_27_clk _0216_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold190 gencon_inst.add_calc.main.in2\[3\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1890_ gencon_inst.operand1\[3\] _0380_ net71 gencon_inst.ALU_out\[3\] VGND VGND
+ VPWR VPWR _0999_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2442_ clknet_leaf_1_clk _0040_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_2511_ clknet_leaf_39_clk _0082_ net123 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2373_ _0516_ _0517_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__nor2_1
X_1255_ gencon_inst.operand1\[7\] _0593_ net75 VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__o21ai_1
X_1324_ gencon_inst.operand2\[4\] net47 _0654_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2709_ clknet_leaf_20_clk _0263_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_45_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1942_ gencon_inst.operand2\[14\] net64 net40 net279 VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_54_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1873_ gencon_inst.operand1\[15\] _0623_ _0986_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__o21a_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2425_ input_ctrl_inst.col_index\[30\] net54 _0553_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__a21o_1
X_2356_ _1192_ _0433_ _0498_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_67_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1238_ gencon_inst.ALU_out\[3\] net71 net51 gencon_inst.mult_calc.out\[3\] net43
+ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a221o_1
X_1307_ _0633_ _0636_ _0638_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a211oi_1
X_2287_ net402 _0471_ _0445_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ input_ctrl_inst.col_index\[17\] input_ctrl_inst.col_index\[16\] input_ctrl_inst.col_index\[19\]
+ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and3_1
X_2072_ input_ctrl_inst.debounce_cnt\[6\] _1136_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__or2_1
XFILLER_38_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2141_ input_ctrl_inst.col_index\[2\] input_ctrl_inst.col_index\[3\] VGND VGND VPWR
+ VPWR _1191_ sky130_fd_sc_hd__nor2_1
XFILLER_61_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1925_ _1022_ net243 net46 VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
X_1856_ gencon_inst.operand1\[13\] net232 net61 VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux2_1
X_1787_ gencon_inst.operand2\[1\] gencon_inst.operand1\[1\] net76 VGND VGND VPWR VPWR
+ _0962_ sky130_fd_sc_hd__mux2_1
XFILLER_57_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2408_ input_ctrl_inst.col_index\[25\] _0537_ input_ctrl_inst.col_index\[26\] VGND
+ VGND VPWR VPWR _0541_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2339_ input_ctrl_inst.col_index\[0\] _0452_ input_ctrl_inst.col_index\[1\] VGND
+ VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a21oi_1
XFILLER_71_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold61 gencon_inst.ALU_in2\[13\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 gencon_inst.ALU_in2\[15\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold50 gencon_inst.ALU_in2\[12\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 gencon_inst.ALU_in2\[7\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 _0327_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2690_ clknet_leaf_18_clk _0244_ net154 VGND VGND VPWR VPWR gencon_inst.ALU_out\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1641_ _0859_ _0861_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__xnor2_1
X_1572_ gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1 _0791_ _0792_ VGND
+ VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nand3_1
X_1710_ net438 _0918_ gencon_inst.add_calc.state\[1\] VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2124_ input_ctrl_inst.debounce_cnt\[18\] _1122_ _1177_ _1121_ _1046_ VGND VGND VPWR
+ VPWR _1178_ sky130_fd_sc_hd__a221o_1
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2055_ input_ctrl_inst.debounce_cnt\[1\] input_ctrl_inst.debounce_cnt\[0\] VGND VGND
+ VPWR VPWR _1126_ sky130_fd_sc_hd__or2_1
XFILLER_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1839_ gencon_inst.operand2\[12\] net207 net62 VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
X_1908_ gencon_inst.ALU_out\[9\] net73 net46 net26 VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a22o_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_25_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_75_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2742_ clknet_leaf_3_clk _0296_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_2811_ clknet_leaf_3_clk _0361_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn2\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1624_ _0789_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__nor2_1
X_2673_ clknet_leaf_9_clk _0232_ net135 VGND VGND VPWR VPWR gencon_inst.add_calc.diffSign
+ sky130_fd_sc_hd__dfrtp_1
X_1555_ net107 gencon_inst.add_calc.main.in2\[14\] VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
X_2107_ input_ctrl_inst.debounce_cnt\[13\] _1157_ input_ctrl_inst.debounce_cnt\[14\]
+ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1486_ _0711_ _0715_ _0712_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o21a_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2038_ gencon_inst.mult_calc.compCount.in2\[12\] _1077_ _1109_ gencon_inst.mult_calc.compCount.in2\[11\]
+ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__a22o_1
XFILLER_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1340_ gencon_inst.mult_calc.out\[8\] net49 _0666_ net55 _0628_ VGND VGND VPWR VPWR
+ _0667_ sky130_fd_sc_hd__a221o_1
X_1271_ gencon_inst.ALU_out\[10\] net73 net52 gencon_inst.mult_calc.out\[10\] net44
+ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__a221o_1
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_2725_ clknet_leaf_17_clk _0279_ net154 VGND VGND VPWR VPWR gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2656_ clknet_leaf_27_clk _0215_ net144 VGND VGND VPWR VPWR gencon_inst.mult_calc.compCount.in2\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_1607_ net105 gencon_inst.add_calc.main.a0.in1 gencon_inst.add_calc.main.in2\[0\]
+ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__mux2_1
Xfanout148 net151 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
Xfanout115 net116 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
X_1469_ gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
+ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nor2_1
X_1538_ _0758_ _0760_ _0759_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__a21boi_1
Xfanout104 gencon_inst.mult_calc.next_finish VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_4
X_2587_ clknet_leaf_30_clk _0146_ net139 VGND VGND VPWR VPWR gencon_inst.mult_calc.countSave\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
Xfanout137 net5 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
XFILLER_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold180 gencon_inst.add_calc.main.in2\[8\] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold191 gencon_inst.add_calc.main.in2\[5\] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2510_ clknet_leaf_39_clk _0081_ net121 VGND VGND VPWR VPWR input_ctrl_inst.col_index\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1323_ gencon_inst.mult_calc.out\[4\] net49 _0652_ _0653_ VGND VGND VPWR VPWR _0654_
+ sky130_fd_sc_hd__a22o_1
X_2441_ clknet_leaf_1_clk _0039_ VGND VGND VPWR VPWR input_ctrl_inst.scan_timer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_2372_ input_ctrl_inst.col_index\[13\] input_ctrl_inst.col_index\[14\] _0515_ VGND
+ VGND VPWR VPWR _0517_ sky130_fd_sc_hd__and3_1
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1254_ gencon_inst.operand1\[7\] _0593_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__and2_1
XFILLER_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2708_ clknet_leaf_20_clk _0262_ net155 VGND VGND VPWR VPWR gencon_inst.add_calc.main.in2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2639_ clknet_leaf_26_clk _0198_ net146 VGND VGND VPWR VPWR gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1872_ gencon_inst.operand1\[15\] _0623_ _0556_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__a21oi_1
X_1941_ gencon_inst.operand2\[13\] net64 net41 net288 VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__a22o_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1306_ gencon_inst.operand2\[2\] gencon_inst.latched_keypad_input\[2\] VGND VGND
+ VPWR VPWR _0639_ sky130_fd_sc_hd__nor2_1
X_2424_ input_ctrl_inst.col_index\[30\] _0550_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__o21a_1
X_2355_ input_ctrl_inst.col_index\[6\] _0506_ net392 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21oi_1
X_2286_ input_ctrl_inst.scan_timer\[15\] _0471_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_67_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1237_ _0582_ _0583_ net75 VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__and3b_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ input_ctrl_inst.decoded_key\[2\] net82 _1181_ _1190_ VGND VGND VPWR VPWR _0029_
+ sky130_fd_sc_hd__a211o_1
X_2071_ net36 _1135_ _1137_ net37 net429 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__a32o_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1855_ gencon_inst.operand1\[12\] net224 net62 VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
X_1924_ gencon_inst.operand1\[14\] _0990_ net58 gencon_inst.mult_calc.out\[14\] _1021_
+ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__a221o_1
XFILLER_39_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1786_ _0961_ net193 net39 VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
X_2269_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__inv_2
X_2407_ net33 _0540_ _0539_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a21o_1
X_2338_ input_ctrl_inst.col_index\[0\] _0451_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 gencon_inst.ALU_in2\[4\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 gencon_inst.ALU_in1\[1\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 gencon_inst.ALU_in1\[5\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 gencon_inst.ALU_in1\[4\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 gencon_inst.ALU_in2\[14\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold95 gencon_inst.mult_calc.countSave\[8\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1640_ _0831_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__xnor2_1
X_1571_ _0791_ _0792_ gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1 VGND
+ VGND VPWR VPWR _0793_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2123_ _1040_ _1163_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__a21oi_1
X_2054_ _1047_ _1048_ _1057_ _1122_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__a22o_1
X_1838_ gencon_inst.operand2\[11\] net206 net62 VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
X_1907_ _1009_ _1010_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__or2_1
X_1769_ net358 _0948_ net112 VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput30 net30 VGND VGND VPWR VPWR key_pressed sky130_fd_sc_hd__buf_2
Xoutput6 net6 VGND VGND VPWR VPWR ColOut[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2810_ clknet_leaf_4_clk gencon_inst.next_state\[3\] net132 VGND VGND VPWR VPWR gencon_inst.gencon_state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_2741_ clknet_leaf_25_clk _0295_ VGND VGND VPWR VPWR gencon_inst.mult_calc.INn1\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_2672_ clknet_leaf_27_clk _0231_ net145 VGND VGND VPWR VPWR gencon_inst.mult_calc.adderSave\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_1623_ _0793_ _0797_ _0842_ _0794_ _0790_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__o311a_1
X_1554_ net107 gencon_inst.add_calc.main.in2\[14\] VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__or2_1
X_1485_ _0717_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nand2_1
.ends

