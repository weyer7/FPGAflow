VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO calculator_top
  CLASS BLOCK ;
  FOREIGN calculator_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 218.215 BY 228.935 ;
  PIN ColOut[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END ColOut[0]
  PIN ColOut[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END ColOut[1]
  PIN ColOut[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END ColOut[2]
  PIN ColOut[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END ColOut[3]
  PIN RowIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END RowIn[0]
  PIN RowIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END RowIn[1]
  PIN RowIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END RowIn[2]
  PIN RowIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END RowIn[3]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 217.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 212.760 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 212.760 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 217.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 212.760 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 212.760 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END clk
  PIN complete
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 224.935 103.410 228.935 ;
    END
  END complete
  PIN display_output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 224.935 87.310 228.935 ;
    END
  END display_output[0]
  PIN display_output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 132.640 218.215 133.240 ;
    END
  END display_output[10]
  PIN display_output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 156.440 218.215 157.040 ;
    END
  END display_output[11]
  PIN display_output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 122.440 218.215 123.040 ;
    END
  END display_output[12]
  PIN display_output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 142.840 218.215 143.440 ;
    END
  END display_output[13]
  PIN display_output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 125.840 218.215 126.440 ;
    END
  END display_output[14]
  PIN display_output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 224.935 100.190 228.935 ;
    END
  END display_output[15]
  PIN display_output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 224.935 96.970 228.935 ;
    END
  END display_output[1]
  PIN display_output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 224.935 113.070 228.935 ;
    END
  END display_output[2]
  PIN display_output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 224.935 116.290 228.935 ;
    END
  END display_output[3]
  PIN display_output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 224.935 125.950 228.935 ;
    END
  END display_output[4]
  PIN display_output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 129.240 218.215 129.840 ;
    END
  END display_output[5]
  PIN display_output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 224.935 145.270 228.935 ;
    END
  END display_output[6]
  PIN display_output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 136.040 218.215 136.640 ;
    END
  END display_output[7]
  PIN display_output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 139.440 218.215 140.040 ;
    END
  END display_output[8]
  PIN display_output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 214.215 146.240 218.215 146.840 ;
    END
  END display_output[9]
  PIN input_state_FPGA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END input_state_FPGA[0]
  PIN input_state_FPGA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END input_state_FPGA[1]
  PIN input_state_FPGA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END input_state_FPGA[2]
  PIN key_pressed
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END key_pressed
  PIN nRST
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 214.215 17.040 218.215 17.640 ;
    END
  END nRST
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 212.710 217.685 ;
      LAYER li1 ;
        RECT 5.520 10.795 212.520 217.685 ;
      LAYER met1 ;
        RECT 4.210 10.640 212.820 217.840 ;
      LAYER met2 ;
        RECT 4.230 224.655 86.750 225.490 ;
        RECT 87.590 224.655 96.410 225.490 ;
        RECT 97.250 224.655 99.630 225.490 ;
        RECT 100.470 224.655 102.850 225.490 ;
        RECT 103.690 224.655 112.510 225.490 ;
        RECT 113.350 224.655 115.730 225.490 ;
        RECT 116.570 224.655 125.390 225.490 ;
        RECT 126.230 224.655 144.710 225.490 ;
        RECT 145.550 224.655 211.050 225.490 ;
        RECT 4.230 4.280 211.050 224.655 ;
        RECT 4.230 4.000 57.770 4.280 ;
        RECT 58.610 4.000 211.050 4.280 ;
      LAYER met3 ;
        RECT 3.990 208.440 214.215 217.765 ;
        RECT 4.400 207.040 214.215 208.440 ;
        RECT 3.990 157.440 214.215 207.040 ;
        RECT 3.990 156.040 213.815 157.440 ;
        RECT 3.990 147.240 214.215 156.040 ;
        RECT 3.990 145.840 213.815 147.240 ;
        RECT 3.990 143.840 214.215 145.840 ;
        RECT 3.990 142.440 213.815 143.840 ;
        RECT 3.990 140.440 214.215 142.440 ;
        RECT 3.990 139.040 213.815 140.440 ;
        RECT 3.990 137.040 214.215 139.040 ;
        RECT 3.990 135.640 213.815 137.040 ;
        RECT 3.990 133.640 214.215 135.640 ;
        RECT 4.400 132.240 213.815 133.640 ;
        RECT 3.990 130.240 214.215 132.240 ;
        RECT 3.990 128.840 213.815 130.240 ;
        RECT 3.990 126.840 214.215 128.840 ;
        RECT 3.990 125.440 213.815 126.840 ;
        RECT 3.990 123.440 214.215 125.440 ;
        RECT 3.990 122.040 213.815 123.440 ;
        RECT 3.990 113.240 214.215 122.040 ;
        RECT 4.400 111.840 214.215 113.240 ;
        RECT 3.990 109.840 214.215 111.840 ;
        RECT 4.400 108.440 214.215 109.840 ;
        RECT 3.990 106.440 214.215 108.440 ;
        RECT 4.400 105.040 214.215 106.440 ;
        RECT 3.990 89.440 214.215 105.040 ;
        RECT 4.400 88.040 214.215 89.440 ;
        RECT 3.990 86.040 214.215 88.040 ;
        RECT 4.400 84.640 214.215 86.040 ;
        RECT 3.990 79.240 214.215 84.640 ;
        RECT 4.400 77.840 214.215 79.240 ;
        RECT 3.990 75.840 214.215 77.840 ;
        RECT 4.400 74.440 214.215 75.840 ;
        RECT 3.990 62.240 214.215 74.440 ;
        RECT 4.400 60.840 214.215 62.240 ;
        RECT 3.990 58.840 214.215 60.840 ;
        RECT 4.400 57.440 214.215 58.840 ;
        RECT 3.990 55.440 214.215 57.440 ;
        RECT 4.400 54.040 214.215 55.440 ;
        RECT 3.990 18.040 214.215 54.040 ;
        RECT 3.990 16.640 213.815 18.040 ;
        RECT 3.990 10.715 214.215 16.640 ;
      LAYER met4 ;
        RECT 26.975 68.175 174.240 214.705 ;
        RECT 176.640 68.175 177.540 214.705 ;
        RECT 179.940 68.175 191.065 214.705 ;
  END
END calculator_top
END LIBRARY

