* NGSPICE file created from outel8227.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

.subckt outel8227 VGND VPWR clk cs dataBusIn[0] dataBusIn[1] dataBusIn[2] dataBusIn[3]
+ dataBusIn[4] dataBusIn[5] dataBusIn[6] dataBusIn[7] dataBusOut[0] dataBusOut[1]
+ dataBusOut[2] dataBusOut[3] dataBusOut[4] dataBusOut[5] dataBusOut[6] dataBusOut[7]
+ dataBusSelect gpio[0] gpio[10] gpio[11] gpio[12] gpio[13] gpio[14] gpio[15] gpio[16]
+ gpio[17] gpio[18] gpio[19] gpio[1] gpio[20] gpio[21] gpio[22] gpio[23] gpio[24]
+ gpio[25] gpio[2] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7] gpio[8] gpio[9] nrst
X_2037_ _1297_ _1302_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__and2_1
XFILLER_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2106_ _1147_ _0145_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__nor2_1
XFILLER_52_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2724_ clknet_4_15_0_clk _0012_ net130 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1606_ net43 _0848_ _0888_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor3_1
X_2655_ _0283_ _0297_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__a21o_1
XFILLER_59_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2586_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0404_ VGND VGND
+ VPWR VPWR _0563_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_57_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1537_ net61 _0835_ net39 net43 VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a211oi_4
Xfanout127 net131 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_2
Xfanout105 net107 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xfanout116 net119 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
X_1468_ _0657_ _0673_ net67 VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__and3_1
X_1399_ _0674_ net69 VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__nor2_4
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2440_ _0440_ _0442_ _0439_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__a21bo_1
X_2371_ _0379_ _0387_ _0378_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__o21a_1
XFILLER_49_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_2569_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] _0403_ _0547_
+ net37 VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__o2bb2a_1
X_2707_ net162 _1265_ _0651_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_1
X_2638_ _0291_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nand2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1940_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] _1211_ _1212_
+ top8227.internalDataflow.accRegToDB\[7\] VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__a22o_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ net60 _0779_ _0818_ _1139_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_16_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2423_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _0438_ _0404_
+ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2354_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] net20 VGND VGND
+ VPWR VPWR _0371_ sky130_fd_sc_hd__nor2_1
XFILLER_49_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2285_ _0323_ top8227.PSRCurrentValue\[1\] _0316_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__and3b_1
XFILLER_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2070_ _1340_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__or2_2
XFILLER_61_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1854_ _1122_ _1125_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__nor3_4
X_1785_ _1056_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__or2_1
X_1923_ net105 _0691_ net67 VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__and3_1
X_2406_ _1313_ _0422_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__nor2_1
X_2337_ _1298_ _0353_ _0739_ _1069_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o211a_1
XFILLER_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2199_ _0238_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__inv_2
X_2268_ _0133_ _0272_ _0302_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__nor3_1
XFILLER_52_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold41 top8227.internalDataflow.addressLowBusModule.busInputs\[39\] VGND VGND VPWR
+ VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 top8227.internalDataflow.accRegToDB\[1\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold30 top8227.internalDataflow.stackBusModule.busInputs\[37\] VGND VGND VPWR VPWR
+ net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_5 _0215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1570_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__inv_2
X_2053_ _1210_ _1325_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__nand2_1
X_2122_ top8227.internalDataflow.stackBusModule.busInputs\[35\] _1204_ _1207_ _0160_
+ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a2111o_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1837_ net94 top8227.demux.state_machine.currentAddress\[12\] _0823_ VGND VGND VPWR
+ VPWR _1110_ sky130_fd_sc_hd__and3_1
X_1906_ net102 _0677_ net55 net93 _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__a221o_1
X_1768_ _1037_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__or2_1
X_1699_ net45 _0897_ _0921_ net33 _0719_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__a32o_1
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1622_ net5 _0850_ _0862_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__and3_2
X_2740_ clknet_4_10_0_clk _0024_ net121 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2671_ _0133_ _0272_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__o21a_1
X_1553_ net133 _0845_ net4 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__or3b_1
X_1484_ net72 _0699_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__nor2_1
X_2036_ top8227.internalDataflow.addressLowBusModule.busInputs\[39\] net24 _1304_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _1306_ VGND VGND VPWR
+ VPWR _1309_ sky130_fd_sc_hd__a221o_1
X_2105_ _0141_ _0144_ _1151_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__o21a_1
XFILLER_39_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2723_ clknet_4_15_0_clk _0011_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2585_ _0392_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__and2b_1
X_1605_ _0848_ _0880_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nor2_4
X_1536_ gpio[19] net61 top8227.pulse_slower.nextEnableState\[0\] VGND VGND VPWR VPWR
+ _0836_ sky130_fd_sc_hd__and3_1
XFILLER_8_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2654_ _0180_ _0610_ _0585_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux2_1
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout128 net130 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
Xfanout117 net118 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_4
Xfanout106 net107 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dlymetal6s2s_1
X_1398_ _0676_ _0699_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nor2_2
X_1467_ _0679_ _0718_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nor2_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2019_ _1077_ _1290_ _1291_ _1246_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__and4bb_1
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2370_ _0380_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and2_1
XFILLER_64_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2706_ net164 _1330_ _0651_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
X_2499_ _0507_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2568_ _0375_ _0376_ _0388_ _0400_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__o31ai_1
X_1519_ top8227.instructionLoader.interruptInjector.resetDetected gpio[21] VGND VGND
+ VPWR VPWR _0819_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2637_ _0283_ _0299_ _0594_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ _0701_ _0711_ _0774_ _0792_ net98 VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__o41a_1
X_2422_ _0433_ _0437_ _0396_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux2_1
X_2353_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] net20 VGND VGND
+ VPWR VPWR _0370_ sky130_fd_sc_hd__and2_1
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2284_ _0790_ _1143_ _1176_ _0322_ net50 VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__o41a_1
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1999_ _1072_ _1271_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__or2_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1922_ net106 _0770_ net60 VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__a21o_1
X_1853_ net41 _1109_ _1119_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__nor3_4
X_1784_ net113 _0739_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__and2_1
X_2405_ _1336_ _0128_ _0420_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__or4_1
X_2336_ _0746_ _0747_ _0749_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a21o_1
XFILLER_6_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2198_ _1152_ _0227_ _0232_ _1148_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__o2bb2a_1
X_2267_ _1344_ _0304_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__xnor2_2
Xhold42 top8227.internalDataflow.addressLowBusModule.busInputs\[35\] VGND VGND VPWR
+ VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 top8227.internalDataflow.stackBusModule.busInputs\[42\] VGND VGND VPWR VPWR
+ net153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 top8227.internalDataflow.stackBusModule.busInputs\[38\] VGND VGND VPWR VPWR
+ net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 top8227.internalDataflow.addressLowBusModule.busInputs\[24\] VGND VGND VPWR
+ VPWR net186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 _0701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ top8227.internalDataflow.stackBusModule.busInputs\[38\] _1204_ _1207_ _1324_
+ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a211o_1
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2121_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\] _1214_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[43\] VGND VGND VPWR VPWR _0161_
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1905_ top8227.demux.state_machine.timeState\[1\] net71 _0691_ VGND VGND VPWR VPWR
+ _1178_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1836_ net58 _1092_ _1097_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a22o_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1698_ net74 net65 net29 _0878_ _0967_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__a32o_1
X_1767_ _0679_ _0710_ _0716_ _0690_ _0656_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__a311oi_4
X_2319_ top8227.PSRCurrentValue\[2\] top8227.demux.setInterruptFlag top8227.instructionLoader.interruptInjector.irqGenerated
+ top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ VGND
+ VGND VPWR VPWR _0345_ sky130_fd_sc_hd__or4b_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR dataBusOut[0] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1552_ net3 net54 VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__nand2_1
X_1621_ net5 _0862_ _0899_ _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__a31o_1
X_2670_ _0133_ _0272_ _0282_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__a21oi_1
X_2104_ net133 _1130_ _1131_ _0143_ _0140_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__a221o_1
X_1483_ net69 _0716_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nor2_2
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2035_ _1261_ _1307_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__nor2_2
X_2799_ clknet_4_15_0_clk _0075_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_1819_ net100 net57 _0693_ net102 _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__a221o_1
XFILLER_60_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2722_ clknet_4_14_0_clk _0010_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_2584_ _0366_ _0367_ _0391_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or3_1
X_1604_ top8227.demux.state_machine.currentAddress\[1\] net36 _0875_ net26 VGND VGND
+ VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
Xfanout129 net130 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_4
X_1535_ _0834_ _0832_ _0827_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__or3b_2
Xfanout107 net108 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout118 net119 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
X_2653_ _0268_ _0587_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_57_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1466_ _0674_ _0718_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__nor2_1
X_1397_ net88 net82 net85 net91 VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__or4b_4
X_2018_ net110 _0696_ top8227.demux.state_machine.currentAddress\[12\] VGND VGND VPWR
+ VPWR _1291_ sky130_fd_sc_hd__or3b_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2705_ net163 _0122_ _0651_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
X_2636_ _0263_ _0581_ _0585_ _0224_ _0282_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__o221a_1
X_2498_ _0497_ _0498_ _0496_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
X_2567_ _0415_ _0545_ _0546_ _0416_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o31a_1
X_1449_ top8227.branchBackward top8227.branchForward VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__or2_1
X_1518_ _0752_ _0817_ net52 VGND VGND VPWR VPWR gpio[21] sky130_fd_sc_hd__o21a_4
XFILLER_55_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2421_ _0435_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__xnor2_1
X_2352_ _0367_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__nor2_1
X_2283_ net108 _0765_ _1177_ _0320_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a211o_1
XFILLER_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1998_ _0707_ _0796_ net109 VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__o21a_1
X_2619_ _1270_ _0577_ _0578_ _1269_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__o31a_1
XFILLER_28_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1852_ _1109_ _1124_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__and2_1
X_1921_ net48 _1188_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__a21o_1
X_1783_ net98 net95 net70 _0691_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__o211a_1
X_2404_ _0153_ _0176_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__or2_1
X_2335_ _0764_ _0821_ _1227_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a21oi_1
X_2266_ _0296_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__xnor2_1
X_2197_ _1154_ _0236_ _0228_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o21bai_4
XFILLER_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold43 top8227.internalDataflow.addressLowBusModule.busInputs\[36\] VGND VGND VPWR
+ VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 top8227.internalDataflow.stackBusModule.busInputs\[35\] VGND VGND VPWR VPWR
+ net154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold32 top8227.internalDataflow.stackBusModule.busInputs\[33\] VGND VGND VPWR VPWR
+ net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 net14 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_60_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2120_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] _1211_ _1212_
+ top8227.internalDataflow.accRegToDB\[3\] VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] _1214_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[46\] _1323_ VGND VGND VPWR VPWR
+ _1324_ sky130_fd_sc_hd__a221o_1
XFILLER_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1904_ _0754_ _0770_ _0775_ _1042_ net96 VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__o41a_1
X_1835_ _1087_ _1104_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__or3_1
XFILLER_22_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1766_ net112 net71 _0709_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__and3_1
X_1697_ _0964_ _0976_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__or2_1
XFILLER_57_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2318_ top8227.demux.nmi _0328_ _0344_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21oi_1
X_2249_ top8227.PSRCurrentValue\[3\] _0283_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__nand2_1
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput11 net11 VGND VGND VPWR VPWR dataBusOut[1] sky130_fd_sc_hd__buf_2
XFILLER_56_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1551_ net8 _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__nor2_1
X_1620_ _0691_ net68 net32 VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__and3_1
X_1482_ _0658_ net69 _0699_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__nor3_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2103_ net103 _0687_ _0142_ _1258_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__a31o_1
X_2034_ net24 _1305_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or2_1
X_2798_ clknet_4_6_0_clk _0074_ net125 VGND VGND VPWR VPWR gpio[15] sky130_fd_sc_hd__dfrtp_4
X_1818_ net113 _0677_ _0687_ net102 VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a22o_1
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1749_ _0979_ _0993_ _0999_ _1011_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__or4_1
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2721_ clknet_4_14_0_clk _0009_ net131 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_2652_ _0791_ _0269_ _0286_ _0608_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a31o_1
X_2583_ net38 _0556_ _0557_ _0560_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a31o_1
X_1603_ net161 net35 _0889_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21bo_1
X_1534_ net94 _0823_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__and3_1
Xfanout108 net109 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
Xfanout119 net9 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__buf_2
X_1465_ _0676_ _0716_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nor2_1
X_1396_ top8227.demux.reset _0696_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__or2_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2017_ _0656_ top8227.demux.state_machine.currentAddress\[1\] _0695_ _0831_ VGND
+ VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a31o_1
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2704_ net168 _0147_ _0651_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
X_2635_ _0262_ _0587_ _0293_ _0193_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o2bb2a_1
X_2566_ _0421_ _0540_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__nor2_1
X_2497_ _1155_ net19 _0506_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__o21ai_2
X_1448_ top8227.branchBackward top8227.branchForward VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__nor2_1
X_1517_ _0705_ net63 net96 net70 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__o211a_1
XFILLER_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1379_ _0657_ net98 _0673_ net76 VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and4_1
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2420_ _0418_ _0424_ _0410_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout90 top8227.demux.state_machine.currentInstruction\[1\] VGND VGND VPWR VPWR
+ net90 sky130_fd_sc_hd__clkbuf_2
X_2351_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] net20 VGND VGND
+ VPWR VPWR _0368_ sky130_fd_sc_hd__nor2_1
X_2282_ _1140_ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or2_1
XFILLER_64_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1997_ _1051_ _1053_ _1073_ _1190_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__or4_2
X_2549_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0384_ _0400_
+ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__o21a_1
X_2618_ _1063_ _1114_ _0276_ _0281_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__or4_2
XFILLER_28_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ net42 _1117_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__nor2_1
X_1920_ gpio[19] _0726_ _1192_ net58 top8227.pulse_slower.nextEnableState\[0\] VGND
+ VGND VPWR VPWR _1193_ sky130_fd_sc_hd__o2111a_1
X_2403_ _0199_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__or2_1
X_1782_ _1044_ _1051_ _1054_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__or3_1
X_2334_ net110 top8227.demux.state_machine.currentAddress\[7\] _0350_ VGND VGND VPWR
+ VPWR _0351_ sky130_fd_sc_hd__a21o_1
X_2196_ _1162_ _0232_ _0235_ _1161_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__o22a_1
X_2265_ _1344_ _0304_ _1340_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a21o_1
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold22 top8227.negEdgeDetector.q1 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 top8227.demux.state_machine.currentAddress\[10\] VGND VGND VPWR VPWR net166
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 top8227.internalDataflow.addressLowBusModule.busInputs\[38\] VGND VGND VPWR
+ VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2050_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] _1211_ _1212_
+ top8227.internalDataflow.accRegToDB\[6\] VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__a22o_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1903_ _0818_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__or2_1
X_1834_ _1045_ _1101_ _1105_ _1106_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__or4_1
X_1765_ net107 _0784_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__and2_1
X_1696_ _0927_ _0972_ _0973_ _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__or4_1
X_2179_ _1148_ _0209_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__nor2_1
X_2317_ _0665_ net144 top8227.demux.nmi VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a21oi_1
X_2248_ _1171_ _0286_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__nand2_1
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput12 net12 VGND VGND VPWR VPWR dataBusOut[2] sky130_fd_sc_hd__buf_2
XFILLER_0_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1550_ net7 net54 VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nand2_2
X_1481_ net69 _0699_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nor2_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2033_ net24 _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__nor2_2
X_2102_ top8227.demux.reset top8227.demux.nmi top8227.demux.setInterruptFlag VGND
+ VGND VPWR VPWR _0142_ sky130_fd_sc_hd__nor3_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2797_ clknet_4_6_0_clk _0073_ net125 VGND VGND VPWR VPWR gpio[14] sky130_fd_sc_hd__dfrtp_4
X_1817_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__inv_2
X_1748_ _1021_ _1022_ _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__or3_1
X_1679_ net57 net30 _0884_ _0919_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_43_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2582_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _0403_ _0558_
+ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a22o_1
X_1602_ _0847_ _0871_ _0888_ _0819_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__a211o_1
X_2720_ clknet_4_14_0_clk _0008_ net131 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2651_ _0148_ _0293_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__nor2_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1533_ top8227.demux.state_machine.currentAddress\[12\] top8227.demux.state_machine.currentAddress\[6\]
+ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__or2_1
X_1395_ net93 _0695_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__or2_1
Xfanout109 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
X_1464_ _0762_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__or2_1
X_2016_ _1138_ _1287_ _1288_ _1181_ _1115_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__a2111o_1
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2565_ _0176_ _0540_ _0155_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o21a_1
X_2703_ net154 _0171_ _0651_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
X_1516_ _0799_ _0812_ _0814_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__or4_1
X_2634_ _0290_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
X_2496_ _1263_ net19 _0408_ _1218_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__o2bb2a_1
X_1447_ net100 _0746_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__and3_1
X_1378_ _0676_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__nor2_1
XFILLER_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout91 net92 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
Xfanout80 top8227.demux.state_machine.currentInstruction\[5\] VGND VGND VPWR VPWR
+ net80 sky130_fd_sc_hd__clkbuf_4
X_2350_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] net20 VGND VGND
+ VPWR VPWR _0367_ sky130_fd_sc_hd__and2_1
X_2281_ _0779_ _1086_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__or2_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1996_ net48 _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__and2_2
X_2548_ _0217_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__xor2_1
X_2617_ net107 _0292_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2_1
X_2479_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] net23 _0476_
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__a21o_1
XFILLER_55_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload0 clknet_4_0_0_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_21_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ _1109_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__and2_1
X_1781_ net60 _1038_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__or3_1
X_2402_ _0217_ _0245_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or2_1
X_2333_ net110 _0825_ _1069_ top8227.demux.state_machine.currentAddress\[6\] _0349_
+ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a221o_1
X_2195_ net1 _1254_ _1256_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__a221oi_2
XFILLER_37_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2264_ _0133_ _0272_ _0303_ _0131_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a211o_1
XFILLER_52_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1979_ net61 _1060_ _1067_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__or4_1
Xhold45 top8227.demux.state_machine.currentAddress\[3\] VGND VGND VPWR VPWR net178
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 top8227.internalDataflow.stackBusModule.busInputs\[43\] VGND VGND VPWR VPWR
+ net156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold34 top8227.internalDataflow.stackBusModule.busInputs\[34\] VGND VGND VPWR VPWR
+ net167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0032_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _0702_ _0735_ net96 net70 VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__o211a_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1833_ net108 _0708_ net60 VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__a21o_1
X_1764_ _0699_ _0710_ _0656_ net72 VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__a211oi_2
X_2316_ _0328_ _0343_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__nor2_1
X_1695_ _0785_ net27 _0855_ net26 _0974_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__a221o_1
X_2178_ _1281_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__nor2_1
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2247_ net108 net50 VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__nand2_1
XFILLER_31_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR dataBusOut[3] sky130_fd_sc_hd__buf_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1480_ net97 net76 _0760_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__and3_1
X_2101_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[4\] _1127_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__a221o_1
X_2032_ _1296_ _1301_ _1286_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2796_ clknet_4_6_0_clk _0072_ net125 VGND VGND VPWR VPWR gpio[13] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1816_ net51 _1088_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__nand2_2
X_1678_ _0806_ net30 _0856_ _0884_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__a22o_1
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1747_ _0974_ _0989_ _1001_ _1004_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2581_ _0391_ _0401_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__nor2_1
X_1601_ _0667_ _0857_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nand2_2
X_1532_ _0829_ _0831_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__or2_1
X_2650_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] _0607_ _0579_
+ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_1
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1394_ net103 net100 net94 VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__nor3_1
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1463_ net70 _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__and2_2
XFILLER_35_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2015_ top8227.demux.state_machine.timeState\[5\] _0695_ net57 VGND VGND VPWR VPWR
+ _1288_ sky130_fd_sc_hd__o21a_1
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2779_ clknet_4_4_0_clk _0055_ net123 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2702_ net167 _0192_ _0651_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
X_2495_ net37 _0503_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__and3_1
X_2564_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _0404_ _0542_
+ net37 _0544_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__o221a_1
X_2633_ _0299_ _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__xnor2_1
X_1515_ net99 _0769_ _0772_ _0807_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__a2111o_1
X_1446_ top8227.PSRCurrentValue\[6\] _0732_ _0740_ _0741_ _0743_ VGND VGND VPWR VPWR
+ _0747_ sky130_fd_sc_hd__o2111a_1
X_1377_ net88 net91 net82 net85 VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__or4b_4
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout92 top8227.demux.state_machine.currentInstruction\[0\] VGND VGND VPWR VPWR
+ net92 sky130_fd_sc_hd__buf_2
Xfanout81 top8227.demux.state_machine.currentInstruction\[4\] VGND VGND VPWR VPWR
+ net81 sky130_fd_sc_hd__buf_2
Xfanout70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_24_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2280_ _1046_ _0313_ _0317_ _0239_ _0319_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2616_ gpio[7] _0575_ _1314_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a21o_1
X_1995_ top8227.demux.state_machine.currentAddress\[12\] _0824_ _1078_ top8227.demux.state_machine.currentAddress\[6\]
+ _1096_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__a221o_1
X_2478_ _0487_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__nor2_1
X_2547_ _0245_ _0412_ net23 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux2_1
X_1429_ _0659_ gpio[22] _0672_ net61 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__a211o_1
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload1 clknet_4_1_0_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_4
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1780_ net107 _0791_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__a21o_1
X_2401_ _1314_ _1335_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or3_1
X_2332_ net101 top8227.demux.state_machine.currentAddress\[7\] net71 _0731_ VGND VGND
+ VPWR VPWR _0349_ sky130_fd_sc_hd__and4_1
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2194_ _1254_ _1256_ _0233_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__nor3_1
X_2263_ _0133_ _0159_ _0297_ _0300_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and4_1
XFILLER_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1978_ net93 _0806_ _1250_ top8227.demux.state_machine.timeState\[1\] _1249_ VGND
+ VGND VPWR VPWR _1251_ sky130_fd_sc_hd__a221o_1
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold46 top8227.internalDataflow.addressLowBusModule.busInputs\[34\] VGND VGND VPWR
+ VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 top8227.internalDataflow.stackBusModule.busInputs\[41\] VGND VGND VPWR VPWR
+ net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 top8227.internalDataflow.stackBusModule.busInputs\[47\] VGND VGND VPWR VPWR
+ net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold35 top8227.internalDataflow.stackBusModule.busInputs\[36\] VGND VGND VPWR VPWR
+ net168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ net41 _1173_ _1170_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__o21ai_4
XFILLER_34_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1832_ _1062_ _1098_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__or2_1
X_1763_ top8227.pulse_slower.currentEnableState\[1\] net137 VGND VGND VPWR VPWR top8227.pulse_slower.nextEnableState\[1\]
+ sky130_fd_sc_hd__and2b_1
X_1694_ _0782_ net27 _0902_ _0914_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__a22o_1
X_2315_ net42 _0842_ top8227.demux.setInterruptFlag VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_27_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2246_ _0656_ net41 VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nor2_4
X_2177_ top8227.demux.reset _0198_ _0216_ _1308_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a211o_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput14 net14 VGND VGND VPWR VPWR dataBusOut[4] sky130_fd_sc_hd__buf_2
X_2100_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] _1109_ _1122_
+ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__and3_1
X_2031_ _1286_ _1296_ _1300_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__and3b_2
X_2795_ clknet_4_7_0_clk _0071_ net125 VGND VGND VPWR VPWR gpio[12] sky130_fd_sc_hd__dfrtp_4
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ net105 _0712_ _1086_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__a211o_1
X_1746_ _0909_ _0915_ _0957_ _0970_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__or4_1
X_1677_ _0770_ net30 _0912_ _0932_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__a22o_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2229_ _0180_ _0268_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__and2b_1
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2580_ _0369_ _0370_ _0390_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__or3_1
X_1600_ _0881_ net26 _0887_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a21o_1
X_1531_ top8227.demux.state_machine.currentAddress\[7\] _0830_ _0828_ VGND VGND VPWR
+ VPWR _0831_ sky130_fd_sc_hd__o21a_1
XFILLER_8_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1462_ net92 net83 net86 net89 VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__and4b_1
X_1393_ net102 net100 VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or2_2
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2014_ top8227.demux.state_machine.timeState\[1\] net56 _0697_ VGND VGND VPWR VPWR
+ _1287_ sky130_fd_sc_hd__a21o_1
X_2778_ clknet_4_7_0_clk _0054_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1729_ _0732_ _0839_ _0879_ _0944_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__o22a_1
XFILLER_58_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2701_ net165 _0212_ _0651_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
X_2632_ _0270_ _0301_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__or2_1
X_2494_ _0487_ _0491_ _0502_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__o21ai_1
X_2563_ _0388_ _0543_ _0400_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__o21ai_1
X_1445_ top8227.PSRCurrentValue\[6\] _0733_ _0742_ _0744_ _0745_ VGND VGND VPWR VPWR
+ _0746_ sky130_fd_sc_hd__a2111oi_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1514_ top8227.demux.state_machine.timeState\[5\] net55 _0779_ _0780_ _0795_ VGND
+ VGND VPWR VPWR _0815_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_2_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376_ net89 top8227.demux.state_machine.currentInstruction\[0\] net84 net87 VGND
+ VGND VPWR VPWR _0678_ sky130_fd_sc_hd__nor4b_2
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout93 net95 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
Xfanout60 _0670_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout82 net83 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout71 _0689_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
XFILLER_64_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1994_ _1148_ _1218_ _1153_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__o21ai_2
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2615_ _1335_ gpio[6] _0575_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_1
X_2477_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] net23 VGND VGND
+ VPWR VPWR _0488_ sky130_fd_sc_hd__nor2_1
X_2546_ _0399_ _0529_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__xnor2_1
X_1428_ gpio[19] _0726_ top8227.pulse_slower.nextEnableState\[0\] net58 VGND VGND
+ VPWR VPWR _0729_ sky130_fd_sc_hd__o211a_1
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1359_ net8 VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__inv_2
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload2 clknet_4_2_0_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_21_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2400_ _0127_ _0416_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2331_ net140 _1267_ _0348_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_1
X_2262_ _0159_ _0297_ _0300_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__and3_1
XFILLER_52_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2193_ _0730_ _1260_ _1261_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__o21ba_1
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1977_ _0693_ net55 VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__or2_1
X_2529_ _0693_ _1228_ _0519_ _0684_ _1056_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__a221oi_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold47 top8227.demux.state_machine.currentAddress\[0\] VGND VGND VPWR VPWR net180
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 top8227.internalDataflow.addressLowBusModule.busInputs\[33\] VGND VGND VPWR
+ VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 top8227.internalDataflow.stackBusModule.busInputs\[45\] VGND VGND VPWR VPWR
+ net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold14 net11 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1900_ _1099_ _1100_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__nor3_1
X_1831_ _1041_ _1100_ _1102_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__or4_1
X_1762_ _0938_ _0947_ _1028_ _1036_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__or4_1
X_1693_ _0700_ net31 _0924_ _0943_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a22o_1
X_2176_ _1306_ _0214_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__nor3_1
X_2314_ gpio[20] net155 net44 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
X_2245_ _0275_ _0282_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__nor3_1
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR dataBusOut[5] sky130_fd_sc_hd__buf_2
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ _1294_ _1301_ _1286_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__and3b_1
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2794_ clknet_4_6_0_clk _0070_ net125 VGND VGND VPWR VPWR gpio[11] sky130_fd_sc_hd__dfrtp_4
X_1745_ _0925_ _0930_ _0969_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__or4_1
X_1814_ _0700_ _0739_ _0765_ net105 VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__o31a_1
X_1676_ _0861_ _0876_ _0952_ _0955_ _0947_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__a311o_1
X_2159_ _1261_ _0198_ _0197_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a21oi_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2228_ _0179_ _0172_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__nand2b_1
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1530_ top8227.demux.state_machine.currentAddress\[3\] top8227.demux.state_machine.currentAddress\[11\]
+ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__or2_1
X_1461_ net76 _0721_ _0760_ net70 VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a22o_1
X_1392_ _0688_ net70 _0691_ net73 net75 VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__a32o_1
X_2013_ _1067_ _1118_ _1178_ _1258_ net51 VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__o41a_2
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2777_ clknet_4_5_0_clk _0053_ net124 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1728_ _1002_ _1004_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__or2_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1659_ _0849_ _0888_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2562_ _0378_ _0379_ _0387_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__nor3_1
X_2700_ net142 _0237_ _0651_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_1
X_2631_ net186 _0590_ _0579_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
X_2493_ _0487_ _0491_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or3_1
X_1444_ top8227.PSRCurrentValue\[1\] net73 net65 VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__and3_1
X_1513_ _0724_ _0759_ _0765_ _0813_ net97 VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__o41a_1
X_1375_ _0674_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__nor2_2
X_2829_ clknet_4_0_0_clk _0105_ net119 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout61 _0670_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
Xfanout94 net95 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout50 net52 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
Xfanout72 _0686_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
Xfanout83 net84 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_64_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ net25 _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__and2_1
XFILLER_20_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2545_ _0662_ _0245_ net38 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux2_1
X_2614_ gpio[5] _0575_ _0127_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__a21o_1
X_2476_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] net23 VGND VGND
+ VPWR VPWR _0487_ sky130_fd_sc_hd__and2_1
X_1427_ _0659_ gpio[22] _0672_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__a21o_1
X_1358_ top8227.internalDataflow.stackBusModule.busInputs\[34\] VGND VGND VPWR VPWR
+ _0663_ sky130_fd_sc_hd__inv_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_4_3_0_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_21_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2192_ _1207_ _0229_ _0230_ _0231_ _1210_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__o41ai_2
X_2330_ net141 _1332_ _0348_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_1
X_2261_ _0297_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1976_ top8227.demux.state_machine.timeState\[5\] net75 net73 VGND VGND VPWR VPWR
+ _1249_ sky130_fd_sc_hd__and3_1
X_2528_ net112 _1228_ net55 VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2459_ _0446_ _0448_ _0458_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__nand3_1
Xhold26 top8227.internalDataflow.stackBusModule.busInputs\[40\] VGND VGND VPWR VPWR
+ net159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold37 top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning VGND
+ VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net10 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 top8227.instructionLoader.interruptInjector.irqGenerated VGND VGND VPWR VPWR
+ net181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1761_ _0908_ _1034_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__or3_1
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1830_ top8227.demux.state_machine.timeState\[1\] net57 _0704_ net107 _1049_ VGND
+ VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a221o_1
X_1692_ _0966_ _0969_ _0970_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__or4_1
X_2313_ top8227.demux.nmi net44 _0342_ _0328_ net170 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_48_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2175_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\] _1297_ _1302_
+ net24 top8227.internalDataflow.addressLowBusModule.busInputs\[33\] VGND VGND VPWR
+ VPWR _0215_ sky130_fd_sc_hd__a32o_1
X_2244_ _1266_ _1315_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__nor2_1
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1959_ net79 _0688_ _0702_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__and3_1
Xoutput16 net16 VGND VGND VPWR VPWR dataBusOut[6] sky130_fd_sc_hd__buf_2
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2793_ clknet_4_7_0_clk _0069_ net126 VGND VGND VPWR VPWR gpio[10] sky130_fd_sc_hd__dfrtp_4
X_1744_ _0902_ _0945_ _1018_ _1019_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__a211o_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1813_ net104 net77 net65 VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__and3_1
X_1675_ _0689_ _0709_ net33 _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2158_ top8227.demux.nmi _1307_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__nor2_1
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2089_ _1283_ _1276_ _0124_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2227_ _0264_ _0266_ _0201_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1391_ net69 _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__nor2_2
X_1460_ _0676_ _0722_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ _1283_ _1276_ _1267_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__mux2_1
X_2776_ clknet_4_6_0_clk _0052_ net124 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_1658_ _0796_ net32 _0906_ _0912_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__a221o_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1727_ _0678_ net74 net29 _0878_ _0897_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_56_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1589_ net39 _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__and2_2
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2492_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] net23 VGND VGND
+ VPWR VPWR _0502_ sky130_fd_sc_hd__xor2_1
X_2561_ _0176_ _0541_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2630_ _0260_ _0283_ _0589_ _0588_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__a31o_1
X_1512_ _0766_ _0784_ _0787_ _0789_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__or4_1
X_1443_ top8227.PSRCurrentValue\[7\] net73 _0705_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__and3_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1374_ net81 net80 VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__nand2b_4
XFILLER_63_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2828_ clknet_4_0_0_clk _0104_ net119 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2759_ clknet_4_3_0_clk _0035_ net114 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_46_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout40 _0820_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
Xfanout62 _0821_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xfanout51 net52 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
Xfanout73 net74 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout95 top8227.demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
Xfanout84 top8227.demux.state_machine.currentInstruction\[3\] VGND VGND VPWR VPWR
+ net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1992_ _1154_ _1264_ _1155_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__o21ai_4
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload10 clknet_4_11_0_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_8
X_2475_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _0403_ _0480_
+ _0400_ _0486_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__a221o_1
X_2544_ _0507_ gpio[15] _0528_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
X_2613_ _0154_ gpio[4] _0575_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_1
X_1357_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] VGND VGND VPWR
+ VPWR _0662_ sky130_fd_sc_hd__inv_2
X_1426_ _0659_ gpio[22] _0672_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload4 clknet_4_5_0_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_21_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2191_ top8227.internalDataflow.stackBusModule.busInputs\[32\] _1204_ VGND VGND VPWR
+ VPWR _0231_ sky130_fd_sc_hd__and2_1
X_2260_ _0298_ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
XFILLER_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1975_ top8227.demux.state_machine.currentAddress\[7\] _0828_ _1110_ _1247_ VGND
+ VGND VPWR VPWR _1248_ sky130_fd_sc_hd__a211o_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2458_ _0446_ _0447_ _0458_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__or3_1
Xhold38 top8227.internalDataflow.addressLowBusModule.busInputs\[32\] VGND VGND VPWR
+ VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 top8227.internalDataflow.stackBusModule.busInputs\[46\] VGND VGND VPWR VPWR
+ net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 top8227.internalDataflow.stackBusModule.busInputs\[44\] VGND VGND VPWR VPWR
+ net160 sky130_fd_sc_hd__dlygate4sd3_1
X_2527_ _1068_ _1228_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or2_1
X_1409_ net72 _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nor2_2
X_2389_ net19 VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__inv_2
Xhold49 _0033_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1691_ _0685_ _0702_ net31 _0877_ _0932_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__a32o_1
X_1760_ _0920_ _0966_ _0973_ _1012_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__or4_1
X_2312_ top8227.PSRCurrentValue\[2\] top8227.demux.setInterruptFlag top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
+ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_48_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _1304_ _1311_
+ net2 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_1
XFILLER_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2243_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1889_ _1154_ _1156_ _1160_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a21o_1
X_1958_ _0806_ _1228_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__a21boi_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput17 net17 VGND VGND VPWR VPWR dataBusOut[7] sky130_fd_sc_hd__buf_2
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ clknet_4_6_0_clk _0068_ net125 VGND VGND VPWR VPWR gpio[9] sky130_fd_sc_hd__dfrtp_4
X_1674_ _0948_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nor2_1
X_1743_ net47 net26 _0897_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__and3_1
X_1812_ net49 _1064_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__and3_1
X_2226_ _0201_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
X_2088_ _0127_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
X_2157_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] _1310_ _1311_
+ net3 _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__a221o_1
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ net88 net91 net82 net85 VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__nand4b_2
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ net41 _1282_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__or2_1
X_2844_ clknet_4_0_0_clk VGND VGND VPWR VPWR gpio[23] sky130_fd_sc_hd__buf_2
X_1588_ net53 _0874_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__nor2_1
X_1726_ _0839_ _0844_ _0851_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__a31o_1
X_2775_ clknet_4_4_0_clk _0051_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_1657_ net68 net64 net32 _0936_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_56_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2209_ net25 _0237_ _0240_ _1281_ _0247_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a221oi_4
XTAP_TAPCELL_ROW_64_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2491_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _0501_ _0404_
+ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux2_1
X_2560_ _0414_ _0540_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nand2_1
X_1442_ top8227.PSRCurrentValue\[1\] net72 _0703_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__or3_1
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1511_ _0802_ _0809_ _0810_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__or4_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1373_ net81 net80 VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__and2b_1
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2758_ clknet_4_3_0_clk _0034_ net115 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
X_2827_ clknet_4_0_0_clk _0103_ net118 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2689_ _0622_ _0640_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__o21ai_1
X_1709_ _0800_ net27 _0902_ _0980_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_18_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_54_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout41 _0730_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_4
Xfanout52 _0729_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout85 net86 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xfanout63 _0755_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_2
Xfanout96 net99 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_2
Xfanout74 _0685_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_63_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload11 clknet_4_12_0_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_6
X_2612_ _0177_ gpio[3] _0575_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
X_1991_ _1160_ _1263_ _1218_ _1162_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2543_ _0496_ gpio[14] _0528_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
X_2474_ net37 _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__nor2_1
X_1425_ _0726_ VGND VGND VPWR VPWR gpio[22] sky130_fd_sc_hd__clkinv_4
X_1356_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] VGND VGND VPWR
+ VPWR _0661_ sky130_fd_sc_hd__inv_2
XFILLER_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload5 clknet_4_6_0_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2190_ top8227.internalDataflow.addressLowBusModule.busInputs\[32\] _1211_ _1212_
+ top8227.internalDataflow.accRegToDB\[0\] VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a22o_1
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ net61 _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__nand2_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold28 top8227.demux.state_machine.currentAddress\[5\] VGND VGND VPWR VPWR net161
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2457_ _0145_ _0444_ _0469_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__a21o_1
Xhold39 top8227.internalDataflow.addressLowBusModule.busInputs\[37\] VGND VGND VPWR
+ VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
X_2526_ net101 _0796_ _1230_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__a21boi_1
X_2388_ net42 _1157_ _1159_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or3_1
Xhold17 top8227.freeCarry VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ net82 net85 net88 net91 VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__or4bb_4
XTAP_TAPCELL_ROW_26_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1690_ _0702_ net68 net30 _0890_ _0919_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__a32o_1
X_2311_ top8227.instructionLoader.interruptInjector.resetDetected net43 VGND VGND
+ VPWR VPWR _0028_ sky130_fd_sc_hd__and2_1
X_2242_ _0276_ _0279_ _0281_ _1269_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__o31ai_4
XTAP_TAPCELL_ROW_48_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2173_ _1085_ _0212_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__nand2_1
X_1957_ top8227.demux.state_machine.timeState\[3\] net57 _1229_ VGND VGND VPWR VPWR
+ _1230_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1888_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__inv_2
X_2509_ net172 _0122_ _0512_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput18 net18 VGND VGND VPWR VPWR dataBusSelect sky130_fd_sc_hd__buf_2
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2791_ clknet_4_7_0_clk _0067_ net126 VGND VGND VPWR VPWR gpio[8] sky130_fd_sc_hd__dfrtp_4
X_1811_ _1076_ _1081_ _1082_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__o2bb2a_1
X_1673_ _0819_ _0843_ net53 _0888_ _0950_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__o41a_1
X_1742_ top8227.demux.state_machine.currentInstruction\[4\] _0721_ net32 _0937_ VGND
+ VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a31o_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2225_ _0193_ _0200_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__and2_1
XFILLER_53_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2156_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\] net24 _1304_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] VGND VGND VPWR VPWR
+ _0196_ sky130_fd_sc_hd__a22o_1
X_2087_ _1306_ _0126_ _1308_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__o21ba_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2010_ net41 _1282_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__nor2_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1725_ _0689_ _0731_ net33 VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__and3_1
X_2774_ clknet_4_4_0_clk _0050_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_2843_ clknet_4_2_0_clk _0117_ net116 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_1587_ _0819_ net53 VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nor2_1
X_1656_ net47 net40 _0890_ _0897_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_56_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2139_ _0177_ _0178_ _1281_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
X_2208_ _1280_ _0240_ _0246_ _0237_ net25 VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_64_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2490_ _0397_ _0500_ _0493_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__o21ai_1
X_1441_ top8227.PSRCurrentValue\[0\] _0678_ net73 VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__and3b_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1510_ _0774_ _0803_ _0804_ net97 VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__o31a_1
X_1372_ net90 net83 net86 net91 VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__or4bb_4
XFILLER_23_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1708_ net56 net31 _0884_ _0945_ _0986_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__a221o_1
X_2757_ clknet_4_2_0_clk top8227.instructionLoader.interruptInjector.nmiSync.in net115
+ VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 sky130_fd_sc_hd__dfrtp_1
X_2688_ _0291_ _0306_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__nor2_1
X_2826_ clknet_4_1_0_clk _0102_ net118 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1639_ _0819_ _0917_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nor2_2
XFILLER_64_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout20 net21 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
Xfanout53 _0849_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
Xfanout42 net44 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
Xfanout64 _0755_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_1
Xfanout31 _0838_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
Xfanout97 net99 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
Xfanout86 net87 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
Xfanout75 _0683_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_2
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1990_ net8 _1254_ _1256_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
+ _1262_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__a221o_1
X_2542_ _0482_ gpio[13] _0528_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
Xclkload12 clknet_4_13_0_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinv_4
XFILLER_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2611_ _1261_ _0198_ _0575_ gpio[2] _0197_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__a221o_1
X_2473_ _0482_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__xnor2_1
X_1355_ top8227.internalDataflow.stackBusModule.busInputs\[33\] VGND VGND VPWR VPWR
+ _0660_ sky130_fd_sc_hd__inv_2
X_1424_ _0714_ _0715_ _0723_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__a31oi_4
Xclkload6 clknet_4_7_0_clk VGND VGND VPWR VPWR clkload6/X sky130_fd_sc_hd__clkbuf_8
XFILLER_59_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2809_ clknet_4_6_0_clk _0085_ net124 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1973_ _1078_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__or2_1
X_2525_ _0697_ _0797_ _1223_ _1258_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__a211oi_1
X_2387_ net38 _0399_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or2_2
X_2456_ _0137_ _0408_ net19 _0138_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold29 top8227.internalDataflow.stackBusModule.busInputs\[39\] VGND VGND VPWR VPWR
+ net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 net12 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ net84 net87 net89 top8227.demux.state_machine.currentInstruction\[0\] VGND
+ VGND VPWR VPWR _0709_ sky130_fd_sc_hd__and4bb_2
XTAP_TAPCELL_ROW_26_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ _1154_ _0211_ _0205_ _1090_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a2bb2o_2
X_2310_ net150 _0313_ _0341_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_1
X_2241_ _1047_ _1058_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__or3_2
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1887_ _1088_ _1157_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__and3b_2
X_1956_ _0705_ net64 net79 _0688_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__o211a_1
XFILLER_33_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2508_ net176 _0147_ _0512_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
X_2439_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] net21 VGND VGND
+ VPWR VPWR _0453_ sky130_fd_sc_hd__xor2_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2790_ clknet_4_14_0_clk _0066_ net128 VGND VGND VPWR VPWR top8227.demux.reset sky130_fd_sc_hd__dfrtp_1
X_1810_ top8227.demux.state_machine.currentAddress\[12\] _0825_ _0830_ net113 VGND
+ VGND VPWR VPWR _1083_ sky130_fd_sc_hd__o31a_1
X_1741_ _0901_ _0935_ _0986_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__or3_1
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1672_ _0916_ _0951_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__nor2_1
XFILLER_53_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2155_ _1284_ _1277_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
X_2224_ _0261_ _0262_ _0223_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a21o_1
X_2086_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\] net24 _1310_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[29\] _0125_ VGND VGND VPWR
+ VPWR _0126_ sky130_fd_sc_hd__a221o_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1939_ _1194_ _1203_ _1174_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__and3b_2
XFILLER_44_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2773_ clknet_4_13_0_clk _0049_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_2842_ clknet_4_15_0_clk _0116_ net130 VGND VGND VPWR VPWR top8227.demux.isAddressing
+ sky130_fd_sc_hd__dfstp_1
X_1724_ _0775_ net29 net26 _0967_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a221o_1
X_1586_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__inv_2
X_1655_ _0689_ net64 net32 _0881_ _0899_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_64_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _1281_ _0245_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__nor2_1
X_2138_ _1283_ _1276_ _0173_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
X_2069_ _1331_ _1339_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__and2_1
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1440_ top8227.PSRCurrentValue\[7\] net72 _0736_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__or3_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1371_ net82 net85 VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__and2b_1
X_2825_ clknet_4_0_0_clk _0101_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1638_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__inv_2
X_1707_ _0793_ net31 _0912_ _0980_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__a221o_1
X_2756_ clknet_4_3_0_clk net135 net115 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ sky130_fd_sc_hd__dfrtp_1
X_2687_ _0631_ _0310_ _0598_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_58_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1569_ net4 net3 net133 net54 VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__o31a_2
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout21 _0362_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout54 _0842_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_4
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xfanout32 net33 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xfanout76 net78 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
Xfanout87 top8227.demux.state_machine.currentInstruction\[2\] VGND VGND VPWR VPWR
+ net87 sky130_fd_sc_hd__buf_2
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout65 _0734_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
Xfanout98 net99 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__buf_2
XFILLER_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2541_ _0470_ gpio[12] _0528_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
X_2472_ _0470_ _0471_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__o21bai_1
X_2610_ _0217_ _0576_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__nand2_1
Xclkload13 clknet_4_14_0_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_6
X_1354_ gpio[19] VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__inv_2
XFILLER_28_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1423_ _0656_ _0724_ net60 VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__a21o_1
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2808_ clknet_4_1_0_clk _0084_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload7 clknet_4_8_0_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_4
XFILLER_59_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2739_ clknet_4_10_0_clk _0023_ net121 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1972_ net101 net94 top8227.demux.state_machine.currentAddress\[6\] VGND VGND VPWR
+ VPWR _1245_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2455_ _0464_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__xor2_1
X_2524_ top8227.instructionLoader.interruptInjector.resetDetected net46 _0516_ top8227.demux.reset
+ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2386_ net38 _0399_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__nor2_2
Xhold19 net15 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
X_1406_ _0657_ net77 _0682_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__and3_1
XFILLER_61_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_334 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2171_ _1160_ _0210_ _0209_ _1162_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__o2bb2a_1
X_2240_ _1067_ _1070_ _1272_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1886_ _1112_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1955_ top8227.demux.state_machine.timeState\[1\] top8227.demux.state_machine.timeState\[5\]
+ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__or2_2
X_2438_ _0450_ _0451_ _0452_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__o21a_1
X_2507_ net175 _0171_ _0512_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
XFILLER_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2369_ _0662_ _0383_ _0382_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__o21ai_1
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1671_ _0844_ _0904_ _0948_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__or3_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ _0972_ _0987_ _1014_ _1016_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__or4_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2085_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _1304_ _1311_
+ net132 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
X_2154_ _0185_ _0191_ _1148_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_2
X_2223_ _0223_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__nand2b_1
XFILLER_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1938_ _1174_ _1193_ _1194_ _1203_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__o211a_2
X_1869_ _0704_ _1042_ net96 VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__o21a_1
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2841_ clknet_4_9_0_clk _0115_ net127 VGND VGND VPWR VPWR top8227.branchBackward
+ sky130_fd_sc_hd__dfrtp_1
X_2772_ clknet_4_13_0_clk _0048_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_1654_ _0930_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__or2_1
X_1723_ net67 net66 net27 _0856_ _0890_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a32o_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1585_ net4 net3 _0667_ _0842_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__or4b_1
X_2206_ _1280_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2137_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
X_2068_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__inv_2
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1370_ _0672_ VGND VGND VPWR VPWR top8227.pulse_slower.nextEnableState\[0\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ clknet_4_1_0_clk _0100_ net118 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1637_ net45 _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__nand2_1
X_1706_ net68 _0735_ net32 _0890_ _0906_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__a32o_1
X_2755_ clknet_4_2_0_clk top8227.instructionLoader.interruptInjector.interruptRequest
+ net115 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqSync.nextQ2
+ sky130_fd_sc_hd__dfrtp_1
X_2686_ _0291_ _0634_ _0639_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__o21ai_1
X_1568_ _0819_ _0848_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__nor2_1
X_1499_ net78 _0763_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__and2_1
Xfanout22 _0362_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xfanout33 net34 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xfanout44 _0728_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_1_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_2
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout99 net101 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_9_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout88 net90 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_2
Xfanout66 _0731_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
Xfanout77 net78 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2540_ _0458_ gpio[11] _0528_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
X_2471_ net21 _0458_ _0459_ _0470_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__and4b_1
Xclkload14 clknet_4_15_0_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinvlp_4
X_1422_ _0710_ _0716_ _0722_ _0718_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__a31oi_2
XPHY_EDGE_ROW_50_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1353_ net96 VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__inv_2
XFILLER_36_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2807_ clknet_4_5_0_clk _0083_ net123 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2738_ clknet_4_10_0_clk _0022_ net121 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload8 clknet_4_9_0_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_8
XFILLER_59_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2669_ _0309_ _0622_ _0291_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1971_ _0659_ gpio[22] _1243_ _0672_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__a211o_2
X_2454_ _0440_ _0465_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__a21oi_1
X_2385_ _0363_ _0364_ _0392_ _0393_ _0400_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__o311a_1
X_2523_ top8227.PSRCurrentValue\[2\] top8227.demux.setInterruptFlag net42 VGND VGND
+ VPWR VPWR _0516_ sky130_fd_sc_hd__or3_1
X_1405_ _0676_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_1
Xinput1 dataBusIn[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ net2 _1254_ _1256_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ _1262_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a221o_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1954_ net62 _1225_ _1226_ _0795_ _0772_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__a2111o_1
XFILLER_21_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1885_ net102 _0739_ _0750_ net61 VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__a31o_1
X_2437_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _0404_ _0443_
+ _0401_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__o22a_1
XFILLER_56_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2368_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _0384_ VGND VGND
+ VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
X_2506_ net179 _0192_ _0512_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_1
X_2299_ _0274_ _0284_ _0275_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o21ba_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1670_ _0819_ _0852_ _0897_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__or4_1
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2222_ net25 _0212_ _0218_ _0222_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a211o_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2084_ _1147_ _1348_ _0121_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__a21oi_2
X_2153_ net25 _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__nand2_1
XFILLER_61_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1937_ _1204_ _1206_ _1208_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__or3_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1799_ top8227.demux.state_machine.timeState\[1\] net57 _0770_ net105 VGND VGND VPWR
+ VPWR _1072_ sky130_fd_sc_hd__a22o_1
X_1868_ _0770_ _0793_ _1074_ net62 VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__o31a_1
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2771_ clknet_4_13_0_clk _0047_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_2840_ clknet_4_1_0_clk _0114_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_1584_ net178 net35 _0867_ _0873_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a22o_1
X_1722_ _0680_ net31 _0912_ _0945_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1653_ _0804_ net28 _0902_ _0932_ _0931_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__a221o_1
X_2205_ _0241_ _0242_ _0244_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_64_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2136_ _1306_ _0175_ _1308_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__o21bai_2
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2067_ _1331_ _1339_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__nor2_1
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2823_ clknet_4_1_0_clk _0099_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_2754_ clknet_4_8_0_clk net134 net120 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ sky130_fd_sc_hd__dfrtp_1
X_1705_ _0977_ _0979_ _0981_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__or4_1
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1567_ net4 net133 _0845_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__a21oi_1
X_1636_ _0843_ _0868_ _0903_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__and3_1
X_2685_ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] _0580_ _0638_
+ _0290_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _0713_ _0798_ net95 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__o21a_1
X_2119_ _0157_ _0158_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__and2b_1
Xfanout23 _0362_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xfanout34 net36 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xfanout45 net46 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xfanout56 _0776_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
Xfanout89 net90 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xfanout78 net79 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xfanout67 _0717_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_2
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2470_ _0120_ _0444_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__a21o_1
X_1421_ _0710_ _0716_ _0722_ _0718_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a31o_1
X_1352_ net88 VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__inv_2
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2806_ clknet_4_13_0_clk _0082_ net126 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_2737_ clknet_4_10_0_clk _0021_ net121 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2668_ _0309_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__or2_1
Xclkload9 clknet_4_10_0_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_6
X_2599_ _1330_ net184 _0568_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_1
X_1619_ net47 _0876_ _0897_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__and3_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1970_ _0825_ _1241_ _1242_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2522_ net157 _1265_ _0515_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
X_2453_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ net20 VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__o41a_1
X_2384_ net37 _0399_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__nand2_2
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1404_ net90 net91 net85 net82 VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__or4b_4
Xinput2 dataBusIn[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1884_ net41 _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__nor2_1
X_1953_ _0700_ _0701_ _0704_ _0688_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__o31a_1
X_2505_ net169 _0212_ _0512_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_1
X_2436_ _0446_ _0447_ _0449_ net37 VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__a31o_1
X_2367_ _0381_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nor2_1
X_2298_ net50 _1105_ _0287_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_24_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2152_ _0187_ _0191_ _1154_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_2
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2221_ _0249_ _0259_ _0248_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o21bai_2
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2083_ net25 _0122_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__and2_1
X_1936_ _1204_ _1206_ _1208_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__nor3_1
XPHY_EDGE_ROW_26_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1867_ net96 _1043_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__and2_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1798_ net60 _1066_ _1067_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_10_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2419_ _1090_ _0205_ _0406_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__a31o_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2770_ clknet_4_13_0_clk _0046_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_1721_ _0773_ net29 _0932_ _0998_ _0996_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__a221o_1
X_1583_ _0819_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__nor2_1
X_1652_ net40 _0923_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__and2_1
XFILLER_58_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2135_ top8227.internalDataflow.addressLowBusModule.busInputs\[35\] net24 _1310_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[27\] _0174_ VGND VGND VPWR
+ VPWR _0175_ sky130_fd_sc_hd__a221o_1
X_2204_ _0730_ _1303_ _1305_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_64_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2066_ _1280_ _1336_ _1337_ _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__a22o_1
X_1919_ _0681_ _1190_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__or3_1
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2822_ clknet_4_7_0_clk _0098_ net124 VGND VGND VPWR VPWR gpio[7] sky130_fd_sc_hd__dfrtp_4
X_2753_ clknet_4_8_0_clk net182 net120 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.irqGenerated
+ sky130_fd_sc_hd__dfrtp_1
X_1704_ _0786_ net27 net26 _0905_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__a221o_1
X_2684_ _0283_ _0635_ _0636_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__a22o_1
X_1566_ net4 _0845_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nor2_1
X_1635_ _0767_ net30 _0912_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__a22o_1
X_1497_ net88 _0673_ net76 VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__and3_1
XFILLER_39_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2049_ _1089_ _1321_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2118_ _0148_ _0156_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__nand2_1
Xfanout35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xfanout24 _1303_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_2
Xfanout46 net47 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xfanout68 _0717_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
Xfanout79 _0675_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_2
Xfanout57 _0687_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1351_ net111 VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__clkinv_4
X_1420_ net88 net91 net82 net85 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__or4_4
X_2805_ clknet_4_7_0_clk _0081_ net126 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_2
X_1618_ net132 _0871_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__or2_1
X_2736_ clknet_4_10_0_clk _0020_ net121 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2667_ _0306_ _0310_ _0312_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or3_1
X_1549_ top8227.instructionLoader.interruptInjector.resetDetected _0841_ VGND VGND
+ VPWR VPWR _0842_ sky130_fd_sc_hd__nor2_2
X_2598_ _0122_ top8227.internalDataflow.accRegToDB\[5\] _0568_ VGND VGND VPWR VPWR
+ _0088_ sky130_fd_sc_hd__mux2_1
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2521_ net149 _1330_ _0515_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
X_2452_ _0364_ _0392_ _0431_ _0453_ _0363_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o2111a_1
X_2383_ net37 _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and2_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1403_ net89 net92 net87 net84 VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor4b_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 dataBusIn[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_2
XFILLER_36_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2719_ clknet_4_15_0_clk _0007_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1883_ _1048_ _1060_ _1067_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor3_1
XFILLER_14_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1952_ net98 _0766_ _0774_ _0791_ _0762_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a2111o_1
X_2435_ _0447_ _0449_ _0446_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_47_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2504_ net171 _0237_ _0512_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_1
X_2366_ _0661_ _0360_ _0361_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__and3_1
X_2297_ _0782_ _1171_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__nor2_1
XFILLER_64_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_56_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2151_ _1127_ _0189_ _0190_ _1151_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__o31a_1
X_2082_ _1350_ _0120_ _1154_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_2
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2220_ _0248_ _0249_ _0259_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or3_1
X_1935_ net51 _1059_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__and2_1
X_1797_ net55 _1069_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__and2_1
X_1866_ net108 _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__and2_1
X_2418_ _0209_ _0408_ net19 _0210_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a2bb2o_1
X_2349_ _0364_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__nor2_1
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1720_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__inv_2
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1651_ net78 _0760_ net28 _0856_ _0902_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a32o_1
X_1582_ net2 _0870_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__nand2_1
X_2134_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _1304_ _1311_
+ net4 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a22o_1
X_2203_ net94 top8227.demux.state_machine.timeState\[1\] _0687_ VGND VGND VPWR VPWR
+ _0243_ sky130_fd_sc_hd__nand3b_1
X_2065_ _1276_ _1332_ _1280_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_64_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1849_ net41 _1120_ _1117_ net48 VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__o211a_2
X_1918_ _0757_ _0796_ _1138_ net109 VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__o31a_1
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ clknet_4_6_0_clk _0097_ net125 VGND VGND VPWR VPWR gpio[6] sky130_fd_sc_hd__dfrtp_4
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1703_ _0685_ _0735_ net30 _0878_ _0918_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__a32o_1
X_1634_ net31 _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__nor2_1
X_2752_ clknet_4_8_0_clk net145 net115 VGND VGND VPWR VPWR top8227.demux.nmi sky130_fd_sc_hd__dfrtp_4
X_2683_ _1343_ _0581_ _0585_ _1341_ _0282_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__o221a_1
X_1565_ top8227.demux.state_machine.currentAddress\[6\] net34 _0851_ _0856_ VGND VGND
+ VPWR VPWR _0009_ sky130_fd_sc_hd__a22o_1
X_1496_ net79 net65 VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__and2_1
X_2048_ _1152_ _1320_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_1_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2117_ _0148_ _0156_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__nor2_1
Xfanout36 _0838_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
Xfanout58 net59 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
Xfanout47 net48 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
Xfanout25 _1085_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout69 _0690_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2804_ clknet_4_7_0_clk _0080_ net126 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1617_ net132 _0871_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__nor2_2
X_2597_ _0147_ top8227.internalDataflow.accRegToDB\[4\] _0568_ VGND VGND VPWR VPWR
+ _0087_ sky130_fd_sc_hd__mux2_1
X_2735_ clknet_4_9_0_clk _0026_ net127 VGND VGND VPWR VPWR top8227.branchForward sky130_fd_sc_hd__dfrtp_1
X_2666_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\] _0580_ _0617_
+ _0621_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__a22o_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ net104 net79 _0678_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and3_1
X_1548_ top8227.demux.nmi top8227.instructionLoader.interruptInjector.irqGenerated
+ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__or2_2
XFILLER_54_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2451_ _0462_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nand2_1
X_2520_ net158 _0122_ _0515_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_1
X_1402_ net69 _0703_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__nor2_4
X_2382_ _0360_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or2_2
Xinput4 dataBusIn[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2718_ clknet_4_15_0_clk _0006_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2649_ _0602_ _0606_ _0291_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux2_1
XFILLER_27_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ _1089_ _1153_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__or2_2
X_1951_ _0688_ _0797_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a21oi_2
X_2434_ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__inv_2
X_2365_ _0360_ _0361_ _0661_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__a21o_1
X_2503_ _1182_ _0511_ net51 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__o21a_4
XFILLER_56_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2296_ _0173_ _0317_ _0332_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ sky130_fd_sc_hd__a21o_1
XFILLER_64_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ net3 _1130_ _1131_ top8227.PSRCurrentValue\[2\] _0188_ VGND VGND VPWR VPWR
+ _0190_ sky130_fd_sc_hd__a221o_1
X_2081_ _1147_ _0120_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__nor2_1
X_1934_ _1204_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nor2_2
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1796_ _0695_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__or2_2
X_1865_ net88 net76 _0682_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__and3_1
X_2417_ _0430_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__xnor2_1
X_2348_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] net20 VGND VGND
+ VPWR VPWR _0365_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2279_ _0315_ _0318_ _0314_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1581_ net7 _0868_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__or2_1
X_1650_ _0924_ _0928_ _0929_ _0886_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a211o_1
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2202_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _1304_ _1311_
+ net1 VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__a22oi_1
XFILLER_3_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _1147_ _0163_ _0170_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__a21oi_2
X_2064_ _1284_ _1332_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__or2_1
XFILLER_19_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1917_ net105 _0675_ net65 VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__and3_1
X_1848_ net41 _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1779_ net106 net70 net63 VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_4_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2820_ clknet_4_7_0_clk _0096_ net124 VGND VGND VPWR VPWR gpio[5] sky130_fd_sc_hd__dfrtp_4
XFILLER_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2751_ clknet_4_8_0_clk _0031_ net115 VGND VGND VPWR VPWR top8227.demux.setInterruptFlag
+ sky130_fd_sc_hd__dfrtp_4
X_1633_ net132 _0870_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__nand2_1
X_1564_ net40 _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and2_2
X_1702_ _0766_ net27 _0890_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__a22o_1
X_2682_ _1266_ _0294_ _0583_ _1342_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1495_ net79 net64 VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__and2_1
Xfanout37 _0397_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
X_2047_ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _1123_ _1318_
+ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__a211o_1
Xfanout26 _0883_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
X_2116_ _0150_ _0155_ _1280_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout59 _0671_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2803_ clknet_4_12_0_clk _0079_ net126 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_2734_ clknet_4_8_0_clk _0019_ net120 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1616_ net8 net40 _0871_ _0891_ _0896_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a41o_1
X_2596_ _0171_ top8227.internalDataflow.accRegToDB\[3\] _0568_ VGND VGND VPWR VPWR
+ _0086_ sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1547_ net95 net44 _0837_ net104 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a22o_1
X_2665_ _0290_ _0620_ _0618_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or3b_1
X_1478_ net98 net77 _0709_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__and3_1
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2450_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] net22 VGND VGND
+ VPWR VPWR _0463_ sky130_fd_sc_hd__or2_1
X_2381_ _0673_ net79 _0286_ _0841_ net40 VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__a32o_1
X_1401_ net88 net85 net82 net91 VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or4bb_4
Xinput5 dataBusIn[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2717_ clknet_4_15_0_clk _0005_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2579_ _0417_ _0555_ _1336_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a21o_1
X_2648_ _0283_ _0298_ _0603_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__a22oi_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1950_ _0805_ _1219_ _1220_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__or4_2
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1881_ _1089_ _1147_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nor2_4
X_2502_ net105 _0705_ net68 _0780_ _1067_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__a311o_1
X_2433_ net21 _0410_ _0423_ _0435_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__and4b_1
X_2364_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] net23 VGND VGND
+ VPWR VPWR _0381_ sky130_fd_sc_hd__and2_1
XFILLER_51_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2295_ _0315_ _0331_ _0330_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_2080_ _1127_ _0119_ _1151_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__o21a_1
X_1933_ _1174_ _1203_ _1194_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__mux2_1
X_1795_ net109 net93 VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__or2_1
X_1864_ _0701_ _0711_ net98 VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__o21a_1
X_2416_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] net22 _0393_
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__a21bo_1
X_2347_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] net20 VGND VGND
+ VPWR VPWR _0364_ sky130_fd_sc_hd__and2_1
X_2278_ _1046_ _0316_ top8227.PSRCurrentValue\[0\] VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__and3b_1
XFILLER_52_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ net7 _0868_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nor2_1
X_2201_ top8227.internalDataflow.addressLowBusModule.busInputs\[24\] _1297_ _1302_
+ net24 top8227.internalDataflow.addressLowBusModule.busInputs\[32\] VGND VGND VPWR
+ VPWR _0241_ sky130_fd_sc_hd__a32o_1
X_2132_ net25 _0171_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__nand2_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2063_ _1335_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__inv_2
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1847_ top8227.branchForward _1047_ _1067_ _1091_ _1118_ VGND VGND VPWR VPWR _1120_
+ sky130_fd_sc_hd__a2111oi_1
X_1916_ net48 _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__and2_1
X_1778_ _0681_ _1037_ _1049_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__or4_1
XFILLER_27_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1701_ net39 _0898_ _0952_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__and3_1
XFILLER_31_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2750_ clknet_4_2_0_clk _0030_ net114 VGND VGND VPWR VPWR top8227.negEdgeDetector.q1
+ sky130_fd_sc_hd__dfrtp_1
X_2681_ _1343_ _0273_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__xnor2_1
X_1632_ net53 _0880_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nor2_2
X_1563_ net132 net47 _0844_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__and3_1
X_1494_ net65 _0735_ net63 net70 net99 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__o311a_1
X_2115_ _1308_ _0153_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__or2_1
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout38 _0396_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
X_2046_ net7 _1130_ _1131_ top8227.PSRCurrentValue\[6\] VGND VGND VPWR VPWR _1319_
+ sky130_fd_sc_hd__a22o_1
Xfanout49 _0727_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_2
Xfanout27 net29 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2802_ clknet_4_12_0_clk _0078_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_2733_ clknet_4_9_0_clk _0018_ net120 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_2664_ _0123_ _0294_ _0587_ _0158_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a221o_1
X_2595_ _0192_ top8227.internalDataflow.accRegToDB\[2\] _0568_ VGND VGND VPWR VPWR
+ _0085_ sky130_fd_sc_hd__mux2_1
X_1615_ _0868_ _0885_ _0894_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__a211o_1
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1546_ top8227.demux.state_machine.timeState\[5\] net44 _0837_ top8227.demux.state_machine.timeState\[1\]
+ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a22o_1
X_1477_ _0676_ _0710_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__nor2_2
XFILLER_54_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2029_ _1294_ _1300_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__or2_1
XFILLER_35_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2380_ _1247_ _0395_ _0394_ net46 _1241_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o2111ai_2
X_1400_ net90 net87 net84 net92 VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__and4bb_4
Xinput6 dataBusIn[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2716_ clknet_4_14_0_clk _0004_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2647_ _0201_ _0265_ _0581_ _0604_ _0282_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__o311a_1
X_2578_ _1336_ _0417_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__nand3_1
X_1529_ net110 top8227.demux.state_machine.currentAddress\[5\] VGND VGND VPWR VPWR
+ _0829_ sky130_fd_sc_hd__and2_1
XFILLER_42_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1880_ _1133_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2501_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] _0404_ _0505_
+ _0510_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__o22a_1
X_2432_ _0410_ _0418_ _0435_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__or3_1
X_2363_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] net22 VGND VGND
+ VPWR VPWR _0380_ sky130_fd_sc_hd__xor2_1
XFILLER_44_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2294_ top8227.PSRCurrentValue\[3\] _0316_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1863_ _1134_ _1135_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nand2_1
X_1932_ _1174_ _1189_ _1203_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__or3_1
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2415_ _0430_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__inv_2
X_1794_ net113 net71 _0691_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__and3_2
X_2346_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] net21 VGND VGND
+ VPWR VPWR _0363_ sky130_fd_sc_hd__xor2_1
X_2277_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__inv_2
XFILLER_52_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2131_ _0165_ _0169_ _1154_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_2
X_2062_ _1333_ _1334_ _1308_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__o21ba_1
X_2200_ _1276_ _1283_ _0238_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1915_ _1158_ _1185_ _1186_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__o31a_1
X_1846_ _1065_ _1067_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__nor3_1
X_1777_ net105 net76 _0709_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2329_ net152 _0124_ _0348_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_1
XFILLER_25_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1631_ _0908_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__or2_1
X_2680_ _0633_ _0307_ _0622_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux2_1
X_1700_ _0784_ net27 net26 _0923_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__a221o_1
X_1562_ top8227.demux.state_machine.currentAddress\[7\] net36 _0853_ _0854_ VGND VGND
+ VPWR VPWR _0010_ sky130_fd_sc_hd__a211o_1
X_1493_ _0792_ _0793_ net98 VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__o21a_1
X_2114_ _1308_ _0153_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__nor2_1
X_2045_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[6\] _1127_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__a221o_1
Xfanout39 net40 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout28 net29 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
X_1829_ net95 net55 _1086_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__a21o_1
XFILLER_38_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2801_ clknet_4_12_0_clk _0077_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_14_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1614_ net45 _0862_ _0876_ net35 top8227.demux.state_machine.currentAddress\[9\]
+ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a32o_1
X_2594_ _0212_ net185 _0568_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
X_2732_ clknet_4_11_0_clk _0017_ net120 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2663_ _0791_ _0159_ _0286_ _0584_ _0157_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__a32o_1
X_1476_ top8227.demux.state_machine.timeState\[5\] net55 VGND VGND VPWR VPWR _0777_
+ sky130_fd_sc_hd__nand2_1
X_1545_ net97 net44 _0837_ top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR
+ VPWR _0017_ sky130_fd_sc_hd__a22o_1
X_2028_ _1224_ _1237_ _1299_ _1244_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_37_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 dataBusIn[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_36_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2715_ clknet_4_15_0_clk _0000_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2577_ _0128_ net21 _0420_ _0421_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__or4_1
X_2646_ _0201_ _0584_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nand2_1
X_1528_ net110 net100 VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__and2b_2
X_1459_ net89 net92 net83 net86 VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__and4_2
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2500_ net38 _0509_ _0403_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__a21o_1
X_2431_ _0191_ _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a21o_1
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2362_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] net22 VGND VGND
+ VPWR VPWR _0379_ sky130_fd_sc_hd__and2_1
XFILLER_37_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2293_ _0800_ _0804_ _0286_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__o21ai_1
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2629_ _0248_ _0249_ _0259_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1862_ top8227.demux.state_machine.currentAddress\[12\] _0828_ net58 VGND VGND VPWR
+ VPWR _1135_ sky130_fd_sc_hd__a21oi_1
X_1931_ _1174_ _1189_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nor3_4
X_1793_ _0806_ _0824_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__and2_1
X_2414_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] net22 VGND VGND
+ VPWR VPWR _0430_ sky130_fd_sc_hd__xnor2_2
XFILLER_6_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2345_ _0360_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__nand2_1
X_2276_ net50 _1098_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_53_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2061_ top8227.internalDataflow.addressLowBusModule.busInputs\[30\] _1310_ _1311_
+ net7 VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a22o_1
X_2130_ _1147_ _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1914_ _0827_ _1135_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__nand2_1
XFILLER_34_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_62_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1845_ net113 net75 net73 VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__and3_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1776_ _0656_ net72 _0716_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__nor3_1
X_2328_ net143 _0149_ _0348_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_1
XFILLER_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2259_ _0261_ _0263_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__xor2_2
XFILLER_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ _0733_ net31 _0856_ _0877_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a221o_1
X_1561_ _0846_ net53 _0839_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__and3b_1
X_1492_ net69 _0736_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__nor2_2
X_2113_ _0151_ _0152_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__nor2_1
X_2044_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__inv_2
Xfanout29 _0838_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_17_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1759_ _1029_ _1031_ _1032_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__or4_1
X_1828_ net104 net77 net75 VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__and3_1
XFILLER_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2800_ clknet_4_13_0_clk _0076_ net130 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_2731_ clknet_4_11_0_clk _0016_ net120 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_14_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1613_ net39 _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__and2_1
X_2593_ _0237_ top8227.internalDataflow.accRegToDB\[0\] _0568_ VGND VGND VPWR VPWR
+ _0083_ sky130_fd_sc_hd__mux2_1
X_1544_ top8227.demux.state_machine.timeState\[3\] net44 _0837_ top8227.demux.state_machine.timeState\[5\]
+ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__a22o_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2662_ _0271_ _0282_ _0615_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_39_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1475_ _0676_ _0736_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nor2_1
X_2027_ _1224_ _1237_ _1299_ _1244_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_37_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 dataBusIn[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2714_ top8227.PSRCurrentValue\[7\] _1267_ _0655_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_1
X_2576_ _0553_ _0554_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__or2_1
X_1527_ net94 top8227.demux.state_machine.currentAddress\[1\] _0823_ _0825_ _0826_
+ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a32oi_4
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2645_ _0172_ _0293_ _0583_ _0265_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o22a_1
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1389_ net89 top8227.demux.state_machine.currentInstruction\[0\] net84 net87 VGND
+ VGND VPWR VPWR _0691_ sky130_fd_sc_hd__and4b_4
X_1458_ _0754_ _0756_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__or3_1
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2361_ _0376_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nor2_1
X_2430_ _0186_ _0408_ net19 _0181_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__a2bb2o_1
X_2292_ _0194_ _0317_ _0328_ _0329_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2559_ net21 _0420_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__or2_1
X_2628_ _0586_ _0582_ _0248_ _0585_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1930_ net42 _1202_ _1170_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__o21a_2
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1861_ _0719_ _0720_ _0832_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__o21ai_1
X_1792_ top8227.branchForward _1047_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__and2_1
X_2413_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _0403_ _0429_
+ net38 _0402_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__a221o_1
X_2344_ top8227.instructionLoader.interruptInjector.resetDetected gpio[21] _0841_
+ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2275_ top8227.demux.setInterruptFlag net59 _1249_ net80 VGND VGND VPWR VPWR _0315_
+ sky130_fd_sc_hd__a31o_1
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2060_ top8227.internalDataflow.addressLowBusModule.busInputs\[38\] net24 _1304_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[22\] _1306_ VGND VGND VPWR
+ VPWR _1333_ sky130_fd_sc_hd__a221o_1
XFILLER_34_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1913_ _0790_ _1143_ _1176_ _1177_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__or4_1
X_1844_ _1115_ _1116_ _1113_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__o21ba_1
X_1775_ top8227.branchBackward _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__and2_1
XFILLER_57_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2327_ net139 _0173_ _0348_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
X_2258_ _0264_ _0266_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__xnor2_2
X_2189_ top8227.internalDataflow.addressLowBusModule.busInputs\[24\] _1214_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[40\] VGND VGND VPWR VPWR _0229_
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1560_ net132 _0844_ _0852_ net36 VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__a211oi_1
X_2112_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\] net24 _1304_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] _1306_ VGND VGND VPWR
+ VPWR _0152_ sky130_fd_sc_hd__a221o_1
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1491_ net71 net65 VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__and2_1
Xfanout19 _0405_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2043_ _1266_ _1315_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1827_ _0778_ _0791_ net107 VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__o21a_1
X_1689_ _0864_ _0952_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__a21o_1
X_1758_ _0970_ _0978_ _0981_ _1027_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_0_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2730_ clknet_4_8_0_clk _0015_ net120 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2661_ _0271_ _0616_ _0290_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__o21ai_1
X_1612_ net133 net45 _0847_ _0862_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__and4_1
X_1543_ _0835_ _0836_ _0839_ _0840_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a211o_1
X_1474_ net78 net66 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__and2_1
X_2592_ _0321_ _0567_ net50 VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_37_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2026_ _0739_ _1238_ _1298_ _0748_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_20_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 nrst VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2713_ _1143_ _0322_ _0654_ net50 VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__o31a_1
X_2644_ _0298_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__xnor2_1
X_2575_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _0403_ _0551_
+ net38 VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__a22o_1
X_1526_ net113 net100 net103 VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__nor3b_1
X_1457_ _0691_ net65 net67 VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__o21a_1
X_1388_ net80 net81 VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__nand2b_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2009_ _1040_ _1045_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__nor2_1
XFILLER_58_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2360_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] net22 VGND VGND
+ VPWR VPWR _0377_ sky130_fd_sc_hd__nor2_1
X_2291_ _0690_ _0722_ _0287_ _0316_ top8227.PSRCurrentValue\[2\] VGND VGND VPWR VPWR
+ _0329_ sky130_fd_sc_hd__o311a_1
XFILLER_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2627_ net107 net52 _0778_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__and3_1
X_2489_ _0496_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__xnor2_1
X_2558_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _0404_ _0539_
+ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__o21a_1
X_1509_ top8227.demux.state_machine.timeState\[3\] net57 _0791_ net99 VGND VGND VPWR
+ VPWR _0810_ sky130_fd_sc_hd__a22o_1
XFILLER_55_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _1123_ _1129_
+ _1132_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__a211o_1
XFILLER_14_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1791_ _1048_ _1055_ _1058_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__or4_1
X_2412_ _0427_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__nor2_1
X_2343_ _0730_ _0359_ _0836_ _0351_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2274_ _0801_ _0286_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nand2_1
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1989_ _1254_ _1256_ _1260_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__and4bb_1
XFILLER_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1912_ _1178_ _1181_ _1183_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__or4_1
X_1843_ net106 _0680_ net57 net98 _1114_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__a221o_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1774_ _0746_ _0747_ _0658_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__a21oi_2
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2326_ net151 _0194_ _0348_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
X_2257_ _0267_ _0269_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_63_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2188_ _1090_ _1152_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__and3_1
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1490_ net69 _0706_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nor2_4
X_2111_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\] _1310_ _1311_
+ net133 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a22o_1
XFILLER_39_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2042_ _1285_ _1314_ _1280_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__mux2_1
Xhold1 top8227.instructionLoader.interruptInjector.irqSync.nextQ2 VGND VGND VPWR VPWR
+ net134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1826_ _1049_ _1062_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__or2_1
X_1688_ _0704_ net34 _0921_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1757_ _0988_ _0996_ _1000_ _1002_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__or4_1
XFILLER_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2309_ net51 _1057_ _0340_ _0836_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ net133 _0862_ _0883_ net35 net166 VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a32o_1
XFILLER_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2660_ _0159_ _0615_ _0301_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__mux2_1
X_1542_ net110 top8227.demux.state_machine.timeState\[3\] net46 VGND VGND VPWR VPWR
+ _0840_ sky130_fd_sc_hd__mux2_1
X_2591_ net96 _0787_ _1165_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a211o_1
X_1473_ _0679_ _0710_ _0690_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__a21oi_2
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2025_ net93 _0822_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_59_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1809_ top8227.demux.state_machine.currentAddress\[1\] _0828_ net58 VGND VGND VPWR
+ VPWR _1082_ sky130_fd_sc_hd__a21o_1
X_2789_ clknet_4_4_0_clk _0065_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2574_ _0372_ _0373_ _0389_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__o31a_1
X_2712_ _0788_ _1105_ _1176_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or3_1
X_2643_ _0599_ _0600_ _0591_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__a21oi_1
X_1525_ top8227.demux.state_machine.currentAddress\[10\] top8227.demux.state_machine.currentAddress\[4\]
+ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__or2_4
X_1456_ net68 net65 VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and2_1
X_1387_ net80 net81 VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__and2b_2
XFILLER_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2008_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__inv_2
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2290_ top8227.demux.setInterruptFlag net59 net49 _1249_ VGND VGND VPWR VPWR _0328_
+ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_22_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2557_ _0396_ _0537_ _0538_ _0403_ _0536_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a311o_1
XFILLER_9_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2626_ _0213_ _0293_ _0583_ _0249_ _0585_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o221a_1
X_2488_ _0497_ _0498_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__nand2_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1439_ net80 _0674_ net81 top8227.PSRCurrentValue\[0\] VGND VGND VPWR VPWR _0740_
+ sky130_fd_sc_hd__or4b_1
X_1508_ net104 _0677_ _0783_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a211o_1
XFILLER_62_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1790_ net107 _0774_ _1059_ _1061_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a2111o_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2411_ _0409_ _0418_ _0424_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and3_1
X_2342_ _0354_ _0358_ _1224_ _0352_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__and4b_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2273_ _0291_ _0311_ _0312_ _0295_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__o31a_1
X_1988_ net94 top8227.demux.state_machine.timeState\[1\] _0687_ net51 VGND VGND VPWR
+ VPWR _1261_ sky130_fd_sc_hd__o211a_2
XFILLER_20_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2609_ gpio[1] _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nand2_1
XFILLER_57_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1842_ net102 _0693_ net60 VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__a21o_1
X_1911_ net102 _0677_ net55 net93 _1180_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a221o_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1773_ _1041_ _1044_ net50 VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__o21a_1
XFILLER_57_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2187_ top8227.internalDataflow.addressLowBusModule.busInputs\[16\] _1123_ _1127_
+ _0225_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__a2111o_1
XPHY_EDGE_ROW_40_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2325_ net147 _0220_ _0348_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
X_2256_ _1316_ _0284_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2041_ _1308_ _1313_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nor2_2
XFILLER_47_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2110_ _1284_ _1277_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_1
Xhold2 top8227.instructionLoader.interruptInjector.nmiSync.nextQ2 VGND VGND VPWR VPWR
+ net135 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1756_ _0876_ _1030_ _1026_ _1019_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a211o_1
X_1825_ _0735_ net63 net104 net76 VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__o211a_1
X_1687_ _0843_ _0903_ _0951_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a21oi_2
X_2308_ net113 _0825_ _0828_ top8227.demux.state_machine.currentAddress\[1\] VGND
+ VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a22o_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ _1073_ _0277_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_23_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1610_ net39 _0867_ _0872_ net35 net173 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a32o_1
X_2590_ net109 _0764_ _0791_ net98 _1196_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a221o_1
X_1541_ net42 _0819_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__nor2_2
X_1472_ _0679_ net69 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__nor2_1
X_2024_ _1286_ _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__nor2_1
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1808_ _0656_ top8227.demux.state_machine.currentAddress\[12\] _0695_ _1080_ VGND
+ VGND VPWR VPWR _1081_ sky130_fd_sc_hd__a31o_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2788_ clknet_4_4_0_clk _0064_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_1739_ _0961_ _1011_ _1012_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__or4_1
XFILLER_18_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2711_ top8227.demux.isAddressing net35 _0653_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2573_ _0390_ _0401_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__nor2_1
X_1524_ net103 net62 VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or2_1
X_2642_ _0299_ _0598_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__nand2_1
X_1386_ net104 net95 VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__or2_2
X_1455_ _0705_ net63 net67 VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__o21a_1
XFILLER_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2007_ _1057_ _1278_ _1279_ net51 VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__o31a_2
XFILLER_23_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2487_ _0482_ _0483_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nand2_1
X_2556_ _0199_ _0534_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__or2_1
X_1507_ net66 _0760_ net97 net78 VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o211a_1
X_2625_ net50 _1099_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nand2_2
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1369_ top8227.pulse_slower.currentEnableState\[1\] top8227.pulse_slower.currentEnableState\[0\]
+ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or2_2
X_1438_ _0737_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__nand2b_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2410_ _0418_ _0424_ _0409_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a21oi_1
X_2341_ _1231_ _1236_ _0355_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__and4_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2272_ _0296_ _0305_ _1316_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a21o_1
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1987_ _1139_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__nor2_1
X_2539_ _0446_ gpio[10] _0528_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_57_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2608_ gpio[0] _0575_ _0245_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_58_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1910_ _0779_ _0780_ _1056_ _1101_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__or4_1
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1772_ net105 net77 net66 VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__and3_1
X_1841_ _0702_ _0735_ net67 net106 VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__o211a_1
X_2324_ net148 _0239_ _0348_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2186_ net1 _1130_ _1131_ top8227.PSRCurrentValue\[0\] VGND VGND VPWR VPWR _0226_
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2255_ _1085_ _0237_ _0294_ _0290_ _0285_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a311o_1
XFILLER_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold3 top8227.demux.state_machine.currentAddress\[8\] VGND VGND VPWR VPWR net136
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _1309_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nor2_1
XFILLER_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1755_ net5 net46 _0857_ _0898_ _0865_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__a41o_1
X_1824_ _0833_ _1078_ _1096_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__a21o_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_30_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1686_ _0855_ _0924_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a21o_1
XFILLER_38_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2307_ top8227.branchForward _0338_ _0339_ _0313_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__a22o_1
X_2238_ _1037_ _1052_ _1059_ _1114_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__or4_1
X_2169_ _0206_ _0207_ _0208_ _1209_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ net45 net40 VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__nand2_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1471_ net99 _0770_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a21o_1
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2023_ net48 _1293_ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__a21oi_2
X_1807_ net111 top8227.demux.state_machine.currentAddress\[7\] _1078_ _1079_ _1077_
+ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__a221o_1
X_1669_ _0844_ _0904_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__or2_1
X_2787_ clknet_4_5_0_clk _0063_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_1738_ net74 _0705_ net27 _0878_ _0905_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_36_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2710_ top8227.demux.isAddressing net43 _0835_ net59 VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2572_ _0127_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__xnor2_1
X_1523_ net111 net103 net100 VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__nor3_1
XFILLER_4_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1454_ net84 net87 net90 net92 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__and4b_1
X_2641_ _0299_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__or2_1
X_1385_ net75 net74 VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__and2_2
XFILLER_50_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2006_ _1059_ _1067_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__or2_1
XFILLER_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2839_ clknet_4_1_0_clk _0113_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2624_ net50 _1099_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__and2_1
XFILLER_20_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2486_ _0470_ _0471_ _0482_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__or3_1
X_2555_ _0199_ _0534_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nand2_1
X_1437_ _0674_ _0679_ _0692_ _0706_ net72 VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__a41o_1
X_1506_ _0693_ _0806_ top8227.demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR
+ _0807_ sky130_fd_sc_hd__o21a_1
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1368_ top8227.demux.state_machine.currentAddress\[2\] top8227.demux.state_machine.currentAddress\[9\]
+ _0669_ top8227.demux.isAddressing VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or4b_1
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2340_ net93 _0806_ _1228_ _1250_ _1249_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a221oi_1
X_2271_ _0306_ _0310_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__nor2_1
X_1986_ net100 _0693_ _1118_ _1181_ _1258_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__a2111o_1
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ _1095_ _0573_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__o21bai_4
X_2538_ _0435_ gpio[9] _0528_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2469_ _1348_ _0408_ _0405_ _1349_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1840_ _0832_ _1110_ _1112_ _1111_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__o31ai_1
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1771_ _1042_ _1043_ net108 VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__o21a_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2323_ _1142_ _0347_ _0346_ net49 VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o211a_2
X_2254_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__inv_2
X_2185_ top8227.internalDataflow.addressHighBusModule.busInputs\[16\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[0\] VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a22o_1
X_1969_ top8227.demux.state_machine.currentAddress\[6\] _1078_ net59 net111 VGND VGND
+ VPWR VPWR _1242_ sky130_fd_sc_hd__a211o_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 top8227.pulse_slower.currentEnableState\[0\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1823_ net58 _1093_ _1094_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__or4_1
XFILLER_30_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1685_ net79 _0702_ net30 VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__and3_1
X_1754_ _0931_ _0958_ _0962_ _0992_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__or4_1
XFILLER_38_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2306_ _0664_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] net51
+ _1057_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__and4_1
X_2237_ net107 _0774_ _1061_ _1190_ _0681_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__a2111o_1
X_2099_ _1162_ _0137_ _0138_ _1160_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__a2bb2o_1
X_2168_ top8227.internalDataflow.addressLowBusModule.busInputs\[33\] _1211_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[41\] VGND VGND VPWR VPWR _0208_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ net109 net70 net66 VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2022_ top8227.demux.state_machine.currentAddress\[5\] top8227.demux.state_machine.currentAddress\[1\]
+ _0836_ net110 VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__o211a_1
X_1806_ top8227.demux.state_machine.currentAddress\[1\] top8227.demux.state_machine.currentAddress\[6\]
+ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__or2_1
X_2786_ clknet_4_4_0_clk _0062_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1599_ top8227.demux.state_machine.currentAddress\[2\] net35 _0869_ _0885_ _0886_
+ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__a221o_1
X_1668_ net45 _0922_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_37_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1737_ _0911_ _0991_ _1006_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__or4_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2640_ _1282_ _0288_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__or2_2
X_2571_ _0155_ _0415_ _0546_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a21oi_1
X_1522_ net109 net102 VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__or2_1
XFILLER_4_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1453_ net75 _0702_ net66 _0735_ net67 VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__o41a_1
X_2005_ net102 net56 _1138_ net100 VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a22o_1
X_1384_ net80 net81 VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__or2_1
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2769_ clknet_4_7_0_clk _0045_ net126 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_2838_ clknet_4_4_0_clk _0112_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2554_ _0387_ net38 _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_30_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2623_ net52 _1050_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__nand2_1
X_2485_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__inv_2
X_1367_ top8227.demux.state_machine.currentAddress\[2\] top8227.demux.state_machine.currentAddress\[9\]
+ _0669_ top8227.demux.isAddressing VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nor4b_2
X_1505_ net79 net75 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__and2_2
X_1436_ _0702_ net66 _0734_ _0735_ net73 VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__o41a_1
XFILLER_62_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2270_ _0307_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__and2_1
XFILLER_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ _0677_ _0680_ net109 VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__o21a_1
X_2537_ _0410_ gpio[8] _0528_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_1
X_2606_ _0352_ _0517_ _0572_ net42 VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a31o_1
X_2468_ _0476_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_58_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2399_ _0155_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__nand2_1
XFILLER_28_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1419_ net89 net92 net83 net86 VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__nor4_2
XFILLER_43_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1770_ _0754_ _0775_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__or2_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2322_ _1115_ _1137_ _1258_ _1279_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or4_1
X_2253_ _0286_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__nand2_2
X_2184_ _0223_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__inv_2
X_1968_ top8227.demux.state_machine.currentAddress\[7\] top8227.demux.state_machine.currentAddress\[6\]
+ net59 VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__or3_1
X_1899_ _0754_ _0769_ _0784_ _1171_ net108 VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__o41a_1
XFILLER_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold5 top8227.pulse_slower.nextEnableState\[1\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1822_ top8227.demux.state_machine.currentAddress\[1\] _0824_ VGND VGND VPWR VPWR
+ _1095_ sky130_fd_sc_hd__and2_1
X_1753_ _0914_ _0998_ _1010_ _0994_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__a211o_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_29_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1684_ _0942_ _0956_ _0961_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__or4_1
X_2167_ top8227.internalDataflow.accRegToDB\[1\] _1212_ _1214_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\]
+ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a22oi_1
X_2305_ net51 _1057_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2236_ net60 _1038_ _1045_ _1066_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__or4_2
X_2098_ net133 _1255_ _1257_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\]
+ _1327_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2021_ net48 _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__and2_1
XFILLER_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1805_ net103 _0658_ net111 VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__a21o_1
X_1736_ _0934_ _0946_ _0982_ _1007_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__or4b_1
X_2785_ clknet_4_4_0_clk _0061_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_1598_ gpio[21] _0847_ _0861_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__and3_1
X_1667_ _0720_ net34 _0858_ _0899_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__a221o_1
XFILLER_53_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2219_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__inv_2
XFILLER_41_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2570_ _0389_ _0548_ _0549_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__o21ai_1
X_1521_ net111 net101 VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__or2_1
X_1383_ net80 net81 VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nor2_2
X_1452_ net75 net66 net67 VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__o21a_1
X_2004_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2768_ clknet_4_7_0_clk _0044_ net126 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_2
X_1719_ _0846_ _0860_ _0888_ net53 VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a31o_1
X_2699_ _0649_ _0650_ net52 VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o21a_4
X_2837_ clknet_4_1_0_clk _0111_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2553_ _0380_ _0386_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__nor2_1
X_1504_ _0803_ _0804_ net97 VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__o21a_1
X_2622_ _0248_ _0249_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__or3_1
X_1366_ top8227.demux.state_machine.currentAddress\[8\] top8227.demux.state_machine.currentAddress\[0\]
+ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__or2_1
X_2484_ _1322_ net19 _0408_ _1326_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__o221a_1
X_1435_ net91 net85 net82 net88 VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__or4bb_2
XFILLER_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1984_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__inv_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2467_ _0477_ _0478_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__nand2_1
X_2536_ net42 _0524_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or3b_4
X_2605_ top8227.demux.state_machine.currentAddress\[6\] _1069_ _1093_ _0526_ VGND
+ VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_58_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2398_ _0177_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__nor2_1
XFILLER_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1418_ _0710_ _0718_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nor2_2
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2321_ _1113_ _1134_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__nand2_1
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2183_ _0218_ _0222_ _0213_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__o21ba_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2252_ net76 _0702_ _0753_ _0700_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a211o_1
XFILLER_33_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ _1224_ _1237_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__and3_1
X_1898_ _0775_ _0785_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__or2_2
X_2519_ net160 _0147_ _0515_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_1
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold6 net13 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1821_ top8227.demux.state_machine.currentAddress\[7\] _0830_ net111 VGND VGND VPWR
+ VPWR _1094_ sky130_fd_sc_hd__o21a_1
X_1752_ net56 net30 _0884_ _0945_ _0985_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a221o_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1683_ _0711_ net27 _0918_ _0924_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__a221o_1
XFILLER_57_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2304_ gpio[18] _0726_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__nand2_1
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2097_ _1210_ _0136_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__nand2_1
X_2166_ _0660_ _1206_ _1205_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _1343_ _0273_ _1317_ _1341_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2020_ _1047_ _1289_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__o21ba_1
XFILLER_35_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1804_ _0825_ _0828_ net59 VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__a21o_1
X_1666_ _0683_ net68 net32 _0890_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__a32o_1
X_2784_ clknet_4_4_0_clk _0060_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_1735_ _0707_ net30 _0905_ _0924_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__a22o_1
X_1597_ net45 net39 _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__and3_1
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2149_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[2\] VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ net49 _0257_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1520_ top8227.instructionLoader.interruptInjector.resetDetected gpio[21] VGND VGND
+ VPWR VPWR _0820_ sky130_fd_sc_hd__or2_1
X_1451_ _0748_ _0751_ _0739_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o21a_1
X_1382_ net81 _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__and2b_1
X_2003_ _1048_ _1065_ _1275_ _1269_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_33_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2836_ clknet_4_4_0_clk _0110_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_2767_ clknet_4_13_0_clk _0043_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_1649_ net71 _0760_ net33 VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__and3_1
X_2698_ _0683_ net63 net70 net100 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__o211a_1
X_1718_ _0768_ net28 _0890_ _0914_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__a22o_1
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2552_ net22 _0419_ _0413_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__o21ba_1
X_2483_ _1328_ net19 VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__nand2_1
X_1503_ net74 _0760_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__and2_1
X_2621_ _0656_ net41 _0791_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__or3b_2
X_1365_ gpio[20] VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__inv_2
X_1434_ top8227.demux.state_machine.currentInstruction\[0\] net87 net84 net89 VGND
+ VGND VPWR VPWR _0735_ sky130_fd_sc_hd__and4bb_4
XFILLER_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2819_ clknet_4_6_0_clk _0095_ net124 VGND VGND VPWR VPWR gpio[4] sky130_fd_sc_hd__dfrtp_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1983_ _1240_ _1244_ _1253_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__nor3_4
X_2604_ _0356_ _0518_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__and3_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2466_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] net23 VGND VGND
+ VPWR VPWR _0478_ sky130_fd_sc_hd__nand2_1
X_2535_ _0825_ _1078_ _1079_ _1069_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a221o_1
X_1417_ _0716_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nor2_1
X_2397_ _0199_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__nand2_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2320_ _0666_ _0328_ _0345_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o21ai_1
X_2251_ _0288_ _0289_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__or2_4
X_2182_ _1283_ _0220_ _0221_ _1281_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1966_ _0751_ net62 _1238_ _0739_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__o22ai_1
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1897_ _0659_ gpio[22] _1169_ _0672_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a211o_1
X_2449_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] net22 VGND VGND
+ VPWR VPWR _0462_ sky130_fd_sc_hd__nand2_1
X_2518_ net156 _0171_ _0515_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold7 net17 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ net62 _0825_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__and2_1
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1751_ _0956_ _1017_ _1024_ _1025_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__or4_1
X_1682_ _0778_ net28 _0882_ _0919_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__a22o_1
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2303_ clknet_4_8_0_clk top8227.pulse_slower.nextEnableState\[0\] VGND VGND VPWR
+ VPWR gpio[24] sky130_fd_sc_hd__and2_2
X_2234_ _1343_ _0273_ _1341_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__o21a_1
X_2165_ _0202_ _0203_ _0204_ _1152_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__o31a_1
X_2096_ top8227.internalDataflow.stackBusModule.busInputs\[36\] _1204_ _1207_ _0135_
+ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ _0688_ _0711_ _0781_ _0783_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__a2111o_1
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2783_ clknet_4_4_0_clk _0059_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_1803_ _1065_ _1071_ _1072_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ net53 _0860_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__nor2_2
X_1665_ net34 _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__nor2_2
X_1734_ _0791_ net31 net26 _0943_ _1010_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a221o_1
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2217_ _0250_ _0252_ _0255_ _0256_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__a22o_1
X_2148_ top8227.internalDataflow.addressLowBusModule.busInputs\[18\] _1109_ _1122_
+ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__and3_1
X_2079_ top8227.internalDataflow.addressLowBusModule.busInputs\[21\] _1123_ _1130_
+ net132 _0118_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ net102 _0749_ net93 VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__a21o_1
X_1381_ net86 net83 net92 net89 VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__and4b_2
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2002_ _1270_ _1272_ _1273_ _1274_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__or4_1
X_2766_ clknet_4_13_0_clk _0042_ net128 VGND VGND VPWR VPWR top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2835_ clknet_4_4_0_clk _0109_ net118 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_1579_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__inv_2
X_1648_ net42 _0913_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nor2_1
X_2697_ _0761_ _0767_ net109 VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__o21a_1
X_1717_ _0964_ _0984_ _0987_ _0995_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__or4_1
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2620_ _1270_ _0577_ _0578_ _1269_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__o31ai_4
X_2482_ net38 _0491_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or3b_1
X_2551_ net38 _0531_ _0533_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a21o_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1502_ net69 _0722_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__nor2_1
X_1433_ net92 net84 net87 net90 VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__and4bb_1
XFILLER_55_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1364_ gpio[16] VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiSync.in
+ sky130_fd_sc_hd__inv_2
XFILLER_11_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2818_ clknet_4_7_0_clk _0094_ net124 VGND VGND VPWR VPWR gpio[3] sky130_fd_sc_hd__dfrtp_4
X_2749_ clknet_4_2_0_clk _0029_ net115 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1982_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__inv_2
X_2534_ _0828_ _0830_ _0525_ _0829_ net58 VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__a2111o_1
X_2603_ _0739_ _1069_ _0570_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__a21oi_1
X_2465_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] net23 VGND VGND
+ VPWR VPWR _0477_ sky130_fd_sc_hd__or2_1
X_2396_ _0217_ net23 _0411_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__and3_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1416_ net80 net81 VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nand2_2
XFILLER_28_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout130 net131 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2250_ _0288_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2181_ _0205_ _0219_ _1277_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__o21ai_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1965_ net74 net63 net62 VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__and3_1
XFILLER_33_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1896_ net58 _1167_ _1168_ _1166_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__o31ai_1
X_2517_ net153 _0192_ _0515_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
X_2448_ _0401_ _0455_ _0461_ net37 _0456_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__o221a_1
X_2379_ _1247_ _0395_ _0394_ net46 _1241_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_3_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold8 net16 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ top8227.demux.state_machine.currentInstruction\[5\] _0721_ net32 VGND VGND
+ VPWR VPWR _1026_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_17_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1681_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__inv_2
X_2164_ net2 _1130_ _1131_ top8227.PSRCurrentValue\[1\] VGND VGND VPWR VPWR _0204_
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2302_ _0668_ net155 net49 _0337_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ sky130_fd_sc_hd__a31o_1
X_2233_ _0133_ _0272_ _0131_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2095_ top8227.internalDataflow.addressLowBusModule.busInputs\[28\] _1214_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[44\] _0134_ VGND VGND VPWR VPWR
+ _0135_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1879_ _1148_ _1151_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__and2_1
X_1948_ _0657_ _0673_ net76 _0695_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__and4_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2782_ clknet_4_4_0_clk _0058_ net122 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_1733_ _0705_ net68 net32 _0894_ _0897_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__a32o_1
X_1802_ _1073_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__or2_1
X_1664_ net6 net8 _0843_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__or3_1
X_1595_ net39 _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__and2_1
X_2147_ _1162_ _0186_ _0181_ _1160_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2216_ top8227.freeCarry _0254_ net59 VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2078_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[5\] _1131_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ net85 net82 VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and2b_1
X_2001_ net60 _1061_ _1062_ _1114_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__or4_1
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2834_ clknet_4_1_0_clk _0108_ net118 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_2765_ clknet_4_2_0_clk _0041_ net114 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_2696_ _0642_ _0648_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
+ _0579_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__o2bb2a_1
X_1716_ _0991_ _0993_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__or3_1
X_1578_ net8 net54 VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nand2_2
X_1647_ _0911_ _0920_ _0925_ _0926_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__or4b_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2550_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _0403_ _0532_
+ _0385_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a22o_1
XFILLER_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2481_ _0477_ _0490_ _0489_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__a21o_1
X_1432_ net72 _0692_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nor2_1
X_1363_ gpio[17] VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.interruptRequest
+ sky130_fd_sc_hd__inv_2
X_1501_ _0800_ _0801_ net97 VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_43_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2748_ clknet_4_12_0_clk _0028_ net128 VGND VGND VPWR VPWR top8227.instructionLoader.interruptInjector.resetDetected
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_52_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2817_ clknet_4_12_0_clk _0093_ net128 VGND VGND VPWR VPWR gpio[2] sky130_fd_sc_hd__dfrtp_4
X_2679_ _0598_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_61_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1981_ _1240_ _1244_ _1253_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__o21a_2
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2533_ top8227.demux.state_machine.currentAddress\[7\] _0821_ _1291_ VGND VGND VPWR
+ VPWR _0525_ sky130_fd_sc_hd__a21bo_1
X_2602_ _0693_ _0519_ _0569_ _1115_ _1118_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a2111o_1
X_2464_ _0464_ _0467_ _0462_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__o21ai_1
X_2395_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__inv_2
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1415_ net80 net81 VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__and2_1
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout131 net9 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__buf_2
Xfanout120 net9 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_57_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2180_ _0205_ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1895_ top8227.demux.state_machine.currentAddress\[11\] top8227.demux.state_machine.currentAddress\[12\]
+ top8227.demux.state_machine.currentAddress\[4\] net110 VGND VGND VPWR VPWR _1168_
+ sky130_fd_sc_hd__o31a_1
X_1964_ _1227_ _1231_ _1235_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__and4b_1
X_2447_ _0458_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__xnor2_1
X_2516_ net146 _0212_ _0515_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2378_ net71 _0731_ _0828_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold9 top8227.internalDataflow.stackBusModule.busInputs\[32\] VGND VGND VPWR VPWR
+ net142 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1680_ _0957_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__nor2_1
X_2301_ _1171_ _0286_ _0289_ _0335_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a41o_1
X_2163_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[1\] _1127_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__a221o_1
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2232_ _0159_ _0270_ _0157_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__a21o_1
X_2094_ top8227.internalDataflow.addressLowBusModule.busInputs\[36\] _1211_ _1212_
+ top8227.internalDataflow.accRegToDB\[4\] VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1878_ _1122_ _1125_ _1126_ _1150_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__or4_2
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1947_ _0724_ _0778_ _0784_ _0787_ net62 VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__o41a_1
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2781_ clknet_4_6_0_clk _0057_ net124 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_1663_ net6 _0844_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__and2b_1
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1732_ _0927_ _0942_ _1009_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__or3_1
X_1801_ net105 _0798_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__and2_1
X_1594_ net2 net1 net54 VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ top8227.demux.state_machine.currentAddress\[1\] _0826_ _1077_ VGND VGND VPWR
+ VPWR _0255_ sky130_fd_sc_hd__a21o_1
X_2077_ _1162_ _1348_ _1349_ _1160_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2146_ _0182_ _0183_ _0184_ _1209_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__a31o_1
XFILLER_41_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2000_ _0806_ _0822_ _1068_ net55 _1056_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a221o_1
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2833_ clknet_4_4_0_clk _0107_ net117 VGND VGND VPWR VPWR top8227.internalDataflow.stackBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_1715_ _0797_ net34 _0856_ _0912_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a22o_1
X_1646_ _0674_ _0686_ _0839_ _0879_ _0913_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__o32a_1
X_2764_ clknet_4_2_0_clk _0040_ net114 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
X_2695_ _0291_ _0647_ _0580_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__a21oi_1
X_1577_ net133 net45 _0857_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__and3_1
X_2129_ _1127_ _0166_ _0167_ _0168_ _1151_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__o41a_1
XFILLER_41_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2480_ _0477_ _0489_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__and3_1
X_1500_ net78 _0691_ _0763_ net74 VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__a22o_1
X_1362_ net133 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__inv_2
X_1431_ _0685_ net66 VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nand2_1
X_2816_ clknet_4_6_0_clk _0092_ net125 VGND VGND VPWR VPWR gpio[1] sky130_fd_sc_hd__dfrtp_4
X_1629_ _0693_ net33 _0885_ _0905_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a22o_1
X_2747_ clknet_4_9_0_clk _0027_ net119 VGND VGND VPWR VPWR top8227.freeCarry sky130_fd_sc_hd__dfrtp_1
X_2678_ _0307_ _0309_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__xor2_1
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ net48 _1248_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__and3_1
XFILLER_20_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2463_ top8227.internalDataflow.addressHighBusModule.busInputs\[20\] _0403_ _0468_
+ _0400_ _0475_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a221o_1
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2532_ _1227_ _1299_ _0517_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__and4b_1
X_2601_ _0684_ net55 _1228_ _0697_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__o22a_1
XFILLER_5_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2394_ _0245_ _0398_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__and2_1
X_1414_ net91 net83 net86 net90 VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__or4b_4
XFILLER_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout110 net111 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xfanout132 net6 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_2
Xfanout121 net9 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1894_ _0829_ _0831_ _0719_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__o21a_1
X_1963_ _0775_ net62 _0802_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__a21oi_1
X_2446_ _0447_ _0449_ _0446_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux2_1
X_2515_ net159 _0237_ _0515_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_1
X_2377_ _0771_ _1047_ _1158_ _1251_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or4_2
XFILLER_24_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2300_ net50 _1105_ _1332_ _0334_ top8227.PSRCurrentValue\[6\] VGND VGND VPWR VPWR
+ _0336_ sky130_fd_sc_hd__a32o_1
X_2231_ _0159_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__and2_1
X_2162_ top8227.internalDataflow.addressLowBusModule.busInputs\[17\] _1109_ _1122_
+ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and3_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2093_ _0131_ _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__and2b_2
XFILLER_61_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1877_ _1048_ _1149_ net51 VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__o21a_1
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1946_ _0754_ _0756_ _0758_ _0769_ net96 VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__o41a_1
X_2429_ _1154_ _0406_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__and2_1
XFILLER_29_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ _0704_ _0793_ net106 VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__o21a_1
X_2780_ clknet_4_5_0_clk _0056_ net123 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_1662_ _0934_ _0935_ _0938_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__or4_1
X_1731_ _0977_ _1005_ _1006_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__or4_1
X_1593_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__inv_2
X_2214_ _0708_ _1171_ _0253_ top8227.PSRCurrentValue\[0\] net108 VGND VGND VPWR VPWR
+ _0254_ sky130_fd_sc_hd__o311a_1
X_2076_ net132 _1255_ _1257_ top8227.internalDataflow.addressHighBusModule.busInputs\[21\]
+ _1327_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__o221a_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2145_ _0182_ _0183_ _0184_ _1209_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a31oi_1
XFILLER_26_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1929_ _1082_ _1201_ _1197_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__o21ai_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2763_ clknet_4_3_0_clk _0039_ net114 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
X_2832_ clknet_4_11_0_clk net138 net120 VGND VGND VPWR VPWR top8227.pulse_slower.currentEnableState\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1576_ _0864_ _0866_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__or2_1
X_1645_ _0701_ net34 _0923_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__a22o_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2694_ _0283_ _0643_ _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__a21o_1
X_1714_ _0792_ net28 _0890_ _0932_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a221o_1
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2128_ net4 _1130_ _1131_ top8227.PSRCurrentValue\[3\] VGND VGND VPWR VPWR _0168_
+ sky130_fd_sc_hd__a22o_1
X_2059_ _1148_ _1326_ _1321_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__o21ai_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1430_ net89 net92 net84 net87 VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__and4bb_2
X_1361_ net181 VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2815_ clknet_4_7_0_clk _0091_ net127 VGND VGND VPWR VPWR gpio[0] sky130_fd_sc_hd__dfrtp_4
X_2746_ clknet_4_3_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ net114 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1559_ _0846_ net53 VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__or2_1
X_1628_ _0901_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__or2_1
X_2677_ _0307_ _0309_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nor2_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2600_ _1265_ top8227.internalDataflow.accRegToDB\[7\] _0568_ VGND VGND VPWR VPWR
+ _0090_ sky130_fd_sc_hd__mux2_1
XFILLER_42_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2462_ _0470_ _0473_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__o21a_1
X_2393_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__inv_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2531_ _1236_ _0518_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__and3_1
X_1413_ _0700_ _0701_ _0704_ _0712_ _0695_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__o41ai_2
X_2729_ clknet_4_9_0_clk _0014_ net120 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout133 net5 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout111 net112 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__buf_2
Xfanout122 net127 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_4
Xfanout100 net101 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ _0777_ _1233_ _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__and3_1
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1893_ net61 _1039_ _1163_ _1164_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__or4_1
X_2376_ _0364_ _0392_ _0363_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__o21ai_1
X_2445_ _0410_ _0426_ _0435_ _0446_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and4_1
X_2514_ net41 _0514_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nor2_4
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_49_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2230_ _0267_ _0269_ _0180_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__a21o_1
X_2161_ _0193_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2092_ _0123_ _0130_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or2_1
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1945_ _1210_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1876_ _0681_ _1052_ _1056_ _1061_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__or4_1
X_2428_ _0440_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__xor2_1
X_2359_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] net22 VGND VGND
+ VPWR VPWR _0376_ sky130_fd_sc_hd__and2_1
XFILLER_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1592_ _0667_ _0862_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nand2_2
X_1661_ _0789_ _0940_ _0839_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__mux2_1
XFILLER_7_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1730_ _0995_ _0999_ _1000_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__or4b_1
X_2144_ top8227.internalDataflow.addressLowBusModule.busInputs\[34\] _1211_ _1212_
+ top8227.internalDataflow.accRegToDB\[2\] VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a22oi_2
X_2213_ net66 _0735_ net67 VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__o21a_1
X_2075_ _1210_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__nand2_1
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1928_ net110 top8227.demux.state_machine.currentAddress\[10\] _0720_ _1199_ _1200_
+ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a221o_1
X_1859_ net8 _1130_ _1131_ top8227.PSRCurrentValue\[7\] VGND VGND VPWR VPWR _1132_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1713_ net39 _0893_ _0898_ net33 _0757_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__a32o_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2831_ clknet_4_8_0_clk top8227.pulse_slower.nextEnableState\[0\] net120 VGND VGND
+ VPWR VPWR top8227.pulse_slower.currentEnableState\[0\] sky130_fd_sc_hd__dfrtp_1
X_2762_ clknet_4_3_0_clk _0038_ net114 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
X_1575_ net39 _0848_ _0865_ net36 top8227.demux.state_machine.currentAddress\[4\]
+ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a32o_1
X_1644_ _0859_ _0860_ _0863_ _0921_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a31o_2
X_2693_ _1316_ _0645_ _0585_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[3\] VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a22o_1
X_2058_ net25 _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__nand2_1
XFILLER_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1360_ top8227.instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning VGND
+ VGND VPWR VPWR _0665_ sky130_fd_sc_hd__inv_2
XFILLER_48_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2814_ clknet_4_5_0_clk _0090_ net124 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2745_ clknet_4_3_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ net114 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[3\] sky130_fd_sc_hd__dfrtp_1
X_2676_ top8227.internalDataflow.addressLowBusModule.busInputs\[29\] _0580_ _0623_
+ _0624_ _0630_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__a221o_1
X_1558_ _0846_ net53 VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nor2_1
X_1627_ net79 _0691_ net32 _0902_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__a32o_1
X_1489_ _0784_ _0787_ _0789_ net96 VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__o31a_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ _1233_ _0520_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__and3_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2461_ _0470_ _0473_ net37 VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a21oi_1
X_2392_ _0235_ _0406_ _0408_ _0232_ _0407_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__o221a_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1412_ _0681_ _0694_ _0698_ net57 VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2728_ clknet_4_14_0_clk _0013_ net131 VGND VGND VPWR VPWR top8227.demux.state_machine.timeState\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_2659_ _0159_ _0270_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__nor2_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout112 net113 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout123 net127 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
Xfanout101 top8227.demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1961_ net93 top8227.demux.state_machine.timeState\[5\] _0693_ VGND VGND VPWR VPWR
+ _1234_ sky130_fd_sc_hd__o21ai_1
X_1892_ net108 net67 net63 VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__and3_1
X_2513_ net109 _0513_ _0794_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__a21oi_2
X_2375_ _0367_ _0391_ _0366_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o21a_1
X_2444_ _0169_ _0444_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_19_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2160_ _0195_ _0199_ _1280_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2091_ _0123_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__and2_1
X_1875_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__inv_2
X_1944_ top8227.internalDataflow.stackBusModule.busInputs\[39\] _1204_ _1207_ _1216_
+ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a211o_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2427_ _0393_ _0430_ _0441_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2358_ _0373_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__nor2_1
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2289_ _0220_ _0317_ _0324_ _0327_ VGND VGND VPWR VPWR top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ net136 net35 _0878_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a21o_1
X_1660_ _0843_ _0868_ _0939_ _0905_ _0851_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__a32o_1
X_2143_ top8227.internalDataflow.addressLowBusModule.busInputs\[26\] _1214_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[42\] VGND VGND VPWR VPWR _0183_
+ sky130_fd_sc_hd__a22oi_1
X_2212_ _1065_ _1278_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__or3_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2074_ top8227.internalDataflow.stackBusModule.busInputs\[37\] _1204_ _1207_ _1346_
+ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__a211o_1
X_1927_ net110 _0720_ net62 top8227.demux.state_machine.currentAddress\[3\] VGND VGND
+ VPWR VPWR _1200_ sky130_fd_sc_hd__o211a_1
X_1858_ _1109_ _1121_ _1124_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__and3_2
X_1789_ net108 net73 net63 VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__and3_1
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2830_ clknet_4_0_0_clk _0106_ net119 VGND VGND VPWR VPWR top8227.internalDataflow.addressLowBusModule.busInputs\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_1643_ net43 _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_1
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2761_ clknet_4_3_0_clk _0037_ net114 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
X_2692_ _0296_ _0581_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__o21ba_1
XANTENNA_1 _0687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1712_ _0988_ _0989_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__or3_1
X_1574_ net4 net3 net45 _0842_ _0863_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__o2111a_1
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2126_ top8227.internalDataflow.addressLowBusModule.busInputs\[19\] _1109_ _1122_
+ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__and3_1
X_2057_ _1154_ _1329_ _1322_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__o21ai_2
XFILLER_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2813_ clknet_4_5_0_clk _0089_ net123 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ net47 net40 _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__and3_1
X_2744_ clknet_4_3_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ net114 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2675_ _0626_ _0629_ _0291_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__o21a_1
X_1557_ net53 VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__inv_2
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1488_ net74 net63 VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__and2_1
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2109_ _1147_ _0137_ _0146_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_52_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2460_ _0471_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__nand2_1
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2391_ net58 _1088_ net19 VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a21o_1
X_1411_ _0700_ _0701_ _0704_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__or4_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2589_ _0401_ _0562_ _0565_ net37 _0563_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__o221a_1
X_2727_ clknet_4_15_0_clk _0003_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_1609_ top8227.demux.state_machine.currentAddress\[12\] net35 _0861_ net26 VGND VGND
+ VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
Xfanout113 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
Xfanout102 net104 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_2
X_2658_ top8227.internalDataflow.addressLowBusModule.busInputs\[27\] _0580_ _0614_
+ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__a21o_1
Xfanout124 net126 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_4
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1891_ net65 _0735_ net112 _0689_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__o211a_1
X_1960_ _0764_ net62 _1232_ net60 VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__a211oi_1
XFILLER_52_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2443_ _0163_ _0408_ net19 _0164_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a2bb2o_1
X_2512_ net71 _0760_ _0768_ _0757_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a211o_1
X_2374_ _0370_ _0390_ _0369_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__o21a_1
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2090_ _0127_ _0129_ _1281_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1874_ net48 _1136_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__and3_4
X_1943_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\] _1214_ _1215_
+ top8227.internalDataflow.stackBusModule.busInputs\[47\] _1213_ VGND VGND VPWR VPWR
+ _1216_ sky130_fd_sc_hd__a221o_1
X_2426_ top8227.internalDataflow.addressHighBusModule.busInputs\[17\] top8227.internalDataflow.addressHighBusModule.busInputs\[16\]
+ net22 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2357_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] net20 VGND VGND
+ VPWR VPWR _0374_ sky130_fd_sc_hd__nor2_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2288_ _1267_ _0239_ _0325_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__nor4_1
XFILLER_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ net40 _0877_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__nand2_1
XFILLER_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2073_ top8227.internalDataflow.accRegToDB\[5\] _1212_ _1215_ top8227.internalDataflow.stackBusModule.busInputs\[45\]
+ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__a221o_1
X_2142_ _0663_ _1206_ _1205_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2211_ _1040_ _1075_ _1139_ _1195_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_28_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1926_ _0828_ _1198_ _0829_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__a21o_1
X_1857_ _1121_ _1124_ _1109_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__and3b_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1788_ _0701_ _0792_ net105 VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__o21a_1
X_2409_ _1314_ _1335_ _0127_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__and4_1
XFILLER_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
X_1642_ net132 _0664_ _0843_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__or3_1
XANTENNA_2 _0701_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2760_ clknet_4_3_0_clk _0036_ net115 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
X_1711_ net74 _0763_ net27 _0902_ _0919_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a32o_1
X_2691_ _0259_ _0293_ _0583_ _0284_ _0581_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__o221a_1
X_1573_ _0859_ _0860_ _0863_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__and3_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2125_ _1162_ _0163_ _0164_ _1160_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__a2bb2o_1
X_2056_ _1162_ _1326_ _1328_ _1160_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a2bb2oi_1
X_1909_ _1101_ _1179_ _1180_ _1181_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__or4_1
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2812_ clknet_4_5_0_clk _0088_ net123 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2743_ clknet_4_3_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ net116 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_16_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1556_ net2 net1 net54 VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__o21a_1
X_1625_ _0664_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__and2_2
X_2674_ _0131_ _0585_ _0627_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__o22a_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1487_ _0784_ _0787_ net96 VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__o21a_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2039_ top8227.internalDataflow.addressLowBusModule.busInputs\[31\] _1310_ _1311_
+ net8 VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__a22o_1
X_2108_ net25 _0147_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__nand2_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1410_ _0657_ net76 _0682_ net73 _0709_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a32o_1
X_2390_ _0228_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nand2_1
XFILLER_36_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2726_ clknet_4_12_0_clk _0002_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
X_2588_ _1314_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__xnor2_1
X_1608_ net180 net35 _0892_ net39 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a22o_1
Xfanout103 net104 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout114 net116 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
X_1539_ net104 net44 _0837_ net97 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a22o_1
X_2657_ _0291_ _0591_ _0613_ _0612_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o31a_1
XFILLER_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1890_ _0705_ net64 net68 net112 VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2442_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\] _0404_ VGND
+ VGND VPWR VPWR _0456_ sky130_fd_sc_hd__or2_1
X_2373_ _0373_ _0389_ _0372_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__o21a_1
X_2511_ net174 _1265_ _0512_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2709_ _0313_ _0652_ _0338_ net183 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_45_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1942_ _1194_ _1203_ _1174_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__nor3b_4
XFILLER_14_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1873_ _0790_ _1143_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__or3_1
X_2425_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] net20 VGND VGND
+ VPWR VPWR _0440_ sky130_fd_sc_hd__xor2_1
X_2356_ top8227.internalDataflow.addressLowBusModule.busInputs\[20\] net20 VGND VGND
+ VPWR VPWR _0373_ sky130_fd_sc_hd__and2_1
XFILLER_56_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2287_ _1332_ _0149_ _0173_ _0194_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or4_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2210_ net113 top8227.demux.state_machine.currentAddress\[1\] _1135_ VGND VGND VPWR
+ VPWR _0250_ sky130_fd_sc_hd__a21bo_1
X_2141_ net3 _1254_ _1256_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\]
+ _1262_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__a221o_1
X_2072_ top8227.internalDataflow.addressLowBusModule.busInputs\[37\] _1211_ _1214_
+ top8227.internalDataflow.addressLowBusModule.busInputs\[29\] VGND VGND VPWR VPWR
+ _1345_ sky130_fd_sc_hd__a22o_1
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1925_ top8227.demux.state_machine.currentAddress\[7\] top8227.demux.state_machine.currentAddress\[11\]
+ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__or2_1
X_1856_ top8227.internalDataflow.addressHighBusModule.busInputs\[23\] _1126_ _1128_
+ top8227.internalDataflow.accRegToDB\[7\] _1127_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a221o_1
X_1787_ net113 _0701_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__and2_1
X_2408_ _0153_ _0176_ _0420_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nor3_1
X_2339_ _1236_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold50 top8227.branchBackward VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1572_ _0858_ _0862_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__nor2_1
X_1641_ gpio[21] _0847_ _0858_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__and3_1
X_1710_ _0764_ net33 net26 _0928_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__a22o_1
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2690_ _0274_ _0296_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__xnor2_1
XANTENNA_3 _0782_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2124_ net4 _1254_ _1256_ top8227.internalDataflow.addressHighBusModule.busInputs\[19\]
+ _1262_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a221o_1
X_2055_ net7 _1255_ _1257_ top8227.internalDataflow.addressHighBusModule.busInputs\[22\]
+ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__o221a_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1839_ net61 _0827_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__nand2_1
X_1908_ net98 _0798_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__and2_1
XFILLER_57_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2811_ clknet_4_5_0_clk _0087_ net123 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2742_ clknet_4_2_0_clk top8227.internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ net116 VGND VGND VPWR VPWR top8227.PSRCurrentValue\[0\] sky130_fd_sc_hd__dfrtp_4
X_1555_ net2 net54 VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nand2_2
X_1624_ net7 _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_1
X_2673_ _0791_ _0133_ _0286_ _0584_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a31o_1
X_2107_ _0139_ _0145_ _1154_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_2
X_1486_ _0699_ _0716_ net72 VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__a21oi_2
X_2038_ _1286_ _1294_ _1296_ _1300_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__nor4_4
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2725_ clknet_4_14_0_clk _0001_ net129 VGND VGND VPWR VPWR top8227.demux.state_machine.currentAddress\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2656_ _0298_ _0599_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nor2_1
XFILLER_59_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2587_ _0417_ _0555_ _1335_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux2_1
Xfanout126 net127 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
X_1607_ net45 _0890_ _0891_ _0664_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__a22o_1
Xfanout115 net116 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__buf_2
X_1538_ top8227.demux.state_machine.timeState\[1\] net44 _0837_ net95 VGND VGND VPWR
+ VPWR _0014_ sky130_fd_sc_hd__a22o_1
Xfanout104 top8227.demux.state_machine.timeState\[2\] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_2
X_1469_ net75 net71 VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__and2_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2510_ net177 _1330_ _0512_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_1
X_2441_ _0453_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__xor2_1
X_2372_ _0376_ _0388_ _0375_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_19_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2708_ _0664_ top8227.internalDataflow.addressLowBusModule.busInputs\[23\] _0338_
+ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
X_2639_ top8227.internalDataflow.addressLowBusModule.busInputs\[25\] _0580_ _0593_
+ _0597_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__a22o_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1941_ _1174_ _1193_ _1203_ _1189_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__and4bb_2
X_1872_ _1140_ _1141_ _1142_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_16_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2424_ top8227.internalDataflow.addressHighBusModule.busInputs\[18\] net21 VGND VGND
+ VPWR VPWR _0439_ sky130_fd_sc_hd__nand2_1
X_2355_ _0370_ _0371_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__nor2_1
X_2286_ _0124_ _0220_ _0323_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or3b_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2140_ net25 _0171_ _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__and3_1
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2071_ _1343_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__inv_2
X_1855_ net42 _1109_ _1117_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nor3b_4
X_1924_ net106 _0773_ _1052_ _1195_ _1196_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__a2111o_1
X_1786_ net57 _0824_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__and2_1
X_2407_ _1313_ net21 _0422_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__or3_1
XFILLER_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2338_ _1232_ _1238_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__nor2_1
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2269_ _0133_ _0272_ _0303_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_64_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 top8227.demux.state_machine.currentAddress\[11\] VGND VGND VPWR VPWR net173
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold51 top8227.internalDataflow.accRegToDB\[6\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1571_ net3 net54 net4 VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__and3b_2
X_1640_ _0677_ net30 _0912_ _0919_ _0915_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__a221o_1
XANTENNA_4 top8227.demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2123_ _1210_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__nand2_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2054_ _1260_ _1261_ _1254_ _1256_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__a211o_1
XFILLER_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ net68 _0721_ net58 VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__a21o_1
X_1907_ net93 net75 net73 VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__and3_1
X_1769_ _0699_ _0703_ _0706_ _0676_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__a31oi_2
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2810_ clknet_4_5_0_clk _0086_ net124 VGND VGND VPWR VPWR top8227.internalDataflow.accRegToDB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2741_ clknet_4_10_0_clk _0025_ net121 VGND VGND VPWR VPWR top8227.demux.state_machine.currentInstruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2672_ _1331_ _0293_ _0587_ _0132_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a2bb2o_1
X_1554_ net2 net54 VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__and2_1
X_1623_ net132 net54 VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nand2_1
X_1485_ net72 _0716_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__nor2_1
.ends

