* NGSPICE file created from fpgacell.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt fpgacell CBeast_in[0] CBeast_in[10] CBeast_in[11] CBeast_in[12] CBeast_in[13]
+ CBeast_in[1] CBeast_in[2] CBeast_in[3] CBeast_in[4] CBeast_in[5] CBeast_in[6] CBeast_in[7]
+ CBeast_in[8] CBeast_in[9] CBeast_out[0] CBeast_out[10] CBeast_out[11] CBeast_out[12]
+ CBeast_out[13] CBeast_out[1] CBeast_out[2] CBeast_out[3] CBeast_out[4] CBeast_out[5]
+ CBeast_out[6] CBeast_out[7] CBeast_out[8] CBeast_out[9] CBnorth_in[0] CBnorth_in[10]
+ CBnorth_in[11] CBnorth_in[12] CBnorth_in[13] CBnorth_in[1] CBnorth_in[2] CBnorth_in[3]
+ CBnorth_in[4] CBnorth_in[5] CBnorth_in[6] CBnorth_in[7] CBnorth_in[8] CBnorth_in[9]
+ CBnorth_out[0] CBnorth_out[10] CBnorth_out[11] CBnorth_out[12] CBnorth_out[13] CBnorth_out[1]
+ CBnorth_out[2] CBnorth_out[3] CBnorth_out[4] CBnorth_out[5] CBnorth_out[6] CBnorth_out[7]
+ CBnorth_out[8] CBnorth_out[9] SBsouth_in[0] SBsouth_in[10] SBsouth_in[11] SBsouth_in[12]
+ SBsouth_in[13] SBsouth_in[1] SBsouth_in[2] SBsouth_in[3] SBsouth_in[4] SBsouth_in[5]
+ SBsouth_in[6] SBsouth_in[7] SBsouth_in[8] SBsouth_in[9] SBsouth_out[0] SBsouth_out[10]
+ SBsouth_out[11] SBsouth_out[12] SBsouth_out[13] SBsouth_out[1] SBsouth_out[2] SBsouth_out[3]
+ SBsouth_out[4] SBsouth_out[5] SBsouth_out[6] SBsouth_out[7] SBsouth_out[8] SBsouth_out[9]
+ SBwest_in[0] SBwest_in[10] SBwest_in[11] SBwest_in[12] SBwest_in[13] SBwest_in[1]
+ SBwest_in[2] SBwest_in[3] SBwest_in[4] SBwest_in[5] SBwest_in[6] SBwest_in[7] SBwest_in[8]
+ SBwest_in[9] SBwest_out[0] SBwest_out[10] SBwest_out[11] SBwest_out[12] SBwest_out[13]
+ SBwest_out[1] SBwest_out[2] SBwest_out[3] SBwest_out[4] SBwest_out[5] SBwest_out[6]
+ SBwest_out[7] SBwest_out[8] SBwest_out[9] clk config_data_in config_data_out config_en
+ le_clk le_en le_nrst nrst vccd1 vssd1
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2037_ CB_1.config_dataA\[1\] CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0822_
+ sky130_fd_sc_hd__nand2_1
X_2106_ _0879_ _0889_ _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__o21a_1
X_2939_ clknet_leaf_27_clk _0201_ net209 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[65\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1606_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] CB_0.config_dataA\[19\] CB_0.config_dataA\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__or4_1
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2724_ net286 LE_1B.config_data\[5\] net257 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__mux2_1
X_2655_ SB0.route_sel\[109\] SB0.route_sel\[108\] net251 vssd1 vssd1 vccd1 vccd1 _0245_
+ sky130_fd_sc_hd__mux2_1
Xfanout149 CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
Xfanout127 _1219_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_2
X_1399_ CB_0.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__inv_2
X_1537_ _1325_ _1326_ _1329_ CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 _1331_
+ sky130_fd_sc_hd__o31a_1
Xfanout138 CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
X_2586_ SB0.route_sel\[40\] SB0.route_sel\[39\] net231 vssd1 vssd1 vccd1 vccd1 _0176_
+ sky130_fd_sc_hd__mux2_1
X_1468_ SB0.route_sel\[58\] SB0.route_sel\[59\] vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__nor2_1
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2440_ net373 net370 net268 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__mux2_1
X_2371_ _1099_ _1100_ _0428_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__o21a_1
X_2707_ CB_1.config_dataA\[9\] net141 net265 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__mux2_1
X_2638_ SB0.route_sel\[92\] SB0.route_sel\[91\] net246 vssd1 vssd1 vccd1 vccd1 _0228_
+ sky130_fd_sc_hd__mux2_1
X_2569_ SB0.route_sel\[23\] SB0.route_sel\[22\] net227 vssd1 vssd1 vccd1 vccd1 _0159_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1871_ net132 net127 net123 net120 LEI0.config_data\[3\] LEI0.config_data\[4\] vssd1
+ vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__mux4_1
X_1940_ net154 net156 net153 _0492_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_16_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2423_ LEI0.config_data\[14\] LEI0.config_data\[13\] net267 vssd1 vssd1 vccd1 vccd1
+ _0015_ sky130_fd_sc_hd__mux2_1
X_2285_ _1299_ _1307_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__nand2_1
X_2354_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__and2b_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2070_ net132 net127 net123 net120 LEI0.config_data\[30\] LEI0.config_data\[31\]
+ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__mux4_1
X_2972_ clknet_leaf_10_clk _0234_ net203 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[98\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1785_ _0453_ _0473_ _0517_ _0492_ CB_0.config_dataA\[8\] net166 vssd1 vssd1 vccd1
+ vccd1 _0574_ sky130_fd_sc_hd__mux4_1
X_1923_ net23 net24 net25 net26 net155 net154 vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__mux4_1
X_1854_ _0636_ _0637_ _0640_ _0627_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__o31a_1
X_2406_ SB0.route_sel\[81\] _1174_ _1172_ _1173_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__a2bb2o_1
X_2268_ _1310_ _1040_ _1314_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__o21ai_1
X_2199_ _1218_ _1219_ net123 _1221_ LEI0.config_data\[33\] LEI0.config_data\[34\]
+ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__mux4_1
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2337_ SB0.route_sel\[57\] SB0.route_sel\[56\] SB0.route_sel\[58\] _1156_ vssd1 vssd1
+ vccd1 vccd1 _1078_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_27_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold30 LEI0.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 LE_0A.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 LE_0A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 LE_0A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 LE_0B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 LEI0.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 LEI0.config_data\[26\] vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_41_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1570_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] CB_0.config_dataA\[17\] CB_0.config_dataA\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__or4bb_1
XANTENNA_5 LEI0.config_data\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2053_ net4 net5 CB_1.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__mux2_1
X_2122_ _0906_ _0899_ _0895_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ clknet_leaf_2_clk _0217_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[81\]
+ sky130_fd_sc_hd__dfstp_1
X_1906_ net15 net20 net21 net22 net157 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _0693_ sky130_fd_sc_hd__mux4_1
X_1768_ _1192_ net167 vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
X_1837_ CB_0.config_dataB\[7\] _0622_ _0623_ _0620_ vssd1 vssd1 vccd1 vccd1 _0624_
+ sky130_fd_sc_hd__o22ai_1
X_2886_ clknet_leaf_29_clk _0148_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_1699_ _0483_ _0486_ _0487_ SB0.route_sel\[89\] SB0.route_sel\[88\] vssd1 vssd1 vccd1
+ vccd1 _0488_ sky130_fd_sc_hd__o311a_1
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 CBeast_out[10] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 CBeast_out[8] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 CBnorth_out[5] sky130_fd_sc_hd__buf_2
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 SBsouth_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2671_ CB_0.config_dataA\[13\] CB_0.config_dataA\[12\] net248 vssd1 vssd1 vccd1 vccd1
+ _0261_ sky130_fd_sc_hd__mux2_1
X_2740_ clknet_leaf_16_clk _0002_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1622_ SB0.route_sel\[3\] SB0.route_sel\[2\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__nor2_1
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1553_ _0338_ _0340_ _0341_ _0329_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__a31oi_1
X_1484_ net123 _1273_ _1275_ _1276_ _1277_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__o221ai_4
X_2036_ _0469_ _0791_ _1203_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__a21o_1
X_2105_ CB_1.config_dataA\[15\] _0887_ _0888_ _0873_ vssd1 vssd1 vccd1 vccd1 _0890_
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2938_ clknet_leaf_27_clk _0200_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[64\]
+ sky130_fd_sc_hd__dfstp_1
X_2869_ clknet_leaf_21_clk _0131_ net215 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2723_ net310 LE_1B.config_data\[4\] net252 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__mux2_1
X_1536_ _1325_ _1326_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__or3_4
X_1605_ SB0.route_sel\[0\] SB0.route_sel\[1\] vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__nand2_1
X_2654_ SB0.route_sel\[108\] SB0.route_sel\[107\] net251 vssd1 vssd1 vccd1 vccd1 _0244_
+ sky130_fd_sc_hd__mux2_1
X_2585_ SB0.route_sel\[39\] SB0.route_sel\[38\] net232 vssd1 vssd1 vccd1 vccd1 _0175_
+ sky130_fd_sc_hd__mux2_1
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_2
X_1398_ net166 vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__inv_2
Xfanout139 CB_1.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_1467_ _1256_ _1260_ _1246_ _1250_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2019_ _0514_ _0803_ vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__and2_2
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2370_ _1136_ SB0.route_sel\[18\] SB0.route_sel\[23\] SB0.route_sel\[22\] vssd1 vssd1
+ vccd1 vccd1 _1100_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_19_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2706_ net141 CB_1.config_dataA\[7\] net265 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__mux2_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1519_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__inv_2
X_2637_ SB0.route_sel\[91\] SB0.route_sel\[90\] net246 vssd1 vssd1 vccd1 vccd1 _0227_
+ sky130_fd_sc_hd__mux2_1
X_2568_ SB0.route_sel\[22\] SB0.route_sel\[21\] net227 vssd1 vssd1 vccd1 vccd1 _0158_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2499_ LE_0B.edge_mode LE_0B.config_data\[16\] net231 vssd1 vssd1 vccd1 vccd1 _0090_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ _0648_ _0653_ _0655_ _0656_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1
+ _0657_ sky130_fd_sc_hd__o311ai_4
XFILLER_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2422_ LEI0.config_data\[13\] LEI0.config_data\[12\] net267 vssd1 vssd1 vccd1 vccd1
+ _0014_ sky130_fd_sc_hd__mux2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2353_ _1282_ _1088_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__nor2_1
X_2284_ net136 _1048_ _1270_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__mux2_1
X_1999_ _0782_ _0783_ _0410_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__a21bo_2
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1922_ net155 _0346_ _0706_ _0708_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__o211a_1
XFILLER_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ clknet_leaf_11_clk _0233_ net203 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[97\]
+ sky130_fd_sc_hd__dfstp_1
X_1784_ net15 net20 net21 net22 net167 net166 vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__mux4_1
X_1853_ CB_0.config_dataB\[7\] _0628_ _0630_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_
+ sky130_fd_sc_hd__o211a_1
X_2336_ SB0.route_sel\[60\] _1157_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nor2_1
X_2405_ SB0.route_sel\[82\] _1170_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nor2_1
X_2267_ _1330_ net127 _1311_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__mux2_1
X_2198_ net180 _1214_ CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_27_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 _0008_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 _0013_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 _0062_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 LE_0A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 LEI0.config_data\[22\] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 LE_1B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 LE_1A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 LE_0B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 LEI0.config_data\[31\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2052_ net9 net10 net11 net12 net144 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0837_ sky130_fd_sc_hd__mux4_1
X_2121_ _0904_ _0905_ _0868_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__mux2_1
X_1905_ CB_0.config_dataB\[9\] net157 CB_0.config_dataB\[11\] _0492_ vssd1 vssd1 vccd1
+ vccd1 _0692_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_32_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2885_ clknet_leaf_28_clk _0147_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_2954_ clknet_leaf_3_clk _0216_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[80\]
+ sky130_fd_sc_hd__dfstp_1
X_1767_ LE_0A.config_data\[7\] LE_0A.config_data\[6\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0556_ sky130_fd_sc_hd__mux2_1
X_1836_ net18 net19 net159 vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__mux2_1
X_1698_ SB0.route_sel\[92\] SB0.route_sel\[93\] net31 vssd1 vssd1 vccd1 vccd1 _0487_
+ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2319_ _0420_ _1066_ _0422_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__a21o_1
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 CBnorth_out[6] sky130_fd_sc_hd__buf_2
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 CBeast_out[11] sky130_fd_sc_hd__buf_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 SBsouth_out[3] sky130_fd_sc_hd__buf_2
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 CBeast_out[9] sky130_fd_sc_hd__buf_2
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2670_ net165 CB_0.config_dataA\[11\] net248 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__mux2_1
X_1552_ SB0.route_sel\[100\] SB0.route_sel\[101\] net32 vssd1 vssd1 vccd1 vccd1 _0341_
+ sky130_fd_sc_hd__a21bo_1
X_1621_ _0405_ _0409_ _0394_ _0400_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__a2bb2o_2
X_2104_ net2 net3 net139 vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__mux2_1
X_1483_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__nand2_2
X_2035_ CB_1.config_dataA\[1\] CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0820_
+ sky130_fd_sc_hd__nand2b_1
X_2937_ clknet_leaf_28_clk _0199_ net193 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[63\]
+ sky130_fd_sc_hd__dfstp_1
X_2868_ clknet_leaf_21_clk _0130_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2799_ clknet_leaf_6_clk net300 net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_1819_ LE_0A.config_data\[15\] LE_0A.config_data\[14\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0608_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_37_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2722_ net315 net294 net251 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__mux2_1
Xfanout129 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_1
X_1604_ _0391_ _0392_ _0390_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__a21bo_2
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2653_ SB0.route_sel\[107\] SB0.route_sel\[106\] net253 vssd1 vssd1 vccd1 vccd1 _0243_
+ sky130_fd_sc_hd__mux2_1
X_1535_ SB0.route_sel\[106\] SB0.route_sel\[107\] _1187_ SB0.route_sel\[109\] _1328_
+ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__o221a_1
X_2584_ SB0.route_sel\[38\] SB0.route_sel\[37\] net232 vssd1 vssd1 vccd1 vccd1 _0174_
+ sky130_fd_sc_hd__mux2_1
X_1397_ LEI0.config_data\[26\] vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__inv_2
XFILLER_27_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1466_ SB0.route_sel\[58\] SB0.route_sel\[59\] _1258_ _1259_ _1246_ vssd1 vssd1 vccd1
+ vccd1 _1260_ sky130_fd_sc_hd__a41o_1
X_2018_ _1172_ SB0.route_sel\[86\] SB0.route_sel\[81\] _1174_ _0802_ vssd1 vssd1 vccd1
+ vccd1 _0803_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2705_ CB_1.config_dataA\[7\] CB_1.config_dataA\[6\] net265 vssd1 vssd1 vccd1 vccd1
+ _0295_ sky130_fd_sc_hd__mux2_1
X_2636_ SB0.route_sel\[90\] SB0.route_sel\[89\] net246 vssd1 vssd1 vccd1 vccd1 _0226_
+ sky130_fd_sc_hd__mux2_1
X_1518_ net19 net131 _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__mux2_1
X_2567_ SB0.route_sel\[21\] SB0.route_sel\[20\] net229 vssd1 vssd1 vccd1 vccd1 _0157_
+ sky130_fd_sc_hd__mux2_1
X_1449_ SB0.route_sel\[52\] _1153_ SB0.route_sel\[55\] _1154_ _1242_ vssd1 vssd1 vccd1
+ vccd1 _1243_ sky130_fd_sc_hd__a221o_1
X_2498_ LE_0B.config_data\[16\] net333 net233 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2421_ LEI0.config_data\[12\] net301 net267 vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__mux2_1
X_2283_ _1286_ net128 _1267_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__mux2_1
X_2352_ _1148_ SB0.route_sel\[42\] SB0.route_sel\[47\] SB0.route_sel\[46\] _1087_
+ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_24_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1998_ SB0.route_sel\[4\] SB0.route_sel\[5\] SB0.route_sel\[7\] _1129_ vssd1 vssd1
+ vccd1 vccd1 _0783_ sky130_fd_sc_hd__o22a_1
X_2619_ SB0.route_sel\[73\] SB0.route_sel\[72\] net238 vssd1 vssd1 vccd1 vccd1 _0209_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1921_ net155 _1330_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__nand2_1
X_1852_ CB_0.config_dataB\[5\] CB_0.config_dataB\[7\] _0638_ _0635_ CB_0.config_dataB\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__a311oi_1
X_2970_ clknet_leaf_11_clk _0232_ net203 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[96\]
+ sky130_fd_sc_hd__dfstp_1
X_1783_ _1192_ _0569_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__a21oi_1
X_2404_ _1121_ _1122_ _0514_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__o21a_1
X_2266_ net59 LE_1B.edge_mode vssd1 vssd1 vccd1 vccd1 LE_1B.sel_clk sky130_fd_sc_hd__xnor2_1
X_2335_ _1075_ _1076_ _0450_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__o21a_1
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2197_ _0973_ _0975_ _0977_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__a22o_1
Xhold98 LEI0.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 LE_0A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 LEI0.config_data\[25\] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _0064_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _0024_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 LE_0B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 LE_0B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold32 LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0109_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 LE_1B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2120_ _0903_ _0902_ _0814_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__mux2_1
X_2051_ _0343_ _0762_ net144 vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1904_ net157 _0472_ _0677_ _0690_ vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__a211o_1
X_1835_ net23 net24 net25 net26 net159 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1
+ _0622_ sky130_fd_sc_hd__mux4_1
X_2884_ clknet_leaf_29_clk _0146_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_2953_ clknet_leaf_3_clk _0215_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[79\]
+ sky130_fd_sc_hd__dfstp_1
X_1766_ _0551_ _0552_ _0554_ _0539_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__a31oi_4
X_1697_ _1177_ _1178_ net45 SB0.route_sel\[93\] SB0.route_sel\[92\] vssd1 vssd1 vccd1
+ vccd1 _0486_ sky130_fd_sc_hd__o2111a_1
X_2318_ _0419_ _0787_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__nand2_1
X_2249_ _0936_ LE_1B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__and2b_1
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 CBnorth_out[0] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 CBnorth_out[7] sky130_fd_sc_hd__buf_2
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 CBeast_out[12] sky130_fd_sc_hd__buf_2
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 SBsouth_out[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1551_ _1182_ _1183_ net46 SB0.route_sel\[101\] SB0.route_sel\[100\] vssd1 vssd1
+ vccd1 vccd1 _0340_ sky130_fd_sc_hd__o2111ai_1
X_1620_ SB0.route_sel\[3\] SB0.route_sel\[2\] _0407_ _0408_ _0394_ vssd1 vssd1 vccd1
+ vccd1 _0409_ sky130_fd_sc_hd__a41o_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1482_ net10 _1274_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__and2b_1
X_2103_ net13 net14 net139 vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__mux2_1
X_2034_ CB_1.config_dataA\[1\] CB_1.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0819_
+ sky130_fd_sc_hd__and2b_1
XFILLER_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1818_ _0606_ _0581_ _0579_ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__mux2_1
X_2798_ clknet_leaf_6_clk _0060_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2936_ clknet_leaf_28_clk _0198_ net193 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[62\]
+ sky130_fd_sc_hd__dfstp_1
X_2867_ clknet_leaf_21_clk _0129_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_2
X_1749_ net132 net127 net123 net120 LEI0.config_data\[12\] LEI0.config_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_51_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2721_ net294 LE_1B.config_data\[2\] net251 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__mux2_1
X_2652_ SB0.route_sel\[106\] SB0.route_sel\[105\] net253 vssd1 vssd1 vccd1 vccd1 _0242_
+ sky130_fd_sc_hd__mux2_1
X_1603_ SB0.route_sel\[11\] SB0.route_sel\[10\] _1132_ SB0.route_sel\[13\] vssd1 vssd1
+ vccd1 vccd1 _0392_ sky130_fd_sc_hd__o22a_1
X_1465_ SB0.route_sel\[60\] SB0.route_sel\[61\] net40 vssd1 vssd1 vccd1 vccd1 _1259_
+ sky130_fd_sc_hd__a21bo_1
X_1534_ SB0.route_sel\[110\] net119 vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__nand2b_1
X_2583_ SB0.route_sel\[37\] SB0.route_sel\[36\] net232 vssd1 vssd1 vccd1 vccd1 _0173_
+ sky130_fd_sc_hd__mux2_1
X_1396_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__inv_2
X_2017_ SB0.route_sel\[84\] SB0.route_sel\[85\] vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__nor2_1
X_2919_ clknet_leaf_31_clk _0181_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[45\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2704_ CB_1.config_dataA\[6\] CB_1.config_dataA\[5\] net265 vssd1 vssd1 vccd1 vccd1
+ _0294_ sky130_fd_sc_hd__mux2_1
X_2635_ SB0.route_sel\[89\] SB0.route_sel\[88\] net246 vssd1 vssd1 vccd1 vccd1 _0225_
+ sky130_fd_sc_hd__mux2_1
X_1517_ net150 net152 net146 net148 vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__and4b_1
XFILLER_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2566_ SB0.route_sel\[20\] SB0.route_sel\[19\] net229 vssd1 vssd1 vccd1 vccd1 _0156_
+ sky130_fd_sc_hd__mux2_1
X_1448_ SB0.route_sel\[51\] SB0.route_sel\[50\] vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__nor2_1
X_2497_ net333 net306 net231 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__mux2_1
X_1379_ SB0.route_sel\[86\] vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__inv_2
X_3049_ clknet_leaf_24_clk net295 net206 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2420_ net301 net316 net267 vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2282_ net133 _1047_ _1228_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__mux2_1
X_2351_ SB0.route_sel\[41\] SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__nand2b_1
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1997_ SB0.route_sel\[0\] _1130_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__or2_1
X_2549_ SB0.route_sel\[3\] SB0.route_sel\[2\] net250 vssd1 vssd1 vccd1 vccd1 _0139_
+ sky130_fd_sc_hd__mux2_1
X_2618_ SB0.route_sel\[72\] SB0.route_sel\[71\] net237 vssd1 vssd1 vccd1 vccd1 _0208_
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1920_ net154 net153 vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__nand2b_1
X_1851_ _0517_ _0492_ net160 vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__mux2_1
X_1782_ _0431_ _0557_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__a21o_1
X_2403_ SB0.route_sel\[81\] SB0.route_sel\[80\] SB0.route_sel\[82\] _1170_ vssd1 vssd1
+ vccd1 vccd1 _1122_ sky130_fd_sc_hd__a2bb2o_1
X_2196_ CB_1.config_dataB\[9\] _1214_ _0978_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or3_1
X_2265_ net184 LE_1B.reset_mode vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__xor2_2
X_2334_ _1159_ SB0.route_sel\[66\] _1161_ _1162_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold22 _0083_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 LE_1B.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 LEI0.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 _0026_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 LE_0A.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold99 LEI0.config_data\[30\] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold33 _0317_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 LE_1B.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 LE_1B.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ _1325_ _1326_ _0767_ net144 vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__o31a_1
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2952_ clknet_leaf_3_clk _0214_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[78\]
+ sky130_fd_sc_hd__dfstp_1
X_1765_ _0536_ _0537_ _0553_ _0532_ CB_0.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1
+ _0554_ sky130_fd_sc_hd__o311ai_4
X_1903_ net157 _0453_ vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1834_ net159 _1330_ _0619_ _0620_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__a211o_1
X_2883_ clknet_leaf_29_clk _0145_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_1696_ _0481_ _0482_ _0483_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__o211ai_1
X_2179_ net181 _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__o21a_1
X_2248_ LE_1B.config_data\[7\] LE_1B.config_data\[6\] _0936_ vssd1 vssd1 vccd1 vccd1
+ _1031_ sky130_fd_sc_hd__mux2_1
X_2317_ net124 _1251_ _0361_ _1065_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__a31o_1
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 CBnorth_out[10] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 CBnorth_out[8] sky130_fd_sc_hd__buf_2
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 CBeast_out[13] sky130_fd_sc_hd__buf_2
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1550_ _0334_ _0336_ _0337_ _0338_ vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__a211o_1
X_1481_ net121 _1274_ _1272_ net137 vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__a2bb2o_1
X_2033_ _0450_ _0795_ net144 vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__a21o_1
X_2102_ net1 net6 net7 net8 net139 CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1
+ _0887_ sky130_fd_sc_hd__mux4_1
X_2935_ clknet_leaf_28_clk _0197_ net193 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[61\]
+ sky130_fd_sc_hd__dfstp_1
X_1748_ _1244_ _0523_ _0526_ _1264_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__a22o_1
X_1817_ _0604_ _0605_ _0555_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__mux2_1
X_2797_ clknet_leaf_6_clk _0059_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2866_ clknet_leaf_21_clk _0128_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_2
X_1679_ SB0.route_sel\[74\] SB0.route_sel\[75\] _0466_ _0467_ _0455_ vssd1 vssd1 vccd1
+ vccd1 _0468_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_51_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1602_ SB0.route_sel\[15\] _1133_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__nand2_1
X_2720_ LE_1B.config_data\[2\] net276 net251 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__mux2_1
X_2651_ SB0.route_sel\[105\] SB0.route_sel\[104\] net253 vssd1 vssd1 vccd1 vccd1 _0241_
+ sky130_fd_sc_hd__mux2_1
X_2582_ SB0.route_sel\[36\] SB0.route_sel\[35\] net232 vssd1 vssd1 vccd1 vccd1 _0172_
+ sky130_fd_sc_hd__mux2_1
X_1395_ CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__inv_2
X_1464_ SB0.route_sel\[63\] SB0.route_sel\[62\] _1257_ vssd1 vssd1 vccd1 vccd1 _1258_
+ sky130_fd_sc_hd__a21bo_1
X_1533_ _1325_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__or2_1
X_2016_ _0489_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__and2_2
X_3065_ clknet_leaf_31_clk _0327_ net184 vssd1 vssd1 vccd1 vccd1 LE_1B.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_30_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2918_ clknet_leaf_31_clk _0180_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[44\]
+ sky130_fd_sc_hd__dfstp_1
X_2849_ clknet_leaf_22_clk _0111_ net212 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1516_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1269_ vssd1 vssd1 vccd1 vccd1
+ _1310_ sky130_fd_sc_hd__and3_1
X_2703_ CB_1.config_dataA\[5\] net143 net265 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__mux2_1
X_2634_ SB0.route_sel\[88\] SB0.route_sel\[87\] net246 vssd1 vssd1 vccd1 vccd1 _0224_
+ sky130_fd_sc_hd__mux2_1
X_2565_ SB0.route_sel\[19\] SB0.route_sel\[18\] net229 vssd1 vssd1 vccd1 vccd1 _0155_
+ sky130_fd_sc_hd__mux2_1
X_1378_ SB0.route_sel\[87\] vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1447_ _1236_ _1240_ _1223_ _1229_ vssd1 vssd1 vccd1 vccd1 _1241_ sky130_fd_sc_hd__a2bb2o_1
X_2496_ net306 net291 net231 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__mux2_1
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3048_ clknet_leaf_24_clk net277 net206 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2281_ _1245_ net128 _1224_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__mux2_1
X_2350_ _1282_ _1086_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1996_ _0779_ _0780_ _0390_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__a21bo_2
X_2548_ SB0.route_sel\[2\] SB0.route_sel\[1\] net250 vssd1 vssd1 vccd1 vccd1 _0138_
+ sky130_fd_sc_hd__mux2_1
X_2617_ SB0.route_sel\[71\] SB0.route_sel\[70\] net237 vssd1 vssd1 vccd1 vccd1 _0207_
+ sky130_fd_sc_hd__mux2_1
X_2479_ LE_0A.reset_mode LE_0A.reset_val net227 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__mux2_1
XFILLER_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
Xfanout270 net271 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ CB_0.config_dataA\[9\] net167 _0374_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__and3_1
X_1850_ CB_0.config_dataB\[7\] _0618_ _0621_ _0624_ CB_0.config_dataB\[6\] vssd1 vssd1
+ vccd1 vccd1 _0637_ sky130_fd_sc_hd__o2111a_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2402_ SB0.route_sel\[84\] _1171_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__nor2_1
X_2333_ SB0.route_sel\[65\] _1164_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__nor2_1
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2264_ net59 LE_1A.edge_mode vssd1 vssd1 vccd1 vccd1 LE_1A.sel_clk sky130_fd_sc_hd__xnor2_1
X_2195_ net4 net5 net180 vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__mux2_1
X_1979_ _0343_ _0762_ net143 vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__a21oi_1
Xhold45 LEI0.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 LE_0A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 _0315_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 LE_1B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 LE_1A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 LE_0A.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold89 LE_1B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 LE_0B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _0317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1902_ CB_0.config_dataB\[11\] _0688_ vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__or2_1
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2951_ clknet_leaf_3_clk _0213_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[77\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_19_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1764_ _0533_ _0534_ _1190_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a21oi_1
X_1833_ CB_0.config_dataB\[5\] CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0620_
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_40_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2882_ clknet_leaf_29_clk _0144_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_1695_ net125 _1251_ _0440_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__nand3_1
X_2316_ _0362_ _0778_ _0363_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__a21oi_1
X_2178_ net3 _0943_ _0945_ net2 CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0961_
+ sky130_fd_sc_hd__o221a_1
X_2247_ _0998_ _1000_ _1024_ _1029_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a211o_1
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 CBnorth_out[11] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 CBeast_out[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1480_ net175 net171 net173 net177 vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__or4bb_1
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2032_ _0781_ _0784_ _0778_ _0787_ _1203_ CB_1.config_dataA\[1\] vssd1 vssd1 vccd1
+ vccd1 _0817_ sky130_fd_sc_hd__mux4_1
X_2101_ CB_1.config_dataA\[13\] net138 CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1
+ _0886_ sky130_fd_sc_hd__and3_1
X_2934_ clknet_leaf_25_clk _0196_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[60\]
+ sky130_fd_sc_hd__dfstp_1
X_2865_ clknet_leaf_21_clk _0127_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_1747_ _1189_ _1190_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__and3_1
X_1816_ LE_0A.config_data\[1\] LE_0A.config_data\[0\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0605_ sky130_fd_sc_hd__mux2_1
X_2796_ clknet_leaf_6_clk _0058_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1678_ SB0.route_sel\[76\] SB0.route_sel\[77\] net42 vssd1 vssd1 vccd1 vccd1 _0467_
+ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2650_ SB0.route_sel\[104\] SB0.route_sel\[103\] net253 vssd1 vssd1 vccd1 vccd1 _0240_
+ sky130_fd_sc_hd__mux2_1
X_1601_ _0376_ _0380_ _0385_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__a22o_1
X_2581_ SB0.route_sel\[35\] SB0.route_sel\[34\] net237 vssd1 vssd1 vccd1 vccd1 _0171_
+ sky130_fd_sc_hd__mux2_1
X_1532_ _1320_ _1324_ _1309_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__a21oi_2
X_1463_ SB0.route_sel\[60\] SB0.route_sel\[61\] net54 vssd1 vssd1 vccd1 vccd1 _1257_
+ sky130_fd_sc_hd__and3_1
X_1394_ SB0.route_sel\[105\] vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__inv_2
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2015_ _1177_ SB0.route_sel\[94\] _1179_ SB0.route_sel\[89\] _0799_ vssd1 vssd1 vccd1
+ vccd1 _0800_ sky130_fd_sc_hd__a221o_1
X_3064_ clknet_leaf_25_clk _0326_ net206 vssd1 vssd1 vccd1 vccd1 LE_1B.reset_val sky130_fd_sc_hd__dfrtp_2
X_2917_ clknet_leaf_31_clk _0179_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[43\]
+ sky130_fd_sc_hd__dfstp_1
X_2848_ clknet_leaf_22_clk net280 net212 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2779_ clknet_leaf_11_clk net366 net219 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2702_ net143 CB_1.config_dataA\[3\] net264 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__mux2_1
X_2633_ SB0.route_sel\[87\] SB0.route_sel\[86\] net233 vssd1 vssd1 vccd1 vccd1 _0223_
+ sky130_fd_sc_hd__mux2_1
X_2564_ SB0.route_sel\[18\] SB0.route_sel\[17\] net229 vssd1 vssd1 vccd1 vccd1 _0154_
+ sky130_fd_sc_hd__mux2_1
X_1515_ SB0.route_sel\[104\] SB0.route_sel\[105\] vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nand2_1
X_2495_ net291 net272 net232 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__mux2_1
X_1377_ SB0.route_sel\[85\] vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__inv_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1446_ SB0.route_sel\[51\] SB0.route_sel\[50\] _1238_ _1239_ _1223_ vssd1 vssd1 vccd1
+ vccd1 _1240_ sky130_fd_sc_hd__a41o_1
X_3047_ clknet_leaf_25_clk _0309_ net206 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2280_ _1046_ net133 _1249_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__mux2_1
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ SB0.route_sel\[12\] SB0.route_sel\[13\] SB0.route_sel\[15\] _1133_ vssd1 vssd1
+ vccd1 vccd1 _0780_ sky130_fd_sc_hd__o22a_1
X_2616_ SB0.route_sel\[70\] SB0.route_sel\[69\] net237 vssd1 vssd1 vccd1 vccd1 _0206_
+ sky130_fd_sc_hd__mux2_1
X_2547_ SB0.route_sel\[1\] SB0.route_sel\[0\] net250 vssd1 vssd1 vccd1 vccd1 _0137_
+ sky130_fd_sc_hd__mux2_1
X_1429_ SB0.route_sel\[49\] SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__nand2_1
X_2478_ LE_0A.reset_val LE_0A.edge_mode net231 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload1 clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout271 net58 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout260 net264 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1780_ _0413_ _0393_ net167 vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__mux2_1
X_2401_ _1119_ _1120_ _0489_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__o21a_1
X_2332_ _1073_ _1074_ _0450_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__o21a_1
X_2263_ net210 LE_1A.reset_mode vssd1 vssd1 vccd1 vccd1 _2263_/X sky130_fd_sc_hd__xor2_2
X_2194_ CB_1.config_dataB\[11\] _0976_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__or2_1
X_1978_ _0343_ _0762_ vssd1 vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__and2_1
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold68 _0055_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 LE_0A.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 LE_0A.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 LE_0B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 LE_1B.config_data\[14\] vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _0311_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _0074_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1901_ _0413_ _0431_ _0393_ _0374_ CB_0.config_dataB\[9\] net158 vssd1 vssd1 vccd1
+ vccd1 _0688_ sky130_fd_sc_hd__mux4_1
X_1832_ net159 _0346_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__nor2_1
X_2950_ clknet_leaf_4_clk _0212_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[76\]
+ sky130_fd_sc_hd__dfstp_1
X_2881_ clknet_leaf_29_clk _0143_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_1763_ _1189_ _1190_ net168 CB_0.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 _0552_
+ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_40_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1694_ SB0.route_sel\[90\] SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__nand2_1
X_2246_ _0966_ _1026_ _1027_ _1028_ _0997_ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__o221a_1
X_2315_ _1289_ _1064_ _1291_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__a21o_1
X_2177_ net13 net14 net182 vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__mux2_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 CBeast_out[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2100_ net138 _0793_ _0873_ _0884_ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__a211o_1
X_2031_ _0815_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__inv_2
XFILLER_22_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1815_ LE_0A.config_data\[3\] LE_0A.config_data\[2\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0604_ sky130_fd_sc_hd__mux2_1
X_2795_ clknet_leaf_7_clk _0057_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2933_ clknet_leaf_26_clk _0195_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[59\]
+ sky130_fd_sc_hd__dfstp_1
X_2864_ clknet_leaf_20_clk _0126_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_1746_ _1307_ _1285_ net168 vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1677_ _1167_ _1168_ net56 SB0.route_sel\[77\] SB0.route_sel\[76\] vssd1 vssd1 vccd1
+ vccd1 _0466_ sky130_fd_sc_hd__o2111ai_1
X_2229_ _0792_ _0796_ _0801_ _0804_ _1215_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1
+ vccd1 _1012_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_51_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1531_ _1310_ _1313_ _1314_ _1309_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__o211a_2
X_1600_ SB0.route_sel\[11\] SB0.route_sel\[10\] _0388_ _0376_ vssd1 vssd1 vccd1 vccd1
+ _0389_ sky130_fd_sc_hd__a31oi_1
X_1462_ _1253_ _1254_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__a21oi_1
X_2580_ SB0.route_sel\[34\] SB0.route_sel\[33\] net232 vssd1 vssd1 vccd1 vccd1 _0170_
+ sky130_fd_sc_hd__mux2_1
X_3063_ clknet_leaf_25_clk _0325_ net208 vssd1 vssd1 vccd1 vccd1 LE_1B.edge_mode sky130_fd_sc_hd__dfstp_1
X_1393_ SB0.route_sel\[108\] vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__inv_2
X_2014_ SB0.route_sel\[92\] SB0.route_sel\[93\] vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nor2_1
X_2778_ clknet_leaf_12_clk _0040_ net219 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_2916_ clknet_leaf_31_clk _0178_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[42\]
+ sky130_fd_sc_hd__dfstp_1
X_2847_ clknet_leaf_22_clk net336 net214 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold110 LE_1A.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _0514_ _0516_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ CB_1.config_dataA\[3\] CB_1.config_dataA\[2\] net264 vssd1 vssd1 vccd1 vccd1
+ _0291_ sky130_fd_sc_hd__mux2_1
X_2632_ SB0.route_sel\[86\] SB0.route_sel\[85\] net233 vssd1 vssd1 vccd1 vccd1 _0222_
+ sky130_fd_sc_hd__mux2_1
X_1514_ _1307_ _1285_ _1244_ _1264_ net170 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1
+ vccd1 _1308_ sky130_fd_sc_hd__mux4_1
X_2494_ net272 LE_0B.config_data\[11\] net232 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__mux2_1
X_2563_ SB0.route_sel\[17\] SB0.route_sel\[16\] net229 vssd1 vssd1 vccd1 vccd1 _0153_
+ sky130_fd_sc_hd__mux2_1
X_1445_ SB0.route_sel\[52\] SB0.route_sel\[53\] net39 vssd1 vssd1 vccd1 vccd1 _1239_
+ sky130_fd_sc_hd__a21bo_1
X_3046_ clknet_leaf_31_clk _0308_ net184 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1376_ SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__inv_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ SB0.route_sel\[8\] SB0.route_sel\[9\] vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__nand2b_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload30 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_8
X_2615_ SB0.route_sel\[69\] SB0.route_sel\[68\] net238 vssd1 vssd1 vccd1 vccd1 _0205_
+ sky130_fd_sc_hd__mux2_1
X_1428_ net132 net127 net123 net120 LEI0.config_data\[0\] LEI0.config_data\[1\] vssd1
+ vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__mux4_2
X_2546_ SB0.route_sel\[0\] net171 net250 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__mux2_1
X_2477_ LE_0A.edge_mode LE_0A.config_data\[16\] net231 vssd1 vssd1 vccd1 vccd1 _0068_
+ sky130_fd_sc_hd__mux2_1
X_3029_ clknet_leaf_12_clk _0291_ net220 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1359_ SB0.route_sel\[53\] vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__inv_2
Xclkload2 clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
Xfanout261 net263 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout250 net252 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2400_ _1179_ SB0.route_sel\[89\] _1177_ _1178_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2262_ net59 LE_0B.edge_mode vssd1 vssd1 vccd1 vccd1 LE_0B.sel_clk sky130_fd_sc_hd__xnor2_1
X_2331_ SB0.route_sel\[65\] SB0.route_sel\[64\] _1159_ SB0.route_sel\[66\] vssd1 vssd1
+ vccd1 vccd1 _1074_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2193_ net9 net10 net11 net12 net180 net179 vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__mux4_1
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1977_ _1182_ SB0.route_sel\[102\] _1184_ SB0.route_sel\[97\] _0761_ vssd1 vssd1
+ vccd1 vccd1 _0762_ sky130_fd_sc_hd__a221o_1
X_2529_ CB_1.config_dataB\[3\] CB_1.config_dataB\[2\] net260 vssd1 vssd1 vccd1 vccd1
+ _0119_ sky130_fd_sc_hd__mux2_1
Xhold58 LE_0A.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 LE_0B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 LE_0B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 _0323_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 LE_1B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 LE_1B.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1900_ _0686_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__inv_2
X_1831_ _1307_ _1285_ _1244_ _1264_ net159 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1
+ vccd1 _0618_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2880_ clknet_leaf_29_clk _0142_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_1762_ _0544_ _0545_ _0550_ _0542_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_40_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1693_ net3 _0480_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__nor2_1
X_2176_ _0801_ _0943_ _0945_ _0804_ CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1
+ _0959_ sky130_fd_sc_hd__o221ai_1
X_2245_ LE_1B.config_data\[8\] _0936_ _0966_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a21bo_1
X_2314_ _1288_ _0756_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2030_ net135 net131 net126 net122 LEI0.config_data\[6\] LEI0.config_data\[7\] vssd1
+ vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__mux4_1
X_2932_ clknet_leaf_28_clk _0194_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[58\]
+ sky130_fd_sc_hd__dfstp_1
X_1745_ net168 _0346_ _1189_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__o21a_1
X_2794_ clknet_leaf_7_clk _0056_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1814_ LEI0.config_data\[38\] _0595_ _0602_ _0593_ vssd1 vssd1 vccd1 vccd1 _0603_
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2863_ clknet_leaf_20_clk _0125_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_1676_ _0462_ _0463_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__o21ba_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2159_ _1209_ _0753_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__o21bai_1
X_2228_ CB_1.config_dataB\[13\] _1215_ CB_1.config_dataB\[15\] _1010_ vssd1 vssd1
+ vccd1 vccd1 _1011_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_51_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_24_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1461_ net124 net137 _1251_ SB0.route_sel\[59\] SB0.route_sel\[58\] vssd1 vssd1 vccd1
+ vccd1 _1255_ sky130_fd_sc_hd__a32o_1
X_1530_ _1322_ _1323_ _1319_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__or3b_1
X_1392_ SB0.route_sel\[106\] vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__inv_2
X_2013_ net142 _0796_ _0797_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__o21a_1
X_3062_ clknet_leaf_25_clk _0324_ net206 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_15_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2915_ clknet_leaf_0_clk _0177_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[41\]
+ sky130_fd_sc_hd__dfstp_1
X_2777_ clknet_leaf_12_clk _0039_ net219 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[38\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold111 LEI0.config_data\[45\] vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
X_1728_ _0514_ _0516_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__and2_1
X_2846_ clknet_leaf_22_clk net378 net212 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold100 LE_1A.config_data\[10\] vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
X_1659_ _0447_ _1163_ _0446_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__mux2_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ CB_1.config_dataA\[2\] CB_1.config_dataA\[1\] net264 vssd1 vssd1 vccd1 vccd1
+ _0290_ sky130_fd_sc_hd__mux2_1
X_2562_ SB0.route_sel\[16\] SB0.route_sel\[15\] net229 vssd1 vssd1 vccd1 vccd1 _0152_
+ sky130_fd_sc_hd__mux2_1
X_2631_ SB0.route_sel\[85\] SB0.route_sel\[84\] net233 vssd1 vssd1 vccd1 vccd1 _0221_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_4_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1513_ _1304_ _1306_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__nand2_2
X_2493_ net322 net292 net242 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__mux2_1
X_1444_ SB0.route_sel\[55\] SB0.route_sel\[54\] _1237_ vssd1 vssd1 vccd1 vccd1 _1238_
+ sky130_fd_sc_hd__a21bo_1
X_1375_ SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__inv_2
X_3045_ clknet_leaf_26_clk _0307_ net207 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_2
X_2829_ clknet_leaf_0_clk _0091_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.reset_val sky130_fd_sc_hd__dfrtp_1
X_1993_ _0776_ _0777_ _0371_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__a21bo_2
XTAP_TAPCELL_ROW_15_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload20 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_12
X_2545_ net171 net173 net250 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__mux2_1
X_2614_ SB0.route_sel\[68\] SB0.route_sel\[67\] net238 vssd1 vssd1 vccd1 vccd1 _0204_
+ sky130_fd_sc_hd__mux2_1
X_1427_ net122 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__inv_2
X_2476_ LE_0A.config_data\[16\] net345 net241 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__mux2_1
X_1358_ SB0.route_sel\[51\] vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__inv_2
X_3028_ clknet_leaf_12_clk _0290_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_38_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload3 clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout240 net242 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2261_ net184 LE_0B.reset_mode vssd1 vssd1 vccd1 vccd1 _2261_/X sky130_fd_sc_hd__xor2_2
X_2330_ SB0.route_sel\[68\] _1160_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__nor2_1
X_2192_ net179 _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__nand2_1
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1976_ SB0.route_sel\[100\] SB0.route_sel\[101\] vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nor2_1
X_2528_ CB_1.config_dataB\[2\] CB_1.config_dataB\[1\] net260 vssd1 vssd1 vccd1 vccd1
+ _0118_ sky130_fd_sc_hd__mux2_1
Xhold48 LE_0A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 LEI0.config_data\[43\] vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold26 _0082_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 _0079_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 LE_1B.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ LE_0B.dff1_out _1217_ _1125_ vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__a21o_1
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1761_ CB_0.config_dataA\[7\] _0546_ _0549_ CB_0.config_dataA\[6\] vssd1 vssd1 vccd1
+ vccd1 _0550_ sky130_fd_sc_hd__a211o_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ LE_0A.config_data\[16\] _0615_ _0616_ _0617_ vssd1 vssd1 vccd1 vccd1 CB_0.le_outA
+ sky130_fd_sc_hd__o211a_1
X_1692_ _1251_ _0440_ _0480_ net120 vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__a22o_1
X_2313_ net124 net137 _1272_ _1063_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__a31o_1
X_2175_ net182 _0792_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__a21oi_1
X_2244_ _0936_ LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__and2b_1
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1959_ _1202_ LE_0B.dff_out vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2931_ clknet_leaf_28_clk _0193_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[57\]
+ sky130_fd_sc_hd__dfstp_1
X_2793_ clknet_leaf_7_clk net339 net200 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1744_ net169 _1330_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__nand2_1
X_1813_ _0596_ _0598_ _0601_ CB_0.config_dataA\[15\] CB_0.config_dataA\[14\] vssd1
+ vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a221o_1
X_2862_ clknet_leaf_20_clk _0124_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1675_ net125 _1272_ _0440_ SB0.route_sel\[75\] SB0.route_sel\[74\] vssd1 vssd1 vccd1
+ vccd1 _0464_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2158_ _1209_ _1304_ _0755_ CB_1.config_dataB\[7\] net181 vssd1 vssd1 vccd1 vccd1
+ _0941_ sky130_fd_sc_hd__a311o_1
X_2089_ net4 net5 net138 vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__mux2_1
X_2227_ _1002_ _1004_ _1009_ CB_1.config_dataB\[15\] _1008_ vssd1 vssd1 vccd1 vccd1
+ _1010_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1391_ net18 vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__inv_2
X_1460_ net12 _1252_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2012_ net142 _0793_ _0765_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__a21oi_1
X_3061_ clknet_leaf_24_clk net285 net206 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2845_ clknet_leaf_22_clk _0107_ net212 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2914_ clknet_leaf_0_clk _0176_ net188 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[40\]
+ sky130_fd_sc_hd__dfstp_1
X_2776_ clknet_leaf_12_clk _0038_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_1727_ SB0.route_sel\[84\] _1171_ SB0.route_sel\[87\] _1173_ _0515_ vssd1 vssd1 vccd1
+ vccd1 _0516_ sky130_fd_sc_hd__a221o_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 LE_1A.reset_val vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
X_1658_ SB0.route_sel\[71\] SB0.route_sel\[70\] net55 vssd1 vssd1 vccd1 vccd1 _0447_
+ sky130_fd_sc_hd__a21bo_1
X_1589_ net130 net20 _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__mux2_1
XFILLER_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2492_ net292 LE_0B.config_data\[9\] net240 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__mux2_1
X_2561_ SB0.route_sel\[15\] SB0.route_sel\[14\] net234 vssd1 vssd1 vccd1 vccd1 _0151_
+ sky130_fd_sc_hd__mux2_1
X_1512_ SB0.route_sel\[36\] _1143_ SB0.route_sel\[39\] _1145_ _1305_ vssd1 vssd1 vccd1
+ vccd1 _1306_ sky130_fd_sc_hd__a221o_1
X_2630_ SB0.route_sel\[84\] SB0.route_sel\[83\] net233 vssd1 vssd1 vccd1 vccd1 _0220_
+ sky130_fd_sc_hd__mux2_1
X_1374_ SB0.route_sel\[78\] vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__inv_2
X_1443_ SB0.route_sel\[52\] SB0.route_sel\[53\] net53 vssd1 vssd1 vccd1 vccd1 _1237_
+ sky130_fd_sc_hd__and3_1
X_3044_ clknet_leaf_26_clk _0306_ net207 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_18_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2828_ clknet_leaf_1_clk _0090_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.edge_mode sky130_fd_sc_hd__dfstp_1
X_2759_ clknet_leaf_16_clk _0021_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload10 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__clkinvlp_4
X_1992_ SB0.route_sel\[28\] SB0.route_sel\[29\] SB0.route_sel\[31\] _1142_ vssd1 vssd1
+ vccd1 vccd1 _0777_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_15_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload21 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_12
X_2475_ net345 net317 net241 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__mux2_1
X_2544_ net173 net175 net250 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__mux2_1
X_2613_ SB0.route_sel\[67\] SB0.route_sel\[66\] net238 vssd1 vssd1 vccd1 vccd1 _0203_
+ sky130_fd_sc_hd__mux2_1
X_1426_ net126 vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__inv_2
X_1357_ SB0.route_sel\[46\] vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__inv_2
X_3027_ clknet_leaf_11_clk _0289_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_38_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload4 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__bufinv_16
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
Xfanout252 net253 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_2
Xfanout230 net239 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2260_ LE_0A.edge_mode net59 vssd1 vssd1 vccd1 vccd1 LE_0A.sel_clk sky130_fd_sc_hd__xnor2_1
X_2191_ _0750_ _0759_ _1212_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1975_ _0756_ _0759_ _0753_ _0750_ CB_1.config_dataA\[5\] net142 vssd1 vssd1 vccd1
+ vccd1 _0760_ sky130_fd_sc_hd__mux4_1
X_1409_ net144 vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__inv_2
Xhold38 LE_0B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
X_2458_ _0703_ _0734_ _0738_ _0743_ net60 vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__o221a_1
X_2527_ CB_1.config_dataB\[1\] net183 net253 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__mux2_1
Xhold27 LE_1A.config_data\[8\] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 _0314_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 LE_0A.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_26_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ _1327_ _1112_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__and2b_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1760_ CB_0.config_dataA\[5\] _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_40_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1691_ net174 net172 net178 net176 vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__and4b_1
X_2312_ _1274_ _0753_ _1275_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__a21oi_1
X_2174_ _1209_ _0450_ _0795_ net181 vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__a31o_1
X_2243_ LE_1B.config_data\[11\] LE_1B.config_data\[10\] _0936_ vssd1 vssd1 vccd1 vccd1
+ _1026_ sky130_fd_sc_hd__mux2_1
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1889_ net157 _0346_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__nor2_1
X_1958_ LE_0B.dff0_out LE_0B.dff1_out LE_0B.reset_val vssd1 vssd1 vccd1 vccd1 LE_0B.dff_out
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2861_ clknet_leaf_17_clk _0123_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_2
X_2930_ clknet_leaf_28_clk _0192_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[56\]
+ sky130_fd_sc_hd__dfstp_1
X_1743_ CB_0.config_dataA\[7\] _0527_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__o21ai_1
X_2792_ clknet_leaf_7_clk _0054_ net200 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1812_ _0599_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__nor2_1
XFILLER_30_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1674_ net14 _0461_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__and2b_1
X_2226_ _0753_ _0756_ _0750_ _0759_ _1215_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1
+ vccd1 _1009_ sky130_fd_sc_hd__mux4_1
X_2157_ _1208_ _0938_ _0939_ _1211_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__a31o_1
X_2088_ CB_1.config_dataA\[13\] CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0873_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1390_ SB0.route_sel\[96\] vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__inv_2
X_3060_ clknet_leaf_23_clk _0322_ net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2011_ _0450_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__and2_1
X_2844_ clknet_leaf_22_clk _0106_ net212 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2913_ clknet_leaf_0_clk _0175_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[39\]
+ sky130_fd_sc_hd__dfstp_1
X_1588_ net150 net145 net147 net152 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__or4b_1
Xhold102 LEI0.config_data\[31\] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
X_2775_ clknet_leaf_16_clk _0037_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_1657_ SB0.route_sel\[68\] SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__nand2_1
X_1726_ SB0.route_sel\[82\] SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__nor2_1
X_2209_ net2 _0981_ _0988_ net3 vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o22a_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2491_ LE_0B.config_data\[9\] net296 net240 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__mux2_1
X_2560_ SB0.route_sel\[14\] SB0.route_sel\[13\] net234 vssd1 vssd1 vccd1 vccd1 _0150_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1442_ _1233_ _1234_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__a21oi_1
X_1511_ SB0.route_sel\[35\] SB0.route_sel\[34\] vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nor2_1
X_3043_ clknet_leaf_26_clk _0305_ net207 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1373_ SB0.route_sel\[79\] vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2758_ clknet_leaf_16_clk _0020_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_2827_ clknet_leaf_1_clk _0089_ net190 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2689_ CB_0.config_dataB\[11\] CB_0.config_dataB\[10\] net249 vssd1 vssd1 vccd1 vccd1
+ _0279_ sky130_fd_sc_hd__mux2_1
X_1709_ net170 net16 _0352_ _0497_ _1332_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__o32a_1
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload22 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__inv_12
XPHY_EDGE_ROW_41_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1991_ SB0.route_sel\[24\] SB0.route_sel\[25\] vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__nand2b_1
X_2612_ SB0.route_sel\[66\] SB0.route_sel\[65\] net253 vssd1 vssd1 vccd1 vccd1 _0202_
+ sky130_fd_sc_hd__mux2_1
Xclkload11 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_6
X_1425_ net130 vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__inv_2
X_2474_ net317 net313 net241 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__mux2_1
X_2543_ net175 net177 net250 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3026_ clknet_leaf_12_clk _0288_ net218 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_38_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1356_ SB0.route_sel\[47\] vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__inv_2
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload5 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout264 net271 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_2
Xfanout220 net62 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout242 net245 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_2
Xfanout253 net271 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_4
Xfanout231 net233 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2190_ _0970_ _0971_ _0972_ _0969_ _1214_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__a32o_1
X_1974_ _0757_ _0758_ _1241_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__a21bo_2
Xhold28 LE_0A.config_data\[9\] vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
X_2526_ net183 CB_1.config_dataA\[19\] net253 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__mux2_1
Xhold17 LE_1A.config_data\[7\] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 LE_1B.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ LE_0B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__inv_2
X_2388_ _1186_ SB0.route_sel\[107\] SB0.route_sel\[104\] _1188_ _1111_ vssd1 vssd1
+ vccd1 vccd1 _1112_ sky130_fd_sc_hd__a221o_1
X_2457_ LE_0A.dff0_out _0615_ net60 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__mux2_1
X_3009_ clknet_leaf_5_clk _0271_ net198 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_26_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1339_ SB0.route_sel\[14\] vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_7_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1690_ _0477_ net135 _0478_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ net124 net137 _1231_ _1233_ _1062_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__a32o_1
X_2242_ CB_0.config_data_inA _1001_ _1023_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__o21ai_1
X_2173_ _0778_ _0781_ _0787_ _0784_ _1208_ _1209_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__mux4_1
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1957_ _0703_ _0734_ _0738_ _0743_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__o22a_1
X_1888_ _1307_ _1285_ _1244_ _1264_ net157 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1
+ vccd1 _0675_ sky130_fd_sc_hd__mux4_1
X_2509_ LE_1A.config_data\[4\] LE_1A.config_data\[3\] net255 vssd1 vssd1 vccd1 vccd1
+ _0099_ sky130_fd_sc_hd__mux2_1
XFILLER_11_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2791_ clknet_leaf_7_clk _0053_ net200 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1811_ net27 net28 net16 net17 net165 net164 vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__mux4_1
X_2860_ clknet_leaf_18_clk _0122_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1742_ CB_0.config_dataA\[5\] CB_0.config_dataA\[7\] _0528_ _0530_ vssd1 vssd1 vccd1
+ vccd1 _0531_ sky130_fd_sc_hd__o31a_1
X_1673_ net122 _0461_ _0440_ _1272_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__a2bb2o_1
X_2225_ CB_1.config_dataB\[15\] _1005_ _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__o21ai_1
XFILLER_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2156_ _0343_ _0762_ net182 vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2087_ net9 net10 net11 net12 net138 CB_1.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1
+ _0872_ sky130_fd_sc_hd__mux4_1
X_2989_ clknet_leaf_4_clk _0251_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2010_ _1161_ SB0.route_sel\[70\] SB0.route_sel\[65\] _1164_ _0794_ vssd1 vssd1 vccd1
+ vccd1 _0795_ sky130_fd_sc_hd__a221o_2
X_2912_ clknet_leaf_0_clk _0174_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[38\]
+ sky130_fd_sc_hd__dfstp_1
X_2774_ clknet_leaf_14_clk _0036_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_1725_ _0500_ _0504_ _0510_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__a22o_2
X_2843_ clknet_leaf_22_clk _0105_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
Xhold103 LEI0.config_data\[27\] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
X_1587_ SB0.route_sel\[9\] SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__nand2_1
X_1656_ SB0.route_sel\[67\] SB0.route_sel\[66\] _0442_ _0443_ _0444_ vssd1 vssd1 vccd1
+ vccd1 _0445_ sky130_fd_sc_hd__a221o_1
X_2139_ LEI0.config_data\[11\] _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__or2_1
X_2208_ net13 net14 net180 vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_36_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2490_ net296 net312 net240 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1441_ net124 net137 _1231_ SB0.route_sel\[50\] SB0.route_sel\[51\] vssd1 vssd1 vccd1
+ vccd1 _1235_ sky130_fd_sc_hd__a32o_1
X_1510_ _1292_ _1297_ _1303_ _1293_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__a22o_2
X_1372_ SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__inv_2
X_3042_ clknet_leaf_21_clk _0304_ net215 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2688_ CB_0.config_dataB\[10\] CB_0.config_dataB\[9\] net248 vssd1 vssd1 vccd1 vccd1
+ _0278_ sky130_fd_sc_hd__mux2_1
X_2757_ clknet_leaf_15_clk _0019_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_1708_ net27 net28 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__mux2_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2826_ clknet_leaf_1_clk _0088_ net190 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1639_ _0414_ _0418_ _0423_ _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ _0747_ _0774_ CB_1.config_dataA\[6\] vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__clkinv_8
X_2542_ net177 CB_1.config_dataB\[15\] net258 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__mux2_1
Xclkload12 clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinvlp_4
X_2611_ SB0.route_sel\[65\] SB0.route_sel\[64\] net238 vssd1 vssd1 vccd1 vccd1 _0201_
+ sky130_fd_sc_hd__mux2_1
X_1424_ net134 vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__inv_2
X_2473_ net313 LE_0A.config_data\[12\] net240 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__mux2_1
X_1355_ SB0.route_sel\[44\] vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__inv_2
X_3025_ clknet_leaf_13_clk _0287_ net220 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__bufinv_16
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2809_ LE_0B.sel_clk _0071_ net61 vssd1 vssd1 vccd1 vccd1 LE_0B.dff0_out sky130_fd_sc_hd__dfrtp_1
Xfanout243 net245 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
Xfanout221 net226 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__clkbuf_4
Xfanout265 net270 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net257 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net213 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_12_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1973_ SB0.route_sel\[52\] SB0.route_sel\[53\] SB0.route_sel\[55\] _1154_ vssd1 vssd1
+ vccd1 vccd1 _0758_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_23_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2525_ LE_1B.dff0_out _1217_ _1126_ vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__a21o_1
Xhold29 _0061_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
X_2456_ CB_0.config_data_inA net351 net266 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__mux2_1
X_1407_ CB_0.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__inv_2
X_1338_ SB0.route_sel\[12\] vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__inv_2
Xhold18 _0102_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
X_2387_ net119 SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nor2_1
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3008_ clknet_leaf_5_clk _0270_ net198 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_3_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2172_ CB_1.config_dataB\[6\] CB_1.config_dataB\[7\] _0946_ vssd1 vssd1 vccd1 vccd1
+ _0955_ sky130_fd_sc_hd__and3_1
X_2310_ _1232_ _0759_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2241_ CB_0.config_data_inA _1001_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_48_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1956_ _0701_ _0740_ _0742_ _0729_ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__o31ai_1
X_1887_ LE_0B.config_data\[5\] _0672_ _0642_ vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a21o_1
X_2508_ LE_1A.config_data\[3\] LE_1A.config_data\[2\] net255 vssd1 vssd1 vccd1 vccd1
+ _0098_ sky130_fd_sc_hd__mux2_1
X_2439_ net370 LEI0.config_data\[29\] net269 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__mux2_1
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ clknet_leaf_7_clk net321 net200 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1741_ net19 net169 _0529_ CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _0530_
+ sky130_fd_sc_hd__a211o_1
X_1810_ _0453_ _0473_ _0517_ _0492_ net165 net164 vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__mux4_1
X_1672_ net176 net174 net172 net178 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__or4bb_1
X_2155_ _1325_ _1326_ _0767_ net182 vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o31ai_1
X_2224_ net4 _1215_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__a211o_1
X_2086_ _0756_ _0759_ _0753_ _0750_ CB_1.config_dataA\[13\] net138 vssd1 vssd1 vccd1
+ vccd1 _0871_ sky130_fd_sc_hd__mux4_1
X_1939_ _0707_ _0723_ _0725_ _0722_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__o211a_1
X_2988_ clknet_leaf_4_clk _0250_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[2\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_59_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ clknet_leaf_0_clk _0173_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[37\]
+ sky130_fd_sc_hd__dfstp_1
X_2773_ clknet_leaf_15_clk _0035_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[34\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold104 LEI0.config_data\[35\] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
X_2842_ clknet_leaf_22_clk _0104_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1724_ _0508_ _0511_ _0512_ SB0.route_sel\[80\] SB0.route_sel\[81\] vssd1 vssd1 vccd1
+ vccd1 _0513_ sky130_fd_sc_hd__o311a_1
X_1586_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
X_1655_ net125 _1287_ _0440_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__and3_1
X_2138_ net132 net127 net123 net120 LEI0.config_data\[9\] LEI0.config_data\[10\] vssd1
+ vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__mux4_1
X_2069_ net140 _0853_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__nor2_1
X_2207_ CB_1.config_dataB\[11\] _0989_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1440_ net11 _1232_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__nand2b_1
X_1371_ SB0.route_sel\[74\] vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__inv_2
X_3041_ clknet_leaf_21_clk _0303_ net215 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_61_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2825_ clknet_leaf_1_clk _0087_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2687_ CB_0.config_dataB\[9\] net158 net245 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__mux2_1
X_2756_ clknet_leaf_15_clk _0018_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1707_ _1135_ net17 _0352_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__or3_1
X_1638_ SB0.route_sel\[19\] SB0.route_sel\[18\] _0426_ _0414_ vssd1 vssd1 vccd1 vccd1
+ _0427_ sky130_fd_sc_hd__a31oi_1
X_1569_ net22 net128 _0357_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__mux2_1
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload24 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload24/X sky130_fd_sc_hd__clkbuf_4
X_2472_ net326 net323 net240 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__mux2_1
Xclkload13 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload13/X sky130_fd_sc_hd__clkbuf_8
X_2610_ SB0.route_sel\[64\] SB0.route_sel\[63\] net238 vssd1 vssd1 vccd1 vccd1 _0200_
+ sky130_fd_sc_hd__mux2_1
X_2541_ CB_1.config_dataB\[15\] CB_1.config_dataB\[14\] net259 vssd1 vssd1 vccd1 vccd1
+ _0131_ sky130_fd_sc_hd__mux2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1423_ net60 vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__inv_2
X_1354_ SB0.route_sel\[43\] vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__inv_2
X_3024_ clknet_leaf_13_clk _0286_ net220 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2808_ clknet_leaf_31_clk _0070_ net184 vssd1 vssd1 vccd1 vccd1 LE_0A.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
Xclkload7 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__inv_6
Xfanout222 net226 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_4
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
Xfanout211 net213 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
X_2739_ clknet_leaf_22_clk _0001_ net214 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout244 net245 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
Xfanout266 net270 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout233 net239 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net257 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1972_ _1155_ SB0.route_sel\[48\] vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2455_ net351 LEI0.config_data\[45\] net266 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__mux2_1
X_2524_ LE_1A.reset_mode net372 net254 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1406_ LEI0.config_data\[41\] vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__inv_2
X_1337_ SB0.route_sel\[11\] vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__inv_2
Xhold19 LE_1B.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ _1327_ _1110_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__nor2_2
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3007_ clknet_leaf_5_clk _0269_ net198 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_34_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2171_ _0940_ _0942_ _0947_ _0953_ _1210_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__a311oi_1
XFILLER_32_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2240_ _1022_ _1011_ CB_1.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_38_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1955_ LE_0B.config_data\[11\] _0672_ _0741_ _0641_ vssd1 vssd1 vccd1 vccd1 _0742_
+ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_31_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1886_ LE_0B.config_data\[4\] _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0673_
+ sky130_fd_sc_hd__and4_1
X_2438_ LEI0.config_data\[29\] net354 net267 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__mux2_1
X_2507_ LE_1A.config_data\[2\] LE_1A.config_data\[1\] net255 vssd1 vssd1 vccd1 vccd1
+ _0097_ sky130_fd_sc_hd__mux2_1
X_2369_ SB0.route_sel\[17\] SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__and2b_1
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1740_ _1185_ net169 CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__o21ai_1
X_1671_ _0457_ _0458_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__a21o_1
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2154_ net132 net127 net123 _1221_ LEI0.config_data\[21\] LEI0.config_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__mux4_1
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2085_ _0844_ _0869_ _0814_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__mux2_1
X_2223_ net5 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__and2_1
X_2987_ clknet_leaf_4_clk _0249_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_1938_ net16 _0713_ _0724_ net17 vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__o22a_1
X_1869_ _1199_ _0645_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2841_ clknet_leaf_22_clk _0103_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2910_ clknet_leaf_2_clk _0172_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[36\]
+ sky130_fd_sc_hd__dfstp_1
X_2772_ clknet_leaf_15_clk _0034_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold105 LEI0.config_data\[39\] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
X_1654_ net13 _0441_ vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__nand2b_1
X_1723_ SB0.route_sel\[84\] SB0.route_sel\[85\] net30 vssd1 vssd1 vccd1 vccd1 _0512_
+ sky130_fd_sc_hd__a21boi_1
X_1585_ _0372_ _0373_ _0371_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__a21bo_4
X_2206_ net1 net6 net7 net8 net180 net179 vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__mux4_1
X_2137_ net183 _0919_ CB_1.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__o21ai_1
X_2068_ CB_1.config_dataA\[9\] CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0853_
+ sky130_fd_sc_hd__nand2_1
XFILLER_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1370_ SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__inv_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3040_ clknet_leaf_21_clk _0302_ net215 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_61_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2824_ clknet_leaf_1_clk _0086_ net189 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2755_ clknet_leaf_15_clk _0017_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2686_ net158 CB_0.config_dataB\[7\] net241 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__mux2_1
X_1706_ CB_0.config_dataA\[3\] _0494_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__or2_1
X_1637_ _0425_ _1139_ _0424_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__mux2_1
X_1568_ net145 net147 net149 net151 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__and4bb_1
X_1499_ SB0.route_sel\[33\] SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nand2_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload25 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__clkinv_4
X_2471_ net323 LE_0A.config_data\[10\] net240 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__mux2_1
X_1422_ LE_1B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__inv_2
Xclkload14 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__bufinv_16
X_2540_ CB_1.config_dataB\[14\] CB_1.config_dataB\[13\] net258 vssd1 vssd1 vccd1 vccd1
+ _0130_ sky130_fd_sc_hd__mux2_1
X_3023_ clknet_leaf_13_clk _0285_ net220 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1353_ SB0.route_sel\[32\] vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__inv_2
Xclkload8 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__clkinv_2
X_2807_ clknet_leaf_1_clk _0069_ net188 vssd1 vssd1 vccd1 vccd1 LE_0A.reset_val sky130_fd_sc_hd__dfrtp_1
X_2738_ LE_0A.sel_clk _0000_ net61 vssd1 vssd1 vccd1 vccd1 LE_0A.dff1_out sky130_fd_sc_hd__dfstp_1
Xfanout245 net249 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout201 net205 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
Xfanout223 net226 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_2
X_2669_ CB_0.config_dataA\[11\] CB_0.config_dataA\[10\] net243 vssd1 vssd1 vccd1 vccd1
+ _0259_ sky130_fd_sc_hd__mux2_1
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_2
Xfanout267 net270 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
XFILLER_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _1304_ _0755_ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__nand2_2
X_2454_ net382 LEI0.config_data\[44\] net266 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__mux2_1
X_1405_ CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__inv_2
X_2523_ net372 LE_1A.edge_mode net254 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__mux2_1
X_2385_ _1186_ SB0.route_sel\[107\] SB0.route_sel\[104\] SB0.route_sel\[105\] _1109_
+ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__o221a_1
X_3006_ clknet_leaf_9_clk _0268_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xinput1 CBeast_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1336_ SB0.route_sel\[1\] vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__inv_2
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ CB_1.config_dataB\[7\] _0948_ _0950_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_
+ sky130_fd_sc_hd__o211a_1
X_1954_ LE_0B.config_data\[10\] _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0741_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_31_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1885_ _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__nand3_4
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2437_ net354 LEI0.config_data\[27\] net267 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__mux2_1
X_2506_ LE_1A.config_data\[1\] LE_1A.config_data\[0\] net255 vssd1 vssd1 vccd1 vccd1
+ _0096_ sky130_fd_sc_hd__mux2_1
X_2368_ _0428_ _1098_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__and2_1
X_2299_ _0334_ _1056_ _0337_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__a21o_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ net136 _1269_ _0437_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__and3_1
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2222_ net9 net10 net11 net12 CB_1.config_dataB\[12\] CB_1.config_dataB\[13\] vssd1
+ vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__mux4_1
X_2153_ _0918_ _0920_ _0935_ CB_1.config_dataB\[2\] _0922_ vssd1 vssd1 vccd1 vccd1
+ _0936_ sky130_fd_sc_hd__o221a_4
X_2084_ LE_1A.config_data\[7\] LE_1A.config_data\[6\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0869_ sky130_fd_sc_hd__mux2_1
X_1937_ CB_0.config_dataB\[13\] net156 net153 vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__nand3_1
X_2986_ clknet_leaf_17_clk _0248_ net221 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1799_ _1195_ _0587_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__a21o_1
X_1868_ net162 _0346_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_59_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2771_ clknet_leaf_16_clk _0033_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_2840_ clknet_leaf_24_clk net289 net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1722_ _1172_ _1173_ net44 SB0.route_sel\[85\] SB0.route_sel\[84\] vssd1 vssd1 vccd1
+ vccd1 _0511_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1584_ SB0.route_sel\[26\] SB0.route_sel\[27\] _1141_ SB0.route_sel\[29\] vssd1 vssd1
+ vccd1 vccd1 _0373_ sky130_fd_sc_hd__o22a_1
Xhold106 LE_1A.config_data\[13\] vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
X_1653_ _1287_ _0440_ _0441_ net121 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__o2bb2a_1
X_2205_ net179 net180 CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__nand3_1
X_2067_ CB_1.config_dataA\[11\] _0845_ _0848_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_
+ sky130_fd_sc_hd__o211a_1
X_2136_ CB_1.config_dataB\[1\] CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0919_
+ sky130_fd_sc_hd__nand2_1
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2969_ clknet_leaf_4_clk _0231_ net203 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[95\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2754_ clknet_leaf_15_clk _0016_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_1705_ net15 net20 net21 net22 net170 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0494_ sky130_fd_sc_hd__mux4_1
X_2823_ clknet_leaf_2_clk net273 net189 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2685_ CB_0.config_dataB\[7\] CB_0.config_dataB\[6\] net241 vssd1 vssd1 vccd1 vccd1
+ _0275_ sky130_fd_sc_hd__mux2_1
X_1636_ SB0.route_sel\[23\] SB0.route_sel\[22\] net49 vssd1 vssd1 vccd1 vccd1 _0425_
+ sky130_fd_sc_hd__a21bo_1
X_1567_ SB0.route_sel\[25\] SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__nand2_1
X_2119_ _0900_ _0901_ _0814_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__mux2_1
X_1498_ SB0.route_sel\[35\] SB0.route_sel\[34\] _1289_ _1290_ _1291_ vssd1 vssd1 vccd1
+ vccd1 _1292_ sky130_fd_sc_hd__a221o_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload26 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__clkinv_2
Xclkload15 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload15/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_23_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2470_ LE_0A.config_data\[10\] net299 net243 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__mux2_1
X_1421_ CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__inv_2
X_3022_ clknet_leaf_12_clk _0284_ net219 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1352_ net37 vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__inv_2
X_2668_ CB_0.config_dataA\[10\] net166 net243 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__mux2_1
X_2737_ LE_1B.reset_mode LE_1B.reset_val net227 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__mux2_1
Xclkload9 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__clkinv_2
X_2806_ clknet_leaf_1_clk _0068_ net188 vssd1 vssd1 vccd1 vccd1 LE_0A.edge_mode sky130_fd_sc_hd__dfstp_1
Xfanout268 net270 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
Xfanout224 net226 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net248 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_4
X_1619_ SB0.route_sel\[4\] SB0.route_sel\[5\] net29 vssd1 vssd1 vccd1 vccd1 _0408_
+ sky130_fd_sc_hd__a21bo_1
X_2599_ SB0.route_sel\[53\] SB0.route_sel\[52\] net236 vssd1 vssd1 vccd1 vccd1 _0189_
+ sky130_fd_sc_hd__mux2_1
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
Xfanout213 net216 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
Xfanout257 net271 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_37_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1970_ _1144_ SB0.route_sel\[38\] SB0.route_sel\[33\] _1147_ _0754_ vssd1 vssd1 vccd1
+ vccd1 _0755_ sky130_fd_sc_hd__a221o_2
X_2522_ LE_1A.edge_mode LE_1A.config_data\[16\] net254 vssd1 vssd1 vccd1 vccd1 _0112_
+ sky130_fd_sc_hd__mux2_1
X_2453_ LEI0.config_data\[44\] net330 net261 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__mux2_1
X_1335_ SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__inv_2
X_2384_ _1187_ SB0.route_sel\[109\] vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__nand2_1
X_1404_ LE_0A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__inv_2
X_3005_ clknet_leaf_13_clk _0267_ net219 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[19\]
+ sky130_fd_sc_hd__dfstp_2
Xinput2 CBeast_in[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_34_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_27_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1884_ _0663_ _0665_ _0670_ CB_0.config_dataB\[2\] vssd1 vssd1 vccd1 vccd1 _0671_
+ sky130_fd_sc_hd__a31o_2
X_1953_ LE_0B.config_data\[9\] _0672_ _0739_ _0642_ vssd1 vssd1 vccd1 vccd1 _0740_
+ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_31_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2505_ LE_1A.config_data\[0\] LE_0B.reset_mode net227 vssd1 vssd1 vccd1 vccd1 _0095_
+ sky130_fd_sc_hd__mux2_1
X_2436_ net374 net367 net266 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__mux2_1
X_2298_ _0763_ net121 _0335_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__mux2_1
X_2367_ _1136_ SB0.route_sel\[18\] _1137_ SB0.route_sel\[21\] _1097_ vssd1 vssd1 vccd1
+ vccd1 _1098_ sky130_fd_sc_hd__a221o_1
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2152_ CB_1.config_dataB\[3\] _0923_ _0934_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__o21ba_1
X_2221_ CB_1.config_dataB\[12\] _0768_ _1003_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__a21o_1
X_2083_ _1204_ _0852_ _0854_ _0867_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__o31a_1
X_1936_ net27 net28 net156 vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__mux2_1
X_1867_ net162 _1330_ _0652_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__a21oi_1
X_2985_ clknet_leaf_24_clk _0247_ net207 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfstp_1
X_1798_ _1307_ _1285_ net165 vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__mux2_1
Xinput60 le_en vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
X_2419_ net316 net337 net262 vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2770_ clknet_leaf_15_clk _0032_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_1721_ _0506_ _0507_ _0508_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__o211ai_1
X_1583_ SB0.route_sel\[31\] _1142_ vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__nand2_1
Xhold107 _0108_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
X_1652_ net176 net178 net173 net171 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__or4b_1
X_2135_ CB_1.config_dataB\[3\] _0909_ _0913_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_
+ sky130_fd_sc_hd__o211a_1
X_2204_ CB_1.config_dataB\[8\] _0796_ _0972_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_
+ sky130_fd_sc_hd__o211a_1
X_2066_ CB_1.config_dataA\[11\] _0849_ _0850_ _0846_ vssd1 vssd1 vccd1 vccd1 _0851_
+ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_14_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1919_ net154 net153 vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__and2b_1
X_2968_ clknet_leaf_4_clk _0230_ net203 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[94\]
+ sky130_fd_sc_hd__dfstp_1
X_2899_ clknet_leaf_30_clk _0161_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_27_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2753_ clknet_leaf_15_clk _0015_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2684_ CB_0.config_dataB\[6\] CB_0.config_dataB\[5\] net241 vssd1 vssd1 vccd1 vccd1
+ _0274_ sky130_fd_sc_hd__mux2_1
X_1704_ _1135_ _0352_ _0489_ _0491_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__and4bb_1
X_2822_ clknet_leaf_5_clk _0084_ net198 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1566_ CB_0.config_dataA\[2\] _0353_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__and2_1
X_1635_ SB0.route_sel\[20\] SB0.route_sel\[21\] vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__nand2_1
X_1497_ net125 net137 _1287_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__and3_1
X_2049_ _0753_ _0756_ _0750_ _0759_ _1203_ CB_1.config_dataA\[1\] vssd1 vssd1 vccd1
+ vccd1 _0834_ sky130_fd_sc_hd__mux4_1
X_2118_ LE_1A.config_data\[9\] LE_1A.config_data\[8\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0903_ sky130_fd_sc_hd__mux2_1
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload27 clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__bufinv_16
Xclkload16 clknet_leaf_26_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_23_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1351_ SB0.route_sel\[38\] vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__inv_2
X_1420_ CB_1.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__inv_2
X_3021_ clknet_leaf_12_clk _0283_ net219 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2805_ clknet_leaf_6_clk _0067_ net196 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_2667_ net166 net167 net243 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__mux2_1
X_1618_ SB0.route_sel\[7\] SB0.route_sel\[6\] _0406_ vssd1 vssd1 vccd1 vccd1 _0407_
+ sky130_fd_sc_hd__a21bo_1
X_2736_ LE_1B.reset_val LE_1B.edge_mode net250 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__mux2_1
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_2
Xfanout225 net226 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_2
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
X_1549_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__and2_1
Xfanout247 net248 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_2
Xfanout258 net271 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
Xfanout214 net216 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
Xfanout236 net239 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_2
X_2598_ SB0.route_sel\[52\] SB0.route_sel\[51\] net237 vssd1 vssd1 vccd1 vccd1 _0188_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2521_ LE_1A.config_data\[16\] net279 net256 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__mux2_1
X_1403_ CB_0.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__inv_2
X_2452_ net330 net353 net261 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__mux2_1
X_2383_ _0410_ _1108_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__and2_1
X_1334_ SB0.route_sel\[5\] vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3004_ clknet_leaf_13_clk _0266_ net219 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[18\]
+ sky130_fd_sc_hd__dfstp_1
Xinput3 CBeast_in[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2719_ net276 LE_1B.config_data\[0\] net251 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__mux2_1
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1883_ _0518_ _0656_ _0669_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__o21ba_1
X_1952_ LE_0B.config_data\[8\] _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0739_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_31_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2435_ net367 net358 net261 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__mux2_1
X_2504_ LE_1B.dff1_out _1217_ _1126_ vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__a21o_1
X_2366_ SB0.route_sel\[17\] SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__nor2_1
X_2297_ _1315_ _1055_ _1318_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__a21o_1
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2082_ LEI0.config_data\[32\] _0855_ _0866_ CB_1.config_dataA\[10\] vssd1 vssd1 vccd1
+ vccd1 _0867_ sky130_fd_sc_hd__o22a_1
X_2151_ _0912_ _0924_ _0925_ _0926_ _0933_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__a311o_1
X_2220_ CB_1.config_dataB\[13\] CB_1.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 _1003_
+ sky130_fd_sc_hd__nand2b_1
X_2984_ clknet_leaf_26_clk _0246_ net206 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[110\]
+ sky130_fd_sc_hd__dfstp_1
X_1797_ CB_0.config_dataA\[15\] _0583_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__o21ai_1
X_1935_ net153 _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__or2_1
X_1866_ _0650_ _0651_ _0652_ _0649_ CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1
+ _0653_ sky130_fd_sc_hd__o32a_1
Xinput61 le_nrst vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_4
Xinput50 SBwest_in[3] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2418_ net337 LEI0.config_data\[8\] net262 vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__mux2_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2349_ _1148_ SB0.route_sel\[42\] _1149_ SB0.route_sel\[45\] _1085_ vssd1 vssd1 vccd1
+ vccd1 _1086_ sky130_fd_sc_hd__a221o_1
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold108 LEI0.config_data\[23\] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
X_1720_ net125 _1231_ _0440_ vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__nand3_1
X_1651_ CB_1.config_dataA\[18\] CB_1.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 _0440_
+ sky130_fd_sc_hd__and2b_2
X_1582_ _0366_ _0370_ _0356_ _0360_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__a2bb2o_1
X_2065_ net4 net5 net140 vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__mux2_1
X_2134_ _0916_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__inv_2
X_2203_ CB_1.config_dataB\[8\] _0793_ vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__nand2_1
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2967_ clknet_leaf_4_clk _0229_ net203 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[93\]
+ sky130_fd_sc_hd__dfstp_1
X_1918_ net153 _0704_ vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__nor2_1
X_1849_ net160 CB_0.config_dataB\[6\] CB_0.config_dataB\[7\] CB_0.config_dataB\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__and4b_1
X_2898_ clknet_leaf_30_clk _0160_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[24\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2821_ clknet_leaf_5_clk net293 net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2752_ clknet_leaf_14_clk _0014_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2683_ CB_0.config_dataB\[5\] net160 net241 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1703_ _0489_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__and2_2
X_1634_ SB0.route_sel\[19\] SB0.route_sel\[18\] _0420_ _0421_ _0422_ vssd1 vssd1 vccd1
+ vccd1 _0423_ sky130_fd_sc_hd__a221o_1
X_1565_ CB_0.config_dataA\[3\] _1308_ _0351_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1
+ vccd1 _0354_ sky130_fd_sc_hd__o211a_1
X_1496_ net9 _1288_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nand2b_1
X_2048_ CB_1.config_dataA\[3\] _0817_ _0832_ vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__o21ba_1
X_2117_ LE_1A.config_data\[11\] LE_1A.config_data\[10\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0902_ sky130_fd_sc_hd__mux2_1
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload28 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload17 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_23_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1350_ SB0.route_sel\[39\] vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__inv_2
X_3020_ clknet_leaf_10_clk _0282_ net217 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2804_ clknet_leaf_6_clk _0066_ net197 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout204 net205 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
X_2666_ net167 CB_0.config_dataA\[7\] net244 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__mux2_1
X_1617_ SB0.route_sel\[4\] SB0.route_sel\[5\] net43 vssd1 vssd1 vccd1 vccd1 _0406_
+ sky130_fd_sc_hd__and3_1
X_2735_ LE_1B.edge_mode LE_1B.config_data\[16\] net250 vssd1 vssd1 vccd1 vccd1 _0325_
+ sky130_fd_sc_hd__mux2_1
X_2597_ SB0.route_sel\[51\] SB0.route_sel\[50\] net238 vssd1 vssd1 vccd1 vccd1 _0187_
+ sky130_fd_sc_hd__mux2_1
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net62 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout259 net271 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_2
X_1479_ _1230_ _1272_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__nand2_1
X_1548_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] net125 _1287_ vssd1 vssd1
+ vccd1 vccd1 _0337_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_37_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1402_ CB_0.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__inv_2
X_2451_ net353 LEI0.config_data\[41\] net261 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__mux2_1
X_2520_ net279 LE_1A.config_data\[14\] net256 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__mux2_1
Xinput4 CBeast_in[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_4
X_3003_ clknet_leaf_9_clk _0265_ net219 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2382_ SB0.route_sel\[3\] _1127_ SB0.route_sel\[0\] _1130_ _1107_ vssd1 vssd1 vccd1
+ vccd1 _1108_ sky130_fd_sc_hd__a221o_1
X_1333_ SB0.route_sel\[2\] vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__inv_2
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2718_ LE_1B.config_data\[0\] LE_0A.reset_mode net227 vssd1 vssd1 vccd1 vccd1 _0308_
+ sky130_fd_sc_hd__mux2_1
X_2649_ SB0.route_sel\[103\] SB0.route_sel\[102\] net260 vssd1 vssd1 vccd1 vccd1 _0239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1882_ CB_0.config_dataB\[1\] net163 CB_0.config_dataB\[3\] _0492_ _0668_ vssd1 vssd1
+ vccd1 vccd1 _0669_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_31_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ _0735_ _0736_ _0737_ _0641_ _0701_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__o221a_1
X_2434_ net358 LEI0.config_data\[24\] net261 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__mux2_1
X_2503_ net60 _1030_ _1038_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__and3_1
X_2365_ _1095_ _1096_ _0371_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__o21a_1
X_2296_ _0769_ net122 _1316_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__mux2_1
XANTENNA_31 CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2081_ CB_1.config_dataA\[11\] _0856_ _0858_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_
+ sky130_fd_sc_hd__o211a_1
X_2150_ _0489_ _0800_ _0928_ _0932_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__a31o_1
X_1934_ net15 net20 net21 net22 net155 net154 vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__mux4_1
X_2983_ clknet_leaf_22_clk _0245_ net213 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[109\]
+ sky130_fd_sc_hd__dfstp_1
Xinput62 nrst vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_2
X_1796_ net164 _1197_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or3_1
X_1865_ net161 _1199_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__or2_1
Xinput40 SBsouth_in[7] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_1
Xinput51 SBwest_in[4] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
X_2417_ LEI0.config_data\[8\] net356 net261 vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__mux2_1
X_2348_ SB0.route_sel\[41\] SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__nor2_1
X_2279_ _1265_ net128 _1247_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1650_ net134 _0436_ _0438_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold109 LE_1A.config_data\[6\] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1581_ SB0.route_sel\[26\] SB0.route_sel\[27\] _0368_ _0369_ _0356_ vssd1 vssd1 vccd1
+ vccd1 _0370_ sky130_fd_sc_hd__a41o_1
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2202_ CB_1.config_dataB\[11\] _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_53_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2064_ net9 net10 net11 net12 net140 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0849_ sky130_fd_sc_hd__mux4_1
X_2133_ CB_1.config_dataB\[3\] _0914_ _0915_ _0911_ vssd1 vssd1 vccd1 vccd1 _0916_
+ sky130_fd_sc_hd__o22a_1
X_1917_ _1307_ _1285_ _1244_ _1264_ net155 net154 vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__mux4_1
X_2966_ clknet_leaf_4_clk _0228_ net202 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[92\]
+ sky130_fd_sc_hd__dfstp_1
X_2897_ clknet_leaf_31_clk _0159_ net184 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[23\]
+ sky130_fd_sc_hd__dfstp_1
X_1779_ CB_0.config_dataA\[11\] _0557_ _0561_ _0567_ _1193_ vssd1 vssd1 vccd1 vccd1
+ _0568_ sky130_fd_sc_hd__a221oi_1
X_1848_ _0625_ _0632_ _0634_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_4_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2751_ clknet_leaf_14_clk net302 net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_2820_ clknet_leaf_6_clk net297 net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1564_ net170 _0352_ vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__nor2_1
X_2682_ net159 CB_0.config_dataB\[3\] net242 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__mux2_1
X_1702_ SB0.route_sel\[92\] _1176_ SB0.route_sel\[95\] _1178_ _0490_ vssd1 vssd1 vccd1
+ vccd1 _0491_ sky130_fd_sc_hd__a221o_1
X_1633_ net124 _1231_ _0361_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__and3_1
X_1495_ net137 _1287_ _1288_ net121 vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__o2bb2a_1
X_2047_ _0818_ _0819_ _0821_ _0823_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_1_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2116_ LE_1A.config_data\[15\] LE_1A.config_data\[14\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0901_ sky130_fd_sc_hd__mux2_1
XFILLER_22_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2949_ clknet_leaf_27_clk _0211_ net209 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[75\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload29 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__clkinv_8
Xclkload18 clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_23_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2803_ clknet_leaf_6_clk _0065_ net197 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2734_ LE_1B.config_data\[16\] net368 net251 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__mux2_1
Xfanout205 net62 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
X_2665_ CB_0.config_dataA\[7\] CB_0.config_dataA\[6\] net244 vssd1 vssd1 vccd1 vccd1
+ _0255_ sky130_fd_sc_hd__mux2_1
X_1547_ net4 CB_1.le_outB _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__mux2_1
Xfanout216 net62 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
X_1616_ _0402_ _0403_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__o21ba_1
Xfanout227 net230 vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_4
X_2596_ SB0.route_sel\[50\] SB0.route_sel\[49\] net237 vssd1 vssd1 vccd1 vccd1 _0186_
+ sky130_fd_sc_hd__mux2_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
Xfanout249 net58 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_2
X_1478_ CB_1.config_dataA\[17\] CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1272_
+ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_37_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1401_ net164 vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__inv_2
X_2450_ LEI0.config_data\[41\] net365 net263 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__mux2_1
X_2381_ SB0.route_sel\[7\] SB0.route_sel\[6\] vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nor2_1
Xinput5 CBeast_in[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_4
X_3002_ clknet_leaf_9_clk _0264_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2717_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] net252 vssd1 vssd1 vccd1 vccd1
+ _0307_ sky130_fd_sc_hd__mux2_1
X_2648_ SB0.route_sel\[102\] SB0.route_sel\[101\] net260 vssd1 vssd1 vccd1 vccd1 _0238_
+ sky130_fd_sc_hd__mux2_1
X_2579_ SB0.route_sel\[33\] SB0.route_sel\[32\] net232 vssd1 vssd1 vccd1 vccd1 _0169_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1950_ LE_0B.config_data\[14\] LE_0B.config_data\[15\] _0672_ vssd1 vssd1 vccd1 vccd1
+ _0737_ sky130_fd_sc_hd__mux2_1
X_1881_ _0666_ _0667_ _1199_ vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2502_ LE_1A.dff0_out _0907_ net60 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__mux2_1
X_2433_ LEI0.config_data\[24\] net379 net266 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__mux2_1
X_2364_ SB0.route_sel\[26\] _1140_ SB0.route_sel\[31\] SB0.route_sel\[30\] vssd1 vssd1
+ vccd1 vccd1 _1096_ sky130_fd_sc_hd__o22ai_1
X_2295_ _0397_ _1054_ _0399_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__a21o_1
XANTENNA_10 _0687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_32 LE_1B.config_data\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2080_ _0804_ _0854_ _0859_ _0801_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__a221oi_1
X_1933_ _0518_ _0713_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__nor2_1
X_2982_ clknet_leaf_26_clk _0244_ net206 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[108\]
+ sky130_fd_sc_hd__dfstp_1
X_1795_ net18 net19 net165 vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__mux2_1
X_1864_ _1185_ net163 vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__nor2_1
Xinput30 SBsouth_in[10] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 SBsouth_in[8] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_1
Xinput52 SBwest_in[5] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
X_2416_ net356 LEI0.config_data\[6\] net261 vssd1 vssd1 vccd1 vccd1 _0008_ sky130_fd_sc_hd__mux2_1
X_2278_ net135 _1045_ _0438_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__mux2_1
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2347_ _1083_ _1084_ _1241_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_58_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ SB0.route_sel\[28\] SB0.route_sel\[29\] net36 vssd1 vssd1 vccd1 vccd1 _0369_
+ sky130_fd_sc_hd__a21bo_1
X_2132_ net4 net5 net183 vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__mux2_1
X_2201_ _0781_ _0784_ _0778_ _0787_ _1212_ net179 vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__mux4_1
X_2063_ net140 _0763_ _0847_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1847_ CB_0.config_dataB\[7\] _0631_ _0633_ _0620_ vssd1 vssd1 vccd1 vccd1 _0634_
+ sky130_fd_sc_hd__o22a_1
X_2965_ clknet_leaf_4_clk _0227_ net202 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[91\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1916_ _0673_ _0674_ _0702_ _0641_ _0701_ vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__o221a_1
X_2896_ clknet_leaf_31_clk _0158_ net184 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[22\]
+ sky130_fd_sc_hd__dfstp_1
X_1778_ _1244_ _0557_ _0563_ _0565_ _0566_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ clknet_leaf_14_clk _0012_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2681_ CB_0.config_dataB\[3\] CB_0.config_dataB\[2\] net242 vssd1 vssd1 vccd1 vccd1
+ _0271_ sky130_fd_sc_hd__mux2_1
X_1701_ SB0.route_sel\[90\] SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__nor2_1
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1563_ CB_0.config_dataA\[1\] CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _0352_
+ sky130_fd_sc_hd__nand2_1
X_1632_ net7 _0419_ vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__nand2b_1
X_1494_ net176 net177 net172 net173 vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_1_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ LE_1A.config_data\[13\] LE_1A.config_data\[12\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0900_ sky130_fd_sc_hd__mux2_1
X_2046_ _0489_ _0800_ _0826_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__a31o_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2948_ clknet_leaf_27_clk _0210_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[74\]
+ sky130_fd_sc_hd__dfstp_1
X_2879_ clknet_leaf_29_clk _0141_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[5\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_15_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload19 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_6
XFILLER_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2664_ CB_0.config_dataA\[6\] CB_0.config_dataA\[5\] net244 vssd1 vssd1 vccd1 vccd1
+ _0254_ sky130_fd_sc_hd__mux2_1
X_2802_ clknet_leaf_6_clk net314 net197 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2733_ LE_1B.config_data\[15\] net284 net251 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__mux2_1
X_1477_ net133 _1268_ _1270_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__mux2_2
Xfanout217 net220 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_4
Xfanout239 net249 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
X_1615_ net124 _1287_ _0361_ SB0.route_sel\[2\] SB0.route_sel\[3\] vssd1 vssd1 vccd1
+ vccd1 _0404_ sky130_fd_sc_hd__a32o_1
X_2595_ SB0.route_sel\[49\] SB0.route_sel\[48\] net236 vssd1 vssd1 vccd1 vccd1 _0185_
+ sky130_fd_sc_hd__mux2_1
Xfanout228 net230 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_2
Xfanout206 net209 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
X_1546_ net176 net177 net171 net174 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__and4bb_1
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2029_ _0775_ _0812_ _0813_ LEI0.config_data\[20\] vssd1 vssd1 vccd1 vccd1 _0814_
+ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_20_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1400_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__inv_2
X_2380_ _1105_ _1106_ _0410_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__a21boi_2
X_3001_ clknet_leaf_9_clk _0263_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[15\]
+ sky130_fd_sc_hd__dfstp_2
Xinput6 CBeast_in[1] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_34_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2647_ SB0.route_sel\[101\] SB0.route_sel\[100\] net260 vssd1 vssd1 vccd1 vccd1 _0237_
+ sky130_fd_sc_hd__mux2_1
X_2716_ CB_1.config_dataA\[18\] CB_1.config_dataA\[17\] net252 vssd1 vssd1 vccd1 vccd1
+ _0306_ sky130_fd_sc_hd__mux2_1
X_2578_ SB0.route_sel\[32\] SB0.route_sel\[31\] net230 vssd1 vssd1 vccd1 vccd1 _0168_
+ sky130_fd_sc_hd__mux2_1
X_1529_ SB0.route_sel\[108\] SB0.route_sel\[109\] net33 vssd1 vssd1 vccd1 vccd1 _1323_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ net15 net20 net21 net22 net163 net161 vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2501_ LE_0B.reset_mode LE_0B.reset_val net227 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__mux2_1
X_2294_ _0396_ _0413_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__nand2_1
X_2432_ LEI0.config_data\[23\] net346 net268 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2363_ SB0.route_sel\[25\] SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_33 _0578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 _0781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput20 CBnorth_in[1] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
X_1932_ net155 _0453_ _0706_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__o211a_1
X_1863_ net19 net162 vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__and2_1
Xinput31 SBsouth_in[11] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dlymetal6s2s_1
X_2981_ clknet_leaf_26_clk _0243_ net206 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[107\]
+ sky130_fd_sc_hd__dfstp_1
X_2415_ LEI0.config_data\[6\] net341 net267 vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__mux2_1
X_1794_ net23 net24 net25 net26 net165 net164 vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__mux4_1
Xinput42 SBsouth_in[9] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_1
Xinput53 SBwest_in[6] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
X_2277_ net131 _0453_ _0435_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__mux2_1
X_2346_ SB0.route_sel\[55\] SB0.route_sel\[54\] _1155_ SB0.route_sel\[48\] vssd1 vssd1
+ vccd1 vccd1 _1084_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_50_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2200_ LEI0.config_data\[35\] _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nor2_1
X_2062_ net140 _0768_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__a21oi_1
X_2131_ net9 net10 net11 net12 net183 CB_1.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1
+ _0914_ sky130_fd_sc_hd__mux4_1
X_2964_ clknet_leaf_4_clk _0226_ net202 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[90\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_14_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1777_ net166 net167 _1264_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__and3_1
X_1846_ net27 net28 net160 vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__mux2_1
X_1915_ LE_0B.config_data\[6\] LE_0B.config_data\[7\] _0672_ vssd1 vssd1 vccd1 vccd1
+ _0702_ sky130_fd_sc_hd__mux2_1
X_2895_ clknet_leaf_31_clk _0157_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[21\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _1071_ _1072_ _0469_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__o21a_1
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ CB_0.config_dataB\[2\] net161 net242 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__mux2_1
X_1700_ _0475_ _0479_ _0485_ _0488_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__a22o_2
X_1631_ _1231_ _0361_ _0419_ net121 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__o2bb2a_1
X_1562_ _1331_ _1332_ _0347_ _0350_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__o31a_1
X_1493_ CB_1.config_dataA\[17\] CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1287_
+ sky130_fd_sc_hd__nor2_2
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2045_ _0825_ _0827_ _0829_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0830_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _0870_ _0898_ _0868_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__mux2_1
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2947_ clknet_leaf_3_clk _0209_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[73\]
+ sky130_fd_sc_hd__dfstp_1
X_2878_ clknet_leaf_29_clk _0140_ net192 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_1829_ _1198_ LE_0A.dff_out vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__or2_1
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_35_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2801_ clknet_leaf_6_clk _0063_ net196 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2663_ CB_0.config_dataA\[5\] net168 net245 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__mux2_1
X_1614_ net1 _0401_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__and2b_1
X_2732_ net284 net290 net254 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__mux2_1
X_2594_ SB0.route_sel\[48\] SB0.route_sel\[47\] net230 vssd1 vssd1 vccd1 vccd1 _0184_
+ sky130_fd_sc_hd__mux2_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_4
X_1476_ _1226_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__nand2_1
Xfanout229 net230 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_4
Xfanout207 net209 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_1545_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] _1287_ vssd1 vssd1 vccd1 vccd1
+ _0334_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_59_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2028_ net132 net127 net123 net120 LEI0.config_data\[18\] LEI0.config_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__mux4_1
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3000_ clknet_leaf_8_clk _0262_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xinput7 CBeast_in[2] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2646_ SB0.route_sel\[100\] SB0.route_sel\[99\] net260 vssd1 vssd1 vccd1 vccd1 _0236_
+ sky130_fd_sc_hd__mux2_1
X_2715_ CB_1.config_dataA\[17\] CB_1.config_dataA\[16\] net252 vssd1 vssd1 vccd1 vccd1
+ _0305_ sky130_fd_sc_hd__mux2_1
X_2577_ SB0.route_sel\[31\] SB0.route_sel\[30\] net230 vssd1 vssd1 vccd1 vccd1 _0167_
+ sky130_fd_sc_hd__mux2_1
X_1528_ SB0.route_sel\[108\] SB0.route_sel\[109\] net47 _1321_ vssd1 vssd1 vccd1 vccd1
+ _1322_ sky130_fd_sc_hd__and4_1
X_1459_ net137 _1251_ _1252_ net120 vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__a22oi_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2431_ net346 LEI0.config_data\[21\] net268 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__mux2_1
X_2500_ LE_0B.reset_val LE_0B.edge_mode net231 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__mux2_1
X_2293_ net135 _1053_ _0379_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__mux2_1
X_2362_ _0371_ _1094_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_23 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _1219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2629_ SB0.route_sel\[83\] SB0.route_sel\[82\] net232 vssd1 vssd1 vccd1 vccd1 _0219_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ clknet_leaf_26_clk _0242_ net216 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[106\]
+ sky130_fd_sc_hd__dfstp_1
Xinput21 CBnorth_in[2] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
X_1793_ _1195_ net165 vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__nor2_1
Xinput10 CBeast_in[5] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_2
X_1931_ net155 _0472_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__nand2_1
X_1862_ net23 net24 net25 net26 net163 net161 vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__mux4_1
Xinput43 SBwest_in[0] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_1
Xinput32 SBsouth_in[12] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_1
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput54 SBwest_in[7] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
X_2414_ net341 net331 net266 vssd1 vssd1 vccd1 vccd1 _0006_ sky130_fd_sc_hd__mux2_1
X_2276_ _0457_ _1044_ _0459_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__a21o_1
XFILLER_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2345_ _1152_ SB0.route_sel\[50\] vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2061_ CB_1.config_dataA\[9\] CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0846_
+ sky130_fd_sc_hd__nand2b_1
X_2130_ net183 _0768_ _0910_ _0911_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__a211o_1
XFILLER_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2963_ clknet_leaf_4_clk _0225_ net202 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[89\]
+ sky130_fd_sc_hd__dfstp_1
X_1914_ _0700_ vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__inv_2
X_1776_ net167 _1330_ _0564_ _1194_ net166 vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__a2111o_1
X_1845_ net16 net17 net159 vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__mux2_1
X_2894_ clknet_leaf_31_clk _0156_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2328_ _1165_ SB0.route_sel\[75\] _1167_ _1168_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_40_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2259_ net184 LE_0A.reset_mode vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_4_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1630_ net177 net171 net173 net175 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__or4b_1
X_1492_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__inv_2
X_1561_ CB_0.config_dataA\[3\] _0348_ _0349_ _1332_ vssd1 vssd1 vccd1 vccd1 _0350_
+ sky130_fd_sc_hd__o22ai_1
X_2044_ net2 net144 _0822_ _0828_ _0820_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__o32a_1
X_2113_ _0896_ _0897_ _0814_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__mux2_1
X_2877_ clknet_leaf_25_clk _0139_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_2946_ clknet_leaf_3_clk _0208_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[72\]
+ sky130_fd_sc_hd__dfstp_1
X_1759_ net21 _0524_ _0525_ net22 _1190_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__o221a_1
X_1828_ LE_0A.dff0_out LE_0A.dff1_out LE_0A.reset_val vssd1 vssd1 vccd1 vccd1 LE_0A.dff_out
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2800_ clknet_leaf_6_clk net324 net196 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2731_ net290 net340 net254 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__mux2_1
X_1544_ net134 _0331_ _0332_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__mux2_1
X_2662_ net169 CB_0.config_dataA\[3\] net246 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__mux2_1
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1613_ net121 _0401_ _0361_ _1287_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__a2bb2o_1
X_2593_ SB0.route_sel\[47\] SB0.route_sel\[46\] net228 vssd1 vssd1 vccd1 vccd1 _0183_
+ sky130_fd_sc_hd__mux2_1
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_4
X_1475_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1269_
+ sky130_fd_sc_hd__and2b_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2027_ CB_1.config_dataA\[6\] _0789_ _0798_ _0811_ vssd1 vssd1 vccd1 vccd1 _0812_
+ sky130_fd_sc_hd__nor4_1
X_2929_ clknet_leaf_28_clk _0191_ net193 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[55\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 CBeast_in[3] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_2
X_2714_ CB_1.config_dataA\[16\] CB_1.config_dataA\[15\] net259 vssd1 vssd1 vccd1 vccd1
+ _0304_ sky130_fd_sc_hd__mux2_1
X_2645_ SB0.route_sel\[99\] SB0.route_sel\[98\] net260 vssd1 vssd1 vccd1 vccd1 _0235_
+ sky130_fd_sc_hd__mux2_1
X_2576_ SB0.route_sel\[30\] SB0.route_sel\[29\] net229 vssd1 vssd1 vccd1 vccd1 _0166_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1527_ net119 SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__nand2_1
X_1389_ SB0.route_sel\[102\] vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__inv_2
X_1458_ net171 net173 net175 net178 vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__and4b_1
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3059_ clknet_leaf_24_clk _0321_ net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_56_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2430_ LEI0.config_data\[21\] LEI0.config_data\[20\] net268 vssd1 vssd1 vccd1 vccd1
+ _0022_ sky130_fd_sc_hd__mux2_1
XFILLER_41_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2361_ SB0.route_sel\[26\] _1140_ _1141_ SB0.route_sel\[29\] _1093_ vssd1 vssd1 vccd1
+ vccd1 _1094_ sky130_fd_sc_hd__a221o_1
X_2292_ net127 _0377_ _1052_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_47_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_13 net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_24 net108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _1244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2559_ SB0.route_sel\[13\] SB0.route_sel\[12\] net234 vssd1 vssd1 vccd1 vccd1 _0149_
+ sky130_fd_sc_hd__mux2_1
X_2628_ SB0.route_sel\[82\] SB0.route_sel\[81\] net232 vssd1 vssd1 vccd1 vccd1 _0218_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1930_ net153 _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput22 CBnorth_in[3] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_2
X_1792_ _0556_ _0580_ _0555_ vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__mux2_1
Xinput11 CBeast_in[6] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_2
X_1861_ _0644_ _0647_ CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__a21oi_1
Xinput44 SBwest_in[10] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
Xinput33 SBsouth_in[13] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_1
XFILLER_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput55 SBwest_in[8] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
X_2413_ net331 LEI0.config_data\[3\] net266 vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__mux2_1
X_2344_ _1081_ _1082_ _1241_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__o21a_1
X_2275_ _0456_ _0472_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2060_ _0756_ _0759_ _0753_ _0750_ CB_1.config_dataA\[9\] net140 vssd1 vssd1 vccd1
+ vccd1 _0845_ sky130_fd_sc_hd__mux4_1
X_1913_ _0682_ _0685_ _0687_ LEI0.config_data\[29\] _0699_ vssd1 vssd1 vccd1 vccd1
+ _0700_ sky130_fd_sc_hd__o221a_1
X_2962_ clknet_leaf_5_clk _0224_ net202 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[88\]
+ sky130_fd_sc_hd__dfstp_1
X_2893_ clknet_leaf_30_clk _0155_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_1775_ net167 _0346_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__nor2_1
X_1844_ net15 net20 net21 net22 net160 CB_0.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1
+ _0631_ sky130_fd_sc_hd__mux4_1
X_2327_ SB0.route_sel\[73\] _1169_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__nor2_1
X_2258_ _1216_ LE_1B.dff_out _1039_ _0616_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outB sky130_fd_sc_hd__o211a_1
X_2189_ net179 _1214_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nor2_1
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ net18 net19 net170 vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__mux2_1
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2112_ LE_1A.config_data\[3\] LE_1A.config_data\[2\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0897_ sky130_fd_sc_hd__mux2_1
X_1491_ _1282_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__or2_4
X_2043_ net13 net14 net144 vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__mux2_1
X_2876_ clknet_leaf_25_clk _0138_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_1827_ net227 net185 vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__and2b_2
X_2945_ clknet_leaf_3_clk _0207_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[71\]
+ sky130_fd_sc_hd__dfstp_1
X_1758_ net15 net20 net168 vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__mux2_1
X_1689_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] _0437_ vssd1 vssd1 vccd1 vccd1
+ _0478_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2661_ CB_0.config_dataA\[3\] CB_0.config_dataA\[2\] net246 vssd1 vssd1 vccd1 vccd1
+ _0251_ sky130_fd_sc_hd__mux2_1
X_2730_ net340 net360 net254 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1543_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1298_ vssd1 vssd1 vccd1 vccd1
+ _0332_ sky130_fd_sc_hd__nand3_1
X_1474_ net24 net128 _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__mux2_1
Xfanout209 net216 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_4
X_1612_ net175 net177 net171 net173 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__or4_1
X_2592_ SB0.route_sel\[46\] SB0.route_sel\[45\] net227 vssd1 vssd1 vccd1 vccd1 _0182_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2026_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\] _0810_ _0809_ vssd1 vssd1 vccd1
+ vccd1 _0811_ sky130_fd_sc_hd__a31o_1
X_2859_ clknet_leaf_19_clk _0121_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2928_ clknet_leaf_30_clk _0190_ net193 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[54\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_28_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 CBeast_in[4] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_2
X_2644_ SB0.route_sel\[98\] SB0.route_sel\[97\] net260 vssd1 vssd1 vccd1 vccd1 _0234_
+ sky130_fd_sc_hd__mux2_1
X_2713_ CB_1.config_dataA\[15\] CB_1.config_dataA\[14\] net259 vssd1 vssd1 vccd1 vccd1
+ _0303_ sky130_fd_sc_hd__mux2_1
X_2575_ SB0.route_sel\[29\] SB0.route_sel\[28\] net229 vssd1 vssd1 vccd1 vccd1 _0165_
+ sky130_fd_sc_hd__mux2_1
X_1457_ CB_1.config_dataA\[17\] CB_1.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1251_
+ sky130_fd_sc_hd__and2_2
X_1526_ _1315_ _1317_ _1318_ _1319_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__a211o_1
X_1388_ SB0.route_sel\[103\] vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__inv_2
X_3058_ clknet_leaf_23_clk _0320_ net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2009_ SB0.route_sel\[68\] SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2291_ _0393_ _0377_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__nand2b_1
X_2360_ SB0.route_sel\[25\] SB0.route_sel\[24\] vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nor2_1
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_14 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_25 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_36 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 SBwest_out[1] sky130_fd_sc_hd__buf_2
X_2627_ SB0.route_sel\[81\] SB0.route_sel\[80\] net238 vssd1 vssd1 vccd1 vccd1 _0217_
+ sky130_fd_sc_hd__mux2_1
X_1509_ _1300_ _1301_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__a21o_1
X_2489_ net312 net307 net240 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__mux2_1
X_2558_ SB0.route_sel\[12\] SB0.route_sel\[11\] net234 vssd1 vssd1 vccd1 vccd1 _0148_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ _1244_ _0645_ _0646_ _1264_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_26_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
Xinput23 CBnorth_in[4] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_2
X_1791_ LE_0A.config_data\[5\] LE_0A.config_data\[4\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0580_ sky130_fd_sc_hd__mux2_1
Xinput12 CBeast_in[7] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_2
Xinput45 SBwest_in[11] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_1
Xinput34 SBsouth_in[1] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
Xinput56 SBwest_in[9] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
X_2412_ net369 LEI0.config_data\[2\] net266 vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__mux2_1
X_2274_ net133 _1043_ _0503_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__mux2_1
X_2343_ SB0.route_sel\[49\] SB0.route_sel\[48\] _1152_ SB0.route_sel\[50\] vssd1 vssd1
+ vccd1 vccd1 _1082_ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_50_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1989_ CB_1.config_dataA\[7\] _0760_ _0770_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1912_ _0689_ _0691_ _0698_ CB_0.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _0699_
+ sky130_fd_sc_hd__a31o_1
X_1843_ net159 _0472_ _0620_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a211o_1
X_2961_ clknet_leaf_5_clk _0223_ net198 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[87\]
+ sky130_fd_sc_hd__dfstp_1
X_2892_ clknet_leaf_30_clk _0154_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_1774_ _1192_ _0562_ CB_0.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2326_ _1069_ _1070_ _0469_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__o21a_1
X_2257_ LE_1B.dff0_out LE_1B.dff1_out LE_1B.reset_val vssd1 vssd1 vccd1 vccd1 LE_1B.dff_out
+ sky130_fd_sc_hd__mux2_1
X_2188_ net180 _0768_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1490_ _1149_ SB0.route_sel\[45\] _1150_ SB0.route_sel\[46\] _1283_ vssd1 vssd1 vccd1
+ vccd1 _1284_ sky130_fd_sc_hd__o221a_1
X_2042_ net3 _1203_ _0822_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__or3_1
Xhold1 LE_0B.config_data\[12\] vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ LE_1A.config_data\[1\] LE_1A.config_data\[0\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0896_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1826_ _0614_ _0607_ _0603_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__mux2_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2875_ clknet_leaf_25_clk _0137_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2944_ clknet_leaf_3_clk _0206_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[70\]
+ sky130_fd_sc_hd__dfstp_1
X_1757_ net27 net28 net16 net17 net168 CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0546_ sky130_fd_sc_hd__mux4_1
X_1688_ net17 net131 _0476_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ net125 net137 _1251_ _1253_ _1061_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1611_ _0397_ _0398_ _0399_ vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__a21o_1
X_2660_ CB_0.config_dataA\[2\] CB_0.config_dataA\[1\] net246 vssd1 vssd1 vccd1 vccd1
+ _0250_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1473_ net149 net145 net147 net151 vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__and4bb_1
X_1542_ net18 net130 _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__mux2_1
X_2591_ SB0.route_sel\[45\] SB0.route_sel\[44\] net227 vssd1 vssd1 vccd1 vccd1 _0181_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2025_ _0804_ _0801_ net142 vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__mux2_1
X_2927_ clknet_leaf_28_clk _0189_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[53\]
+ sky130_fd_sc_hd__dfstp_1
X_2789_ clknet_leaf_7_clk _0051_ net199 vssd1 vssd1 vccd1 vccd1 LE_0A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1809_ CB_0.config_dataA\[15\] _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__nor2_1
X_2858_ clknet_leaf_19_clk _0120_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2643_ SB0.route_sel\[97\] SB0.route_sel\[96\] net247 vssd1 vssd1 vccd1 vccd1 _0233_
+ sky130_fd_sc_hd__mux2_1
X_2574_ SB0.route_sel\[28\] SB0.route_sel\[27\] net234 vssd1 vssd1 vccd1 vccd1 _0164_
+ sky130_fd_sc_hd__mux2_1
X_2712_ CB_1.config_dataA\[14\] CB_1.config_dataA\[13\] net259 vssd1 vssd1 vccd1 vccd1
+ _0302_ sky130_fd_sc_hd__mux2_1
X_1456_ _1248_ net133 _1249_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__mux2_1
X_1387_ SB0.route_sel\[101\] vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__inv_2
X_1525_ SB0.route_sel\[106\] SB0.route_sel\[107\] vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__and2_1
X_2008_ _0469_ _0791_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__nand2_2
X_3057_ clknet_leaf_23_clk _0319_ net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2290_ net133 _1051_ _0417_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__mux2_1
XANTENNA_37 net89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 SBwest_out[2] sky130_fd_sc_hd__buf_2
X_2557_ SB0.route_sel\[11\] SB0.route_sel\[10\] net234 vssd1 vssd1 vccd1 vccd1 _0147_
+ sky130_fd_sc_hd__mux2_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 SBsouth_out[5] sky130_fd_sc_hd__buf_2
X_2626_ SB0.route_sel\[80\] SB0.route_sel\[79\] net238 vssd1 vssd1 vccd1 vccd1 _0216_
+ sky130_fd_sc_hd__mux2_1
X_1508_ net135 _1226_ _1298_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__and3_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2488_ net307 LE_0B.config_data\[5\] net240 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__mux2_1
X_1439_ net137 _1231_ _1232_ net121 vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_53_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1790_ _1191_ _0578_ _0577_ _0568_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a211o_1
Xinput13 CBeast_in[8] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_2
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput24 CBnorth_in[5] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_2
Xinput57 config_data_in vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
X_2411_ LEI0.config_data\[2\] net363 net266 vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__mux2_1
Xinput46 SBwest_in[12] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
Xinput35 SBsouth_in[2] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_1
X_2273_ _0517_ net129 _0501_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2342_ SB0.route_sel\[52\] _1153_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1988_ CB_1.config_dataA\[7\] _0771_ _0772_ _0765_ vssd1 vssd1 vccd1 vccd1 _0773_
+ sky130_fd_sc_hd__o22ai_1
X_2609_ SB0.route_sel\[63\] SB0.route_sel\[62\] net236 vssd1 vssd1 vccd1 vccd1 _0199_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout190 net205 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2960_ clknet_leaf_2_clk _0222_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[86\]
+ sky130_fd_sc_hd__dfstp_1
X_1911_ _0518_ _0684_ _0692_ _0697_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__o211a_1
X_1773_ _1307_ _1285_ net167 vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__mux2_1
X_1842_ net159 _0453_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__nor2_1
X_2891_ clknet_leaf_30_clk _0153_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_2325_ SB0.route_sel\[76\] _1166_ SB0.route_sel\[73\] SB0.route_sel\[72\] vssd1 vssd1
+ vccd1 vccd1 _1070_ sky130_fd_sc_hd__o22ai_1
X_2187_ net180 _0763_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__or2_1
X_2256_ _1030_ _1038_ LE_1B.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__a21o_1
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2041_ _1203_ _0822_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__nor2_1
Xhold2 _0085_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
X_2110_ _1205_ _0878_ _0880_ _0894_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_60_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2943_ clknet_leaf_28_clk _0205_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[69\]
+ sky130_fd_sc_hd__dfstp_1
X_1756_ _0517_ _0524_ _0525_ _0492_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1
+ _0545_ sky130_fd_sc_hd__o221a_1
X_1825_ _0613_ _0610_ _0579_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__mux2_1
XFILLER_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2874_ clknet_leaf_25_clk _0136_ net208 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_1687_ net148 net146 net152 net150 vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_13_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2308_ _1252_ _0750_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__nand2b_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2239_ CB_1.config_dataB\[15\] _1014_ _1021_ _1013_ vssd1 vssd1 vccd1 vccd1 _1022_
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1610_ net132 _0395_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__nor2_1
X_2590_ SB0.route_sel\[44\] SB0.route_sel\[43\] net228 vssd1 vssd1 vccd1 vccd1 _0180_
+ sky130_fd_sc_hd__mux2_1
X_1541_ net150 net152 net146 net148 vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and4bb_1
XFILLER_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1472_ SB0.route_sel\[41\] SB0.route_sel\[40\] vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__nand2_1
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ _0765_ _0806_ _0808_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__o21a_1
X_2857_ clknet_leaf_19_clk _0119_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[3\]
+ sky130_fd_sc_hd__dfstp_2
X_2926_ clknet_leaf_3_clk _0188_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[52\]
+ sky130_fd_sc_hd__dfstp_1
X_1739_ net23 net24 net168 vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__mux2_1
X_1808_ net15 net20 net21 net22 net165 net164 vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__mux4_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2788_ LE_0B.sel_clk _0050_ net61 vssd1 vssd1 vccd1 vccd1 LE_0B.dff1_out sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_36_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2711_ CB_1.config_dataA\[13\] net138 net259 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__mux2_1
X_2642_ SB0.route_sel\[96\] SB0.route_sel\[95\] net247 vssd1 vssd1 vccd1 vccd1 _0232_
+ sky130_fd_sc_hd__mux2_1
X_2573_ SB0.route_sel\[27\] SB0.route_sel\[26\] net234 vssd1 vssd1 vccd1 vccd1 _0163_
+ sky130_fd_sc_hd__mux2_1
X_1524_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] net125 _1272_ vssd1 vssd1
+ vccd1 vccd1 _1318_ sky130_fd_sc_hd__and4_1
X_1455_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] _1226_ vssd1 vssd1 vccd1 vccd1
+ _1249_ sky130_fd_sc_hd__and3_1
X_1386_ SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__inv_2
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2007_ _0469_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__and2_1
X_3056_ clknet_leaf_24_clk _0318_ net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ clknet_leaf_3_clk _0171_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_47_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_38 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1507_ net23 _1299_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__nand2b_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 SBwest_out[3] sky130_fd_sc_hd__buf_2
X_2487_ net309 net281 net240 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__mux2_1
X_2556_ SB0.route_sel\[10\] SB0.route_sel\[9\] net234 vssd1 vssd1 vccd1 vccd1 _0146_
+ sky130_fd_sc_hd__mux2_1
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 SBsouth_out[6] sky130_fd_sc_hd__buf_2
X_2625_ SB0.route_sel\[79\] SB0.route_sel\[78\] net237 vssd1 vssd1 vccd1 vccd1 _0215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1369_ net41 vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__inv_2
X_1438_ net177 net172 net174 net175 vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__or4bb_1
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ clknet_leaf_21_clk _0301_ net215 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput25 CBnorth_in[6] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
Xinput14 CBeast_in[9] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_2
Xinput36 SBsouth_in[3] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
Xinput58 config_en vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
X_2410_ net363 LEI0.config_data\[0\] net266 vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__mux2_1
Xinput47 SBwest_in[13] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__dlymetal6s2s_1
X_2341_ _1079_ _1080_ _1261_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__o21a_1
X_2272_ _1042_ net135 _0478_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1987_ net4 net5 net142 vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__mux2_1
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2608_ SB0.route_sel\[62\] SB0.route_sel\[61\] net235 vssd1 vssd1 vccd1 vccd1 _0198_
+ sky130_fd_sc_hd__mux2_1
X_2539_ CB_1.config_dataB\[13\] CB_1.config_dataB\[12\] net258 vssd1 vssd1 vccd1 vccd1
+ _0129_ sky130_fd_sc_hd__mux2_1
XFILLER_11_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout180 CB_1.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout191 net193 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1910_ _0677_ _0694_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o21ai_1
X_2890_ clknet_leaf_29_clk _0152_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_1772_ CB_0.config_dataA\[11\] _0558_ _0560_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__o21ai_1
X_1841_ _0413_ _0431_ _0393_ _0374_ CB_0.config_dataB\[5\] net159 vssd1 vssd1 vccd1
+ vccd1 _0628_ sky130_fd_sc_hd__mux4_1
X_2324_ _1165_ SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__nor2_1
X_2255_ _0997_ _1037_ _1034_ _1025_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__a211o_1
X_2186_ _1212_ _0753_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_3_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2040_ CB_1.config_dataA\[3\] _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__or2_1
Xhold3 LE_0B.config_data\[2\] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2873_ clknet_leaf_25_clk _0135_ net208 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[19\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_17_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2942_ clknet_leaf_28_clk _0204_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[68\]
+ sky130_fd_sc_hd__dfstp_1
X_1755_ net169 _0473_ _0543_ CB_0.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1 _0544_
+ sky130_fd_sc_hd__a211o_1
X_1824_ _0611_ _0612_ _0555_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__mux2_1
X_1686_ SB0.route_sel\[88\] SB0.route_sel\[89\] vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__nand2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2307_ _0442_ _1060_ _0444_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__a21o_1
X_2238_ CB_1.config_dataB\[13\] CB_1.config_dataB\[15\] _1020_ _1018_ _1016_ vssd1
+ vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__a311o_1
X_2169_ net4 _1209_ _1211_ _0951_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1540_ SB0.route_sel\[96\] SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_30_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1471_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__inv_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2023_ CB_1.config_dataA\[7\] _0805_ _0807_ _0746_ vssd1 vssd1 vccd1 vccd1 _0808_
+ sky130_fd_sc_hd__o22a_1
X_1807_ _0413_ _0431_ _0393_ _0374_ net164 net165 vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__mux4_1
X_2856_ clknet_leaf_19_clk _0118_ net217 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_2925_ clknet_leaf_28_clk _0187_ net195 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[51\]
+ sky130_fd_sc_hd__dfstp_1
X_1738_ net25 _0524_ _0525_ net26 vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__o22a_1
X_1669_ net28 _0456_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__nand2b_1
X_2787_ LE_0A.sel_clk _0049_ net61 vssd1 vssd1 vccd1 vccd1 LE_0A.dff0_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2710_ net139 CB_1.config_dataA\[11\] net270 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__mux2_1
X_1454_ net26 net128 _1247_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__mux2_1
X_2641_ SB0.route_sel\[95\] SB0.route_sel\[94\] net247 vssd1 vssd1 vccd1 vccd1 _0231_
+ sky130_fd_sc_hd__mux2_1
X_2572_ SB0.route_sel\[26\] SB0.route_sel\[25\] net234 vssd1 vssd1 vccd1 vccd1 _0162_
+ sky130_fd_sc_hd__mux2_1
X_1523_ net5 net121 _1316_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__mux2_1
X_1385_ SB0.route_sel\[88\] vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__inv_2
X_3055_ clknet_leaf_24_clk net304 net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2006_ _1167_ SB0.route_sel\[78\] SB0.route_sel\[73\] _1169_ _0790_ vssd1 vssd1 vccd1
+ vccd1 _0791_ sky130_fd_sc_hd__a221o_2
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2839_ clknet_leaf_23_clk _0101_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2908_ clknet_leaf_2_clk _0170_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_29_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_39 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2624_ SB0.route_sel\[78\] SB0.route_sel\[77\] net237 vssd1 vssd1 vccd1 vccd1 _0214_
+ sky130_fd_sc_hd__mux2_1
X_1506_ _1226_ _1298_ _1299_ net131 vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__o2bb2a_1
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 SBwest_out[4] sky130_fd_sc_hd__buf_2
X_2486_ net281 net278 net240 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__mux2_1
X_2555_ SB0.route_sel\[9\] SB0.route_sel\[8\] net234 vssd1 vssd1 vccd1 vccd1 _0145_
+ sky130_fd_sc_hd__mux2_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 SBsouth_out[7] sky130_fd_sc_hd__buf_2
X_1437_ CB_1.config_dataA\[16\] CB_1.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1231_
+ sky130_fd_sc_hd__and2b_2
X_3038_ clknet_leaf_18_clk _0300_ net226 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_1368_ SB0.route_sel\[70\] vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__inv_2
Xinput26 CBnorth_in[7] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_2
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 CBnorth_in[0] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_2
Xinput59 le_clk vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_4
Xinput37 SBsouth_in[4] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_1
Xinput48 SBwest_in[1] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_2271_ _0492_ net130 _0476_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2340_ SB0.route_sel\[58\] _1156_ SB0.route_sel\[63\] SB0.route_sel\[62\] vssd1 vssd1
+ vccd1 vccd1 _1080_ sky130_fd_sc_hd__o22ai_1
X_1986_ net9 net10 net11 net12 net142 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0771_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2607_ SB0.route_sel\[61\] SB0.route_sel\[60\] net235 vssd1 vssd1 vccd1 vccd1 _0197_
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2469_ net299 net305 net243 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__mux2_1
X_2538_ CB_1.config_dataB\[12\] CB_1.config_dataB\[11\] net258 vssd1 vssd1 vccd1 vccd1
+ _0128_ sky130_fd_sc_hd__mux2_1
XFILLER_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout181 CB_1.config_dataB\[5\] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout170 CB_0.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
X_1840_ LEI0.config_data\[17\] _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__or2_2
X_1771_ net166 _1194_ _0559_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__or3_1
XFILLER_6_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2254_ _1035_ _1036_ _0966_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__mux2_1
X_2323_ net124 _1287_ _0361_ _1068_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__a31o_1
X_2185_ _1212_ _1304_ _0755_ net179 vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__a31o_1
X_1969_ SB0.route_sel\[36\] SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_3_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 _0075_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1823_ LE_0A.config_data\[9\] LE_0A.config_data\[8\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0612_ sky130_fd_sc_hd__mux2_1
X_2872_ clknet_leaf_25_clk _0134_ net208 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[18\]
+ sky130_fd_sc_hd__dfstp_1
X_2941_ clknet_leaf_27_clk _0203_ net209 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[67\]
+ sky130_fd_sc_hd__dfstp_1
X_1754_ net169 _0453_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and2b_1
X_1685_ _0469_ _0471_ _1135_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__a21o_1
XFILLER_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2306_ _0450_ _0795_ _0441_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__a21bo_1
X_2237_ _1019_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__inv_2
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2168_ net5 net182 net181 vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__a21o_1
X_2099_ net138 _0796_ vssd1 vssd1 vccd1 vccd1 _0884_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1470_ _1261_ _1263_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2022_ net2 net3 net143 vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__mux2_1
X_1806_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__inv_2
X_2786_ clknet_leaf_14_clk _0048_ net222 vssd1 vssd1 vccd1 vccd1 CB_0.config_data_inA
+ sky130_fd_sc_hd__dfrtp_1
X_2855_ clknet_leaf_20_clk _0117_ net209 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2924_ clknet_leaf_3_clk _0186_ net194 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[50\]
+ sky130_fd_sc_hd__dfstp_1
X_1668_ _1269_ _0437_ _0456_ net129 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__o2bb2a_1
X_1737_ _0525_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__inv_2
X_1599_ _0387_ _1134_ _0386_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ SB0.route_sel\[94\] SB0.route_sel\[93\] net247 vssd1 vssd1 vccd1 vccd1 _0230_
+ sky130_fd_sc_hd__mux2_1
X_1453_ net145 net147 net149 net151 vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__and4b_1
X_2571_ SB0.route_sel\[25\] SB0.route_sel\[24\] net229 vssd1 vssd1 vccd1 vccd1 _0161_
+ sky130_fd_sc_hd__mux2_1
X_1522_ net175 net178 net172 net174 vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__and4b_1
X_1384_ SB0.route_sel\[94\] vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__inv_2
X_2005_ SB0.route_sel\[76\] SB0.route_sel\[77\] vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__nor2_1
X_3054_ clknet_leaf_23_clk _0316_ net210 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2907_ clknet_leaf_0_clk _0169_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[33\]
+ sky130_fd_sc_hd__dfstp_1
X_2769_ clknet_leaf_15_clk _0031_ net225 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_2838_ clknet_leaf_23_clk _0100_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_29 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 SBwest_out[5] sky130_fd_sc_hd__buf_2
X_2623_ SB0.route_sel\[77\] SB0.route_sel\[76\] net237 vssd1 vssd1 vccd1 vccd1 _0213_
+ sky130_fd_sc_hd__mux2_1
X_2554_ SB0.route_sel\[8\] SB0.route_sel\[7\] net235 vssd1 vssd1 vccd1 vccd1 _0144_
+ sky130_fd_sc_hd__mux2_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 SBsouth_out[8] sky130_fd_sc_hd__buf_2
X_1505_ net149 net151 net146 net148 vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__or4b_1
X_2485_ net278 net274 net231 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__mux2_1
X_1436_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _1230_
+ sky130_fd_sc_hd__and2b_1
X_1367_ SB0.route_sel\[71\] vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__inv_2
X_3037_ clknet_leaf_17_clk _0299_ net226 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_52_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 CBnorth_in[10] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_2
Xinput27 CBnorth_in[8] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_2
Xinput38 SBsouth_in[5] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
Xinput49 SBwest_in[2] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
X_2270_ net134 _1041_ _0332_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1985_ net142 _0768_ _0765_ _0764_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__a211o_1
X_2606_ SB0.route_sel\[60\] SB0.route_sel\[59\] net235 vssd1 vssd1 vccd1 vccd1 _0196_
+ sky130_fd_sc_hd__mux2_1
X_2537_ CB_1.config_dataB\[11\] CB_1.config_dataB\[10\] net258 vssd1 vssd1 vccd1 vccd1
+ _0127_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2468_ net305 net319 net243 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__mux2_1
X_2399_ SB0.route_sel\[90\] _1175_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nor2_1
X_1419_ CB_1.config_dataB\[10\] vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__inv_2
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout182 CB_1.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout160 CB_0.config_dataB\[4\] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_2
Xfanout171 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout193 net205 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ net18 net19 CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__mux2_1
X_2253_ LE_1B.config_data\[1\] LE_1B.config_data\[0\] _0936_ vssd1 vssd1 vccd1 vccd1
+ _1036_ sky130_fd_sc_hd__mux2_1
X_2184_ LE_1B.config_data\[15\] LE_1B.config_data\[14\] _0936_ vssd1 vssd1 vccd1 vccd1
+ _0967_ sky130_fd_sc_hd__mux2_1
X_2322_ _0401_ _0784_ _0402_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__a21oi_1
X_1899_ net134 net131 net126 net122 LEI0.config_data\[27\] LEI0.config_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__mux4_1
XFILLER_33_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1968_ _1282_ _0752_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_3_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold5 LE_1B.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_17_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2940_ clknet_leaf_26_clk _0202_ net209 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[66\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_60_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1753_ _1189_ _0540_ _0541_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__a21oi_1
X_1822_ LE_0A.config_data\[11\] LE_0A.config_data\[10\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0611_ sky130_fd_sc_hd__mux2_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2871_ clknet_leaf_25_clk _0133_ net208 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_1684_ _0472_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__inv_2
X_2167_ net9 _1209_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__a21o_1
X_2305_ net125 _1272_ _0440_ _1059_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ net2 net3 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__mux2_1
X_2098_ _0784_ _0787_ _0781_ _0778_ CB_1.config_dataA\[13\] net138 vssd1 vssd1 vccd1
+ vccd1 _0883_ sky130_fd_sc_hd__mux4_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2021_ net13 net14 net142 vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__mux2_1
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2923_ clknet_leaf_0_clk _0185_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[49\]
+ sky130_fd_sc_hd__dfstp_1
X_1805_ net134 net130 net126 net122 LEI0.config_data\[36\] LEI0.config_data\[37\]
+ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__mux4_1
X_2785_ clknet_leaf_14_clk net352 net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_1736_ CB_0.config_dataA\[5\] net168 vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__nand2_1
X_2854_ clknet_leaf_20_clk _0116_ net209 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[0\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_17_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1667_ net149 net147 net145 net151 vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__or4bb_1
X_1598_ SB0.route_sel\[15\] SB0.route_sel\[14\] net48 vssd1 vssd1 vccd1 vccd1 _0387_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ CB_1.config_dataB\[12\] _0763_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2570_ SB0.route_sel\[24\] SB0.route_sel\[23\] net229 vssd1 vssd1 vccd1 vccd1 _0160_
+ sky130_fd_sc_hd__mux2_1
X_1383_ SB0.route_sel\[95\] vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__inv_2
X_1452_ SB0.route_sel\[57\] SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__nand2_1
X_1521_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] _1272_ vssd1 vssd1 vccd1 vccd1
+ _1315_ sky130_fd_sc_hd__nand3_1
X_2004_ CB_1.config_dataA\[7\] _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__nor2_1
X_3053_ clknet_leaf_24_clk net283 net213 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2906_ clknet_leaf_0_clk _0168_ net187 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2768_ clknet_leaf_14_clk _0030_ net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_2699_ CB_1.config_dataA\[1\] net144 net260 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__mux2_1
X_2837_ clknet_leaf_23_clk _0099_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1719_ SB0.route_sel\[82\] SB0.route_sel\[83\] vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__nand2_1
XFILLER_41_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_19 net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1504_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] vssd1 vssd1 vccd1 vccd1 _1298_
+ sky130_fd_sc_hd__nor2_1
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 SBwest_out[6] sky130_fd_sc_hd__buf_2
X_2622_ SB0.route_sel\[76\] SB0.route_sel\[75\] net237 vssd1 vssd1 vccd1 vccd1 _0212_
+ sky130_fd_sc_hd__mux2_1
X_2553_ SB0.route_sel\[7\] SB0.route_sel\[6\] net235 vssd1 vssd1 vccd1 vccd1 _0143_
+ sky130_fd_sc_hd__mux2_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 SBsouth_out[9] sky130_fd_sc_hd__buf_2
X_1435_ net133 _1225_ _1228_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__mux2_1
X_1366_ SB0.route_sel\[69\] vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__inv_2
X_2484_ net274 LE_0B.config_data\[1\] net231 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__mux2_1
X_3036_ clknet_leaf_17_clk _0298_ net226 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_43_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_52_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 CBnorth_in[11] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
Xinput28 CBnorth_in[9] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_2
Xinput39 SBsouth_in[6] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_9_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1984_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__inv_2
X_2467_ net319 net325 net243 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__mux2_1
X_2605_ SB0.route_sel\[59\] SB0.route_sel\[58\] net252 vssd1 vssd1 vccd1 vccd1 _0195_
+ sky130_fd_sc_hd__mux2_1
X_2536_ CB_1.config_dataB\[10\] net179 net258 vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2398_ _1117_ _1118_ _0489_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__o21a_1
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1349_ SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__inv_2
X_1418_ net180 vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__inv_2
X_3019_ clknet_leaf_10_clk _0281_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[13\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_5_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout150 CB_0.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_1
Xfanout161 CB_0.config_dataB\[1\] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout183 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout172 CB_1.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_1
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2321_ _0382_ _1067_ _0384_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__a21o_1
X_2183_ _0954_ _0955_ _0965_ _0937_ LEI0.config_data\[23\] vssd1 vssd1 vccd1 vccd1
+ _0966_ sky130_fd_sc_hd__o32a_2
X_2252_ LE_1B.config_data\[3\] LE_1B.config_data\[2\] _0936_ vssd1 vssd1 vccd1 vccd1
+ _1035_ sky130_fd_sc_hd__mux2_1
XFILLER_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1898_ CB_0.config_dataB\[10\] _0684_ vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__nand2_1
X_1967_ SB0.route_sel\[44\] SB0.route_sel\[45\] SB0.route_sel\[47\] _1151_ _0751_
+ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__o221a_1
X_2519_ net335 LE_1A.config_data\[13\] net258 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold6 _0310_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2870_ clknet_leaf_20_clk _0132_ net214 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataB\[16\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_17_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1752_ _0431_ _0523_ _0526_ _0374_ CB_0.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1
+ _0541_ sky130_fd_sc_hd__a221o_1
X_1821_ _0608_ _0609_ _0555_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1683_ _0469_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__nand2_2
X_2304_ _0461_ _0793_ _0462_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__a21oi_1
X_2097_ _0881_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__inv_2
X_2166_ net10 net182 CB_1.config_dataB\[7\] net181 vssd1 vssd1 vccd1 vccd1 _0949_
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _1003_ _1017_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__nor2_1
X_2999_ clknet_leaf_8_clk _0261_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[13\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2020_ net1 net6 net7 net8 net143 CB_1.config_dataA\[5\] vssd1 vssd1 vccd1 vccd1
+ _0805_ sky130_fd_sc_hd__mux4_1
X_2853_ LE_1B.sel_clk _0115_ net61 vssd1 vssd1 vccd1 vccd1 LE_1B.dff0_out sky130_fd_sc_hd__dfrtp_1
X_2922_ clknet_leaf_0_clk _0184_ net187 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[48\]
+ sky130_fd_sc_hd__dfstp_1
X_1735_ _1189_ net168 vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__or2_1
X_1804_ CB_0.config_dataA\[15\] _0582_ _0586_ _0592_ _1196_ vssd1 vssd1 vccd1 vccd1
+ _0593_ sky130_fd_sc_hd__a221o_1
X_2784_ clknet_leaf_14_clk _0046_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_1666_ SB0.route_sel\[73\] SB0.route_sel\[72\] vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__nand2_1
X_1597_ SB0.route_sel\[12\] SB0.route_sel\[13\] vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__nand2_1
X_2218_ net132 _1219_ _1220_ _1221_ LEI0.config_data\[45\] LEI0.config_data\[46\]
+ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__mux4_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2149_ _0919_ _0929_ _0931_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__o21a_1
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1520_ net135 _1310_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__nand2_1
X_1451_ _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__inv_2
X_1382_ SB0.route_sel\[93\] vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__inv_2
XFILLER_35_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _0784_ _0787_ _0781_ _0778_ CB_1.config_dataA\[5\] net142 vssd1 vssd1 vccd1
+ vccd1 _0788_ sky130_fd_sc_hd__mux4_1
X_3052_ clknet_leaf_24_clk net287 net213 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2836_ clknet_leaf_23_clk _0098_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2905_ clknet_leaf_0_clk _0167_ net187 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[31\]
+ sky130_fd_sc_hd__dfstp_1
X_1649_ _1298_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__nand2_1
X_2767_ clknet_leaf_14_clk net355 net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_2698_ net144 net146 net261 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__mux2_1
X_1718_ net2 _0505_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__nor2_1
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 SBwest_out[7] sky130_fd_sc_hd__buf_2
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 SBwest_out[0] sky130_fd_sc_hd__buf_2
X_2621_ SB0.route_sel\[75\] SB0.route_sel\[74\] net253 vssd1 vssd1 vccd1 vccd1 _0211_
+ sky130_fd_sc_hd__mux2_1
X_2552_ SB0.route_sel\[6\] SB0.route_sel\[5\] net235 vssd1 vssd1 vccd1 vccd1 _0142_
+ sky130_fd_sc_hd__mux2_1
X_1503_ SB0.route_sel\[35\] SB0.route_sel\[34\] _1296_ _1293_ vssd1 vssd1 vccd1 vccd1
+ _1297_ sky130_fd_sc_hd__a31oi_1
X_2483_ net349 LE_0B.config_data\[0\] net231 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__mux2_1
X_1434_ _1226_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__nand2_1
X_3035_ clknet_leaf_16_clk _0297_ net226 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_1365_ SB0.route_sel\[67\] vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__inv_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2819_ clknet_leaf_6_clk _0081_ net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 CBnorth_in[12] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput29 SBsouth_in[0] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2604_ SB0.route_sel\[58\] SB0.route_sel\[57\] net250 vssd1 vssd1 vccd1 vccd1 _0194_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_21_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1983_ _1325_ _1326_ _0767_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__or3_4
X_2466_ net325 net329 net243 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__mux2_1
X_1417_ CB_1.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__inv_2
X_2535_ net179 net180 net258 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3018_ clknet_leaf_10_clk _0280_ net205 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_2397_ SB0.route_sel\[88\] SB0.route_sel\[89\] SB0.route_sel\[90\] _1175_ vssd1 vssd1
+ vccd1 vccd1 _1118_ sky130_fd_sc_hd__a2bb2o_1
X_1348_ SB0.route_sel\[30\] vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__inv_2
XFILLER_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout151 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_2
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
Xfanout195 net205 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
Xfanout173 CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_4
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2320_ _0381_ _0781_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__nand2_1
X_2251_ _0966_ _1031_ _1032_ _1033_ _0998_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__o221a_1
X_2182_ CB_1.config_dataB\[7\] _0956_ _0958_ _0959_ _0964_ vssd1 vssd1 vccd1 vccd1
+ _0965_ sky130_fd_sc_hd__o221a_1
X_1966_ SB0.route_sel\[40\] SB0.route_sel\[41\] vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__nand2b_1
X_1897_ net157 _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__or2_1
X_2449_ net365 LEI0.config_data\[39\] net263 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__mux2_1
X_2518_ net377 LE_1A.config_data\[12\] net256 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7 LE_0B.config_data\[3\] vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_60_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1820_ LE_0A.config_data\[13\] LE_0A.config_data\[12\] _0522_ vssd1 vssd1 vccd1 vccd1
+ _0609_ sky130_fd_sc_hd__mux2_1
X_1751_ _0413_ _0393_ net169 vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__mux2_1
X_1682_ SB0.route_sel\[76\] _1166_ SB0.route_sel\[79\] _1168_ _0470_ vssd1 vssd1 vccd1
+ vccd1 _0471_ sky130_fd_sc_hd__a221o_1
X_2303_ _0506_ _1058_ _0509_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__o21ai_1
X_2234_ net13 net14 CB_1.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__mux2_1
X_2096_ net134 net130 net126 net122 LEI0.config_data\[42\] LEI0.config_data\[43\]
+ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__mux4_1
X_2165_ net12 _0943_ _0945_ net11 vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2998_ clknet_leaf_8_clk _0260_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_1949_ LE_0B.config_data\[13\] _0672_ _0642_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a21o_1
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1803_ _1244_ _0582_ _0588_ _0590_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__a221o_1
X_2783_ clknet_leaf_12_clk _0045_ net221 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_2921_ clknet_leaf_31_clk _0183_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[47\]
+ sky130_fd_sc_hd__dfstp_1
X_2852_ clknet_leaf_22_clk _0114_ net213 vssd1 vssd1 vccd1 vccd1 LE_1A.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1734_ _1189_ net168 vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__nor2_1
X_1665_ _0450_ _0452_ net170 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__a21o_1
X_1596_ SB0.route_sel\[11\] SB0.route_sel\[10\] _0382_ _0383_ _0384_ vssd1 vssd1 vccd1
+ vccd1 _0385_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2217_ _0967_ _0999_ _0966_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__mux2_1
X_2079_ _0853_ _0862_ _0863_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_36_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2148_ CB_1.config_dataB\[3\] _0927_ _0930_ _0911_ vssd1 vssd1 vccd1 vccd1 _0931_
+ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1450_ _1241_ _1243_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__nand2_4
X_1381_ SB0.route_sel\[91\] vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__inv_2
X_3051_ clknet_leaf_24_clk net311 net207 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2002_ _0785_ _0786_ _0428_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__a21bo_2
X_2766_ clknet_leaf_14_clk _0028_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_2835_ clknet_leaf_23_clk _0097_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2904_ clknet_leaf_0_clk _0166_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_2697_ net146 net148 net262 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__mux2_1
X_1648_ CB_0.config_dataA\[18\] CB_0.config_dataA\[19\] vssd1 vssd1 vccd1 vccd1 _0437_
+ sky130_fd_sc_hd__and2b_1
X_1717_ _1231_ _0440_ _0505_ net120 vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__a22o_1
X_1579_ SB0.route_sel\[31\] SB0.route_sel\[30\] _0367_ vssd1 vssd1 vccd1 vccd1 _0368_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2620_ SB0.route_sel\[74\] SB0.route_sel\[73\] net239 vssd1 vssd1 vccd1 vccd1 _0210_
+ sky130_fd_sc_hd__mux2_1
X_1433_ CB_0.config_dataA\[16\] CB_0.config_dataA\[17\] vssd1 vssd1 vccd1 vccd1 _1227_
+ sky130_fd_sc_hd__and2b_1
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 SBwest_out[8] sky130_fd_sc_hd__buf_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 SBwest_out[10] sky130_fd_sc_hd__buf_2
X_2551_ SB0.route_sel\[5\] SB0.route_sel\[4\] net235 vssd1 vssd1 vccd1 vccd1 _0141_
+ sky130_fd_sc_hd__mux2_1
X_2482_ net364 LE_1B.reset_mode net228 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__mux2_1
X_1502_ _1295_ _1146_ _1294_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__mux2_1
X_3034_ clknet_leaf_17_clk _0296_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_1364_ SB0.route_sel\[62\] vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__inv_2
X_2749_ clknet_leaf_14_clk _0011_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2818_ clknet_leaf_5_clk _0080_ net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 CBnorth_in[13] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1982_ SB0.route_sel\[108\] SB0.route_sel\[109\] SB0.route_sel\[104\] _1188_ _0766_
+ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o221a_1
X_2534_ CB_1.config_dataB\[8\] CB_1.config_dataB\[7\] net258 vssd1 vssd1 vccd1 vccd1
+ _0124_ sky130_fd_sc_hd__mux2_1
X_2603_ SB0.route_sel\[57\] SB0.route_sel\[56\] net235 vssd1 vssd1 vccd1 vccd1 _0193_
+ sky130_fd_sc_hd__mux2_1
X_2465_ net329 net343 net243 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__mux2_1
X_1416_ CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__inv_2
X_2396_ SB0.route_sel\[92\] _1176_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__nor2_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1347_ SB0.route_sel\[28\] vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__inv_2
X_3017_ clknet_leaf_8_clk _0279_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[11\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout152 CB_0.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_1
Xfanout163 CB_0.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout130 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xfanout141 CB_1.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_2
Xfanout174 CB_1.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ LE_1B.config_data\[4\] _0936_ _0966_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a21bo_1
X_2181_ _1211_ _0963_ _0962_ CB_1.config_dataB\[6\] vssd1 vssd1 vccd1 vccd1 _0964_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1965_ _0748_ _0749_ _1261_ vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__a21bo_2
X_1896_ CB_0.config_dataB\[9\] CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0683_
+ sky130_fd_sc_hd__nand2_1
X_2517_ LE_1A.config_data\[12\] LE_1A.config_data\[11\] net256 vssd1 vssd1 vccd1 vccd1
+ _0107_ sky130_fd_sc_hd__mux2_1
X_2448_ net376 net361 net263 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__mux2_1
X_2379_ SB0.route_sel\[3\] _1127_ SB0.route_sel\[4\] _1128_ vssd1 vssd1 vccd1 vccd1
+ _1106_ sky130_fd_sc_hd__o22a_1
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold8 LE_1A.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
X_1750_ LEI0.config_data\[14\] _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__nor2_2
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1681_ SB0.route_sel\[74\] SB0.route_sel\[75\] vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__nor2_1
X_2164_ _0750_ _0944_ _0946_ _0759_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__a22oi_1
X_2302_ _0505_ _0804_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__nor2_1
X_2233_ CB_1.config_dataB\[15\] _1015_ vssd1 vssd1 vccd1 vccd1 _1016_ sky130_fd_sc_hd__nor2_1
X_2095_ net139 _0879_ vssd1 vssd1 vccd1 vccd1 _0880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2997_ clknet_leaf_6_clk _0259_ net199 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_1879_ net27 net28 net16 net17 net163 net161 vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__mux4_1
X_1948_ LE_0B.config_data\[12\] _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0735_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_39_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2920_ clknet_leaf_31_clk _0182_ net185 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_1802_ net164 CB_0.config_dataA\[12\] _1264_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__and3_1
X_2782_ clknet_leaf_12_clk _0044_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_1733_ _0354_ _0355_ _0521_ _1222_ LEI0.config_data\[2\] vssd1 vssd1 vccd1 vccd1
+ _0522_ sky130_fd_sc_hd__o32a_4
X_2851_ clknet_leaf_24_clk _0113_ net210 vssd1 vssd1 vccd1 vccd1 LE_1A.reset_val sky130_fd_sc_hd__dfrtp_1
X_1664_ _0450_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__and2_2
X_1595_ net124 _1272_ _0361_ vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__and3_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ net13 net14 net183 vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux2_1
X_2216_ LE_1B.config_data\[13\] LE_1B.config_data\[12\] _0936_ vssd1 vssd1 vccd1 vccd1
+ _0999_ sky130_fd_sc_hd__mux2_1
X_2078_ CB_1.config_dataA\[11\] _0860_ _0861_ _0846_ vssd1 vssd1 vccd1 vccd1 _0863_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1380_ SB0.route_sel\[80\] vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__inv_2
X_2001_ SB0.route_sel\[20\] SB0.route_sel\[21\] SB0.route_sel\[23\] _1138_ vssd1 vssd1
+ vccd1 vccd1 _0786_ sky130_fd_sc_hd__o22a_1
X_3050_ clknet_leaf_24_clk _0312_ net206 vssd1 vssd1 vccd1 vccd1 LE_1B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2903_ clknet_leaf_30_clk _0165_ net186 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[29\]
+ sky130_fd_sc_hd__dfstp_1
X_2696_ net148 net150 net262 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__mux2_1
X_2765_ clknet_leaf_14_clk _0027_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_2834_ clknet_leaf_23_clk _0096_ net211 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1716_ net178 net174 net172 net176 vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__and4bb_1
X_1647_ net130 net27 _0435_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__mux2_1
X_1578_ SB0.route_sel\[28\] SB0.route_sel\[29\] net50 vssd1 vssd1 vccd1 vccd1 _0367_
+ sky130_fd_sc_hd__and3_1
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 SBwest_out[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_30_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2550_ SB0.route_sel\[4\] SB0.route_sel\[3\] net235 vssd1 vssd1 vccd1 vccd1 _0140_
+ sky130_fd_sc_hd__mux2_1
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 SBwest_out[9] sky130_fd_sc_hd__buf_2
X_1432_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _1226_
+ sky130_fd_sc_hd__and2b_1
X_2481_ LE_1A.dff1_out _0907_ net60 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__mux2_1
X_1363_ SB0.route_sel\[61\] vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__inv_2
X_1501_ SB0.route_sel\[39\] SB0.route_sel\[38\] net51 vssd1 vssd1 vccd1 vccd1 _1295_
+ sky130_fd_sc_hd__a21bo_1
X_3033_ clknet_leaf_17_clk _0295_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_2
X_2748_ clknet_leaf_13_clk _0010_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_2679_ net161 net162 net242 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__mux2_1
X_2817_ clknet_leaf_5_clk net308 net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_44_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1981_ net119 SB0.route_sel\[110\] vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__nand2b_1
X_2533_ CB_1.config_dataB\[7\] CB_1.config_dataB\[6\] net265 vssd1 vssd1 vccd1 vccd1
+ _0123_ sky130_fd_sc_hd__mux2_1
X_2602_ SB0.route_sel\[56\] SB0.route_sel\[55\] net235 vssd1 vssd1 vccd1 vccd1 _0192_
+ sky130_fd_sc_hd__mux2_1
X_2464_ LE_0A.config_data\[4\] net338 net244 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__mux2_1
X_1415_ net182 vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__inv_2
X_2395_ _1115_ _1116_ _0343_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__o21a_1
X_1346_ SB0.route_sel\[27\] vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__inv_2
X_3016_ clknet_leaf_9_clk _0278_ net204 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[10\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_31_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout131 CB_0.le_outB vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_1
Xfanout120 _1221_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
Xfanout164 CB_0.config_dataA\[13\] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_2
Xfanout153 CB_0.config_dataB\[15\] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
Xfanout175 CB_1.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_22_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ net1 net6 net7 net8 CB_1.config_dataB\[4\] net181 vssd1 vssd1 vccd1 vccd1
+ _0963_ sky130_fd_sc_hd__mux4_1
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_1895_ CB_0.config_dataB\[11\] _0675_ _0678_ _0681_ vssd1 vssd1 vccd1 vccd1 _0682_
+ sky130_fd_sc_hd__o211a_1
X_1964_ SB0.route_sel\[60\] SB0.route_sel\[61\] SB0.route_sel\[63\] _1158_ vssd1 vssd1
+ vccd1 vccd1 _0749_ sky130_fd_sc_hd__o22a_1
X_2447_ net361 net344 net261 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__mux2_1
X_2516_ net381 net371 net256 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__mux2_1
X_2378_ SB0.route_sel\[0\] SB0.route_sel\[1\] vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__or2_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold9 _0110_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _0481_ _1057_ _0484_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__o21ai_1
X_1680_ _0465_ _0468_ _0455_ _0460_ vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__a2bb2o_2
X_2163_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__inv_2
X_2232_ net1 net6 net7 net8 CB_1.config_dataB\[12\] CB_1.config_dataB\[13\] vssd1
+ vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2094_ CB_1.config_dataA\[13\] CB_1.config_dataA\[15\] vssd1 vssd1 vccd1 vccd1 _0879_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2996_ clknet_leaf_6_clk _0258_ net199 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_1878_ net162 _0472_ _0652_ _0664_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__a211o_1
X_1947_ _0700_ _0731_ _0733_ _0729_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__a31o_1
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2850_ clknet_leaf_24_clk _0112_ net210 vssd1 vssd1 vccd1 vccd1 LE_1A.edge_mode sky130_fd_sc_hd__dfstp_1
X_1801_ net165 _1330_ _0589_ _1197_ net164 vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__a2111o_1
X_2781_ clknet_leaf_12_clk _0043_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_1732_ CB_0.config_dataA\[3\] _0433_ _0520_ vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__o21ba_1
X_1663_ SB0.route_sel\[68\] _1160_ SB0.route_sel\[71\] _1162_ _0451_ vssd1 vssd1 vccd1
+ vccd1 _0452_ sky130_fd_sc_hd__a221o_1
X_1594_ net6 _0381_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2077_ net2 net3 net140 vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__mux2_1
X_2146_ net2 net3 CB_1.config_dataB\[0\] vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__mux2_1
X_2215_ CB_1.config_dataB\[10\] _0980_ _0981_ _0983_ _0996_ vssd1 vssd1 vccd1 vccd1
+ _0998_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_36_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2979_ clknet_leaf_26_clk _0241_ net216 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[105\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2000_ SB0.route_sel\[16\] SB0.route_sel\[17\] vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__nand2b_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2833_ clknet_leaf_31_clk _0095_ net184 vssd1 vssd1 vccd1 vccd1 LE_1A.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2902_ clknet_leaf_30_clk _0164_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_2695_ net150 net152 net262 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__mux2_1
X_1646_ net149 net152 net147 net145 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__or4b_1
X_2764_ clknet_leaf_12_clk net359 net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_1715_ net136 _0502_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__mux2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1577_ _0363_ _0364_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__o21ba_1
X_2129_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__inv_2
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 SBwest_out[12] sky130_fd_sc_hd__buf_2
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 config_data_out sky130_fd_sc_hd__buf_2
X_2480_ LE_0B.dff0_out _1217_ _1125_ vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__a21o_1
X_1500_ SB0.route_sel\[36\] SB0.route_sel\[37\] vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__nand2_1
X_1431_ net25 net128 _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__mux2_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 CBnorth_out[9] sky130_fd_sc_hd__buf_2
X_1362_ SB0.route_sel\[59\] vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__inv_2
X_3032_ clknet_leaf_17_clk _0294_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_2816_ clknet_leaf_5_clk _0078_ net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1629_ net133 _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__mux2_1
X_2747_ clknet_leaf_13_clk _0009_ net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2678_ net163 CB_0.config_dataA\[19\] net248 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__mux2_1
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1980_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0765_
+ sky130_fd_sc_hd__nand2b_1
X_2463_ net338 net334 net244 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__mux2_1
X_2532_ CB_1.config_dataB\[6\] net181 net265 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__mux2_1
X_2601_ SB0.route_sel\[55\] SB0.route_sel\[54\] net236 vssd1 vssd1 vccd1 vccd1 _0191_
+ sky130_fd_sc_hd__mux2_1
X_3015_ clknet_leaf_7_clk _0277_ net201 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_2394_ SB0.route_sel\[98\] _1180_ _1182_ _1183_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__a2bb2o_1
X_1414_ net181 vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__inv_2
X_1345_ net35 vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__inv_2
Xfanout165 CB_0.config_dataA\[12\] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout132 _1218_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
Xfanout154 CB_0.config_dataB\[13\] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout143 CB_1.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_2
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout198 net201 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout187 net205 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout176 CB_1.config_dataB\[17\] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_25_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1894_ CB_0.config_dataB\[11\] _0679_ _0680_ _0677_ vssd1 vssd1 vccd1 vccd1 _0681_
+ sky130_fd_sc_hd__o22ai_1
X_1963_ SB0.route_sel\[56\] SB0.route_sel\[57\] vssd1 vssd1 vccd1 vccd1 _0748_ sky130_fd_sc_hd__nand2b_1
X_2446_ net344 LEI0.config_data\[36\] net261 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__mux2_1
X_2515_ net371 net327 net255 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__mux2_1
X_2377_ _1103_ _1104_ _0390_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__o21a_1
XFILLER_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ _0480_ _0801_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__nor2_1
X_2231_ _0781_ _0784_ _0778_ _0787_ _1215_ CB_1.config_dataB\[13\] vssd1 vssd1 vccd1
+ vccd1 _1014_ sky130_fd_sc_hd__mux4_1
X_2162_ CB_1.config_dataB\[5\] _1209_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nand2_1
X_2093_ CB_1.config_dataA\[15\] _0871_ _0876_ _0877_ _0875_ vssd1 vssd1 vccd1 vccd1
+ _0878_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2995_ clknet_leaf_6_clk _0257_ net199 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_1877_ net163 _0453_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nor2_1
X_1946_ LE_0B.config_data\[1\] _0672_ _0732_ _0642_ vssd1 vssd1 vccd1 vccd1 _0733_
+ sky130_fd_sc_hd__a211o_1
X_2429_ LEI0.config_data\[20\] net362 net268 vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__mux2_1
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1800_ CB_0.config_dataA\[12\] _0346_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ clknet_leaf_12_clk _0042_ net219 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_1731_ _0328_ _0454_ _0474_ _0493_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__a311o_1
X_1662_ SB0.route_sel\[67\] SB0.route_sel\[66\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__nor2_1
X_2214_ CB_1.config_dataB\[10\] _0980_ _0981_ _0983_ _0996_ vssd1 vssd1 vccd1 vccd1
+ _0997_ sky130_fd_sc_hd__a311oi_2
X_1593_ _1272_ _0361_ _0381_ net121 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2076_ net13 net14 net141 vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _1207_ _0919_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_28_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1929_ _0413_ _0431_ _0393_ _0374_ net154 net155 vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__mux4_1
X_2978_ clknet_leaf_27_clk _0240_ net209 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[104\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_12_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold90 LEI0.config_data\[38\] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__dlygate4sd3_1
X_2763_ clknet_leaf_16_clk _0025_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2832_ LE_1B.sel_clk _0094_ net61 vssd1 vssd1 vccd1 vccd1 LE_1B.dff1_out sky130_fd_sc_hd__dfstp_1
X_2901_ clknet_leaf_29_clk _0163_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_1714_ _1227_ _0437_ vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__nand2_1
X_2694_ net151 net153 net263 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__mux2_1
X_1576_ net124 _1251_ _0361_ SB0.route_sel\[27\] SB0.route_sel\[26\] vssd1 vssd1 vccd1
+ vccd1 _0365_ sky130_fd_sc_hd__a32o_1
X_1645_ SB0.route_sel\[65\] SB0.route_sel\[64\] vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__nand2_1
X_2128_ CB_1.config_dataB\[1\] CB_1.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0911_
+ sky130_fd_sc_hd__nand2b_1
X_2059_ LE_1A.config_data\[5\] LE_1A.config_data\[4\] _0843_ vssd1 vssd1 vccd1 vccd1
+ _0844_ sky130_fd_sc_hd__mux2_1
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1430_ net151 net145 net147 net149 vssd1 vssd1 vccd1 vccd1 _1224_ sky130_fd_sc_hd__and4bb_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 SBwest_out[13] sky130_fd_sc_hd__buf_2
X_3031_ clknet_leaf_17_clk _0293_ net221 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_2
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 CBnorth_out[12] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 SBsouth_out[0] sky130_fd_sc_hd__buf_2
X_1361_ SB0.route_sel\[49\] vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__inv_2
X_2746_ clknet_leaf_13_clk net357 net218 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2815_ clknet_leaf_5_clk _0077_ net196 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_2677_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] net263 vssd1 vssd1 vccd1 vccd1
+ _0267_ sky130_fd_sc_hd__mux2_1
X_1628_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1227_ vssd1 vssd1 vccd1 vccd1
+ _0417_ sky130_fd_sc_hd__or3b_1
X_1559_ net23 net24 net25 net26 net170 CB_0.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0348_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_43_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2600_ SB0.route_sel\[54\] SB0.route_sel\[53\] net236 vssd1 vssd1 vccd1 vccd1 _0190_
+ sky130_fd_sc_hd__mux2_1
X_2462_ net334 net320 net244 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__mux2_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2531_ net181 net182 net265 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__mux2_1
X_2393_ _1184_ SB0.route_sel\[97\] vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nor2_1
X_1413_ net183 vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__inv_2
X_3014_ clknet_leaf_6_clk _0276_ net197 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1344_ SB0.route_sel\[22\] vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__inv_2
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2729_ net360 net348 net254 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__mux2_1
Xfanout199 net201 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_57_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout133 net136 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_2
Xfanout144 CB_1.config_dataA\[0\] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
Xfanout166 CB_0.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout155 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout122 CB_1.le_outB vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout177 CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net190 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1962_ net142 _0746_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__nor2_1
X_1893_ net18 net19 net157 vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__mux2_1
X_2445_ LEI0.config_data\[36\] net375 net268 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__mux2_1
X_2514_ net327 net298 net255 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__mux2_1
X_2376_ _1131_ SB0.route_sel\[10\] SB0.route_sel\[15\] SB0.route_sel\[14\] vssd1 vssd1
+ vccd1 vccd1 _1104_ sky130_fd_sc_hd__o22ai_1
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ CB_1.config_dataB\[15\] _1012_ vssd1 vssd1 vccd1 vccd1 _1013_ sky130_fd_sc_hd__nand2_1
X_2161_ _0943_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__inv_2
X_2092_ net138 _0768_ _0873_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__a21o_1
X_2994_ clknet_leaf_7_clk _0256_ net200 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[8\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_16_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1945_ LE_0B.config_data\[0\] _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0732_
+ sky130_fd_sc_hd__and4_1
X_1876_ _0661_ _0662_ CB_0.config_dataB\[3\] vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__a21o_1
X_2428_ net362 LEI0.config_data\[18\] net268 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__mux2_1
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2359_ _1091_ _1092_ _1304_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__o21a_1
XFILLER_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1730_ _0353_ _0514_ _0516_ _0499_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__a31o_1
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1592_ net175 net171 net173 net177 vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__or4b_1
X_1661_ _0434_ _0439_ _0445_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__a22o_2
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2144_ net1 net6 net7 net8 CB_1.config_dataB\[0\] CB_1.config_dataB\[1\] vssd1 vssd1
+ vccd1 vccd1 _0927_ sky130_fd_sc_hd__mux4_1
X_2213_ _0985_ _0987_ _0994_ _0995_ _1213_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__o41a_1
X_2075_ net1 net6 net7 net8 net141 CB_1.config_dataA\[9\] vssd1 vssd1 vccd1 vccd1
+ _0860_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_36_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1928_ net134 net130 net126 net122 LEI0.config_data\[39\] LEI0.config_data\[40\]
+ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__mux4_1
X_1859_ net161 net162 vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__nand2_1
X_2977_ clknet_leaf_27_clk _0239_ net217 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[103\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold80 LEI0.config_data\[46\] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 LEI0.config_data\[19\] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
X_2900_ clknet_leaf_30_clk _0162_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_1713_ net16 net129 _0501_ vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__mux2_1
X_2762_ clknet_leaf_16_clk net347 net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2831_ LE_1A.sel_clk _0093_ net61 vssd1 vssd1 vccd1 vccd1 LE_1A.dff0_out sky130_fd_sc_hd__dfrtp_1
X_2693_ net153 CB_0.config_dataB\[14\] net263 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__mux2_1
X_1644_ _0393_ _0413_ _0374_ _0431_ _1135_ CB_0.config_dataA\[1\] vssd1 vssd1 vccd1
+ vccd1 _0433_ sky130_fd_sc_hd__mux4_1
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1575_ net8 _0362_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__and2b_1
X_2127_ _0343_ _0762_ net183 vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2058_ _0833_ _0841_ _0842_ _0816_ LEI0.config_data\[8\] vssd1 vssd1 vccd1 vccd1
+ _0843_ sky130_fd_sc_hd__o32a_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ SB0.route_sel\[54\] vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__inv_2
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 CBeast_out[3] sky130_fd_sc_hd__buf_2
X_3030_ clknet_leaf_19_clk _0292_ net220 vssd1 vssd1 vccd1 vccd1 CB_1.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 CBnorth_out[13] sky130_fd_sc_hd__buf_2
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 SBsouth_out[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2676_ CB_0.config_dataA\[18\] CB_0.config_dataA\[17\] net263 vssd1 vssd1 vccd1 vccd1
+ _0266_ sky130_fd_sc_hd__mux2_1
X_2745_ clknet_leaf_15_clk net342 net223 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2814_ clknet_leaf_1_clk _0076_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1627_ net128 net21 _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__mux2_1
X_1558_ _0343_ _0345_ net170 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__a21oi_1
X_1489_ SB0.route_sel\[43\] SB0.route_sel\[42\] vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__or2_1
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_2_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2530_ net182 CB_1.config_dataB\[3\] net264 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__mux2_1
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2461_ net320 LE_0A.config_data\[0\] net244 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__mux2_1
X_2392_ _1113_ _1114_ _0343_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__o21a_1
X_1343_ SB0.route_sel\[20\] vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__inv_2
X_1412_ LE_1A.config_data\[16\] vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__inv_2
X_3013_ clknet_leaf_6_clk _0275_ net197 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[7\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2659_ CB_0.config_dataA\[1\] net170 net246 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__mux2_1
X_2728_ net348 net303 net254 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout145 CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_2
Xfanout167 CB_0.config_dataA\[8\] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
Xfanout123 _1220_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
Xfanout134 net136 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_2
Xfanout156 CB_0.config_dataB\[12\] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_1
Xfanout189 net190 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout178 CB_1.config_dataB\[16\] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_1
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1892_ net23 net24 net25 net26 net157 CB_0.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1
+ _0679_ sky130_fd_sc_hd__mux4_1
X_1961_ CB_1.config_dataA\[5\] CB_1.config_dataA\[7\] vssd1 vssd1 vccd1 vccd1 _0746_
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2513_ net298 net288 net255 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__mux2_1
X_2444_ net375 LEI0.config_data\[34\] net269 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2375_ SB0.route_sel\[9\] SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__and2b_1
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2160_ net181 net182 vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2_1
X_2091_ net138 _0763_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2993_ clknet_leaf_7_clk _0255_ net200 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[7\]
+ sky130_fd_sc_hd__dfstp_2
X_1875_ _0431_ _0645_ _0646_ _0374_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__o22a_1
X_1944_ LE_0B.config_data\[3\] _0672_ _0730_ _0641_ vssd1 vssd1 vccd1 vccd1 _0731_
+ sky130_fd_sc_hd__a211o_1
X_2427_ LEI0.config_data\[18\] LEI0.config_data\[17\] net269 vssd1 vssd1 vccd1 vccd1
+ _0019_ sky130_fd_sc_hd__mux2_1
X_2289_ net128 _0432_ _0415_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__mux2_1
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2358_ SB0.route_sel\[33\] _1147_ _1144_ _1145_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_39_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1591_ net134 _0378_ _0379_ vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__mux2_1
X_1660_ SB0.route_sel\[67\] SB0.route_sel\[66\] _0448_ _0434_ vssd1 vssd1 vccd1 vccd1
+ _0449_ sky130_fd_sc_hd__a31oi_1
XFILLER_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2143_ _0919_ _0803_ _0514_ _1207_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__and4b_1
X_2212_ CB_1.config_dataB\[9\] CB_1.config_dataB\[8\] CB_1.config_dataB\[11\] _0801_
+ _0993_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__a41o_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_46_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2074_ CB_1.config_dataA\[9\] net141 CB_1.config_dataA\[11\] vssd1 vssd1 vccd1 vccd1
+ _0859_ sky130_fd_sc_hd__and3_1
X_1927_ _0705_ _0709_ _0712_ _0713_ CB_0.config_dataB\[14\] vssd1 vssd1 vccd1 vccd1
+ _0714_ sky130_fd_sc_hd__o311a_1
X_1858_ net162 net161 vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__nand2b_1
X_2976_ clknet_leaf_11_clk _0238_ net217 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[102\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_55_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1789_ net134 net130 net126 net122 LEI0.config_data\[24\] LEI0.config_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__mux4_2
XFILLER_39_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold70 LEI0.config_data\[5\] vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 LEI0.config_data\[1\] vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 _0047_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ clknet_leaf_31_clk _0092_ net184 vssd1 vssd1 vccd1 vccd1 LE_0B.reset_mode
+ sky130_fd_sc_hd__dfrtp_1
X_1643_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
X_1712_ net151 net147 net145 net149 vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__and4bb_1
X_2761_ clknet_leaf_16_clk _0023_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_1 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2692_ CB_0.config_dataB\[14\] net154 net260 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__mux2_1
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1574_ net121 _0362_ _0361_ _1251_ vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_49_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ CB_1.config_dataA\[3\] _0834_ _0840_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1
+ vccd1 _0842_ sky130_fd_sc_hd__o211a_1
X_2126_ _0753_ _0756_ _0750_ _0759_ _1207_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1
+ vccd1 _0909_ sky130_fd_sc_hd__mux4_1
X_2959_ clknet_leaf_2_clk _0221_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[85\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 CBnorth_out[1] sky130_fd_sc_hd__buf_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 SBsouth_out[11] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 CBeast_out[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2813_ clknet_leaf_1_clk net275 net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2675_ CB_0.config_dataA\[17\] CB_0.config_dataA\[16\] net248 vssd1 vssd1 vccd1 vccd1
+ _0265_ sky130_fd_sc_hd__mux2_1
X_2744_ clknet_leaf_15_clk _0006_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1626_ net151 net145 net147 net149 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__or4b_1
X_1557_ _0343_ _0345_ vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__and2_2
X_1488_ _1266_ _1271_ _1278_ _1281_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__a22oi_2
XFILLER_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2109_ LEI0.config_data\[44\] _0882_ _0893_ CB_1.config_dataA\[14\] vssd1 vssd1 vccd1
+ vccd1 _0894_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_9_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2460_ net328 net57 net243 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__mux2_1
X_2391_ SB0.route_sel\[96\] SB0.route_sel\[97\] SB0.route_sel\[98\] _1180_ vssd1 vssd1
+ vccd1 vccd1 _1114_ sky130_fd_sc_hd__a2bb2o_1
X_1411_ CB_1.config_dataA\[14\] vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__inv_2
X_1342_ SB0.route_sel\[19\] vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__inv_2
X_3012_ clknet_leaf_6_clk _0274_ net197 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_1609_ net15 _0396_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__nand2b_1
X_2658_ CB_0.config_dataA\[0\] CB_0.config_data_inA net265 vssd1 vssd1 vccd1 vccd1
+ _0248_ sky130_fd_sc_hd__mux2_1
X_2727_ net303 LE_1B.config_data\[8\] net254 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__mux2_1
X_2589_ SB0.route_sel\[43\] SB0.route_sel\[42\] net228 vssd1 vssd1 vccd1 vccd1 _0179_
+ sky130_fd_sc_hd__mux2_1
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout146 CB_0.config_dataB\[19\] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_1
Xfanout124 net126 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
Xfanout179 CB_1.config_dataB\[9\] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ net157 _1330_ _0676_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a211o_1
X_1960_ LE_0B.config_data\[16\] _0744_ _0745_ _0616_ vssd1 vssd1 vccd1 vccd1 CB_0.le_outB
+ sky130_fd_sc_hd__o211a_1
X_2443_ LEI0.config_data\[34\] LEI0.config_data\[33\] net269 vssd1 vssd1 vccd1 vccd1
+ _0035_ sky130_fd_sc_hd__mux2_1
X_2512_ net288 LE_1A.config_data\[6\] net255 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__mux2_1
X_2374_ _0390_ _1102_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__and2_1
XFILLER_30_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2090_ CB_1.config_dataA\[15\] _0872_ _0873_ _0874_ vssd1 vssd1 vccd1 vccd1 _0875_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_17_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ clknet_leaf_7_clk _0254_ net200 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[6\]
+ sky130_fd_sc_hd__dfstp_1
X_1874_ net162 _0393_ _0660_ net161 vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__a211o_1
X_1943_ LE_0B.config_data\[2\] _0657_ _0659_ _0671_ vssd1 vssd1 vccd1 vccd1 _0730_
+ sky130_fd_sc_hd__and4_1
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2426_ LEI0.config_data\[17\] LEI0.config_data\[16\] net269 vssd1 vssd1 vccd1 vccd1
+ _0018_ sky130_fd_sc_hd__mux2_1
X_2288_ net133 _1050_ _0359_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2357_ SB0.route_sel\[34\] SB0.route_sel\[35\] vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__and2b_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1590_ CB_0.config_dataA\[19\] CB_0.config_dataA\[18\] _1269_ vssd1 vssd1 vccd1 vccd1
+ _0379_ sky130_fd_sc_hd__or3b_1
X_2073_ net140 _0793_ _0846_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__a211o_1
X_2142_ _0469_ _0791_ _1207_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__a21o_1
X_2211_ _0981_ _0803_ _0514_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__and3b_1
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2975_ clknet_leaf_12_clk _0237_ net217 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[101\]
+ sky130_fd_sc_hd__dfstp_1
X_1788_ CB_0.config_dataA\[11\] _0572_ _0573_ _0576_ _1193_ vssd1 vssd1 vccd1 vccd1
+ _0577_ sky130_fd_sc_hd__o311a_1
X_1926_ net156 CB_0.config_dataB\[15\] net154 vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__nand3b_1
X_1857_ net162 _1285_ _0643_ net161 vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__a211o_1
X_2409_ LEI0.config_data\[0\] LE_1A.reset_mode net258 vssd1 vssd1 vccd1 vccd1 _0001_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold71 _0007_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 LEI0.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 LEI0.config_data\[42\] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 LE_0B.config_data\[0\] vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
X_2760_ clknet_leaf_16_clk _0022_ net224 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 CBeast_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2691_ net154 net155 net246 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__mux2_1
X_1642_ _0429_ _0430_ _0428_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__a21bo_4
X_1711_ SB0.route_sel\[81\] SB0.route_sel\[80\] vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__nand2_1
X_1573_ net171 net173 net175 net177 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_49_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2056_ _0822_ _1203_ CB_1.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__and3b_1
X_2125_ LE_1A.config_data\[16\] _0907_ _0908_ _0616_ vssd1 vssd1 vccd1 vccd1 CB_1.le_outA
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_16_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1909_ CB_0.config_dataB\[11\] _0693_ _0695_ _0683_ vssd1 vssd1 vccd1 vccd1 _0696_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_32_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2958_ clknet_leaf_1_clk _0220_ net190 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[84\]
+ sky130_fd_sc_hd__dfstp_1
X_2889_ clknet_leaf_29_clk _0151_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[15\]
+ sky130_fd_sc_hd__dfstp_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 CBnorth_out[2] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 SBsouth_out[12] sky130_fd_sc_hd__buf_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 CBeast_out[5] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2743_ clknet_leaf_14_clk net332 net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2812_ clknet_leaf_1_clk net350 net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2674_ CB_0.config_dataA\[16\] CB_0.config_dataA\[15\] net248 vssd1 vssd1 vccd1 vccd1
+ _0264_ sky130_fd_sc_hd__mux2_1
X_1556_ SB0.route_sel\[100\] _1181_ SB0.route_sel\[103\] _1183_ _0344_ vssd1 vssd1
+ vccd1 vccd1 _0345_ sky130_fd_sc_hd__a221o_1
X_1625_ SB0.route_sel\[17\] SB0.route_sel\[16\] vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__nand2_1
X_1487_ _1277_ _1279_ _1280_ SB0.route_sel\[40\] SB0.route_sel\[41\] vssd1 vssd1 vccd1
+ vccd1 _1281_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_52_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2039_ net1 net6 net7 net8 net144 CB_1.config_dataA\[1\] vssd1 vssd1 vccd1 vccd1
+ _0824_ sky130_fd_sc_hd__mux4_1
X_2108_ CB_1.config_dataA\[15\] _0883_ _0885_ _0892_ vssd1 vssd1 vccd1 vccd1 _0893_
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1410_ CB_1.config_dataA\[10\] vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__inv_2
X_3011_ clknet_leaf_6_clk _0273_ net197 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[5\]
+ sky130_fd_sc_hd__dfstp_2
X_2390_ SB0.route_sel\[100\] _1181_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__nor2_1
X_1341_ net170 vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__inv_2
X_2726_ net318 net282 net254 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__mux2_1
Xfanout147 CB_0.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__clkbuf_2
X_1608_ net129 _0396_ _0395_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__o21a_1
Xfanout136 CB_0.le_outA vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_2
X_1539_ _1332_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
X_2657_ net119 SB0.route_sel\[110\] net251 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__mux2_1
X_2588_ SB0.route_sel\[42\] SB0.route_sel\[41\] net228 vssd1 vssd1 vccd1 vccd1 _0178_
+ sky130_fd_sc_hd__mux2_1
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout169 CB_0.config_dataA\[4\] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 CB_0.config_dataB\[8\] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_19_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ CB_0.config_dataB\[9\] CB_0.config_dataB\[11\] vssd1 vssd1 vccd1 vccd1 _0677_
+ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2442_ LEI0.config_data\[33\] LEI0.config_data\[32\] net268 vssd1 vssd1 vccd1 vccd1
+ _0034_ sky130_fd_sc_hd__mux2_1
X_2373_ _1131_ SB0.route_sel\[10\] _1132_ SB0.route_sel\[13\] _1101_ vssd1 vssd1 vccd1
+ vccd1 _1102_ sky130_fd_sc_hd__a221o_1
X_2511_ net380 LE_1A.config_data\[5\] net255 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2709_ CB_1.config_dataA\[11\] CB_1.config_dataA\[10\] net270 vssd1 vssd1 vccd1 vccd1
+ _0299_ sky130_fd_sc_hd__mux2_1
XFILLER_3_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2991_ clknet_leaf_7_clk _0253_ net201 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[5\]
+ sky130_fd_sc_hd__dfstp_2
X_1942_ _1200_ _0715_ _0728_ _1201_ _0714_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__a221o_1
XFILLER_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1873_ _0410_ _0412_ net163 vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__a21oi_1
X_2425_ LEI0.config_data\[16\] LEI0.config_data\[15\] net269 vssd1 vssd1 vccd1 vccd1
+ _0017_ sky130_fd_sc_hd__mux2_1
XFILLER_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2356_ _1089_ _1090_ _1304_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__o21a_1
X_2287_ _0375_ net128 _0357_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2210_ net179 _1214_ _0991_ _0992_ _0990_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__o311a_1
XFILLER_46_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2072_ net140 _0796_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nor2_1
X_2141_ _0450_ _0795_ net183 vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__a21o_1
X_1925_ net153 _0710_ _0711_ _0707_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__o22a_1
X_2974_ clknet_leaf_11_clk _0236_ net217 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[100\]
+ sky130_fd_sc_hd__dfstp_1
X_1787_ _1194_ _0574_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__or3_1
X_1856_ _1304_ _1306_ net162 vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2339_ SB0.route_sel\[57\] SB0.route_sel\[56\] vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__and2b_1
X_2408_ LE_0A.dff1_out _0615_ net60 vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold50 _0052_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 LEI0.config_data\[28\] vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 LE_0A.config_data\[4\] vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 _0005_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 LEI0.config_data\[40\] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_31_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_3 CBeast_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2690_ net155 CB_0.config_dataB\[11\] net249 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__mux2_1
X_1710_ _0495_ _0496_ _0498_ CB_0.config_dataA\[2\] vssd1 vssd1 vccd1 vccd1 _0499_
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1641_ SB0.route_sel\[19\] SB0.route_sel\[18\] _1137_ SB0.route_sel\[21\] vssd1 vssd1
+ vccd1 vccd1 _0430_ sky130_fd_sc_hd__o22a_1
X_1572_ CB_1.config_dataA\[19\] CB_1.config_dataA\[18\] vssd1 vssd1 vccd1 vccd1 _0361_
+ sky130_fd_sc_hd__nor2_2
X_2124_ _1206_ LE_1A.dff_out vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _0820_ _0835_ _0836_ _0839_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__o31a_1
X_1839_ net132 net127 net123 net120 LEI0.config_data\[15\] LEI0.config_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__mux4_1
X_1908_ net16 net17 net158 vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2888_ clknet_leaf_30_clk _0150_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_2957_ clknet_leaf_2_clk _0219_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[83\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_55_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 CBnorth_out[3] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 SBsouth_out[13] sky130_fd_sc_hd__buf_2
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 CBeast_out[6] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_2_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2742_ clknet_leaf_14_clk _0004_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2811_ clknet_leaf_0_clk _0073_ net188 vssd1 vssd1 vccd1 vccd1 LE_0B.config_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2673_ CB_0.config_dataA\[15\] CB_0.config_dataA\[14\] net248 vssd1 vssd1 vccd1 vccd1
+ _0263_ sky130_fd_sc_hd__mux2_1
X_1555_ SB0.route_sel\[98\] SB0.route_sel\[99\] vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__nor2_1
X_1624_ _0410_ _0412_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2107_ _0804_ _0880_ _0886_ _0801_ _0891_ vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__a221oi_1
X_1486_ SB0.route_sel\[44\] SB0.route_sel\[45\] net38 vssd1 vssd1 vccd1 vccd1 _1280_
+ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_52_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _0822_ _0803_ _0514_ _1203_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__and4b_1
XFILLER_7_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1340_ net34 vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__inv_2
X_3010_ clknet_leaf_5_clk _0272_ net198 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataB\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
X_2725_ net282 LE_1B.config_data\[6\] net257 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__mux2_1
X_2656_ SB0.route_sel\[110\] SB0.route_sel\[109\] net251 vssd1 vssd1 vccd1 vccd1 _0246_
+ sky130_fd_sc_hd__mux2_1
X_1607_ net149 net151 net145 net147 vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__or4_1
Xfanout148 CB_0.config_dataB\[18\] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_1
X_1538_ CB_0.config_dataA\[1\] CB_0.config_dataA\[3\] vssd1 vssd1 vccd1 vccd1 _1332_
+ sky130_fd_sc_hd__nand2b_1
Xfanout159 net160 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
Xfanout126 CB_1.le_outA vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
X_2587_ SB0.route_sel\[41\] SB0.route_sel\[40\] net228 vssd1 vssd1 vccd1 vccd1 _0177_
+ sky130_fd_sc_hd__mux2_1
X_1469_ SB0.route_sel\[60\] _1157_ SB0.route_sel\[63\] _1158_ _1262_ vssd1 vssd1 vccd1
+ vccd1 _1263_ sky130_fd_sc_hd__a221o_1
Xfanout137 _1230_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_57_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2510_ LE_1A.config_data\[5\] LE_1A.config_data\[4\] net255 vssd1 vssd1 vccd1 vccd1
+ _0100_ sky130_fd_sc_hd__mux2_1
X_2441_ LEI0.config_data\[32\] net373 net268 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__mux2_1
X_2372_ SB0.route_sel\[9\] SB0.route_sel\[8\] vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_20_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2708_ CB_1.config_dataA\[10\] CB_1.config_dataA\[9\] net265 vssd1 vssd1 vccd1 vccd1
+ _0298_ sky130_fd_sc_hd__mux2_1
X_2639_ SB0.route_sel\[93\] SB0.route_sel\[92\] net247 vssd1 vssd1 vccd1 vccd1 _0229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1872_ LEI0.config_data\[5\] _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__or2_4
X_1941_ _0717_ _0719_ _0720_ _0727_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__or4_1
X_2990_ clknet_leaf_10_clk _0252_ net202 vssd1 vssd1 vccd1 vccd1 CB_0.config_dataA\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2424_ LEI0.config_data\[15\] LEI0.config_data\[14\] net268 vssd1 vssd1 vccd1 vccd1
+ _0016_ sky130_fd_sc_hd__mux2_1
X_2286_ _1300_ _1049_ _1302_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__a21o_1
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2355_ SB0.route_sel\[36\] _1143_ SB0.route_sel\[33\] SB0.route_sel\[32\] vssd1 vssd1
+ vccd1 vccd1 _1090_ sky130_fd_sc_hd__o22ai_1
XFILLER_28_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2140_ _0781_ _0784_ _0778_ _0787_ _1207_ CB_1.config_dataB\[1\] vssd1 vssd1 vccd1
+ vccd1 _0923_ sky130_fd_sc_hd__mux4_1
X_2071_ _0784_ _0787_ _0781_ _0778_ CB_1.config_dataA\[9\] net140 vssd1 vssd1 vccd1
+ vccd1 _0856_ sky130_fd_sc_hd__mux4_1
X_1924_ net18 net19 net156 vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__mux2_1
X_2973_ clknet_leaf_10_clk _0235_ net217 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[99\]
+ sky130_fd_sc_hd__dfstp_1
X_1855_ _0636_ _0637_ _0640_ _0627_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o31ai_4
X_1786_ net27 net28 net16 net17 CB_0.config_dataA\[8\] net166 vssd1 vssd1 vccd1 vccd1
+ _0575_ sky130_fd_sc_hd__mux4_1
X_2269_ _0346_ net130 _0330_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__mux2_1
X_2407_ _1123_ _1124_ _0514_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__o21a_1
X_2338_ _1077_ _1078_ _1261_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 _0313_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold73 LEI0.config_data\[37\] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _0029_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0041_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 LE_0B.config_data\[11\] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 LE_0B.config_data\[15\] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ net133 _0358_ _0359_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_4 LEI0.config_data\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1640_ SB0.route_sel\[23\] _1138_ vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__nand2_1
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ LE_1A.dff0_out LE_1A.dff1_out LE_1A.reset_val vssd1 vssd1 vccd1 vccd1 LE_1A.dff_out
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2054_ CB_1.config_dataA\[3\] _0837_ _0838_ _0820_ vssd1 vssd1 vccd1 vccd1 _0839_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1907_ net27 net28 net158 vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__mux2_1
X_1838_ CB_0.config_dataB\[5\] CB_0.config_dataB\[7\] vssd1 vssd1 vccd1 vccd1 _0625_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2887_ clknet_leaf_29_clk _0149_ net191 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_2956_ clknet_leaf_2_clk _0218_ net189 vssd1 vssd1 vccd1 vccd1 SB0.route_sel\[82\]
+ sky130_fd_sc_hd__dfstp_1
X_1769_ net23 net24 net25 net26 CB_0.config_dataA\[8\] net166 vssd1 vssd1 vccd1 vccd1
+ _0558_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_55_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 CBnorth_out[4] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 SBsouth_out[1] sky130_fd_sc_hd__buf_2
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 CBeast_out[0] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 CBeast_out[7] sky130_fd_sc_hd__buf_2
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2672_ CB_0.config_dataA\[14\] net164 net248 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__mux2_1
X_2741_ clknet_leaf_17_clk _0003_ net222 vssd1 vssd1 vccd1 vccd1 LEI0.config_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2810_ LE_1A.sel_clk _0072_ net61 vssd1 vssd1 vccd1 vccd1 LE_1A.dff1_out sky130_fd_sc_hd__dfstp_1
X_1554_ _0329_ _0333_ _0339_ _0342_ vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__a22o_2
X_1623_ SB0.route_sel\[4\] _1128_ SB0.route_sel\[7\] _1129_ _0411_ vssd1 vssd1 vccd1
+ vccd1 _0412_ sky130_fd_sc_hd__a221o_1
X_1485_ _1150_ _1151_ net52 SB0.route_sel\[45\] SB0.route_sel\[44\] vssd1 vssd1 vccd1
+ vccd1 _1279_ sky130_fd_sc_hd__o2111a_1
.ends

