magic
tech sky130A
magscale 1 2
timestamp 1748220643
<< viali >>
rect 17693 43401 17727 43435
rect 19533 43401 19567 43435
rect 20269 43401 20303 43435
rect 20821 43401 20855 43435
rect 22845 43401 22879 43435
rect 23397 43401 23431 43435
rect 25329 43401 25363 43435
rect 29193 43401 29227 43435
rect 24685 43333 24719 43367
rect 28181 43333 28215 43367
rect 17509 43265 17543 43299
rect 19717 43265 19751 43299
rect 20085 43265 20119 43299
rect 21005 43265 21039 43299
rect 22661 43265 22695 43299
rect 23581 43265 23615 43299
rect 24593 43265 24627 43299
rect 24777 43265 24811 43299
rect 24961 43265 24995 43299
rect 25513 43265 25547 43299
rect 28365 43265 28399 43299
rect 29377 43265 29411 43299
rect 24409 43061 24443 43095
rect 28549 43061 28583 43095
rect 17417 42857 17451 42891
rect 26157 42857 26191 42891
rect 28457 42857 28491 42891
rect 24409 42721 24443 42755
rect 26341 42721 26375 42755
rect 35173 42721 35207 42755
rect 15669 42653 15703 42687
rect 18337 42653 18371 42687
rect 19441 42653 19475 42687
rect 19809 42653 19843 42687
rect 21005 42653 21039 42687
rect 24041 42653 24075 42687
rect 28641 42653 28675 42687
rect 29009 42653 29043 42687
rect 15945 42585 15979 42619
rect 18521 42585 18555 42619
rect 19533 42585 19567 42619
rect 19625 42585 19659 42619
rect 21281 42585 21315 42619
rect 23857 42585 23891 42619
rect 24225 42585 24259 42619
rect 24685 42585 24719 42619
rect 26617 42585 26651 42619
rect 28733 42585 28767 42619
rect 28825 42585 28859 42619
rect 35449 42585 35483 42619
rect 18705 42517 18739 42551
rect 19257 42517 19291 42551
rect 22753 42517 22787 42551
rect 28089 42517 28123 42551
rect 36921 42517 36955 42551
rect 16865 42313 16899 42347
rect 26985 42313 27019 42347
rect 29561 42313 29595 42347
rect 35357 42313 35391 42347
rect 39037 42313 39071 42347
rect 16313 42245 16347 42279
rect 17141 42245 17175 42279
rect 18153 42245 18187 42279
rect 27629 42245 27663 42279
rect 28089 42245 28123 42279
rect 16129 42177 16163 42211
rect 16497 42177 16531 42211
rect 17049 42177 17083 42211
rect 17233 42177 17267 42211
rect 17417 42177 17451 42211
rect 17877 42177 17911 42211
rect 19901 42177 19935 42211
rect 27261 42177 27295 42211
rect 32413 42177 32447 42211
rect 35633 42177 35667 42211
rect 36277 42177 36311 42211
rect 36737 42177 36771 42211
rect 37289 42177 37323 42211
rect 19625 42109 19659 42143
rect 20177 42109 20211 42143
rect 22385 42109 22419 42143
rect 22661 42109 22695 42143
rect 22937 42109 22971 42143
rect 27169 42109 27203 42143
rect 27537 42109 27571 42143
rect 27813 42109 27847 42143
rect 30205 42109 30239 42143
rect 30481 42109 30515 42143
rect 35541 42109 35575 42143
rect 35909 42109 35943 42143
rect 36001 42109 36035 42143
rect 36553 42109 36587 42143
rect 36645 42109 36679 42143
rect 37565 42109 37599 42143
rect 32229 42041 32263 42075
rect 37105 42041 37139 42075
rect 21649 41973 21683 42007
rect 21833 41973 21867 42007
rect 24409 41973 24443 42007
rect 31953 41973 31987 42007
rect 36093 41973 36127 42007
rect 20453 41769 20487 41803
rect 21741 41769 21775 41803
rect 23305 41769 23339 41803
rect 27353 41769 27387 41803
rect 28457 41769 28491 41803
rect 28917 41769 28951 41803
rect 30849 41769 30883 41803
rect 33149 41769 33183 41803
rect 34805 41769 34839 41803
rect 35357 41769 35391 41803
rect 36461 41769 36495 41803
rect 30757 41701 30791 41735
rect 35265 41701 35299 41735
rect 14841 41633 14875 41667
rect 17141 41633 17175 41667
rect 20085 41633 20119 41667
rect 21097 41633 21131 41667
rect 23949 41633 23983 41667
rect 26157 41633 26191 41667
rect 26893 41633 26927 41667
rect 27629 41633 27663 41667
rect 29101 41633 29135 41667
rect 36277 41633 36311 41667
rect 36645 41633 36679 41667
rect 19993 41565 20027 41599
rect 20821 41565 20855 41599
rect 22017 41565 22051 41599
rect 22109 41565 22143 41599
rect 22385 41565 22419 41599
rect 23673 41565 23707 41599
rect 25881 41565 25915 41599
rect 25973 41565 26007 41599
rect 26065 41565 26099 41599
rect 26985 41565 27019 41599
rect 27077 41565 27111 41599
rect 27169 41565 27203 41599
rect 28365 41565 28399 41599
rect 28733 41565 28767 41599
rect 28825 41565 28859 41599
rect 30481 41565 30515 41599
rect 30573 41565 30607 41599
rect 31033 41565 31067 41599
rect 31125 41565 31159 41599
rect 31493 41565 31527 41599
rect 31769 41565 31803 41599
rect 31861 41565 31895 41599
rect 31953 41565 31987 41599
rect 32045 41565 32079 41599
rect 32689 41565 32723 41599
rect 32781 41565 32815 41599
rect 32873 41565 32907 41599
rect 32965 41565 32999 41599
rect 33149 41565 33183 41599
rect 33241 41565 33275 41599
rect 34713 41565 34747 41599
rect 34989 41565 35023 41599
rect 35541 41565 35575 41599
rect 35633 41565 35667 41599
rect 35725 41565 35759 41599
rect 35817 41565 35851 41599
rect 36185 41565 36219 41599
rect 36829 41565 36863 41599
rect 36921 41565 36955 41599
rect 15117 41497 15151 41531
rect 17417 41497 17451 41531
rect 20913 41497 20947 41531
rect 21373 41497 21407 41531
rect 21557 41497 21591 41531
rect 22201 41497 22235 41531
rect 28457 41497 28491 41531
rect 30757 41497 30791 41531
rect 31401 41497 31435 41531
rect 35265 41497 35299 41531
rect 36645 41497 36679 41531
rect 16589 41429 16623 41463
rect 18889 41429 18923 41463
rect 20361 41429 20395 41463
rect 21833 41429 21867 41463
rect 23765 41429 23799 41463
rect 25697 41429 25731 41463
rect 28641 41429 28675 41463
rect 29101 41429 29135 41463
rect 31585 41429 31619 41463
rect 32505 41429 32539 41463
rect 33517 41429 33551 41463
rect 35081 41429 35115 41463
rect 15577 41225 15611 41259
rect 19993 41225 20027 41259
rect 23489 41225 23523 41259
rect 27353 41225 27387 41259
rect 28825 41225 28859 41259
rect 16037 41157 16071 41191
rect 17417 41157 17451 41191
rect 17617 41157 17651 41191
rect 19330 41157 19364 41191
rect 26985 41157 27019 41191
rect 29193 41157 29227 41191
rect 31769 41157 31803 41191
rect 31953 41157 31987 41191
rect 15945 41089 15979 41123
rect 16681 41089 16715 41123
rect 17969 41089 18003 41123
rect 19157 41089 19191 41123
rect 19441 41089 19475 41123
rect 19534 41089 19568 41123
rect 19901 41089 19935 41123
rect 20085 41089 20119 41123
rect 22661 41089 22695 41123
rect 22845 41089 22879 41123
rect 23121 41089 23155 41123
rect 23581 41089 23615 41123
rect 23765 41089 23799 41123
rect 24777 41089 24811 41123
rect 27169 41089 27203 41123
rect 27905 41089 27939 41123
rect 28457 41089 28491 41123
rect 31585 41089 31619 41123
rect 32137 41089 32171 41123
rect 32229 41089 32263 41123
rect 32413 41089 32447 41123
rect 36093 41089 36127 41123
rect 38209 41089 38243 41123
rect 16221 41021 16255 41055
rect 17233 41021 17267 41055
rect 18705 41021 18739 41055
rect 22753 41021 22787 41055
rect 23213 41021 23247 41055
rect 25053 41021 25087 41055
rect 28273 41021 28307 41055
rect 28365 41021 28399 41055
rect 28917 41021 28951 41055
rect 32505 41021 32539 41055
rect 32781 41021 32815 41055
rect 36001 41021 36035 41055
rect 19809 40953 19843 40987
rect 17601 40885 17635 40919
rect 17785 40885 17819 40919
rect 18981 40885 19015 40919
rect 23949 40885 23983 40919
rect 26525 40885 26559 40919
rect 30665 40885 30699 40919
rect 32413 40885 32447 40919
rect 34253 40885 34287 40919
rect 35725 40885 35759 40919
rect 36093 40885 36127 40919
rect 17325 40681 17359 40715
rect 20545 40681 20579 40715
rect 20913 40681 20947 40715
rect 21005 40681 21039 40715
rect 25329 40681 25363 40715
rect 27445 40681 27479 40715
rect 28457 40681 28491 40715
rect 32505 40681 32539 40715
rect 35541 40681 35575 40715
rect 17233 40613 17267 40647
rect 17693 40613 17727 40647
rect 20453 40613 20487 40647
rect 26065 40613 26099 40647
rect 27905 40613 27939 40647
rect 31125 40613 31159 40647
rect 34989 40613 35023 40647
rect 35817 40613 35851 40647
rect 37473 40613 37507 40647
rect 17601 40545 17635 40579
rect 20637 40545 20671 40579
rect 21189 40545 21223 40579
rect 21741 40545 21775 40579
rect 22017 40545 22051 40579
rect 22109 40545 22143 40579
rect 25513 40545 25547 40579
rect 25973 40545 26007 40579
rect 27629 40545 27663 40579
rect 28273 40545 28307 40579
rect 30665 40545 30699 40579
rect 32689 40545 32723 40579
rect 33057 40545 33091 40579
rect 37933 40545 37967 40579
rect 38853 40545 38887 40579
rect 16957 40477 16991 40511
rect 17049 40477 17083 40511
rect 17509 40477 17543 40511
rect 17785 40477 17819 40511
rect 18153 40477 18187 40511
rect 20269 40477 20303 40511
rect 20545 40477 20579 40511
rect 21281 40477 21315 40511
rect 21925 40477 21959 40511
rect 22201 40477 22235 40511
rect 25605 40477 25639 40511
rect 26341 40477 26375 40511
rect 27721 40477 27755 40511
rect 28181 40477 28215 40511
rect 30757 40477 30791 40511
rect 32781 40477 32815 40511
rect 35173 40477 35207 40511
rect 35265 40477 35299 40511
rect 35357 40477 35391 40511
rect 36001 40477 36035 40511
rect 37841 40477 37875 40511
rect 42165 40477 42199 40511
rect 17233 40409 17267 40443
rect 20085 40409 20119 40443
rect 21557 40409 21591 40443
rect 21649 40409 21683 40443
rect 25881 40409 25915 40443
rect 26065 40409 26099 40443
rect 27445 40409 27479 40443
rect 33149 40409 33183 40443
rect 34989 40409 35023 40443
rect 38117 40409 38151 40443
rect 26249 40341 26283 40375
rect 41521 40341 41555 40375
rect 17509 40137 17543 40171
rect 19441 40137 19475 40171
rect 20998 40137 21032 40171
rect 23489 40137 23523 40171
rect 25421 40137 25455 40171
rect 30757 40137 30791 40171
rect 32689 40137 32723 40171
rect 37013 40137 37047 40171
rect 21097 40069 21131 40103
rect 16037 40001 16071 40035
rect 17141 40001 17175 40035
rect 19073 40001 19107 40035
rect 20824 40023 20858 40057
rect 20913 40001 20947 40035
rect 23121 40001 23155 40035
rect 25053 40001 25087 40035
rect 27169 40001 27203 40035
rect 30665 40001 30699 40035
rect 30849 40001 30883 40035
rect 32321 40001 32355 40035
rect 35909 40001 35943 40035
rect 36001 40001 36035 40035
rect 36921 40001 36955 40035
rect 37105 40001 37139 40035
rect 38393 40001 38427 40035
rect 38669 40001 38703 40035
rect 38865 40001 38899 40035
rect 39129 40001 39163 40035
rect 39588 40001 39622 40035
rect 39681 40001 39715 40035
rect 40049 40001 40083 40035
rect 13277 39933 13311 39967
rect 13553 39933 13587 39967
rect 15669 39933 15703 39967
rect 15945 39933 15979 39967
rect 16405 39933 16439 39967
rect 17233 39933 17267 39967
rect 18981 39933 19015 39967
rect 23213 39933 23247 39967
rect 25145 39933 25179 39967
rect 27077 39933 27111 39967
rect 32229 39933 32263 39967
rect 33793 39933 33827 39967
rect 34069 39933 34103 39967
rect 35817 39933 35851 39967
rect 36093 39933 36127 39967
rect 37289 39933 37323 39967
rect 38485 39933 38519 39967
rect 39313 39933 39347 39967
rect 40325 39933 40359 39967
rect 27537 39865 27571 39899
rect 38025 39865 38059 39899
rect 38945 39865 38979 39899
rect 39037 39865 39071 39899
rect 15025 39797 15059 39831
rect 15117 39797 15151 39831
rect 35541 39797 35575 39831
rect 35633 39797 35667 39831
rect 37933 39797 37967 39831
rect 41797 39797 41831 39831
rect 13185 39593 13219 39627
rect 23121 39593 23155 39627
rect 24225 39593 24259 39627
rect 25145 39593 25179 39627
rect 26525 39593 26559 39627
rect 26801 39593 26835 39627
rect 28181 39593 28215 39627
rect 30573 39593 30607 39627
rect 32137 39593 32171 39627
rect 32229 39593 32263 39627
rect 34713 39593 34747 39627
rect 39589 39593 39623 39627
rect 42165 39593 42199 39627
rect 17325 39525 17359 39559
rect 18245 39525 18279 39559
rect 18613 39525 18647 39559
rect 18705 39525 18739 39559
rect 20545 39525 20579 39559
rect 23213 39525 23247 39559
rect 23857 39525 23891 39559
rect 24777 39525 24811 39559
rect 25237 39525 25271 39559
rect 27261 39525 27295 39559
rect 28549 39525 28583 39559
rect 31125 39525 31159 39559
rect 31861 39525 31895 39559
rect 32321 39525 32355 39559
rect 38577 39525 38611 39559
rect 13737 39457 13771 39491
rect 14841 39457 14875 39491
rect 15485 39457 15519 39491
rect 17601 39457 17635 39491
rect 19625 39457 19659 39491
rect 20269 39457 20303 39491
rect 20821 39457 20855 39491
rect 21097 39457 21131 39491
rect 22569 39457 22603 39491
rect 23949 39457 23983 39491
rect 27353 39457 27387 39491
rect 27997 39457 28031 39491
rect 28365 39457 28399 39491
rect 30849 39457 30883 39491
rect 31217 39457 31251 39491
rect 32689 39457 32723 39491
rect 35265 39457 35299 39491
rect 35725 39457 35759 39491
rect 38025 39457 38059 39491
rect 38669 39457 38703 39491
rect 40417 39457 40451 39491
rect 13553 39389 13587 39423
rect 17693 39389 17727 39423
rect 17969 39389 18003 39423
rect 18245 39389 18279 39423
rect 18429 39389 18463 39423
rect 18613 39389 18647 39423
rect 18980 39389 19014 39423
rect 19073 39389 19107 39423
rect 19441 39389 19475 39423
rect 19533 39389 19567 39423
rect 19717 39389 19751 39423
rect 19901 39389 19935 39423
rect 20177 39389 20211 39423
rect 22937 39389 22971 39423
rect 23121 39389 23155 39423
rect 23488 39389 23522 39423
rect 23581 39389 23615 39423
rect 23765 39389 23799 39423
rect 24041 39389 24075 39423
rect 24409 39389 24443 39423
rect 24593 39389 24627 39423
rect 24685 39389 24719 39423
rect 24869 39389 24903 39423
rect 25053 39389 25087 39423
rect 26341 39389 26375 39423
rect 26525 39389 26559 39423
rect 26892 39389 26926 39423
rect 26985 39389 27019 39423
rect 27169 39389 27203 39423
rect 27445 39389 27479 39423
rect 27629 39389 27663 39423
rect 27905 39389 27939 39423
rect 30664 39389 30698 39423
rect 30757 39389 30791 39423
rect 31033 39389 31067 39423
rect 31309 39389 31343 39423
rect 31493 39389 31527 39423
rect 31677 39389 31711 39423
rect 31769 39389 31803 39423
rect 31953 39389 31987 39423
rect 34897 39389 34931 39423
rect 34989 39389 35023 39423
rect 35817 39389 35851 39423
rect 38485 39389 38519 39423
rect 38761 39389 38795 39423
rect 38945 39389 38979 39423
rect 39405 39389 39439 39423
rect 39497 39389 39531 39423
rect 39957 39389 39991 39423
rect 40325 39389 40359 39423
rect 14933 39321 14967 39355
rect 15761 39321 15795 39355
rect 18061 39321 18095 39355
rect 25605 39321 25639 39355
rect 28825 39321 28859 39355
rect 35357 39321 35391 39355
rect 37749 39321 37783 39355
rect 39681 39321 39715 39355
rect 40141 39321 40175 39355
rect 40693 39321 40727 39355
rect 13645 39253 13679 39287
rect 15025 39253 15059 39287
rect 15393 39253 15427 39287
rect 17233 39253 17267 39287
rect 19257 39253 19291 39287
rect 36185 39253 36219 39287
rect 36277 39253 36311 39287
rect 38301 39253 38335 39287
rect 16681 39049 16715 39083
rect 17601 39049 17635 39083
rect 19625 39049 19659 39083
rect 20821 39049 20855 39083
rect 24225 39049 24259 39083
rect 25237 39049 25271 39083
rect 31677 39049 31711 39083
rect 32505 39049 32539 39083
rect 32781 39049 32815 39083
rect 35817 39049 35851 39083
rect 35909 39049 35943 39083
rect 37289 39049 37323 39083
rect 37657 39049 37691 39083
rect 38669 39049 38703 39083
rect 39957 39049 39991 39083
rect 40141 39049 40175 39083
rect 40693 39049 40727 39083
rect 41061 39049 41095 39083
rect 24133 38981 24167 39015
rect 30665 38981 30699 39015
rect 30849 38981 30883 39015
rect 37749 38981 37783 39015
rect 3617 38913 3651 38947
rect 15669 38913 15703 38947
rect 17049 38913 17083 38947
rect 17509 38913 17543 38947
rect 17693 38913 17727 38947
rect 19165 38913 19199 38947
rect 19257 38913 19291 38947
rect 19349 38913 19383 38947
rect 19441 38913 19475 38947
rect 21035 38913 21069 38947
rect 21189 38913 21223 38947
rect 23581 38913 23615 38947
rect 23765 38913 23799 38947
rect 23857 38913 23891 38947
rect 23949 38913 23983 38947
rect 24225 38913 24259 38947
rect 25145 38913 25179 38947
rect 25237 38913 25271 38947
rect 25421 38913 25455 38947
rect 27353 38913 27387 38947
rect 27629 38913 27663 38947
rect 27813 38913 27847 38947
rect 30297 38913 30331 38947
rect 30481 38913 30515 38947
rect 30757 38913 30791 38947
rect 31033 38913 31067 38947
rect 31401 38913 31435 38947
rect 31585 38913 31619 38947
rect 31677 38913 31711 38947
rect 32137 38913 32171 38947
rect 32505 38913 32539 38947
rect 32781 38903 32815 38937
rect 32873 38913 32907 38947
rect 33057 38913 33091 38947
rect 35357 38913 35391 38947
rect 35633 38913 35667 38947
rect 36185 38913 36219 38947
rect 39773 38913 39807 38947
rect 40049 38913 40083 38947
rect 40141 38913 40175 38947
rect 40325 38913 40359 38947
rect 42073 38913 42107 38947
rect 13185 38845 13219 38879
rect 13461 38845 13495 38879
rect 14933 38845 14967 38879
rect 17141 38845 17175 38879
rect 17325 38845 17359 38879
rect 27445 38845 27479 38879
rect 32689 38845 32723 38879
rect 35449 38845 35483 38879
rect 35909 38845 35943 38879
rect 37841 38845 37875 38879
rect 39129 38845 39163 38879
rect 41153 38845 41187 38879
rect 41245 38845 41279 38879
rect 23581 38777 23615 38811
rect 27537 38777 27571 38811
rect 31033 38777 31067 38811
rect 35541 38777 35575 38811
rect 38853 38777 38887 38811
rect 39773 38777 39807 38811
rect 3525 38709 3559 38743
rect 15025 38709 15059 38743
rect 27169 38709 27203 38743
rect 36093 38709 36127 38743
rect 41521 38709 41555 38743
rect 14105 38505 14139 38539
rect 19533 38505 19567 38539
rect 19717 38505 19751 38539
rect 21189 38505 21223 38539
rect 21557 38505 21591 38539
rect 22017 38505 22051 38539
rect 23581 38505 23615 38539
rect 24133 38505 24167 38539
rect 25237 38505 25271 38539
rect 26157 38505 26191 38539
rect 28549 38505 28583 38539
rect 29193 38505 29227 38539
rect 31309 38505 31343 38539
rect 40509 38505 40543 38539
rect 13553 38437 13587 38471
rect 22477 38437 22511 38471
rect 25973 38437 26007 38471
rect 38577 38437 38611 38471
rect 1685 38369 1719 38403
rect 6561 38369 6595 38403
rect 8585 38369 8619 38403
rect 9505 38369 9539 38403
rect 14749 38369 14783 38403
rect 29561 38369 29595 38403
rect 32045 38369 32079 38403
rect 35725 38369 35759 38403
rect 37381 38369 37415 38403
rect 41061 38369 41095 38403
rect 4353 38301 4387 38335
rect 4721 38301 4755 38335
rect 4997 38301 5031 38335
rect 6101 38301 6135 38335
rect 6285 38301 6319 38335
rect 6837 38301 6871 38335
rect 11805 38301 11839 38335
rect 14473 38301 14507 38335
rect 19257 38301 19291 38335
rect 19349 38301 19383 38335
rect 19809 38301 19843 38335
rect 19901 38301 19935 38335
rect 21189 38301 21223 38335
rect 21281 38301 21315 38335
rect 21465 38301 21499 38335
rect 22017 38301 22051 38335
rect 22201 38301 22235 38335
rect 22293 38301 22327 38335
rect 22385 38301 22419 38335
rect 22569 38301 22603 38335
rect 23765 38301 23799 38335
rect 24041 38301 24075 38335
rect 24225 38301 24259 38335
rect 25421 38301 25455 38335
rect 25697 38301 25731 38335
rect 25789 38301 25823 38335
rect 26065 38301 26099 38335
rect 26249 38301 26283 38335
rect 28549 38301 28583 38335
rect 28825 38301 28859 38335
rect 28917 38301 28951 38335
rect 32413 38301 32447 38335
rect 35265 38301 35299 38335
rect 35817 38301 35851 38335
rect 37933 38301 37967 38335
rect 38209 38301 38243 38335
rect 38577 38301 38611 38335
rect 38761 38301 38795 38335
rect 40877 38301 40911 38335
rect 41889 38301 41923 38335
rect 1961 38233 1995 38267
rect 4537 38233 4571 38267
rect 5089 38233 5123 38267
rect 5273 38233 5307 38267
rect 5457 38233 5491 38267
rect 6193 38233 6227 38267
rect 6423 38233 6457 38267
rect 7113 38233 7147 38267
rect 12081 38233 12115 38267
rect 19533 38233 19567 38267
rect 19625 38233 19659 38267
rect 21741 38233 21775 38267
rect 21925 38233 21959 38267
rect 23949 38233 23983 38267
rect 25605 38233 25639 38267
rect 25983 38233 26017 38267
rect 28641 38233 28675 38267
rect 29193 38233 29227 38267
rect 29837 38233 29871 38267
rect 32689 38233 32723 38267
rect 41337 38233 41371 38267
rect 3433 38165 3467 38199
rect 3801 38165 3835 38199
rect 4905 38165 4939 38199
rect 5917 38165 5951 38199
rect 8953 38165 8987 38199
rect 14565 38165 14599 38199
rect 29009 38165 29043 38199
rect 31401 38165 31435 38199
rect 34161 38165 34195 38199
rect 34713 38165 34747 38199
rect 35449 38165 35483 38199
rect 40969 38165 41003 38199
rect 2329 37961 2363 37995
rect 6377 37961 6411 37995
rect 7021 37961 7055 37995
rect 15577 37961 15611 37995
rect 18981 37961 19015 37995
rect 19533 37961 19567 37995
rect 27635 37961 27669 37995
rect 27997 37961 28031 37995
rect 28641 37961 28675 37995
rect 29101 37961 29135 37995
rect 29561 37961 29595 37995
rect 29929 37961 29963 37995
rect 33425 37961 33459 37995
rect 33793 37961 33827 37995
rect 34805 37961 34839 37995
rect 36001 37961 36035 37995
rect 38025 37961 38059 37995
rect 40509 37961 40543 37995
rect 2835 37893 2869 37927
rect 7757 37893 7791 37927
rect 19165 37893 19199 37927
rect 22293 37893 22327 37927
rect 27445 37893 27479 37927
rect 27721 37893 27755 37927
rect 28089 37893 28123 37927
rect 29009 37893 29043 37927
rect 30481 37893 30515 37927
rect 32873 37893 32907 37927
rect 33241 37893 33275 37927
rect 33885 37893 33919 37927
rect 40417 37893 40451 37927
rect 1777 37825 1811 37859
rect 1869 37825 1903 37859
rect 2053 37825 2087 37859
rect 2513 37825 2547 37859
rect 2605 37825 2639 37859
rect 2697 37825 2731 37859
rect 2973 37825 3007 37859
rect 6745 37825 6779 37859
rect 7205 37825 7239 37859
rect 7297 37825 7331 37859
rect 7389 37825 7423 37859
rect 7507 37825 7541 37859
rect 7665 37825 7699 37859
rect 7941 37825 7975 37859
rect 8125 37825 8159 37859
rect 8217 37825 8251 37859
rect 12817 37825 12851 37859
rect 15117 37825 15151 37859
rect 15393 37825 15427 37859
rect 16865 37825 16899 37859
rect 18429 37825 18463 37859
rect 18889 37825 18923 37859
rect 19073 37825 19107 37859
rect 19349 37825 19383 37859
rect 21649 37825 21683 37859
rect 22201 37825 22235 37859
rect 23029 37825 23063 37859
rect 24133 37825 24167 37859
rect 27077 37825 27111 37859
rect 27261 37825 27295 37859
rect 27537 37825 27571 37859
rect 27813 37825 27847 37859
rect 27905 37825 27939 37859
rect 28181 37825 28215 37859
rect 28825 37825 28859 37859
rect 29101 37825 29135 37859
rect 29285 37825 29319 37859
rect 30389 37825 30423 37859
rect 30573 37825 30607 37859
rect 31677 37825 31711 37859
rect 32137 37825 32171 37859
rect 33149 37825 33183 37859
rect 33333 37825 33367 37859
rect 34437 37825 34471 37859
rect 36369 37825 36403 37859
rect 37381 37825 37415 37859
rect 37565 37825 37599 37859
rect 37841 37825 37875 37859
rect 38239 37825 38273 37859
rect 38393 37825 38427 37859
rect 39957 37825 39991 37859
rect 40141 37825 40175 37859
rect 40601 37825 40635 37859
rect 40693 37825 40727 37859
rect 40969 37825 41003 37859
rect 41889 37825 41923 37859
rect 1685 37757 1719 37791
rect 3709 37757 3743 37791
rect 3801 37757 3835 37791
rect 4077 37757 4111 37791
rect 6561 37757 6595 37791
rect 6653 37757 6687 37791
rect 6837 37757 6871 37791
rect 13093 37757 13127 37791
rect 13369 37757 13403 37791
rect 14841 37757 14875 37791
rect 16957 37757 16991 37791
rect 17233 37757 17267 37791
rect 20361 37757 20395 37791
rect 21005 37757 21039 37791
rect 22477 37757 22511 37791
rect 30021 37757 30055 37791
rect 30113 37757 30147 37791
rect 33977 37757 34011 37791
rect 34345 37757 34379 37791
rect 36461 37757 36495 37791
rect 15301 37689 15335 37723
rect 37657 37689 37691 37723
rect 37749 37689 37783 37723
rect 41705 37689 41739 37723
rect 2237 37621 2271 37655
rect 3065 37621 3099 37655
rect 5549 37621 5583 37655
rect 18521 37621 18555 37655
rect 19809 37621 19843 37655
rect 21833 37621 21867 37655
rect 23581 37621 23615 37655
rect 40325 37621 40359 37655
rect 3249 37417 3283 37451
rect 3433 37417 3467 37451
rect 5536 37417 5570 37451
rect 7021 37417 7055 37451
rect 8493 37417 8527 37451
rect 12081 37417 12115 37451
rect 14105 37417 14139 37451
rect 15577 37417 15611 37451
rect 20637 37417 20671 37451
rect 24225 37417 24259 37451
rect 26157 37417 26191 37451
rect 27997 37417 28031 37451
rect 34253 37417 34287 37451
rect 36461 37417 36495 37451
rect 39405 37417 39439 37451
rect 39957 37417 39991 37451
rect 3157 37349 3191 37383
rect 9045 37349 9079 37383
rect 29101 37349 29135 37383
rect 34897 37349 34931 37383
rect 36369 37349 36403 37383
rect 37473 37349 37507 37383
rect 37565 37349 37599 37383
rect 1409 37281 1443 37315
rect 13369 37281 13403 37315
rect 15301 37281 15335 37315
rect 16037 37281 16071 37315
rect 16313 37281 16347 37315
rect 18613 37281 18647 37315
rect 19809 37281 19843 37315
rect 22109 37281 22143 37315
rect 24685 37281 24719 37315
rect 28641 37281 28675 37315
rect 31769 37281 31803 37315
rect 34069 37281 34103 37315
rect 34989 37281 35023 37315
rect 37197 37281 37231 37315
rect 40141 37281 40175 37315
rect 4721 37213 4755 37247
rect 4997 37213 5031 37247
rect 5181 37213 5215 37247
rect 5273 37213 5307 37247
rect 7113 37213 7147 37247
rect 7665 37213 7699 37247
rect 8125 37213 8159 37247
rect 8217 37213 8251 37247
rect 8493 37213 8527 37247
rect 8585 37213 8619 37247
rect 8769 37213 8803 37247
rect 8953 37213 8987 37247
rect 12265 37213 12299 37247
rect 13553 37213 13587 37247
rect 14289 37213 14323 37247
rect 14473 37213 14507 37247
rect 14565 37213 14599 37247
rect 18429 37213 18463 37247
rect 18797 37213 18831 37247
rect 18981 37213 19015 37247
rect 19073 37213 19107 37247
rect 19625 37213 19659 37247
rect 22385 37213 22419 37247
rect 22477 37213 22511 37247
rect 24409 37213 24443 37247
rect 26249 37213 26283 37247
rect 30205 37213 30239 37247
rect 32597 37213 32631 37247
rect 33149 37213 33183 37247
rect 33977 37213 34011 37247
rect 34161 37213 34195 37247
rect 34253 37213 34287 37247
rect 34437 37213 34471 37247
rect 34805 37213 34839 37247
rect 35081 37213 35115 37247
rect 35265 37213 35299 37247
rect 35357 37213 35391 37247
rect 35449 37213 35483 37247
rect 35541 37213 35575 37247
rect 37381 37213 37415 37247
rect 37657 37213 37691 37247
rect 37841 37213 37875 37247
rect 39681 37213 39715 37247
rect 39865 37213 39899 37247
rect 40049 37213 40083 37247
rect 1685 37145 1719 37179
rect 3617 37145 3651 37179
rect 7849 37145 7883 37179
rect 12357 37145 12391 37179
rect 13093 37145 13127 37179
rect 15853 37145 15887 37179
rect 22753 37145 22787 37179
rect 26525 37145 26559 37179
rect 28917 37145 28951 37179
rect 31585 37145 31619 37179
rect 32045 37145 32079 37179
rect 32965 37145 32999 37179
rect 36001 37145 36035 37179
rect 39405 37145 39439 37179
rect 39589 37145 39623 37179
rect 40417 37145 40451 37179
rect 3417 37077 3451 37111
rect 4997 37077 5031 37111
rect 8033 37077 8067 37111
rect 8401 37077 8435 37111
rect 14657 37077 14691 37111
rect 17785 37077 17819 37111
rect 17877 37077 17911 37111
rect 19257 37077 19291 37111
rect 19717 37077 19751 37111
rect 28089 37077 28123 37111
rect 29653 37077 29687 37111
rect 31217 37077 31251 37111
rect 31677 37077 31711 37111
rect 32781 37077 32815 37111
rect 41889 37077 41923 37111
rect 2513 36873 2547 36907
rect 4261 36873 4295 36907
rect 5181 36873 5215 36907
rect 5365 36873 5399 36907
rect 8585 36873 8619 36907
rect 14657 36873 14691 36907
rect 16497 36873 16531 36907
rect 17417 36873 17451 36907
rect 19901 36873 19935 36907
rect 22477 36873 22511 36907
rect 22845 36873 22879 36907
rect 24869 36873 24903 36907
rect 26985 36873 27019 36907
rect 27905 36873 27939 36907
rect 31953 36873 31987 36907
rect 36921 36873 36955 36907
rect 38025 36873 38059 36907
rect 38951 36873 38985 36907
rect 40141 36873 40175 36907
rect 2789 36805 2823 36839
rect 3019 36805 3053 36839
rect 3433 36805 3467 36839
rect 4169 36805 4203 36839
rect 8677 36805 8711 36839
rect 9045 36805 9079 36839
rect 13185 36805 13219 36839
rect 18429 36805 18463 36839
rect 24041 36805 24075 36839
rect 25329 36805 25363 36839
rect 27353 36805 27387 36839
rect 30481 36805 30515 36839
rect 32873 36805 32907 36839
rect 33793 36805 33827 36839
rect 34009 36805 34043 36839
rect 34713 36805 34747 36839
rect 36001 36805 36035 36839
rect 36645 36805 36679 36839
rect 37013 36805 37047 36839
rect 38117 36805 38151 36839
rect 38393 36805 38427 36839
rect 39037 36805 39071 36839
rect 2697 36737 2731 36771
rect 2881 36737 2915 36771
rect 3157 36737 3191 36771
rect 4445 36737 4479 36771
rect 4537 36737 4571 36771
rect 4629 36737 4663 36771
rect 4767 36737 4801 36771
rect 5273 36737 5307 36771
rect 6561 36737 6595 36771
rect 6745 36737 6779 36771
rect 10333 36737 10367 36771
rect 10517 36737 10551 36771
rect 10609 36737 10643 36771
rect 12449 36737 12483 36771
rect 12633 36737 12667 36771
rect 17233 36737 17267 36771
rect 17601 36737 17635 36771
rect 17693 36737 17727 36771
rect 17969 36737 18003 36771
rect 18153 36737 18187 36771
rect 21925 36737 21959 36771
rect 22109 36737 22143 36771
rect 23305 36737 23339 36771
rect 25237 36737 25271 36771
rect 25789 36737 25823 36771
rect 26341 36737 26375 36771
rect 27445 36737 27479 36771
rect 27813 36737 27847 36771
rect 27997 36737 28031 36771
rect 29653 36737 29687 36771
rect 30205 36737 30239 36771
rect 32597 36737 32631 36771
rect 34253 36737 34287 36771
rect 34345 36737 34379 36771
rect 34529 36737 34563 36771
rect 36185 36737 36219 36771
rect 36369 36737 36403 36771
rect 36461 36737 36495 36771
rect 36737 36737 36771 36771
rect 36829 36737 36863 36771
rect 37105 36737 37139 36771
rect 38025 36737 38059 36771
rect 38301 36737 38335 36771
rect 38577 36737 38611 36771
rect 38761 36737 38795 36771
rect 38853 36737 38887 36771
rect 39129 36737 39163 36771
rect 39497 36737 39531 36771
rect 41889 36737 41923 36771
rect 4905 36669 4939 36703
rect 6837 36669 6871 36703
rect 7113 36669 7147 36703
rect 11345 36669 11379 36703
rect 12081 36669 12115 36703
rect 12909 36669 12943 36703
rect 14749 36669 14783 36703
rect 15025 36669 15059 36703
rect 17877 36669 17911 36703
rect 20545 36669 20579 36703
rect 22937 36669 22971 36703
rect 23121 36669 23155 36703
rect 25513 36669 25547 36703
rect 27537 36669 27571 36703
rect 33149 36669 33183 36703
rect 41613 36669 41647 36703
rect 4997 36601 5031 36635
rect 34161 36601 34195 36635
rect 34529 36601 34563 36635
rect 36461 36601 36495 36635
rect 5549 36533 5583 36567
rect 6653 36533 6687 36567
rect 10149 36533 10183 36567
rect 10701 36533 10735 36567
rect 11529 36533 11563 36567
rect 12265 36533 12299 36567
rect 16681 36533 16715 36567
rect 19993 36533 20027 36567
rect 29101 36533 29135 36567
rect 32321 36533 32355 36567
rect 33977 36533 34011 36567
rect 34805 36533 34839 36567
rect 40049 36533 40083 36567
rect 6929 36329 6963 36363
rect 11345 36329 11379 36363
rect 14105 36329 14139 36363
rect 15761 36329 15795 36363
rect 29377 36329 29411 36363
rect 29561 36329 29595 36363
rect 35449 36329 35483 36363
rect 36829 36329 36863 36363
rect 39313 36329 39347 36363
rect 40785 36329 40819 36363
rect 4077 36261 4111 36295
rect 26709 36261 26743 36295
rect 3433 36193 3467 36227
rect 7573 36193 7607 36227
rect 9873 36193 9907 36227
rect 12265 36193 12299 36227
rect 14565 36193 14599 36227
rect 14657 36193 14691 36227
rect 16405 36193 16439 36227
rect 17141 36193 17175 36227
rect 19809 36193 19843 36227
rect 20361 36193 20395 36227
rect 22201 36193 22235 36227
rect 23949 36193 23983 36227
rect 25697 36193 25731 36227
rect 31309 36193 31343 36227
rect 31861 36193 31895 36227
rect 31953 36193 31987 36227
rect 33517 36193 33551 36227
rect 34345 36193 34379 36227
rect 36001 36193 36035 36227
rect 40141 36193 40175 36227
rect 41613 36193 41647 36227
rect 2973 36125 3007 36159
rect 3065 36125 3099 36159
rect 3893 36125 3927 36159
rect 3985 36125 4019 36159
rect 4169 36125 4203 36159
rect 7113 36125 7147 36159
rect 7297 36125 7331 36159
rect 7849 36125 7883 36159
rect 8033 36125 8067 36159
rect 9597 36125 9631 36159
rect 12081 36125 12115 36159
rect 12173 36125 12207 36159
rect 12817 36125 12851 36159
rect 13829 36125 13863 36159
rect 16129 36125 16163 36159
rect 19625 36125 19659 36159
rect 24961 36125 24995 36159
rect 26433 36125 26467 36159
rect 26985 36125 27019 36159
rect 27629 36125 27663 36159
rect 32781 36125 32815 36159
rect 35265 36125 35299 36159
rect 35817 36125 35851 36159
rect 35909 36125 35943 36159
rect 36093 36125 36127 36159
rect 36369 36125 36403 36159
rect 36737 36125 36771 36159
rect 36921 36125 36955 36159
rect 37381 36125 37415 36159
rect 39221 36125 39255 36159
rect 39405 36125 39439 36159
rect 40877 36125 40911 36159
rect 3157 36057 3191 36091
rect 3295 36057 3329 36091
rect 7205 36057 7239 36091
rect 7435 36057 7469 36091
rect 15577 36057 15611 36091
rect 20637 36057 20671 36091
rect 22477 36057 22511 36091
rect 27905 36057 27939 36091
rect 31033 36057 31067 36091
rect 31769 36057 31803 36091
rect 32229 36057 32263 36091
rect 33333 36057 33367 36091
rect 34161 36057 34195 36091
rect 34713 36057 34747 36091
rect 35633 36057 35667 36091
rect 37657 36057 37691 36091
rect 40417 36057 40451 36091
rect 2789 35989 2823 36023
rect 4353 35989 4387 36023
rect 7665 35989 7699 36023
rect 11713 35989 11747 36023
rect 13369 35989 13403 36023
rect 13737 35989 13771 36023
rect 14473 35989 14507 36023
rect 15485 35989 15519 36023
rect 16221 35989 16255 36023
rect 16589 35989 16623 36023
rect 16957 35989 16991 36023
rect 17049 35989 17083 36023
rect 19257 35989 19291 36023
rect 19717 35989 19751 36023
rect 22109 35989 22143 36023
rect 24409 35989 24443 36023
rect 25145 35989 25179 36023
rect 27537 35989 27571 36023
rect 31401 35989 31435 36023
rect 32965 35989 32999 36023
rect 33425 35989 33459 36023
rect 33793 35989 33827 36023
rect 34253 35989 34287 36023
rect 36553 35989 36587 36023
rect 39129 35989 39163 36023
rect 40325 35989 40359 36023
rect 6101 35785 6135 35819
rect 11023 35785 11057 35819
rect 13553 35785 13587 35819
rect 14657 35785 14691 35819
rect 16957 35785 16991 35819
rect 17417 35785 17451 35819
rect 21833 35785 21867 35819
rect 22937 35785 22971 35819
rect 23305 35785 23339 35819
rect 27353 35785 27387 35819
rect 28273 35785 28307 35819
rect 28641 35785 28675 35819
rect 29745 35785 29779 35819
rect 31953 35785 31987 35819
rect 34253 35785 34287 35819
rect 37933 35785 37967 35819
rect 40233 35785 40267 35819
rect 40601 35785 40635 35819
rect 41061 35785 41095 35819
rect 5733 35717 5767 35751
rect 11805 35717 11839 35751
rect 18245 35717 18279 35751
rect 30481 35717 30515 35751
rect 34345 35717 34379 35751
rect 37381 35717 37415 35751
rect 38393 35717 38427 35751
rect 4261 35649 4295 35683
rect 5181 35649 5215 35683
rect 5273 35649 5307 35683
rect 5365 35649 5399 35683
rect 5503 35649 5537 35683
rect 5917 35649 5951 35683
rect 7573 35649 7607 35683
rect 7757 35649 7791 35683
rect 13828 35649 13862 35683
rect 13921 35649 13955 35683
rect 15025 35649 15059 35683
rect 15485 35649 15519 35683
rect 17049 35649 17083 35683
rect 20177 35649 20211 35683
rect 20269 35649 20303 35683
rect 22201 35649 22235 35683
rect 23397 35649 23431 35683
rect 24133 35649 24167 35683
rect 30205 35649 30239 35683
rect 35909 35649 35943 35683
rect 36369 35649 36403 35683
rect 36921 35649 36955 35683
rect 38301 35649 38335 35683
rect 38761 35649 38795 35683
rect 39313 35649 39347 35683
rect 41429 35649 41463 35683
rect 1409 35581 1443 35615
rect 1685 35581 1719 35615
rect 3341 35581 3375 35615
rect 3617 35581 3651 35615
rect 4905 35581 4939 35615
rect 5641 35581 5675 35615
rect 9229 35581 9263 35615
rect 9597 35581 9631 35615
rect 11529 35581 11563 35615
rect 15117 35581 15151 35615
rect 15301 35581 15335 35615
rect 16497 35581 16531 35615
rect 16865 35581 16899 35615
rect 17969 35581 18003 35615
rect 19717 35581 19751 35615
rect 20453 35581 20487 35615
rect 22293 35581 22327 35615
rect 22477 35581 22511 35615
rect 23489 35581 23523 35615
rect 24409 35581 24443 35615
rect 25881 35581 25915 35615
rect 26525 35581 26559 35615
rect 27445 35581 27479 35615
rect 27629 35581 27663 35615
rect 28733 35581 28767 35615
rect 28917 35581 28951 35615
rect 29561 35581 29595 35615
rect 29653 35581 29687 35615
rect 32505 35581 32539 35615
rect 32781 35581 32815 35615
rect 34897 35581 34931 35615
rect 36001 35581 36035 35615
rect 36093 35581 36127 35615
rect 38485 35581 38519 35615
rect 40693 35581 40727 35615
rect 40785 35581 40819 35615
rect 41521 35581 41555 35615
rect 41613 35581 41647 35615
rect 4997 35513 5031 35547
rect 19809 35513 19843 35547
rect 25973 35513 26007 35547
rect 3157 35445 3191 35479
rect 7757 35445 7791 35479
rect 13277 35445 13311 35479
rect 15669 35445 15703 35479
rect 15853 35445 15887 35479
rect 26985 35445 27019 35479
rect 30113 35445 30147 35479
rect 35541 35445 35575 35479
rect 37473 35445 37507 35479
rect 3617 35241 3651 35275
rect 4537 35241 4571 35275
rect 9873 35241 9907 35275
rect 12357 35241 12391 35275
rect 14197 35241 14231 35275
rect 15945 35241 15979 35275
rect 19349 35241 19383 35275
rect 22477 35241 22511 35275
rect 23489 35241 23523 35275
rect 24777 35241 24811 35275
rect 27629 35241 27663 35275
rect 31401 35241 31435 35275
rect 36737 35241 36771 35275
rect 40417 35241 40451 35275
rect 41245 35241 41279 35275
rect 4261 35173 4295 35207
rect 14657 35173 14691 35207
rect 22385 35173 22419 35207
rect 1869 35105 1903 35139
rect 2145 35105 2179 35139
rect 4813 35105 4847 35139
rect 7021 35105 7055 35139
rect 10609 35105 10643 35139
rect 13645 35105 13679 35139
rect 15301 35105 15335 35139
rect 18429 35105 18463 35139
rect 19993 35105 20027 35139
rect 20361 35105 20395 35139
rect 21833 35105 21867 35139
rect 23029 35105 23063 35139
rect 24087 35105 24121 35139
rect 25329 35105 25363 35139
rect 25881 35105 25915 35139
rect 28825 35105 28859 35139
rect 31953 35105 31987 35139
rect 34989 35105 35023 35139
rect 37381 35105 37415 35139
rect 38485 35105 38519 35139
rect 39313 35105 39347 35139
rect 40969 35105 41003 35139
rect 41797 35105 41831 35139
rect 3801 35037 3835 35071
rect 4077 35037 4111 35071
rect 10057 35037 10091 35071
rect 10333 35037 10367 35071
rect 10517 35037 10551 35071
rect 13553 35037 13587 35071
rect 14105 35037 14139 35071
rect 14289 35037 14323 35071
rect 15025 35037 15059 35071
rect 17325 35037 17359 35071
rect 17417 35037 17451 35071
rect 19809 35037 19843 35071
rect 25145 35037 25179 35071
rect 30113 35037 30147 35071
rect 4353 34969 4387 35003
rect 5096 34969 5130 35003
rect 7297 34969 7331 35003
rect 10885 34969 10919 35003
rect 17058 34969 17092 35003
rect 22017 34969 22051 35003
rect 22937 34969 22971 35003
rect 26157 34969 26191 35003
rect 28549 34969 28583 35003
rect 29561 34969 29595 35003
rect 32229 34969 32263 35003
rect 35265 34969 35299 35003
rect 38301 34969 38335 35003
rect 38761 34969 38795 35003
rect 39957 34969 39991 35003
rect 40785 34969 40819 35003
rect 41705 34969 41739 35003
rect 3893 34901 3927 34935
rect 4553 34901 4587 34935
rect 4721 34901 4755 34935
rect 6561 34901 6595 34935
rect 8769 34901 8803 34935
rect 13921 34901 13955 34935
rect 15117 34901 15151 34935
rect 17877 34901 17911 34935
rect 19717 34901 19751 34935
rect 21005 34901 21039 34935
rect 21925 34901 21959 34935
rect 22845 34901 22879 34935
rect 23857 34901 23891 34935
rect 23949 34901 23983 34935
rect 25237 34901 25271 34935
rect 28181 34901 28215 34935
rect 28641 34901 28675 34935
rect 31769 34901 31803 34935
rect 31861 34901 31895 34935
rect 33517 34901 33551 34935
rect 36829 34901 36863 34935
rect 37933 34901 37967 34935
rect 38393 34901 38427 34935
rect 40049 34901 40083 34935
rect 40877 34901 40911 34935
rect 41613 34901 41647 34935
rect 3433 34697 3467 34731
rect 4353 34697 4387 34731
rect 4813 34697 4847 34731
rect 12541 34697 12575 34731
rect 14013 34697 14047 34731
rect 16037 34697 16071 34731
rect 16497 34697 16531 34731
rect 18061 34697 18095 34731
rect 20085 34697 20119 34731
rect 20177 34697 20211 34731
rect 20637 34697 20671 34731
rect 23489 34697 23523 34731
rect 23857 34697 23891 34731
rect 25237 34697 25271 34731
rect 26065 34697 26099 34731
rect 29193 34697 29227 34731
rect 30021 34697 30055 34731
rect 34161 34697 34195 34731
rect 39129 34697 39163 34731
rect 40785 34697 40819 34731
rect 40969 34697 41003 34731
rect 41429 34697 41463 34731
rect 6653 34629 6687 34663
rect 8553 34629 8587 34663
rect 8769 34629 8803 34663
rect 10977 34629 11011 34663
rect 11529 34629 11563 34663
rect 16129 34629 16163 34663
rect 18972 34629 19006 34663
rect 22201 34629 22235 34663
rect 25605 34629 25639 34663
rect 26525 34629 26559 34663
rect 27721 34629 27755 34663
rect 30389 34629 30423 34663
rect 31309 34629 31343 34663
rect 32689 34629 32723 34663
rect 37657 34629 37691 34663
rect 3433 34561 3467 34595
rect 3617 34561 3651 34595
rect 4445 34561 4479 34595
rect 5089 34561 5123 34595
rect 5365 34561 5399 34595
rect 5457 34561 5491 34595
rect 7849 34561 7883 34595
rect 7941 34561 7975 34595
rect 10609 34561 10643 34595
rect 10793 34561 10827 34595
rect 12909 34561 12943 34595
rect 14105 34561 14139 34595
rect 14372 34561 14406 34595
rect 16681 34561 16715 34595
rect 16948 34561 16982 34595
rect 18705 34561 18739 34595
rect 20545 34561 20579 34595
rect 22293 34561 22327 34595
rect 22661 34561 22695 34595
rect 23213 34561 23247 34595
rect 24869 34561 24903 34595
rect 26433 34561 26467 34595
rect 29377 34561 29411 34595
rect 30481 34561 30515 34595
rect 31217 34561 31251 34595
rect 32413 34561 32447 34595
rect 34805 34561 34839 34595
rect 39405 34561 39439 34595
rect 39672 34561 39706 34595
rect 41337 34561 41371 34595
rect 4997 34493 5031 34527
rect 5549 34493 5583 34527
rect 7389 34493 7423 34527
rect 8217 34493 8251 34527
rect 8309 34493 8343 34527
rect 13001 34493 13035 34527
rect 13185 34493 13219 34527
rect 13461 34493 13495 34527
rect 15853 34493 15887 34527
rect 20821 34493 20855 34527
rect 22385 34493 22419 34527
rect 23949 34493 23983 34527
rect 24041 34493 24075 34527
rect 25697 34493 25731 34527
rect 25789 34493 25823 34527
rect 26617 34493 26651 34527
rect 27445 34493 27479 34527
rect 30665 34493 30699 34527
rect 31493 34493 31527 34527
rect 36553 34493 36587 34527
rect 37381 34493 37415 34527
rect 41521 34493 41555 34527
rect 7665 34425 7699 34459
rect 29653 34425 29687 34459
rect 6193 34357 6227 34391
rect 8401 34357 8435 34391
rect 8585 34357 8619 34391
rect 15485 34357 15519 34391
rect 21833 34357 21867 34391
rect 24317 34357 24351 34391
rect 30849 34357 30883 34391
rect 35062 34357 35096 34391
rect 5273 34153 5307 34187
rect 8033 34153 8067 34187
rect 8125 34153 8159 34187
rect 9689 34153 9723 34187
rect 13185 34153 13219 34187
rect 14197 34153 14231 34187
rect 14933 34153 14967 34187
rect 22293 34153 22327 34187
rect 24225 34153 24259 34187
rect 27813 34153 27847 34187
rect 28641 34153 28675 34187
rect 29561 34153 29595 34187
rect 31493 34153 31527 34187
rect 34161 34153 34195 34187
rect 34989 34153 35023 34187
rect 36645 34153 36679 34187
rect 38209 34153 38243 34187
rect 41981 34153 42015 34187
rect 25973 34085 26007 34119
rect 26985 34085 27019 34119
rect 5457 34017 5491 34051
rect 5825 34017 5859 34051
rect 5917 34017 5951 34051
rect 10701 34017 10735 34051
rect 13093 34017 13127 34051
rect 14381 34017 14415 34051
rect 15485 34017 15519 34051
rect 19257 34017 19291 34051
rect 20913 34017 20947 34051
rect 22845 34017 22879 34051
rect 24593 34017 24627 34051
rect 26617 34017 26651 34051
rect 27537 34017 27571 34051
rect 28365 34017 28399 34051
rect 29285 34017 29319 34051
rect 30205 34017 30239 34051
rect 31953 34017 31987 34051
rect 32137 34017 32171 34051
rect 33609 34017 33643 34051
rect 35633 34017 35667 34051
rect 36461 34017 36495 34051
rect 37197 34017 37231 34051
rect 38853 34017 38887 34051
rect 39129 34017 39163 34051
rect 40509 34017 40543 34051
rect 5549 33949 5583 33983
rect 6009 33949 6043 33983
rect 6285 33949 6319 33983
rect 6469 33949 6503 33983
rect 7297 33949 7331 33983
rect 7481 33949 7515 33983
rect 7757 33949 7791 33983
rect 7849 33949 7883 33983
rect 8401 33949 8435 33983
rect 8585 33949 8619 33983
rect 9505 33949 9539 33983
rect 9965 33949 9999 33983
rect 10149 33949 10183 33983
rect 13829 33949 13863 33983
rect 14473 33949 14507 33983
rect 15761 33949 15795 33983
rect 17049 33949 17083 33983
rect 17969 33949 18003 33983
rect 18521 33949 18555 33983
rect 21180 33949 21214 33983
rect 27353 33949 27387 33983
rect 29009 33949 29043 33983
rect 32413 33949 32447 33983
rect 33701 33949 33735 33983
rect 35357 33949 35391 33983
rect 40601 33949 40635 33983
rect 7665 33881 7699 33915
rect 8953 33881 8987 33915
rect 11345 33881 11379 33915
rect 16497 33881 16531 33915
rect 17233 33881 17267 33915
rect 19073 33881 19107 33915
rect 19502 33881 19536 33915
rect 23112 33881 23146 33915
rect 24860 33881 24894 33915
rect 37013 33881 37047 33915
rect 38577 33881 38611 33915
rect 40868 33881 40902 33915
rect 6193 33813 6227 33847
rect 8309 33813 8343 33847
rect 9873 33813 9907 33847
rect 11253 33813 11287 33847
rect 15301 33813 15335 33847
rect 15393 33813 15427 33847
rect 16405 33813 16439 33847
rect 20637 33813 20671 33847
rect 26065 33813 26099 33847
rect 27445 33813 27479 33847
rect 28181 33813 28215 33847
rect 28273 33813 28307 33847
rect 29101 33813 29135 33847
rect 29929 33813 29963 33847
rect 30021 33813 30055 33847
rect 31861 33813 31895 33847
rect 33057 33813 33091 33847
rect 33793 33813 33827 33847
rect 35449 33813 35483 33847
rect 35817 33813 35851 33847
rect 36185 33813 36219 33847
rect 36277 33813 36311 33847
rect 37105 33813 37139 33847
rect 38669 33813 38703 33847
rect 39681 33813 39715 33847
rect 39865 33813 39899 33847
rect 5273 33609 5307 33643
rect 6377 33609 6411 33643
rect 9873 33609 9907 33643
rect 13369 33609 13403 33643
rect 14197 33609 14231 33643
rect 15669 33609 15703 33643
rect 16129 33609 16163 33643
rect 17141 33609 17175 33643
rect 17601 33609 17635 33643
rect 19993 33609 20027 33643
rect 23397 33609 23431 33643
rect 23857 33609 23891 33643
rect 25053 33609 25087 33643
rect 25513 33609 25547 33643
rect 30849 33609 30883 33643
rect 32597 33609 32631 33643
rect 33425 33609 33459 33643
rect 39497 33609 39531 33643
rect 39589 33609 39623 33643
rect 39957 33609 39991 33643
rect 40417 33609 40451 33643
rect 40785 33609 40819 33643
rect 3985 33541 4019 33575
rect 8033 33541 8067 33575
rect 8401 33541 8435 33575
rect 15332 33541 15366 33575
rect 17509 33541 17543 33575
rect 20361 33541 20395 33575
rect 23765 33541 23799 33575
rect 35817 33541 35851 33575
rect 38669 33541 38703 33575
rect 41245 33541 41279 33575
rect 1409 33473 1443 33507
rect 3433 33473 3467 33507
rect 3893 33473 3927 33507
rect 4169 33473 4203 33507
rect 5089 33473 5123 33507
rect 6561 33473 6595 33507
rect 6653 33473 6687 33507
rect 7021 33473 7055 33507
rect 7297 33473 7331 33507
rect 7757 33473 7791 33507
rect 10232 33473 10266 33507
rect 11989 33473 12023 33507
rect 12256 33473 12290 33507
rect 14013 33473 14047 33507
rect 16037 33473 16071 33507
rect 18153 33473 18187 33507
rect 20453 33473 20487 33507
rect 20821 33473 20855 33507
rect 21373 33473 21407 33507
rect 21833 33473 21867 33507
rect 22100 33473 22134 33507
rect 25421 33473 25455 33507
rect 28733 33473 28767 33507
rect 29736 33473 29770 33507
rect 31493 33473 31527 33507
rect 32505 33473 32539 33507
rect 33793 33473 33827 33507
rect 33885 33473 33919 33507
rect 35909 33473 35943 33507
rect 36277 33473 36311 33507
rect 37289 33473 37323 33507
rect 40325 33473 40359 33507
rect 41153 33473 41187 33507
rect 1685 33405 1719 33439
rect 3525 33405 3559 33439
rect 3617 33405 3651 33439
rect 3709 33405 3743 33439
rect 7113 33405 7147 33439
rect 7389 33405 7423 33439
rect 7849 33405 7883 33439
rect 8125 33405 8159 33439
rect 9965 33405 9999 33439
rect 15577 33405 15611 33439
rect 16221 33405 16255 33439
rect 17693 33405 17727 33439
rect 18429 33405 18463 33439
rect 19901 33405 19935 33439
rect 20637 33405 20671 33439
rect 23949 33405 23983 33439
rect 24777 33405 24811 33439
rect 25697 33405 25731 33439
rect 29469 33405 29503 33439
rect 32781 33405 32815 33439
rect 33977 33405 34011 33439
rect 36001 33405 36035 33439
rect 36829 33405 36863 33439
rect 38025 33405 38059 33439
rect 38761 33405 38795 33439
rect 38945 33405 38979 33439
rect 39773 33405 39807 33439
rect 40509 33405 40543 33439
rect 41337 33405 41371 33439
rect 23213 33337 23247 33371
rect 30941 33337 30975 33371
rect 39129 33337 39163 33371
rect 3157 33269 3191 33303
rect 3249 33269 3283 33303
rect 4169 33269 4203 33303
rect 6837 33269 6871 33303
rect 7113 33269 7147 33303
rect 11345 33269 11379 33303
rect 13461 33269 13495 33303
rect 24225 33269 24259 33303
rect 28641 33269 28675 33303
rect 32137 33269 32171 33303
rect 35449 33269 35483 33303
rect 38301 33269 38335 33303
rect 5917 33065 5951 33099
rect 7389 33065 7423 33099
rect 10241 33065 10275 33099
rect 10333 33065 10367 33099
rect 12817 33065 12851 33099
rect 16681 33065 16715 33099
rect 21741 33065 21775 33099
rect 22753 33065 22787 33099
rect 28365 33065 28399 33099
rect 29929 33065 29963 33099
rect 32229 33065 32263 33099
rect 38761 33065 38795 33099
rect 38853 33065 38887 33099
rect 4721 32997 4755 33031
rect 7113 32997 7147 33031
rect 12449 32997 12483 33031
rect 1685 32929 1719 32963
rect 4353 32929 4387 32963
rect 6009 32929 6043 32963
rect 10057 32929 10091 32963
rect 10977 32929 11011 32963
rect 11069 32929 11103 32963
rect 13369 32929 13403 32963
rect 17049 32929 17083 32963
rect 20085 32929 20119 32963
rect 21097 32929 21131 32963
rect 22385 32929 22419 32963
rect 24961 32929 24995 32963
rect 26341 32929 26375 32963
rect 26709 32929 26743 32963
rect 26801 32929 26835 32963
rect 28917 32929 28951 32963
rect 30481 32929 30515 32963
rect 39405 32929 39439 32963
rect 40969 32929 41003 32963
rect 41889 32929 41923 32963
rect 3985 32861 4019 32895
rect 4261 32861 4295 32895
rect 5181 32861 5215 32895
rect 5365 32861 5399 32895
rect 5457 32861 5491 32895
rect 5733 32861 5767 32895
rect 6837 32861 6871 32895
rect 6929 32861 6963 32895
rect 7113 32861 7147 32895
rect 7573 32861 7607 32895
rect 7665 32861 7699 32895
rect 7849 32861 7883 32895
rect 7941 32861 7975 32895
rect 9965 32861 9999 32895
rect 11325 32861 11359 32895
rect 13277 32861 13311 32895
rect 14105 32861 14139 32895
rect 14933 32861 14967 32895
rect 20913 32861 20947 32895
rect 22201 32861 22235 32895
rect 24133 32861 24167 32895
rect 26893 32861 26927 32895
rect 30389 32861 30423 32895
rect 30849 32861 30883 32895
rect 32597 32861 32631 32895
rect 35081 32861 35115 32895
rect 36921 32861 36955 32895
rect 37381 32861 37415 32895
rect 37648 32861 37682 32895
rect 1961 32793 1995 32827
rect 4169 32793 4203 32827
rect 9597 32793 9631 32827
rect 15209 32793 15243 32827
rect 17325 32793 17359 32827
rect 23866 32793 23900 32827
rect 27353 32793 27387 32827
rect 28181 32793 28215 32827
rect 31116 32793 31150 32827
rect 32864 32793 32898 32827
rect 35348 32793 35382 32827
rect 40785 32793 40819 32827
rect 3433 32725 3467 32759
rect 3801 32725 3835 32759
rect 4813 32725 4847 32759
rect 4997 32725 5031 32759
rect 5549 32725 5583 32759
rect 13185 32725 13219 32759
rect 14749 32725 14783 32759
rect 18797 32725 18831 32759
rect 19533 32725 19567 32759
rect 22109 32725 22143 32759
rect 24409 32725 24443 32759
rect 25789 32725 25823 32759
rect 27261 32725 27295 32759
rect 30297 32725 30331 32759
rect 33977 32725 34011 32759
rect 36461 32725 36495 32759
rect 40417 32725 40451 32759
rect 40877 32725 40911 32759
rect 41337 32725 41371 32759
rect 2145 32521 2179 32555
rect 2789 32521 2823 32555
rect 3433 32521 3467 32555
rect 12633 32521 12667 32555
rect 14105 32521 14139 32555
rect 14565 32521 14599 32555
rect 17785 32521 17819 32555
rect 18153 32521 18187 32555
rect 18613 32521 18647 32555
rect 23397 32521 23431 32555
rect 23857 32521 23891 32555
rect 26157 32521 26191 32555
rect 28365 32521 28399 32555
rect 33149 32521 33183 32555
rect 36461 32521 36495 32555
rect 38761 32521 38795 32555
rect 41705 32521 41739 32555
rect 8125 32453 8159 32487
rect 13768 32453 13802 32487
rect 18981 32453 19015 32487
rect 19349 32453 19383 32487
rect 19717 32453 19751 32487
rect 35348 32453 35382 32487
rect 40592 32453 40626 32487
rect 2329 32385 2363 32419
rect 2513 32385 2547 32419
rect 3341 32385 3375 32419
rect 3617 32385 3651 32419
rect 3801 32385 3835 32419
rect 3893 32385 3927 32419
rect 7297 32385 7331 32419
rect 8401 32385 8435 32419
rect 8953 32385 8987 32419
rect 14013 32385 14047 32419
rect 14473 32385 14507 32419
rect 18751 32385 18785 32419
rect 18889 32385 18923 32419
rect 19164 32385 19198 32419
rect 19257 32385 19291 32419
rect 23765 32385 23799 32419
rect 24777 32385 24811 32419
rect 25044 32385 25078 32419
rect 26985 32385 27019 32419
rect 27252 32385 27286 32419
rect 28713 32385 28747 32419
rect 29929 32385 29963 32419
rect 33517 32385 33551 32419
rect 33609 32385 33643 32419
rect 33977 32385 34011 32419
rect 34529 32385 34563 32419
rect 35081 32385 35115 32419
rect 37648 32385 37682 32419
rect 39405 32385 39439 32419
rect 40325 32385 40359 32419
rect 41889 32385 41923 32419
rect 3065 32317 3099 32351
rect 4261 32317 4295 32351
rect 4537 32317 4571 32351
rect 8033 32317 8067 32351
rect 8493 32317 8527 32351
rect 9137 32317 9171 32351
rect 10057 32317 10091 32351
rect 14657 32317 14691 32351
rect 18245 32317 18279 32351
rect 18337 32317 18371 32351
rect 19901 32317 19935 32351
rect 20177 32317 20211 32351
rect 21649 32317 21683 32351
rect 24041 32317 24075 32351
rect 28457 32317 28491 32351
rect 31217 32317 31251 32351
rect 32137 32317 32171 32351
rect 33793 32317 33827 32351
rect 37381 32317 37415 32351
rect 8769 32249 8803 32283
rect 29837 32249 29871 32283
rect 3249 32181 3283 32215
rect 6009 32181 6043 32215
rect 7941 32181 7975 32215
rect 8677 32181 8711 32215
rect 10609 32181 10643 32215
rect 30573 32181 30607 32215
rect 30665 32181 30699 32215
rect 32781 32181 32815 32215
rect 38853 32181 38887 32215
rect 42073 32181 42107 32215
rect 3157 31977 3191 32011
rect 4721 31977 4755 32011
rect 5641 31977 5675 32011
rect 6377 31977 6411 32011
rect 6653 31977 6687 32011
rect 8677 31977 8711 32011
rect 9321 31977 9355 32011
rect 12357 31977 12391 32011
rect 13553 31977 13587 32011
rect 15669 31977 15703 32011
rect 16129 31977 16163 32011
rect 18061 31977 18095 32011
rect 21833 31977 21867 32011
rect 25237 31977 25271 32011
rect 28549 31977 28583 32011
rect 31033 31977 31067 32011
rect 35449 31977 35483 32011
rect 37841 31977 37875 32011
rect 41337 31977 41371 32011
rect 16313 31909 16347 31943
rect 17049 31909 17083 31943
rect 21281 31909 21315 31943
rect 27813 31909 27847 31943
rect 33977 31909 34011 31943
rect 34253 31909 34287 31943
rect 41245 31909 41279 31943
rect 4997 31841 5031 31875
rect 5089 31841 5123 31875
rect 5457 31841 5491 31875
rect 11161 31841 11195 31875
rect 18889 31841 18923 31875
rect 24041 31841 24075 31875
rect 25697 31841 25731 31875
rect 25789 31841 25823 31875
rect 26433 31841 26467 31875
rect 29009 31841 29043 31875
rect 29101 31841 29135 31875
rect 29561 31841 29595 31875
rect 35265 31841 35299 31875
rect 36001 31841 36035 31875
rect 36829 31841 36863 31875
rect 38301 31841 38335 31875
rect 38393 31841 38427 31875
rect 39037 31841 39071 31875
rect 39221 31841 39255 31875
rect 41889 31841 41923 31875
rect 3341 31773 3375 31807
rect 4905 31773 4939 31807
rect 5181 31773 5215 31807
rect 5549 31773 5583 31807
rect 5641 31773 5675 31807
rect 5825 31773 5859 31807
rect 6653 31773 6687 31807
rect 6837 31773 6871 31807
rect 6929 31773 6963 31807
rect 11069 31773 11103 31807
rect 11713 31773 11747 31807
rect 12173 31773 12207 31807
rect 12357 31773 12391 31807
rect 13829 31773 13863 31807
rect 15853 31773 15887 31807
rect 15945 31773 15979 31807
rect 16221 31773 16255 31807
rect 16497 31773 16531 31807
rect 16589 31773 16623 31807
rect 16681 31773 16715 31807
rect 16865 31773 16899 31807
rect 17233 31773 17267 31807
rect 17325 31773 17359 31807
rect 17509 31773 17543 31807
rect 18199 31773 18233 31807
rect 18337 31773 18371 31807
rect 18429 31773 18463 31807
rect 18612 31773 18646 31807
rect 18705 31773 18739 31807
rect 18797 31773 18831 31807
rect 18981 31773 19015 31807
rect 20729 31773 20763 31807
rect 20913 31773 20947 31807
rect 21005 31773 21039 31807
rect 21097 31773 21131 31807
rect 21373 31773 21407 31807
rect 21557 31773 21591 31807
rect 21649 31773 21683 31807
rect 21925 31773 21959 31807
rect 23765 31773 23799 31807
rect 23857 31773 23891 31807
rect 24133 31773 24167 31807
rect 29828 31773 29862 31807
rect 32413 31773 32447 31807
rect 32597 31773 32631 31807
rect 32864 31773 32898 31807
rect 34069 31773 34103 31807
rect 35909 31773 35943 31807
rect 36277 31773 36311 31807
rect 39865 31773 39899 31807
rect 7205 31705 7239 31739
rect 10793 31705 10827 31739
rect 11897 31705 11931 31739
rect 26678 31705 26712 31739
rect 32146 31705 32180 31739
rect 40110 31705 40144 31739
rect 12541 31637 12575 31671
rect 17417 31637 17451 31671
rect 23581 31637 23615 31671
rect 25605 31637 25639 31671
rect 28917 31637 28951 31671
rect 30941 31637 30975 31671
rect 34713 31637 34747 31671
rect 35817 31637 35851 31671
rect 38209 31637 38243 31671
rect 39313 31637 39347 31671
rect 39681 31637 39715 31671
rect 2605 31433 2639 31467
rect 3919 31433 3953 31467
rect 5181 31433 5215 31467
rect 5349 31433 5383 31467
rect 5825 31433 5859 31467
rect 7573 31433 7607 31467
rect 12357 31433 12391 31467
rect 15485 31433 15519 31467
rect 15945 31433 15979 31467
rect 17049 31433 17083 31467
rect 17141 31433 17175 31467
rect 18061 31433 18095 31467
rect 19625 31433 19659 31467
rect 21373 31433 21407 31467
rect 24777 31433 24811 31467
rect 26157 31433 26191 31467
rect 28273 31433 28307 31467
rect 29745 31433 29779 31467
rect 30573 31433 30607 31467
rect 32597 31433 32631 31467
rect 33333 31433 33367 31467
rect 33793 31433 33827 31467
rect 42165 31433 42199 31467
rect 3709 31365 3743 31399
rect 5549 31365 5583 31399
rect 5641 31365 5675 31399
rect 8125 31365 8159 31399
rect 21005 31365 21039 31399
rect 21097 31365 21131 31399
rect 23213 31365 23247 31399
rect 25053 31365 25087 31399
rect 27353 31365 27387 31399
rect 29408 31365 29442 31399
rect 40049 31365 40083 31399
rect 2513 31297 2547 31331
rect 5917 31297 5951 31331
rect 6469 31297 6503 31331
rect 7757 31297 7791 31331
rect 7849 31297 7883 31331
rect 8217 31297 8251 31331
rect 11529 31297 11563 31331
rect 15025 31297 15059 31331
rect 16129 31297 16163 31331
rect 16221 31297 16255 31331
rect 16313 31297 16347 31331
rect 16497 31297 16531 31331
rect 17509 31297 17543 31331
rect 17693 31297 17727 31331
rect 17785 31297 17819 31331
rect 17877 31297 17911 31331
rect 18337 31297 18371 31331
rect 19717 31297 19751 31331
rect 19993 31297 20027 31331
rect 20085 31297 20119 31331
rect 20269 31297 20303 31331
rect 20361 31297 20395 31331
rect 20729 31297 20763 31331
rect 20877 31297 20911 31331
rect 21235 31297 21269 31331
rect 24961 31297 24995 31331
rect 25145 31297 25179 31331
rect 25329 31297 25363 31331
rect 27445 31297 27479 31331
rect 29653 31297 29687 31331
rect 30113 31297 30147 31331
rect 30205 31297 30239 31331
rect 30941 31297 30975 31331
rect 32505 31297 32539 31331
rect 33701 31297 33735 31331
rect 35081 31297 35115 31331
rect 35173 31297 35207 31331
rect 35449 31297 35483 31331
rect 37289 31297 37323 31331
rect 37565 31297 37599 31331
rect 37657 31297 37691 31331
rect 39957 31297 39991 31331
rect 40141 31297 40175 31331
rect 40325 31297 40359 31331
rect 40417 31297 40451 31331
rect 2789 31229 2823 31263
rect 2973 31229 3007 31263
rect 3525 31229 3559 31263
rect 9321 31229 9355 31263
rect 9597 31229 9631 31263
rect 11069 31229 11103 31263
rect 12081 31229 12115 31263
rect 14749 31229 14783 31263
rect 15209 31229 15243 31263
rect 15393 31229 15427 31263
rect 17233 31229 17267 31263
rect 22937 31229 22971 31263
rect 26801 31229 26835 31263
rect 27537 31229 27571 31263
rect 30297 31229 30331 31263
rect 31033 31229 31067 31263
rect 31125 31229 31159 31263
rect 32689 31229 32723 31263
rect 33977 31229 34011 31263
rect 40693 31229 40727 31263
rect 11897 31161 11931 31195
rect 24685 31161 24719 31195
rect 26985 31161 27019 31195
rect 35357 31161 35391 31195
rect 37381 31161 37415 31195
rect 2145 31093 2179 31127
rect 3893 31093 3927 31127
rect 4077 31093 4111 31127
rect 5365 31093 5399 31127
rect 5641 31093 5675 31127
rect 11989 31093 12023 31127
rect 13277 31093 13311 31127
rect 15853 31093 15887 31127
rect 16681 31093 16715 31127
rect 20545 31093 20579 31127
rect 32137 31093 32171 31127
rect 34897 31093 34931 31127
rect 37841 31093 37875 31127
rect 39773 31093 39807 31127
rect 3157 30889 3191 30923
rect 3249 30889 3283 30923
rect 5273 30889 5307 30923
rect 10793 30889 10827 30923
rect 12633 30889 12667 30923
rect 15025 30889 15059 30923
rect 16129 30889 16163 30923
rect 18061 30889 18095 30923
rect 19441 30889 19475 30923
rect 19901 30889 19935 30923
rect 20637 30889 20671 30923
rect 23581 30889 23615 30923
rect 24409 30889 24443 30923
rect 31033 30889 31067 30923
rect 32229 30889 32263 30923
rect 36461 30889 36495 30923
rect 37289 30889 37323 30923
rect 41061 30889 41095 30923
rect 3801 30821 3835 30855
rect 4721 30821 4755 30855
rect 1409 30753 1443 30787
rect 4813 30753 4847 30787
rect 5181 30753 5215 30787
rect 6929 30753 6963 30787
rect 10517 30753 10551 30787
rect 10885 30753 10919 30787
rect 13277 30753 13311 30787
rect 14381 30753 14415 30787
rect 15853 30753 15887 30787
rect 16589 30753 16623 30787
rect 18889 30753 18923 30787
rect 20821 30753 20855 30787
rect 21005 30753 21039 30787
rect 24777 30753 24811 30787
rect 25145 30753 25179 30787
rect 25329 30753 25363 30787
rect 30481 30753 30515 30787
rect 31585 30753 31619 30787
rect 32781 30753 32815 30787
rect 34713 30753 34747 30787
rect 34989 30753 35023 30787
rect 37657 30753 37691 30787
rect 40417 30753 40451 30787
rect 3433 30685 3467 30719
rect 3525 30685 3559 30719
rect 4077 30685 4111 30719
rect 4537 30685 4571 30719
rect 5641 30685 5675 30719
rect 5917 30685 5951 30719
rect 6101 30685 6135 30719
rect 10609 30685 10643 30719
rect 13461 30685 13495 30719
rect 13645 30685 13679 30719
rect 15577 30685 15611 30719
rect 15761 30685 15795 30719
rect 16313 30685 16347 30719
rect 16405 30685 16439 30719
rect 16681 30685 16715 30719
rect 17601 30663 17635 30697
rect 17693 30685 17727 30719
rect 17877 30685 17911 30719
rect 18153 30685 18187 30719
rect 19257 30685 19291 30719
rect 19441 30685 19475 30719
rect 19993 30685 20027 30719
rect 20177 30685 20211 30719
rect 20269 30685 20303 30719
rect 20381 30685 20415 30719
rect 21557 30685 21591 30719
rect 22017 30685 22051 30719
rect 23765 30685 23799 30719
rect 24133 30685 24167 30719
rect 24593 30685 24627 30719
rect 24685 30685 24719 30719
rect 24869 30685 24903 30719
rect 25053 30685 25087 30719
rect 27307 30685 27341 30719
rect 27445 30685 27479 30719
rect 27665 30685 27699 30719
rect 27813 30685 27847 30719
rect 28917 30685 28951 30719
rect 29837 30685 29871 30719
rect 30021 30685 30055 30719
rect 30573 30685 30607 30719
rect 30757 30685 30791 30719
rect 36645 30685 36679 30719
rect 36793 30685 36827 30719
rect 37013 30685 37047 30719
rect 37110 30685 37144 30719
rect 37381 30685 37415 30719
rect 40325 30685 40359 30719
rect 40877 30685 40911 30719
rect 1685 30617 1719 30651
rect 3801 30617 3835 30651
rect 5089 30617 5123 30651
rect 5549 30617 5583 30651
rect 6193 30617 6227 30651
rect 11161 30617 11195 30651
rect 17141 30617 17175 30651
rect 19533 30617 19567 30651
rect 19717 30617 19751 30651
rect 22201 30617 22235 30651
rect 23857 30617 23891 30651
rect 23949 30617 23983 30651
rect 27537 30617 27571 30651
rect 28733 30617 28767 30651
rect 29193 30617 29227 30651
rect 29561 30617 29595 30651
rect 29929 30617 29963 30651
rect 36921 30617 36955 30651
rect 40693 30617 40727 30651
rect 3985 30549 4019 30583
rect 4353 30549 4387 30583
rect 5457 30549 5491 30583
rect 5825 30549 5859 30583
rect 10149 30549 10183 30583
rect 12725 30549 12759 30583
rect 13553 30549 13587 30583
rect 15393 30549 15427 30583
rect 16865 30549 16899 30583
rect 21097 30549 21131 30583
rect 21465 30549 21499 30583
rect 21649 30549 21683 30583
rect 21833 30549 21867 30583
rect 25329 30549 25363 30583
rect 27169 30549 27203 30583
rect 28457 30549 28491 30583
rect 29101 30549 29135 30583
rect 30941 30549 30975 30583
rect 39129 30549 39163 30583
rect 39865 30549 39899 30583
rect 40233 30549 40267 30583
rect 3065 30345 3099 30379
rect 3249 30345 3283 30379
rect 4169 30345 4203 30379
rect 6377 30345 6411 30379
rect 11069 30345 11103 30379
rect 11529 30345 11563 30379
rect 16221 30345 16255 30379
rect 18705 30345 18739 30379
rect 19717 30345 19751 30379
rect 20637 30345 20671 30379
rect 21005 30345 21039 30379
rect 24317 30345 24351 30379
rect 25237 30345 25271 30379
rect 25329 30345 25363 30379
rect 30481 30345 30515 30379
rect 30849 30345 30883 30379
rect 36277 30345 36311 30379
rect 37841 30345 37875 30379
rect 2881 30277 2915 30311
rect 3617 30277 3651 30311
rect 3801 30277 3835 30311
rect 4353 30277 4387 30311
rect 5758 30277 5792 30311
rect 10149 30277 10183 30311
rect 11897 30277 11931 30311
rect 16405 30277 16439 30311
rect 17325 30277 17359 30311
rect 18153 30277 18187 30311
rect 22753 30277 22787 30311
rect 23581 30277 23615 30311
rect 27261 30277 27295 30311
rect 28825 30277 28859 30311
rect 30113 30277 30147 30311
rect 30313 30277 30347 30311
rect 30941 30277 30975 30311
rect 34069 30277 34103 30311
rect 35336 30277 35370 30311
rect 35541 30277 35575 30311
rect 36645 30277 36679 30311
rect 37657 30277 37691 30311
rect 38301 30277 38335 30311
rect 40601 30277 40635 30311
rect 3157 30209 3191 30243
rect 3433 30209 3467 30243
rect 3541 30209 3575 30243
rect 3985 30209 4019 30243
rect 4169 30209 4203 30243
rect 4261 30209 4295 30243
rect 4445 30209 4479 30243
rect 4537 30209 4571 30243
rect 4721 30209 4755 30243
rect 4813 30209 4847 30243
rect 4905 30209 4939 30243
rect 5641 30209 5675 30243
rect 8125 30209 8159 30243
rect 10425 30209 10459 30243
rect 10885 30209 10919 30243
rect 11069 30209 11103 30243
rect 14841 30209 14875 30243
rect 15025 30209 15059 30243
rect 15209 30209 15243 30243
rect 15301 30209 15335 30243
rect 15945 30209 15979 30243
rect 16129 30209 16163 30243
rect 17509 30209 17543 30243
rect 17693 30209 17727 30243
rect 18245 30209 18279 30243
rect 19073 30209 19107 30243
rect 19349 30209 19383 30243
rect 19533 30209 19567 30243
rect 20269 30209 20303 30243
rect 20913 30209 20947 30243
rect 21097 30209 21131 30243
rect 21465 30209 21499 30243
rect 21649 30209 21683 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 22109 30209 22143 30243
rect 22201 30209 22235 30243
rect 23213 30209 23247 30243
rect 23397 30209 23431 30243
rect 24225 30209 24259 30243
rect 24961 30209 24995 30243
rect 25421 30209 25455 30243
rect 25789 30209 25823 30243
rect 25973 30209 26007 30243
rect 26249 30209 26283 30243
rect 26433 30209 26467 30243
rect 26525 30209 26559 30243
rect 29377 30209 29411 30243
rect 29561 30209 29595 30243
rect 30573 30209 30607 30243
rect 30757 30209 30791 30243
rect 31585 30209 31619 30243
rect 31677 30209 31711 30243
rect 31953 30209 31987 30243
rect 33149 30209 33183 30243
rect 33701 30209 33735 30243
rect 34713 30209 34747 30243
rect 35633 30209 35667 30243
rect 35817 30209 35851 30243
rect 36415 30209 36449 30243
rect 36553 30209 36587 30243
rect 36773 30209 36807 30243
rect 36932 30209 36966 30243
rect 38117 30209 38151 30243
rect 38393 30209 38427 30243
rect 39037 30209 39071 30243
rect 39221 30209 39255 30243
rect 39313 30209 39347 30243
rect 39405 30209 39439 30243
rect 40417 30209 40451 30243
rect 40509 30209 40543 30243
rect 40785 30209 40819 30243
rect 40877 30209 40911 30243
rect 41061 30209 41095 30243
rect 41889 30209 41923 30243
rect 5273 30141 5307 30175
rect 5549 30141 5583 30175
rect 7849 30141 7883 30175
rect 8953 30141 8987 30175
rect 10333 30141 10367 30175
rect 10793 30141 10827 30175
rect 11989 30141 12023 30175
rect 12081 30141 12115 30175
rect 12725 30141 12759 30175
rect 13001 30141 13035 30175
rect 14749 30141 14783 30175
rect 15117 30141 15151 30175
rect 15485 30141 15519 30175
rect 17969 30141 18003 30175
rect 18981 30141 19015 30175
rect 21557 30141 21591 30175
rect 22477 30141 22511 30175
rect 23121 30141 23155 30175
rect 24409 30141 24443 30175
rect 26801 30141 26835 30175
rect 26985 30141 27019 30175
rect 31125 30141 31159 30175
rect 32229 30141 32263 30175
rect 32505 30141 32539 30175
rect 34805 30141 34839 30175
rect 34897 30141 34931 30175
rect 34989 30141 35023 30175
rect 36001 30141 36035 30175
rect 16405 30073 16439 30107
rect 20821 30073 20855 30107
rect 22569 30073 22603 30107
rect 25053 30073 25087 30107
rect 25697 30073 25731 30107
rect 26617 30073 26651 30107
rect 29745 30073 29779 30107
rect 34437 30073 34471 30107
rect 35173 30073 35207 30107
rect 37289 30073 37323 30107
rect 39589 30073 39623 30107
rect 40233 30073 40267 30107
rect 3801 30005 3835 30039
rect 5181 30005 5215 30039
rect 5917 30005 5951 30039
rect 9505 30005 9539 30039
rect 15853 30005 15887 30039
rect 18613 30005 18647 30039
rect 20637 30005 20671 30039
rect 22753 30005 22787 30039
rect 23857 30005 23891 30039
rect 26709 30005 26743 30039
rect 28733 30005 28767 30039
rect 30297 30005 30331 30039
rect 31401 30005 31435 30039
rect 31861 30005 31895 30039
rect 33885 30005 33919 30039
rect 34069 30005 34103 30039
rect 34529 30005 34563 30039
rect 35357 30005 35391 30039
rect 37657 30005 37691 30039
rect 37933 30005 37967 30039
rect 41245 30005 41279 30039
rect 42073 30005 42107 30039
rect 3801 29801 3835 29835
rect 5549 29801 5583 29835
rect 5733 29801 5767 29835
rect 22201 29801 22235 29835
rect 24685 29801 24719 29835
rect 26893 29801 26927 29835
rect 27353 29801 27387 29835
rect 33057 29801 33091 29835
rect 34805 29801 34839 29835
rect 37197 29801 37231 29835
rect 37381 29801 37415 29835
rect 42165 29801 42199 29835
rect 32965 29733 32999 29767
rect 4261 29665 4295 29699
rect 5457 29665 5491 29699
rect 8677 29665 8711 29699
rect 9597 29665 9631 29699
rect 13093 29665 13127 29699
rect 25421 29665 25455 29699
rect 26065 29665 26099 29699
rect 28181 29665 28215 29699
rect 29101 29665 29135 29699
rect 29653 29665 29687 29699
rect 30389 29665 30423 29699
rect 30941 29665 30975 29699
rect 31493 29665 31527 29699
rect 35449 29665 35483 29699
rect 35633 29665 35667 29699
rect 35909 29665 35943 29699
rect 36093 29665 36127 29699
rect 37657 29665 37691 29699
rect 40693 29665 40727 29699
rect 2697 29597 2731 29631
rect 2881 29597 2915 29631
rect 3152 29597 3186 29631
rect 3249 29597 3283 29631
rect 3341 29597 3375 29631
rect 3469 29597 3503 29631
rect 3617 29597 3651 29631
rect 3985 29597 4019 29631
rect 4077 29597 4111 29631
rect 4353 29597 4387 29631
rect 5365 29597 5399 29631
rect 9321 29597 9355 29631
rect 10333 29597 10367 29631
rect 10701 29597 10735 29631
rect 20361 29597 20395 29631
rect 21649 29597 21683 29631
rect 21741 29597 21775 29631
rect 21925 29597 21959 29631
rect 22017 29597 22051 29631
rect 22753 29597 22787 29631
rect 22846 29597 22880 29631
rect 23121 29597 23155 29631
rect 23259 29597 23293 29631
rect 24869 29597 24903 29631
rect 25145 29597 25179 29631
rect 25513 29597 25547 29631
rect 25973 29597 26007 29631
rect 27077 29597 27111 29631
rect 27169 29597 27203 29631
rect 27445 29597 27479 29631
rect 27997 29597 28031 29631
rect 29285 29597 29319 29631
rect 29377 29597 29411 29631
rect 29837 29597 29871 29631
rect 30021 29597 30055 29631
rect 30297 29597 30331 29631
rect 30573 29597 30607 29631
rect 30849 29597 30883 29631
rect 31033 29597 31067 29631
rect 31217 29597 31251 29631
rect 33236 29597 33270 29631
rect 33608 29597 33642 29631
rect 33701 29597 33735 29631
rect 35081 29597 35115 29631
rect 35357 29597 35391 29631
rect 36185 29597 36219 29631
rect 37841 29597 37875 29631
rect 37933 29597 37967 29631
rect 38209 29597 38243 29631
rect 38393 29597 38427 29631
rect 38485 29597 38519 29631
rect 38577 29597 38611 29631
rect 40417 29597 40451 29631
rect 2789 29529 2823 29563
rect 8401 29529 8435 29563
rect 12725 29529 12759 29563
rect 12909 29529 12943 29563
rect 20821 29529 20855 29563
rect 21005 29529 21039 29563
rect 23029 29529 23063 29563
rect 25053 29529 25087 29563
rect 33333 29529 33367 29563
rect 33425 29529 33459 29563
rect 34805 29529 34839 29563
rect 34989 29529 35023 29563
rect 37565 29529 37599 29563
rect 39865 29529 39899 29563
rect 40049 29529 40083 29563
rect 2973 29461 3007 29495
rect 8033 29461 8067 29495
rect 8493 29461 8527 29495
rect 8953 29461 8987 29495
rect 9413 29461 9447 29495
rect 9781 29461 9815 29495
rect 10609 29461 10643 29495
rect 20545 29461 20579 29495
rect 23397 29461 23431 29495
rect 25881 29461 25915 29495
rect 27537 29461 27571 29495
rect 27905 29461 27939 29495
rect 29101 29461 29135 29495
rect 30757 29461 30791 29495
rect 35633 29461 35667 29495
rect 36553 29461 36587 29495
rect 37355 29461 37389 29495
rect 37657 29461 37691 29495
rect 38761 29461 38795 29495
rect 40233 29461 40267 29495
rect 5457 29257 5491 29291
rect 9781 29257 9815 29291
rect 10701 29257 10735 29291
rect 10977 29257 11011 29291
rect 12633 29257 12667 29291
rect 14289 29257 14323 29291
rect 15025 29257 15059 29291
rect 15485 29257 15519 29291
rect 16037 29257 16071 29291
rect 16957 29257 16991 29291
rect 18245 29257 18279 29291
rect 18797 29257 18831 29291
rect 27997 29257 28031 29291
rect 32689 29257 32723 29291
rect 32781 29257 32815 29291
rect 34897 29257 34931 29291
rect 38117 29257 38151 29291
rect 39589 29257 39623 29291
rect 7196 29189 7230 29223
rect 16129 29189 16163 29223
rect 17877 29189 17911 29223
rect 22109 29189 22143 29223
rect 22201 29189 22235 29223
rect 22845 29189 22879 29223
rect 23581 29189 23615 29223
rect 27721 29189 27755 29223
rect 31217 29189 31251 29223
rect 31309 29189 31343 29223
rect 33425 29189 33459 29223
rect 33517 29189 33551 29223
rect 37933 29189 37967 29223
rect 39221 29189 39255 29223
rect 39313 29189 39347 29223
rect 39957 29189 39991 29223
rect 1409 29121 1443 29155
rect 3433 29121 3467 29155
rect 4077 29121 4111 29155
rect 4261 29121 4295 29155
rect 5457 29121 5491 29155
rect 5641 29121 5675 29155
rect 6929 29121 6963 29155
rect 8401 29121 8435 29155
rect 8668 29121 8702 29155
rect 9873 29121 9907 29155
rect 10057 29121 10091 29155
rect 10241 29121 10275 29155
rect 10701 29121 10735 29155
rect 10885 29121 10919 29155
rect 10977 29121 11011 29155
rect 11161 29121 11195 29155
rect 12817 29121 12851 29155
rect 13093 29121 13127 29155
rect 13277 29121 13311 29155
rect 13369 29121 13403 29155
rect 13829 29121 13863 29155
rect 14933 29121 14967 29155
rect 15209 29121 15243 29155
rect 16681 29121 16715 29155
rect 16957 29121 16991 29155
rect 17141 29121 17175 29155
rect 17325 29121 17359 29155
rect 17601 29121 17635 29155
rect 17759 29121 17793 29155
rect 17969 29121 18003 29155
rect 18061 29121 18095 29155
rect 18613 29121 18647 29155
rect 20269 29121 20303 29155
rect 20453 29121 20487 29155
rect 21925 29121 21959 29155
rect 22293 29121 22327 29155
rect 24041 29121 24075 29155
rect 25789 29121 25823 29155
rect 25973 29121 26007 29155
rect 27445 29121 27479 29155
rect 27629 29121 27663 29155
rect 27813 29121 27847 29155
rect 29469 29121 29503 29155
rect 29653 29121 29687 29155
rect 30481 29121 30515 29155
rect 30573 29121 30607 29155
rect 30849 29121 30883 29155
rect 31079 29121 31113 29155
rect 31492 29121 31526 29155
rect 31585 29121 31619 29155
rect 33241 29121 33275 29155
rect 33609 29121 33643 29155
rect 34069 29121 34103 29155
rect 34161 29121 34195 29155
rect 34437 29121 34471 29155
rect 35081 29121 35115 29155
rect 35173 29121 35207 29155
rect 35357 29121 35391 29155
rect 35541 29121 35575 29155
rect 37289 29121 37323 29155
rect 37565 29121 37599 29155
rect 37657 29121 37691 29155
rect 38209 29121 38243 29155
rect 39037 29121 39071 29155
rect 39405 29121 39439 29155
rect 41889 29121 41923 29155
rect 1685 29053 1719 29087
rect 3157 29053 3191 29087
rect 3525 29053 3559 29087
rect 3617 29053 3651 29087
rect 3709 29053 3743 29087
rect 3893 29053 3927 29087
rect 4353 29053 4387 29087
rect 15301 29053 15335 29087
rect 15577 29053 15611 29087
rect 15669 29053 15703 29087
rect 18337 29053 18371 29087
rect 23765 29053 23799 29087
rect 32597 29053 32631 29087
rect 34897 29053 34931 29087
rect 39681 29053 39715 29087
rect 41429 29053 41463 29087
rect 8309 28985 8343 29019
rect 10149 28985 10183 29019
rect 13507 28985 13541 29019
rect 20453 28985 20487 29019
rect 22477 28985 22511 29019
rect 30297 28985 30331 29019
rect 30757 28985 30791 29019
rect 30941 28985 30975 29019
rect 33149 28985 33183 29019
rect 33885 28985 33919 29019
rect 35541 28985 35575 29019
rect 37381 28985 37415 29019
rect 37933 28985 37967 29019
rect 42073 28985 42107 29019
rect 3249 28917 3283 28951
rect 10333 28917 10367 28951
rect 10609 28917 10643 28951
rect 13645 28917 13679 28951
rect 13737 28917 13771 28951
rect 18429 28917 18463 28951
rect 25789 28917 25823 28951
rect 29469 28917 29503 28951
rect 33793 28917 33827 28951
rect 34345 28917 34379 28951
rect 37841 28917 37875 28951
rect 2605 28713 2639 28747
rect 2973 28713 3007 28747
rect 4629 28713 4663 28747
rect 6929 28713 6963 28747
rect 9137 28713 9171 28747
rect 12449 28713 12483 28747
rect 17325 28713 17359 28747
rect 21005 28713 21039 28747
rect 25605 28713 25639 28747
rect 30021 28713 30055 28747
rect 32505 28713 32539 28747
rect 34529 28713 34563 28747
rect 36645 28713 36679 28747
rect 4721 28645 4755 28679
rect 8769 28645 8803 28679
rect 12081 28645 12115 28679
rect 15853 28645 15887 28679
rect 16405 28645 16439 28679
rect 16773 28645 16807 28679
rect 16911 28645 16945 28679
rect 18797 28645 18831 28679
rect 29377 28645 29411 28679
rect 36093 28645 36127 28679
rect 5181 28577 5215 28611
rect 9689 28577 9723 28611
rect 14381 28577 14415 28611
rect 16681 28577 16715 28611
rect 18061 28577 18095 28611
rect 19257 28577 19291 28611
rect 24133 28577 24167 28611
rect 27629 28577 27663 28611
rect 27905 28577 27939 28611
rect 29561 28577 29595 28611
rect 32781 28577 32815 28611
rect 37381 28577 37415 28611
rect 37657 28577 37691 28611
rect 2789 28509 2823 28543
rect 3065 28509 3099 28543
rect 4077 28509 4111 28543
rect 4445 28509 4479 28543
rect 4721 28509 4755 28543
rect 4905 28509 4939 28543
rect 7389 28509 7423 28543
rect 9505 28509 9539 28543
rect 9965 28509 9999 28543
rect 10149 28509 10183 28543
rect 10977 28509 11011 28543
rect 11161 28509 11195 28543
rect 11621 28509 11655 28543
rect 11713 28509 11747 28543
rect 11805 28509 11839 28543
rect 11989 28509 12023 28543
rect 12265 28509 12299 28543
rect 12449 28509 12483 28543
rect 12725 28509 12759 28543
rect 12817 28509 12851 28543
rect 14105 28509 14139 28543
rect 16221 28509 16255 28543
rect 17141 28509 17175 28543
rect 17417 28509 17451 28543
rect 17785 28509 17819 28543
rect 18245 28509 18279 28543
rect 18521 28509 18555 28543
rect 18797 28509 18831 28543
rect 21189 28509 21223 28543
rect 21787 28509 21821 28543
rect 21925 28509 21959 28543
rect 22017 28509 22051 28543
rect 22200 28509 22234 28543
rect 22293 28509 22327 28543
rect 24409 28509 24443 28543
rect 25329 28509 25363 28543
rect 25421 28509 25455 28543
rect 25697 28509 25731 28543
rect 25968 28509 26002 28543
rect 26065 28509 26099 28543
rect 26340 28509 26374 28543
rect 26433 28509 26467 28543
rect 29745 28509 29779 28543
rect 29837 28509 29871 28543
rect 30113 28509 30147 28543
rect 31125 28509 31159 28543
rect 31309 28509 31343 28543
rect 32045 28509 32079 28543
rect 34989 28509 35023 28543
rect 35357 28509 35391 28543
rect 35449 28509 35483 28543
rect 35597 28509 35631 28543
rect 35725 28509 35759 28543
rect 35817 28509 35851 28543
rect 35955 28509 35989 28543
rect 36369 28509 36403 28543
rect 36461 28509 36495 28543
rect 36737 28509 36771 28543
rect 41521 28509 41555 28543
rect 41889 28509 41923 28543
rect 4261 28441 4295 28475
rect 4353 28441 4387 28475
rect 5457 28441 5491 28475
rect 7656 28441 7690 28475
rect 13093 28441 13127 28475
rect 13185 28441 13219 28475
rect 13645 28441 13679 28475
rect 17049 28441 17083 28475
rect 19533 28441 19567 28475
rect 21557 28441 21591 28475
rect 23857 28441 23891 28475
rect 26157 28441 26191 28475
rect 32413 28441 32447 28475
rect 33057 28441 33091 28475
rect 35081 28441 35115 28475
rect 35173 28441 35207 28475
rect 40325 28441 40359 28475
rect 40509 28441 40543 28475
rect 9597 28373 9631 28407
rect 10057 28373 10091 28407
rect 11069 28373 11103 28407
rect 11345 28373 11379 28407
rect 12541 28373 12575 28407
rect 13553 28373 13587 28407
rect 16129 28373 16163 28407
rect 17601 28373 17635 28407
rect 18429 28373 18463 28407
rect 21649 28373 21683 28407
rect 22385 28373 22419 28407
rect 25145 28373 25179 28407
rect 25789 28373 25823 28407
rect 34805 28373 34839 28407
rect 36185 28373 36219 28407
rect 39129 28373 39163 28407
rect 40693 28373 40727 28407
rect 41705 28373 41739 28407
rect 42073 28373 42107 28407
rect 5549 28169 5583 28203
rect 8493 28169 8527 28203
rect 8677 28169 8711 28203
rect 9413 28169 9447 28203
rect 11897 28169 11931 28203
rect 12817 28169 12851 28203
rect 13553 28169 13587 28203
rect 15301 28169 15335 28203
rect 16681 28169 16715 28203
rect 18429 28169 18463 28203
rect 19441 28169 19475 28203
rect 23581 28169 23615 28203
rect 24777 28169 24811 28203
rect 26709 28169 26743 28203
rect 29561 28169 29595 28203
rect 37933 28169 37967 28203
rect 40325 28169 40359 28203
rect 42165 28169 42199 28203
rect 13093 28101 13127 28135
rect 14933 28101 14967 28135
rect 15117 28101 15151 28135
rect 15669 28101 15703 28135
rect 16865 28101 16899 28135
rect 17325 28101 17359 28135
rect 19349 28101 19383 28135
rect 24409 28101 24443 28135
rect 24593 28101 24627 28135
rect 25237 28101 25271 28135
rect 27721 28101 27755 28135
rect 29193 28101 29227 28135
rect 29285 28101 29319 28135
rect 29745 28101 29779 28135
rect 29929 28101 29963 28135
rect 32505 28101 32539 28135
rect 33701 28101 33735 28135
rect 35541 28101 35575 28135
rect 37657 28101 37691 28135
rect 40049 28101 40083 28135
rect 40693 28101 40727 28135
rect 4445 28033 4479 28067
rect 4629 28033 4663 28067
rect 6009 28033 6043 28067
rect 6469 28033 6503 28067
rect 6561 28033 6595 28067
rect 9321 28033 9355 28067
rect 11989 28033 12023 28067
rect 12081 28033 12115 28067
rect 12559 28033 12593 28067
rect 12996 28033 13030 28067
rect 13185 28033 13219 28067
rect 13368 28033 13402 28067
rect 13461 28033 13495 28067
rect 13737 28033 13771 28067
rect 13829 28033 13863 28067
rect 14013 28033 14047 28067
rect 14289 28033 14323 28067
rect 14473 28033 14507 28067
rect 14657 28033 14691 28067
rect 14749 28033 14783 28067
rect 15209 28033 15243 28067
rect 15485 28033 15519 28067
rect 16313 28033 16347 28067
rect 17049 28033 17083 28067
rect 17233 28033 17267 28067
rect 17417 28033 17451 28067
rect 17509 28033 17543 28067
rect 17693 28033 17727 28067
rect 17785 28033 17819 28067
rect 17969 28033 18003 28067
rect 18061 28033 18095 28067
rect 18153 28033 18187 28067
rect 18613 28033 18647 28067
rect 19073 28033 19107 28067
rect 19165 28033 19199 28067
rect 19625 28033 19659 28067
rect 19717 28033 19751 28067
rect 20361 28033 20395 28067
rect 21005 28033 21039 28067
rect 24133 28033 24167 28067
rect 24317 28033 24351 28067
rect 24961 28033 24995 28067
rect 27629 28033 27663 28067
rect 27813 28033 27847 28067
rect 27997 28033 28031 28067
rect 28917 28033 28951 28067
rect 29065 28033 29099 28067
rect 29423 28033 29457 28067
rect 32781 28033 32815 28067
rect 32965 28033 32999 28067
rect 33057 28033 33091 28067
rect 33149 28033 33183 28067
rect 33425 28033 33459 28067
rect 33518 28033 33552 28067
rect 33793 28033 33827 28067
rect 33931 28033 33965 28067
rect 34345 28033 34379 28067
rect 35265 28033 35299 28067
rect 37289 28033 37323 28067
rect 37437 28033 37471 28067
rect 37565 28033 37599 28067
rect 37773 28033 37807 28067
rect 38945 28033 38979 28067
rect 39773 28033 39807 28067
rect 39957 28033 39991 28067
rect 40141 28033 40175 28067
rect 4905 27965 4939 27999
rect 5273 27965 5307 27999
rect 5365 27965 5399 27999
rect 5917 27965 5951 27999
rect 8033 27965 8067 27999
rect 9873 27965 9907 27999
rect 12357 27965 12391 27999
rect 16037 27965 16071 27999
rect 17601 27965 17635 27999
rect 18705 27965 18739 27999
rect 19809 27965 19843 27999
rect 19901 27965 19935 27999
rect 21833 27965 21867 27999
rect 22109 27965 22143 27999
rect 30205 27965 30239 27999
rect 30481 27965 30515 27999
rect 34621 27965 34655 27999
rect 40417 27965 40451 27999
rect 5641 27897 5675 27931
rect 8401 27897 8435 27931
rect 9597 27897 9631 27931
rect 12725 27897 12759 27931
rect 24317 27897 24351 27931
rect 32229 27897 32263 27931
rect 34069 27897 34103 27931
rect 4537 27829 4571 27863
rect 4813 27829 4847 27863
rect 12541 27829 12575 27863
rect 14013 27829 14047 27863
rect 14197 27829 14231 27863
rect 14657 27829 14691 27863
rect 15761 27829 15795 27863
rect 15945 27829 15979 27863
rect 17785 27829 17819 27863
rect 18061 27829 18095 27863
rect 27445 27829 27479 27863
rect 31953 27829 31987 27863
rect 33333 27829 33367 27863
rect 37013 27829 37047 27863
rect 39037 27829 39071 27863
rect 4077 27625 4111 27659
rect 4813 27625 4847 27659
rect 22293 27625 22327 27659
rect 5181 27557 5215 27591
rect 13277 27557 13311 27591
rect 15669 27557 15703 27591
rect 16129 27557 16163 27591
rect 17233 27557 17267 27591
rect 21833 27557 21867 27591
rect 22937 27557 22971 27591
rect 28917 27557 28951 27591
rect 32689 27557 32723 27591
rect 5089 27489 5123 27523
rect 12265 27489 12299 27523
rect 25881 27489 25915 27523
rect 26065 27489 26099 27523
rect 30205 27489 30239 27523
rect 30297 27489 30331 27523
rect 31861 27489 31895 27523
rect 34437 27489 34471 27523
rect 38853 27489 38887 27523
rect 3893 27421 3927 27455
rect 4077 27421 4111 27455
rect 4997 27421 5031 27455
rect 5273 27421 5307 27455
rect 9965 27421 9999 27455
rect 13001 27421 13035 27455
rect 13185 27421 13219 27455
rect 13369 27421 13403 27455
rect 15393 27421 15427 27455
rect 15577 27421 15611 27455
rect 16037 27421 16071 27455
rect 16129 27421 16163 27455
rect 16405 27421 16439 27455
rect 17049 27421 17083 27455
rect 17233 27421 17267 27455
rect 17601 27421 17635 27455
rect 18245 27421 18279 27455
rect 18337 27421 18371 27455
rect 21373 27421 21407 27455
rect 21741 27421 21775 27455
rect 22017 27421 22051 27455
rect 22109 27421 22143 27455
rect 22385 27421 22419 27455
rect 22569 27421 22603 27455
rect 22845 27421 22879 27455
rect 23121 27421 23155 27455
rect 23305 27421 23339 27455
rect 24409 27421 24443 27455
rect 24593 27421 24627 27455
rect 26893 27421 26927 27455
rect 27169 27421 27203 27455
rect 30113 27421 30147 27455
rect 32137 27421 32171 27455
rect 32505 27421 32539 27455
rect 34161 27421 34195 27455
rect 34253 27421 34287 27455
rect 34713 27421 34747 27455
rect 34806 27421 34840 27455
rect 35081 27421 35115 27455
rect 35178 27421 35212 27455
rect 35725 27421 35759 27455
rect 35817 27421 35851 27455
rect 35965 27421 35999 27455
rect 36185 27421 36219 27455
rect 36282 27421 36316 27455
rect 40141 27421 40175 27455
rect 40417 27421 40451 27455
rect 40509 27421 40543 27455
rect 40785 27421 40819 27455
rect 41337 27421 41371 27455
rect 41705 27421 41739 27455
rect 10232 27353 10266 27387
rect 11437 27353 11471 27387
rect 15853 27353 15887 27387
rect 16313 27353 16347 27387
rect 17325 27353 17359 27387
rect 17509 27353 17543 27387
rect 17785 27353 17819 27387
rect 17877 27353 17911 27387
rect 18429 27353 18463 27387
rect 20913 27353 20947 27387
rect 21189 27353 21223 27387
rect 24501 27353 24535 27387
rect 26709 27353 26743 27387
rect 27077 27353 27111 27387
rect 27445 27353 27479 27387
rect 32321 27353 32355 27387
rect 32413 27353 32447 27387
rect 34989 27353 35023 27387
rect 36093 27353 36127 27387
rect 39055 27353 39089 27387
rect 39221 27353 39255 27387
rect 40325 27353 40359 27387
rect 40969 27353 41003 27387
rect 11345 27285 11379 27319
rect 12449 27285 12483 27319
rect 15485 27285 15519 27319
rect 17417 27285 17451 27319
rect 20637 27285 20671 27319
rect 22753 27285 22787 27319
rect 26157 27285 26191 27319
rect 26525 27285 26559 27319
rect 29745 27285 29779 27319
rect 31309 27285 31343 27319
rect 31677 27285 31711 27319
rect 31769 27285 31803 27319
rect 33793 27285 33827 27319
rect 35357 27285 35391 27319
rect 35541 27285 35575 27319
rect 36461 27285 36495 27319
rect 38209 27285 38243 27319
rect 38577 27285 38611 27319
rect 38669 27285 38703 27319
rect 39405 27285 39439 27319
rect 40693 27285 40727 27319
rect 41153 27285 41187 27319
rect 41521 27285 41555 27319
rect 41889 27285 41923 27319
rect 3065 27081 3099 27115
rect 3617 27081 3651 27115
rect 10149 27081 10183 27115
rect 10425 27081 10459 27115
rect 12909 27081 12943 27115
rect 14381 27081 14415 27115
rect 25789 27081 25823 27115
rect 26985 27081 27019 27115
rect 38117 27081 38151 27115
rect 38577 27081 38611 27115
rect 2881 27013 2915 27047
rect 3249 27013 3283 27047
rect 7205 27013 7239 27047
rect 10885 27013 10919 27047
rect 13553 27013 13587 27047
rect 13921 27013 13955 27047
rect 14749 27013 14783 27047
rect 16497 27013 16531 27047
rect 17969 27013 18003 27047
rect 18153 27013 18187 27047
rect 21373 27013 21407 27047
rect 21557 27013 21591 27047
rect 29837 27013 29871 27047
rect 38209 27013 38243 27047
rect 39129 27013 39163 27047
rect 1685 26945 1719 26979
rect 3433 26945 3467 26979
rect 3985 26945 4019 26979
rect 4077 26945 4111 26979
rect 4261 26945 4295 26979
rect 4353 26945 4387 26979
rect 4721 26945 4755 26979
rect 4997 26945 5031 26979
rect 5181 26945 5215 26979
rect 9229 26945 9263 26979
rect 10057 26945 10091 26979
rect 10241 26945 10275 26979
rect 10793 26945 10827 26979
rect 11805 26945 11839 26979
rect 12541 26945 12575 26979
rect 12695 26945 12729 26979
rect 13093 26945 13127 26979
rect 13369 26945 13403 26979
rect 13829 26945 13863 26979
rect 14197 26945 14231 26979
rect 18705 26945 18739 26979
rect 27169 26945 27203 26979
rect 27261 26945 27295 26979
rect 27353 26945 27387 26979
rect 27537 26945 27571 26979
rect 29561 26945 29595 26979
rect 29745 26945 29779 26979
rect 29929 26945 29963 26979
rect 41245 26945 41279 26979
rect 4905 26877 4939 26911
rect 8953 26877 8987 26911
rect 9873 26877 9907 26911
rect 10977 26877 11011 26911
rect 11529 26877 11563 26911
rect 13001 26877 13035 26911
rect 14013 26877 14047 26911
rect 14473 26877 14507 26911
rect 19533 26877 19567 26911
rect 21005 26877 21039 26911
rect 21281 26877 21315 26911
rect 24041 26877 24075 26911
rect 24317 26877 24351 26911
rect 26525 26877 26559 26911
rect 38025 26877 38059 26911
rect 38853 26877 38887 26911
rect 42165 26877 42199 26911
rect 2513 26809 2547 26843
rect 13737 26809 13771 26843
rect 18337 26809 18371 26843
rect 40601 26809 40635 26843
rect 41429 26809 41463 26843
rect 1501 26741 1535 26775
rect 2881 26741 2915 26775
rect 3801 26741 3835 26775
rect 4537 26741 4571 26775
rect 5089 26741 5123 26775
rect 9321 26741 9355 26775
rect 11621 26741 11655 26775
rect 11713 26741 11747 26775
rect 13829 26741 13863 26775
rect 13921 26741 13955 26775
rect 18889 26741 18923 26775
rect 25973 26741 26007 26775
rect 30113 26741 30147 26775
rect 41521 26741 41555 26775
rect 4905 26537 4939 26571
rect 8585 26537 8619 26571
rect 10333 26537 10367 26571
rect 13001 26537 13035 26571
rect 13737 26537 13771 26571
rect 14841 26537 14875 26571
rect 19257 26537 19291 26571
rect 19625 26537 19659 26571
rect 20821 26537 20855 26571
rect 24593 26537 24627 26571
rect 36369 26537 36403 26571
rect 38485 26537 38519 26571
rect 12725 26469 12759 26503
rect 17877 26469 17911 26503
rect 18337 26469 18371 26503
rect 18705 26469 18739 26503
rect 22845 26469 22879 26503
rect 24869 26469 24903 26503
rect 25513 26469 25547 26503
rect 2973 26401 3007 26435
rect 7205 26401 7239 26435
rect 7849 26401 7883 26435
rect 10977 26401 11011 26435
rect 11253 26401 11287 26435
rect 12909 26401 12943 26435
rect 13737 26401 13771 26435
rect 15117 26401 15151 26435
rect 15209 26401 15243 26435
rect 15577 26401 15611 26435
rect 18981 26401 19015 26435
rect 19349 26401 19383 26435
rect 20269 26401 20303 26435
rect 21097 26401 21131 26435
rect 25053 26401 25087 26435
rect 33517 26401 33551 26435
rect 35633 26401 35667 26435
rect 35817 26401 35851 26435
rect 3249 26333 3283 26367
rect 3893 26333 3927 26367
rect 4629 26333 4663 26367
rect 4997 26333 5031 26367
rect 5089 26333 5123 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 5457 26333 5491 26367
rect 8033 26333 8067 26367
rect 8309 26333 8343 26367
rect 8401 26333 8435 26367
rect 8953 26333 8987 26367
rect 13185 26333 13219 26367
rect 13829 26333 13863 26367
rect 14565 26333 14599 26367
rect 14657 26333 14691 26367
rect 15485 26333 15519 26367
rect 17601 26333 17635 26367
rect 17693 26333 17727 26367
rect 17969 26333 18003 26367
rect 18061 26333 18095 26367
rect 19257 26333 19291 26367
rect 23121 26333 23155 26367
rect 23305 26333 23339 26367
rect 24777 26333 24811 26367
rect 24961 26333 24995 26367
rect 25237 26333 25271 26367
rect 25697 26333 25731 26367
rect 25881 26333 25915 26367
rect 29745 26333 29779 26367
rect 33333 26333 33367 26367
rect 35357 26333 35391 26367
rect 35541 26333 35575 26367
rect 37933 26333 37967 26367
rect 38301 26333 38335 26367
rect 38761 26333 38795 26367
rect 39865 26333 39899 26367
rect 5733 26265 5767 26299
rect 8217 26265 8251 26299
rect 9198 26265 9232 26299
rect 13369 26265 13403 26299
rect 18153 26265 18187 26299
rect 18337 26265 18371 26299
rect 20361 26265 20395 26299
rect 21373 26265 21407 26299
rect 23213 26265 23247 26299
rect 29653 26265 29687 26299
rect 35817 26265 35851 26299
rect 36553 26265 36587 26299
rect 38117 26265 38151 26299
rect 38209 26265 38243 26299
rect 39589 26265 39623 26299
rect 1501 26197 1535 26231
rect 7297 26197 7331 26231
rect 13461 26197 13495 26231
rect 14933 26197 14967 26231
rect 15393 26197 15427 26231
rect 17417 26197 17451 26231
rect 18521 26197 18555 26231
rect 20453 26197 20487 26231
rect 32965 26197 32999 26231
rect 33425 26197 33459 26231
rect 36185 26197 36219 26231
rect 36353 26197 36387 26231
rect 3617 25993 3651 26027
rect 6377 25993 6411 26027
rect 7113 25993 7147 26027
rect 8217 25993 8251 26027
rect 14933 25993 14967 26027
rect 20729 25993 20763 26027
rect 21833 25993 21867 26027
rect 22201 25993 22235 26027
rect 25145 25993 25179 26027
rect 27169 25993 27203 26027
rect 31585 25993 31619 26027
rect 38669 25993 38703 26027
rect 42165 25993 42199 26027
rect 3249 25925 3283 25959
rect 4997 25925 5031 25959
rect 7941 25925 7975 25959
rect 8585 25925 8619 25959
rect 8953 25925 8987 25959
rect 13461 25925 13495 25959
rect 17417 25925 17451 25959
rect 20453 25925 20487 25959
rect 25789 25925 25823 25959
rect 32689 25925 32723 25959
rect 37013 25925 37047 25959
rect 37565 25925 37599 25959
rect 37657 25925 37691 25959
rect 38945 25925 38979 25959
rect 2053 25857 2087 25891
rect 2207 25857 2241 25891
rect 2605 25857 2639 25891
rect 2789 25857 2823 25891
rect 2881 25857 2915 25891
rect 3341 25857 3375 25891
rect 3525 25857 3559 25891
rect 4537 25857 4571 25891
rect 4859 25857 4893 25891
rect 5089 25857 5123 25891
rect 5272 25857 5306 25891
rect 5365 25857 5399 25891
rect 6561 25857 6595 25891
rect 6837 25857 6871 25891
rect 7021 25857 7055 25891
rect 7665 25857 7699 25891
rect 7849 25857 7883 25891
rect 8033 25857 8067 25891
rect 8309 25857 8343 25891
rect 8493 25857 8527 25891
rect 8677 25857 8711 25891
rect 9597 25857 9631 25891
rect 9689 25857 9723 25891
rect 9945 25857 9979 25891
rect 20177 25857 20211 25891
rect 20361 25857 20395 25891
rect 20545 25857 20579 25891
rect 23949 25857 23983 25891
rect 24409 25857 24443 25891
rect 24777 25857 24811 25891
rect 24869 25857 24903 25891
rect 25053 25857 25087 25891
rect 25389 25857 25423 25891
rect 25513 25857 25547 25891
rect 25697 25857 25731 25891
rect 25881 25857 25915 25891
rect 25973 25857 26007 25891
rect 26066 25857 26100 25891
rect 26249 25857 26283 25891
rect 26341 25857 26375 25891
rect 26438 25857 26472 25891
rect 26985 25857 27019 25891
rect 28733 25857 28767 25891
rect 28825 25857 28859 25891
rect 28917 25857 28951 25891
rect 29055 25857 29089 25891
rect 29469 25857 29503 25891
rect 30173 25857 30207 25891
rect 30389 25857 30423 25891
rect 31677 25857 31711 25891
rect 32137 25857 32171 25891
rect 32413 25857 32447 25891
rect 34345 25857 34379 25891
rect 36645 25857 36679 25891
rect 36921 25857 36955 25891
rect 37473 25857 37507 25891
rect 37775 25857 37809 25891
rect 38853 25857 38887 25891
rect 39037 25857 39071 25891
rect 39221 25857 39255 25891
rect 40325 25857 40359 25891
rect 2421 25789 2455 25823
rect 6745 25789 6779 25823
rect 13185 25789 13219 25823
rect 17141 25789 17175 25823
rect 19165 25789 19199 25823
rect 22293 25789 22327 25823
rect 22477 25789 22511 25823
rect 23857 25789 23891 25823
rect 25605 25789 25639 25823
rect 29193 25789 29227 25823
rect 29561 25789 29595 25823
rect 31769 25789 31803 25823
rect 34161 25789 34195 25823
rect 34621 25789 34655 25823
rect 36369 25789 36403 25823
rect 37933 25789 37967 25823
rect 40417 25789 40451 25823
rect 40693 25789 40727 25823
rect 25053 25721 25087 25755
rect 29837 25721 29871 25755
rect 4721 25653 4755 25687
rect 8861 25653 8895 25687
rect 11069 25653 11103 25687
rect 23581 25653 23615 25687
rect 23857 25653 23891 25687
rect 24225 25653 24259 25687
rect 26617 25653 26651 25687
rect 28549 25653 28583 25687
rect 29929 25653 29963 25687
rect 30297 25653 30331 25687
rect 31217 25653 31251 25687
rect 32321 25653 32355 25687
rect 36093 25653 36127 25687
rect 36461 25653 36495 25687
rect 36829 25653 36863 25687
rect 37289 25653 37323 25687
rect 40141 25653 40175 25687
rect 7573 25449 7607 25483
rect 10333 25449 10367 25483
rect 17877 25449 17911 25483
rect 20269 25449 20303 25483
rect 21557 25449 21591 25483
rect 23213 25449 23247 25483
rect 25329 25449 25363 25483
rect 25973 25449 26007 25483
rect 28917 25449 28951 25483
rect 30389 25449 30423 25483
rect 32597 25449 32631 25483
rect 33609 25449 33643 25483
rect 39497 25449 39531 25483
rect 42165 25449 42199 25483
rect 17785 25381 17819 25415
rect 23397 25381 23431 25415
rect 3801 25313 3835 25347
rect 6193 25313 6227 25347
rect 12265 25313 12299 25347
rect 15393 25313 15427 25347
rect 16405 25313 16439 25347
rect 17049 25313 17083 25347
rect 17233 25313 17267 25347
rect 18337 25313 18371 25347
rect 23581 25313 23615 25347
rect 24593 25313 24627 25347
rect 28549 25313 28583 25347
rect 28733 25313 28767 25347
rect 30849 25313 30883 25347
rect 32689 25313 32723 25347
rect 34805 25313 34839 25347
rect 35909 25313 35943 25347
rect 36369 25313 36403 25347
rect 37013 25313 37047 25347
rect 37197 25313 37231 25347
rect 38025 25313 38059 25347
rect 3157 25245 3191 25279
rect 3249 25245 3283 25279
rect 3341 25245 3375 25279
rect 3525 25245 3559 25279
rect 8953 25245 8987 25279
rect 15117 25245 15151 25279
rect 15209 25245 15243 25279
rect 15485 25245 15519 25279
rect 16221 25245 16255 25279
rect 16589 25245 16623 25279
rect 16891 25245 16925 25279
rect 17141 25245 17175 25279
rect 17325 25245 17359 25279
rect 17417 25245 17451 25279
rect 17601 25245 17635 25279
rect 18061 25245 18095 25279
rect 18153 25245 18187 25279
rect 18429 25245 18463 25279
rect 20269 25245 20303 25279
rect 20453 25245 20487 25279
rect 21741 25245 21775 25279
rect 21925 25245 21959 25279
rect 22201 25245 22235 25279
rect 22477 25245 22511 25279
rect 22845 25245 22879 25279
rect 23029 25245 23063 25279
rect 23305 25245 23339 25279
rect 23673 25245 23707 25279
rect 23949 25245 23983 25279
rect 24041 25245 24075 25279
rect 24685 25245 24719 25279
rect 25053 25245 25087 25279
rect 25513 25245 25547 25279
rect 25789 25245 25823 25279
rect 26157 25245 26191 25279
rect 29745 25245 29779 25279
rect 29838 25245 29872 25279
rect 30021 25245 30055 25279
rect 30210 25245 30244 25279
rect 30757 25245 30791 25279
rect 32965 25245 32999 25279
rect 33793 25245 33827 25279
rect 33885 25245 33919 25279
rect 34253 25245 34287 25279
rect 35633 25245 35667 25279
rect 36001 25245 36035 25279
rect 37749 25245 37783 25279
rect 40417 25245 40451 25279
rect 4077 25177 4111 25211
rect 6460 25177 6494 25211
rect 9198 25177 9232 25211
rect 11989 25177 12023 25211
rect 15669 25177 15703 25211
rect 16681 25177 16715 25211
rect 16773 25177 16807 25211
rect 21833 25177 21867 25211
rect 22063 25177 22097 25211
rect 23581 25177 23615 25211
rect 23857 25177 23891 25211
rect 24961 25177 24995 25211
rect 25605 25177 25639 25211
rect 26433 25177 26467 25211
rect 28457 25177 28491 25211
rect 29101 25177 29135 25211
rect 29285 25177 29319 25211
rect 30113 25177 30147 25211
rect 31125 25177 31159 25211
rect 34161 25177 34195 25211
rect 36277 25177 36311 25211
rect 40693 25177 40727 25211
rect 2881 25109 2915 25143
rect 5549 25109 5583 25143
rect 11621 25109 11655 25143
rect 12081 25109 12115 25143
rect 14933 25109 14967 25143
rect 22385 25109 22419 25143
rect 24225 25109 24259 25143
rect 24869 25109 24903 25143
rect 27905 25109 27939 25143
rect 28089 25109 28123 25143
rect 30573 25109 30607 25143
rect 35725 25109 35759 25143
rect 37289 25109 37323 25143
rect 37657 25109 37691 25143
rect 3157 24905 3191 24939
rect 3525 24905 3559 24939
rect 6377 24905 6411 24939
rect 7665 24905 7699 24939
rect 16037 24905 16071 24939
rect 16681 24905 16715 24939
rect 18337 24905 18371 24939
rect 19625 24905 19659 24939
rect 20453 24905 20487 24939
rect 21649 24905 21683 24939
rect 22477 24905 22511 24939
rect 26985 24905 27019 24939
rect 33885 24905 33919 24939
rect 34805 24905 34839 24939
rect 35173 24905 35207 24939
rect 35265 24905 35299 24939
rect 35725 24905 35759 24939
rect 40877 24905 40911 24939
rect 41245 24905 41279 24939
rect 7941 24837 7975 24871
rect 11805 24837 11839 24871
rect 14565 24837 14599 24871
rect 16865 24837 16899 24871
rect 21005 24837 21039 24871
rect 27813 24837 27847 24871
rect 29745 24837 29779 24871
rect 32623 24837 32657 24871
rect 37933 24837 37967 24871
rect 3341 24769 3375 24803
rect 3893 24769 3927 24803
rect 4537 24769 4571 24803
rect 4905 24769 4939 24803
rect 6653 24769 6687 24803
rect 6745 24769 6779 24803
rect 6837 24769 6871 24803
rect 7021 24769 7055 24803
rect 7113 24769 7147 24803
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 7573 24769 7607 24803
rect 7665 24769 7699 24803
rect 8033 24769 8067 24803
rect 8217 24769 8251 24803
rect 8953 24769 8987 24803
rect 9137 24769 9171 24803
rect 9229 24769 9263 24803
rect 9321 24769 9355 24803
rect 9597 24769 9631 24803
rect 9781 24769 9815 24803
rect 11529 24769 11563 24803
rect 13829 24769 13863 24803
rect 16221 24769 16255 24803
rect 17049 24769 17083 24803
rect 18153 24769 18187 24803
rect 18429 24769 18463 24803
rect 18521 24769 18555 24803
rect 18613 24769 18647 24803
rect 18797 24769 18831 24803
rect 19533 24769 19567 24803
rect 19717 24769 19751 24803
rect 19809 24769 19843 24803
rect 19993 24769 20027 24803
rect 20085 24769 20119 24803
rect 20177 24769 20211 24803
rect 20545 24769 20579 24803
rect 20729 24769 20763 24803
rect 21097 24769 21131 24803
rect 21189 24769 21223 24803
rect 21373 24769 21407 24803
rect 21465 24769 21499 24803
rect 21833 24769 21867 24803
rect 22017 24769 22051 24803
rect 22109 24769 22143 24803
rect 22201 24769 22235 24803
rect 23673 24769 23707 24803
rect 23949 24769 23983 24803
rect 24317 24769 24351 24803
rect 24501 24769 24535 24803
rect 25513 24769 25547 24803
rect 27169 24769 27203 24803
rect 31493 24769 31527 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32413 24769 32447 24803
rect 32505 24769 32539 24803
rect 33057 24769 33091 24803
rect 33517 24769 33551 24803
rect 33609 24769 33643 24803
rect 34161 24769 34195 24803
rect 34529 24769 34563 24803
rect 35909 24769 35943 24803
rect 36001 24769 36035 24803
rect 36645 24769 36679 24803
rect 36737 24769 36771 24803
rect 36921 24769 36955 24803
rect 37289 24769 37323 24803
rect 37473 24769 37507 24803
rect 38393 24769 38427 24803
rect 40785 24769 40819 24803
rect 41337 24769 41371 24803
rect 41705 24769 41739 24803
rect 42073 24769 42107 24803
rect 1409 24701 1443 24735
rect 1685 24701 1719 24735
rect 4261 24701 4295 24735
rect 4353 24701 4387 24735
rect 14289 24701 14323 24735
rect 20913 24701 20947 24735
rect 23765 24701 23799 24735
rect 24225 24701 24259 24735
rect 24685 24701 24719 24735
rect 27445 24701 27479 24735
rect 27537 24701 27571 24735
rect 29469 24701 29503 24735
rect 31217 24701 31251 24735
rect 31585 24701 31619 24735
rect 31677 24701 31711 24735
rect 31769 24701 31803 24735
rect 31953 24701 31987 24735
rect 32781 24701 32815 24735
rect 33885 24701 33919 24735
rect 34345 24701 34379 24735
rect 34713 24701 34747 24735
rect 35357 24701 35391 24735
rect 36277 24701 36311 24735
rect 36369 24701 36403 24735
rect 37105 24701 37139 24735
rect 37657 24701 37691 24735
rect 37841 24701 37875 24735
rect 38669 24701 38703 24735
rect 40417 24701 40451 24735
rect 41429 24701 41463 24735
rect 4721 24633 4755 24667
rect 7757 24633 7791 24667
rect 8217 24633 8251 24667
rect 9965 24633 9999 24667
rect 18429 24633 18463 24667
rect 24133 24633 24167 24667
rect 27353 24633 27387 24667
rect 29285 24633 29319 24667
rect 32965 24633 32999 24667
rect 34069 24633 34103 24667
rect 38301 24633 38335 24667
rect 9505 24565 9539 24599
rect 13277 24565 13311 24599
rect 13553 24565 13587 24599
rect 16405 24565 16439 24599
rect 18705 24565 18739 24599
rect 20821 24565 20855 24599
rect 25605 24565 25639 24599
rect 33793 24565 33827 24599
rect 37381 24565 37415 24599
rect 40601 24565 40635 24599
rect 1869 24361 1903 24395
rect 3065 24361 3099 24395
rect 7573 24361 7607 24395
rect 10701 24361 10735 24395
rect 16129 24361 16163 24395
rect 19257 24361 19291 24395
rect 20453 24361 20487 24395
rect 21557 24361 21591 24395
rect 21741 24361 21775 24395
rect 29561 24361 29595 24395
rect 31861 24361 31895 24395
rect 35357 24361 35391 24395
rect 36553 24361 36587 24395
rect 36645 24361 36679 24395
rect 37657 24361 37691 24395
rect 42165 24361 42199 24395
rect 7757 24293 7791 24327
rect 25513 24293 25547 24327
rect 31309 24293 31343 24327
rect 35173 24293 35207 24327
rect 3341 24225 3375 24259
rect 6009 24225 6043 24259
rect 7205 24225 7239 24259
rect 8125 24225 8159 24259
rect 8217 24225 8251 24259
rect 8309 24225 8343 24259
rect 9321 24225 9355 24259
rect 10793 24225 10827 24259
rect 11529 24225 11563 24259
rect 14565 24225 14599 24259
rect 15945 24225 15979 24259
rect 17233 24225 17267 24259
rect 36093 24225 36127 24259
rect 36185 24225 36219 24259
rect 36461 24225 36495 24259
rect 1869 24157 1903 24191
rect 2145 24157 2179 24191
rect 2329 24157 2363 24191
rect 2973 24157 3007 24191
rect 3157 24157 3191 24191
rect 3249 24157 3283 24191
rect 3433 24157 3467 24191
rect 4905 24157 4939 24191
rect 5549 24157 5583 24191
rect 5641 24157 5675 24191
rect 6653 24157 6687 24191
rect 8033 24157 8067 24191
rect 13369 24157 13403 24191
rect 13553 24157 13587 24191
rect 13737 24157 13771 24191
rect 15117 24157 15151 24191
rect 17601 24157 17635 24191
rect 18337 24157 18371 24191
rect 18522 24157 18556 24191
rect 18705 24157 18739 24191
rect 18981 24157 19015 24191
rect 19441 24157 19475 24191
rect 19625 24157 19659 24191
rect 19809 24157 19843 24191
rect 20085 24157 20119 24191
rect 20269 24157 20303 24191
rect 21373 24157 21407 24191
rect 21649 24157 21683 24191
rect 21833 24157 21867 24191
rect 24961 24157 24995 24191
rect 25237 24157 25271 24191
rect 25329 24157 25363 24191
rect 25973 24157 26007 24191
rect 26065 24157 26099 24191
rect 26341 24157 26375 24191
rect 28733 24157 28767 24191
rect 29745 24157 29779 24191
rect 29837 24157 29871 24191
rect 31493 24157 31527 24191
rect 36737 24157 36771 24191
rect 37105 24157 37139 24191
rect 37289 24157 37323 24191
rect 37473 24157 37507 24191
rect 40417 24157 40451 24191
rect 7619 24123 7653 24157
rect 6929 24089 6963 24123
rect 7389 24089 7423 24123
rect 9588 24089 9622 24123
rect 11805 24089 11839 24123
rect 13645 24089 13679 24123
rect 15301 24089 15335 24123
rect 16405 24089 16439 24123
rect 17049 24089 17083 24123
rect 18614 24089 18648 24123
rect 18843 24089 18877 24123
rect 19533 24089 19567 24123
rect 21189 24089 21223 24123
rect 25145 24089 25179 24123
rect 26157 24089 26191 24123
rect 31677 24089 31711 24123
rect 35325 24089 35359 24123
rect 35541 24089 35575 24123
rect 37381 24089 37415 24123
rect 40693 24089 40727 24123
rect 2053 24021 2087 24055
rect 2881 24021 2915 24055
rect 6745 24021 6779 24055
rect 8493 24021 8527 24055
rect 11437 24021 11471 24055
rect 13277 24021 13311 24055
rect 13921 24021 13955 24055
rect 16681 24021 16715 24055
rect 17141 24021 17175 24055
rect 25789 24021 25823 24055
rect 28549 24021 28583 24055
rect 31585 24021 31619 24055
rect 35633 24021 35667 24055
rect 36001 24021 36035 24055
rect 3065 23817 3099 23851
rect 6469 23817 6503 23851
rect 6929 23817 6963 23851
rect 7665 23817 7699 23851
rect 9597 23817 9631 23851
rect 11805 23817 11839 23851
rect 12265 23817 12299 23851
rect 16313 23817 16347 23851
rect 18429 23817 18463 23851
rect 18981 23817 19015 23851
rect 22385 23817 22419 23851
rect 26985 23817 27019 23851
rect 29653 23817 29687 23851
rect 38393 23817 38427 23851
rect 40969 23817 41003 23851
rect 41337 23817 41371 23851
rect 9111 23749 9145 23783
rect 9321 23749 9355 23783
rect 16957 23749 16991 23783
rect 20085 23749 20119 23783
rect 24685 23749 24719 23783
rect 35081 23749 35115 23783
rect 2605 23681 2639 23715
rect 2697 23681 2731 23715
rect 2789 23681 2823 23715
rect 3617 23681 3651 23715
rect 4905 23681 4939 23715
rect 5089 23681 5123 23715
rect 6469 23681 6503 23715
rect 6745 23681 6779 23715
rect 6837 23681 6871 23715
rect 7481 23681 7515 23715
rect 7757 23681 7791 23715
rect 9229 23681 9263 23715
rect 9413 23681 9447 23715
rect 9781 23681 9815 23715
rect 10037 23681 10071 23715
rect 12173 23681 12207 23715
rect 13737 23681 13771 23715
rect 14004 23681 14038 23715
rect 15577 23681 15611 23715
rect 16405 23681 16439 23715
rect 16688 23681 16722 23715
rect 18613 23681 18647 23715
rect 18797 23681 18831 23715
rect 19993 23681 20027 23715
rect 20177 23681 20211 23715
rect 20361 23681 20395 23715
rect 24961 23681 24995 23715
rect 28109 23681 28143 23715
rect 29009 23681 29043 23715
rect 32137 23681 32171 23715
rect 32321 23681 32355 23715
rect 32413 23681 32447 23715
rect 32505 23681 32539 23715
rect 34897 23681 34931 23715
rect 34989 23681 35023 23715
rect 35265 23681 35299 23715
rect 39405 23681 39439 23715
rect 39672 23681 39706 23715
rect 6561 23613 6595 23647
rect 7205 23613 7239 23647
rect 8953 23613 8987 23647
rect 12449 23613 12483 23647
rect 15669 23613 15703 23647
rect 15761 23613 15795 23647
rect 21373 23613 21407 23647
rect 22477 23613 22511 23647
rect 22569 23613 22603 23647
rect 25697 23613 25731 23647
rect 25881 23613 25915 23647
rect 28365 23613 28399 23647
rect 29377 23613 29411 23647
rect 29561 23613 29595 23647
rect 30941 23613 30975 23647
rect 33425 23613 33459 23647
rect 34069 23613 34103 23647
rect 38485 23613 38519 23647
rect 38577 23613 38611 23647
rect 41429 23613 41463 23647
rect 41521 23613 41555 23647
rect 2973 23545 3007 23579
rect 23213 23545 23247 23579
rect 30297 23545 30331 23579
rect 4997 23477 5031 23511
rect 7389 23477 7423 23511
rect 11161 23477 11195 23511
rect 15117 23477 15151 23511
rect 15209 23477 15243 23511
rect 19809 23477 19843 23511
rect 20821 23477 20855 23511
rect 22017 23477 22051 23511
rect 25053 23477 25087 23511
rect 26525 23477 26559 23511
rect 28457 23477 28491 23511
rect 30021 23477 30055 23511
rect 32689 23477 32723 23511
rect 34713 23477 34747 23511
rect 38025 23477 38059 23511
rect 40785 23477 40819 23511
rect 3341 23273 3375 23307
rect 7481 23273 7515 23307
rect 9781 23273 9815 23307
rect 11069 23273 11103 23307
rect 15577 23273 15611 23307
rect 23213 23273 23247 23307
rect 28365 23273 28399 23307
rect 30941 23273 30975 23307
rect 37197 23273 37231 23307
rect 39865 23273 39899 23307
rect 41521 23273 41555 23307
rect 2881 23205 2915 23239
rect 4353 23137 4387 23171
rect 4721 23137 4755 23171
rect 6377 23137 6411 23171
rect 10517 23137 10551 23171
rect 12541 23137 12575 23171
rect 15485 23137 15519 23171
rect 18245 23137 18279 23171
rect 27261 23137 27295 23171
rect 27445 23137 27479 23171
rect 31677 23137 31711 23171
rect 33149 23137 33183 23171
rect 35449 23137 35483 23171
rect 37657 23137 37691 23171
rect 40417 23137 40451 23171
rect 40785 23137 40819 23171
rect 42073 23137 42107 23171
rect 1409 23069 1443 23103
rect 2513 23069 2547 23103
rect 2605 23069 2639 23103
rect 2697 23069 2731 23103
rect 3617 23069 3651 23103
rect 3801 23069 3835 23103
rect 6285 23069 6319 23103
rect 6469 23069 6503 23103
rect 6837 23069 6871 23103
rect 7665 23069 7699 23103
rect 7941 23069 7975 23103
rect 8125 23069 8159 23103
rect 8217 23069 8251 23103
rect 8493 23069 8527 23103
rect 8585 23069 8619 23103
rect 9229 23069 9263 23103
rect 9413 23069 9447 23103
rect 9597 23069 9631 23103
rect 11161 23069 11195 23103
rect 15218 23069 15252 23103
rect 16129 23069 16163 23103
rect 17509 23069 17543 23103
rect 19809 23069 19843 23103
rect 20453 23069 20487 23103
rect 21925 23069 21959 23103
rect 24409 23069 24443 23103
rect 26994 23069 27028 23103
rect 28549 23069 28583 23103
rect 28641 23069 28675 23103
rect 28917 23069 28951 23103
rect 29561 23069 29595 23103
rect 31033 23069 31067 23103
rect 31401 23069 31435 23103
rect 33416 23069 33450 23103
rect 34713 23069 34747 23103
rect 37924 23069 37958 23103
rect 40233 23069 40267 23103
rect 2973 23001 3007 23035
rect 3350 23001 3384 23035
rect 6147 23001 6181 23035
rect 7113 23001 7147 23035
rect 7297 23001 7331 23035
rect 8401 23001 8435 23035
rect 9505 23001 9539 23035
rect 12265 23001 12299 23035
rect 20720 23001 20754 23035
rect 24654 23001 24688 23035
rect 28273 23001 28307 23035
rect 28733 23001 28767 23035
rect 29828 23001 29862 23035
rect 31217 23001 31251 23035
rect 31309 23001 31343 23035
rect 31922 23001 31956 23035
rect 35725 23001 35759 23035
rect 1593 22933 1627 22967
rect 3985 22933 4019 22967
rect 6653 22933 6687 22967
rect 7757 22933 7791 22967
rect 8769 22933 8803 22967
rect 11805 22933 11839 22967
rect 11897 22933 11931 22967
rect 12357 22933 12391 22967
rect 14105 22933 14139 22967
rect 19257 22933 19291 22967
rect 21833 22933 21867 22967
rect 25789 22933 25823 22967
rect 25881 22933 25915 22967
rect 31585 22933 31619 22967
rect 33057 22933 33091 22967
rect 34529 22933 34563 22967
rect 35357 22933 35391 22967
rect 39037 22933 39071 22967
rect 40325 22933 40359 22967
rect 41429 22933 41463 22967
rect 1409 22729 1443 22763
rect 5181 22729 5215 22763
rect 9689 22729 9723 22763
rect 13277 22729 13311 22763
rect 18245 22729 18279 22763
rect 19717 22729 19751 22763
rect 21189 22729 21223 22763
rect 32137 22729 32171 22763
rect 33425 22729 33459 22763
rect 41061 22729 41095 22763
rect 41889 22729 41923 22763
rect 2881 22661 2915 22695
rect 6745 22661 6779 22695
rect 9321 22661 9355 22695
rect 9413 22661 9447 22695
rect 10026 22661 10060 22695
rect 11805 22661 11839 22695
rect 17877 22661 17911 22695
rect 17969 22661 18003 22695
rect 23305 22661 23339 22695
rect 23673 22661 23707 22695
rect 26004 22661 26038 22695
rect 34560 22661 34594 22695
rect 41797 22661 41831 22695
rect 4537 22593 4571 22627
rect 4721 22593 4755 22627
rect 4813 22593 4847 22627
rect 4905 22593 4939 22627
rect 5273 22593 5307 22627
rect 6653 22593 6687 22627
rect 6837 22593 6871 22627
rect 6929 22593 6963 22627
rect 7113 22593 7147 22627
rect 7389 22593 7423 22627
rect 7849 22593 7883 22627
rect 8309 22593 8343 22627
rect 8493 22593 8527 22627
rect 8585 22593 8619 22627
rect 8677 22593 8711 22627
rect 9137 22593 9171 22627
rect 9505 22593 9539 22627
rect 11529 22593 11563 22627
rect 14749 22593 14783 22627
rect 17325 22593 17359 22627
rect 17693 22593 17727 22627
rect 18061 22593 18095 22627
rect 18593 22593 18627 22627
rect 20076 22593 20110 22627
rect 26249 22593 26283 22627
rect 26985 22593 27019 22627
rect 27252 22593 27286 22627
rect 30564 22593 30598 22627
rect 34805 22593 34839 22627
rect 36021 22593 36055 22627
rect 36277 22593 36311 22627
rect 37289 22593 37323 22627
rect 37556 22593 37590 22627
rect 39313 22593 39347 22627
rect 39580 22593 39614 22627
rect 41153 22593 41187 22627
rect 3157 22525 3191 22559
rect 5181 22525 5215 22559
rect 7573 22525 7607 22559
rect 7665 22525 7699 22559
rect 7757 22525 7791 22559
rect 8033 22525 8067 22559
rect 9781 22525 9815 22559
rect 14841 22525 14875 22559
rect 18337 22525 18371 22559
rect 19809 22525 19843 22559
rect 23581 22525 23615 22559
rect 24225 22525 24259 22559
rect 28457 22525 28491 22559
rect 28733 22525 28767 22559
rect 30297 22525 30331 22559
rect 32781 22525 32815 22559
rect 36369 22525 36403 22559
rect 36921 22525 36955 22559
rect 40877 22525 40911 22559
rect 8861 22457 8895 22491
rect 4537 22389 4571 22423
rect 4997 22389 5031 22423
rect 5365 22389 5399 22423
rect 7297 22389 7331 22423
rect 11161 22389 11195 22423
rect 15117 22389 15151 22423
rect 16681 22389 16715 22423
rect 21833 22389 21867 22423
rect 24869 22389 24903 22423
rect 28365 22389 28399 22423
rect 30205 22389 30239 22423
rect 31677 22389 31711 22423
rect 34897 22389 34931 22423
rect 38669 22389 38703 22423
rect 40693 22389 40727 22423
rect 41521 22389 41555 22423
rect 2899 22185 2933 22219
rect 27353 22185 27387 22219
rect 29561 22185 29595 22219
rect 30941 22185 30975 22219
rect 37749 22185 37783 22219
rect 5733 22117 5767 22151
rect 7113 22049 7147 22083
rect 7297 22049 7331 22083
rect 8033 22049 8067 22083
rect 15301 22049 15335 22083
rect 15485 22049 15519 22083
rect 16313 22049 16347 22083
rect 18889 22049 18923 22083
rect 19809 22049 19843 22083
rect 21925 22049 21959 22083
rect 22385 22049 22419 22083
rect 23581 22049 23615 22083
rect 26433 22049 26467 22083
rect 26985 22049 27019 22083
rect 27997 22049 28031 22083
rect 28733 22049 28767 22083
rect 30021 22049 30055 22083
rect 30205 22049 30239 22083
rect 31585 22049 31619 22083
rect 32321 22049 32355 22083
rect 33241 22049 33275 22083
rect 38301 22049 38335 22083
rect 39129 22049 39163 22083
rect 40509 22049 40543 22083
rect 41981 22049 42015 22083
rect 3157 21981 3191 22015
rect 3985 21981 4019 22015
rect 6837 21981 6871 22015
rect 7021 21981 7055 22015
rect 7389 21981 7423 22015
rect 7757 21981 7791 22015
rect 7849 21981 7883 22015
rect 8125 21981 8159 22015
rect 8217 21981 8251 22015
rect 8401 21981 8435 22015
rect 8585 21981 8619 22015
rect 9137 21981 9171 22015
rect 11897 21981 11931 22015
rect 16037 21981 16071 22015
rect 16773 21981 16807 22015
rect 18613 21981 18647 22015
rect 21649 21981 21683 22015
rect 22477 21981 22511 22015
rect 23029 21981 23063 22015
rect 25605 21981 25639 22015
rect 26249 21981 26283 22015
rect 27721 21981 27755 22015
rect 31309 21981 31343 22015
rect 32965 21981 32999 22015
rect 33977 21981 34011 22015
rect 34989 21981 35023 22015
rect 37013 21981 37047 22015
rect 38117 21981 38151 22015
rect 40233 21981 40267 22015
rect 4261 21913 4295 21947
rect 6929 21913 6963 21947
rect 8493 21913 8527 21947
rect 9382 21913 9416 21947
rect 12173 21913 12207 21947
rect 13921 21913 13955 21947
rect 15209 21913 15243 21947
rect 17040 21913 17074 21947
rect 20076 21913 20110 21947
rect 22569 21913 22603 21947
rect 35256 21913 35290 21947
rect 1409 21845 1443 21879
rect 7389 21845 7423 21879
rect 7573 21845 7607 21879
rect 8769 21845 8803 21879
rect 10517 21845 10551 21879
rect 14841 21845 14875 21879
rect 15669 21845 15703 21879
rect 16129 21845 16163 21879
rect 18153 21845 18187 21879
rect 18245 21845 18279 21879
rect 18705 21845 18739 21879
rect 21189 21845 21223 21879
rect 21281 21845 21315 21879
rect 21741 21845 21775 21879
rect 22937 21845 22971 21879
rect 24961 21845 24995 21879
rect 25697 21845 25731 21879
rect 27813 21845 27847 21879
rect 28181 21845 28215 21879
rect 29929 21845 29963 21879
rect 31401 21845 31435 21879
rect 31769 21845 31803 21879
rect 32597 21845 32631 21879
rect 33057 21845 33091 21879
rect 33425 21845 33459 21879
rect 36369 21845 36403 21879
rect 36461 21845 36495 21879
rect 38209 21845 38243 21879
rect 38577 21845 38611 21879
rect 1593 21641 1627 21675
rect 4353 21641 4387 21675
rect 7757 21641 7791 21675
rect 12357 21641 12391 21675
rect 12817 21641 12851 21675
rect 16497 21641 16531 21675
rect 24317 21641 24351 21675
rect 24409 21641 24443 21675
rect 28181 21641 28215 21675
rect 30113 21641 30147 21675
rect 31309 21641 31343 21675
rect 33517 21641 33551 21675
rect 35265 21641 35299 21675
rect 39497 21641 39531 21675
rect 39865 21641 39899 21675
rect 4521 21573 4555 21607
rect 4721 21573 4755 21607
rect 9597 21573 9631 21607
rect 12725 21573 12759 21607
rect 14105 21573 14139 21607
rect 14381 21573 14415 21607
rect 15025 21573 15059 21607
rect 32404 21573 32438 21607
rect 34069 21573 34103 21607
rect 34161 21573 34195 21607
rect 35541 21573 35575 21607
rect 1409 21505 1443 21539
rect 1777 21505 1811 21539
rect 4813 21505 4847 21539
rect 4997 21505 5031 21539
rect 7481 21505 7515 21539
rect 10149 21505 10183 21539
rect 14565 21505 14599 21539
rect 22937 21505 22971 21539
rect 23204 21505 23238 21539
rect 24593 21505 24627 21539
rect 24685 21505 24719 21539
rect 24777 21505 24811 21539
rect 24961 21505 24995 21539
rect 25320 21505 25354 21539
rect 28089 21505 28123 21539
rect 28549 21505 28583 21539
rect 30665 21505 30699 21539
rect 31217 21505 31251 21539
rect 33885 21505 33919 21539
rect 34253 21505 34287 21539
rect 35449 21505 35483 21539
rect 35633 21505 35667 21539
rect 35817 21505 35851 21539
rect 39957 21505 39991 21539
rect 7757 21437 7791 21471
rect 13001 21437 13035 21471
rect 14749 21437 14783 21471
rect 17141 21437 17175 21471
rect 17417 21437 17451 21471
rect 19533 21437 19567 21471
rect 20269 21437 20303 21471
rect 21649 21437 21683 21471
rect 22385 21437 22419 21471
rect 25053 21437 25087 21471
rect 26985 21437 27019 21471
rect 28273 21437 28307 21471
rect 29101 21437 29135 21471
rect 31401 21437 31435 21471
rect 32137 21437 32171 21471
rect 35081 21437 35115 21471
rect 37289 21437 37323 21471
rect 37565 21437 37599 21471
rect 40049 21437 40083 21471
rect 40325 21437 40359 21471
rect 40601 21437 40635 21471
rect 1961 21369 1995 21403
rect 4813 21369 4847 21403
rect 18889 21369 18923 21403
rect 26433 21369 26467 21403
rect 34437 21369 34471 21403
rect 4537 21301 4571 21335
rect 7573 21301 7607 21335
rect 14197 21301 14231 21335
rect 18981 21301 19015 21335
rect 19717 21301 19751 21335
rect 21005 21301 21039 21335
rect 21833 21301 21867 21335
rect 27629 21301 27663 21335
rect 27721 21301 27755 21335
rect 30849 21301 30883 21335
rect 34529 21301 34563 21335
rect 39037 21301 39071 21335
rect 42073 21301 42107 21335
rect 1409 21097 1443 21131
rect 11161 21097 11195 21131
rect 16589 21097 16623 21131
rect 17693 21097 17727 21131
rect 23029 21097 23063 21131
rect 23489 21097 23523 21131
rect 28917 21097 28951 21131
rect 31953 21097 31987 21131
rect 37197 21097 37231 21131
rect 40509 21097 40543 21131
rect 41337 21097 41371 21131
rect 35265 21029 35299 21063
rect 2881 20961 2915 20995
rect 5549 20961 5583 20995
rect 14105 20961 14139 20995
rect 14381 20961 14415 20995
rect 15853 20961 15887 20995
rect 15945 20961 15979 20995
rect 18153 20961 18187 20995
rect 18245 20961 18279 20995
rect 18613 20961 18647 20995
rect 20913 20961 20947 20995
rect 21005 20961 21039 20995
rect 21281 20961 21315 20995
rect 23949 20961 23983 20995
rect 24041 20961 24075 20995
rect 24869 20961 24903 20995
rect 25053 20961 25087 20995
rect 26157 20961 26191 20995
rect 27169 20961 27203 20995
rect 30113 20961 30147 20995
rect 30389 20961 30423 20995
rect 37657 20961 37691 20995
rect 37841 20961 37875 20995
rect 39589 20961 39623 20995
rect 41061 20961 41095 20995
rect 41889 20961 41923 20995
rect 3157 20893 3191 20927
rect 3985 20893 4019 20927
rect 4077 20893 4111 20927
rect 4261 20893 4295 20927
rect 4353 20893 4387 20927
rect 4905 20893 4939 20927
rect 4997 20893 5031 20927
rect 5181 20893 5215 20927
rect 5273 20893 5307 20927
rect 5457 20893 5491 20927
rect 5917 20893 5951 20927
rect 16773 20893 16807 20927
rect 18521 20893 18555 20927
rect 18797 20893 18831 20927
rect 18889 20893 18923 20927
rect 19073 20893 19107 20927
rect 19349 20893 19383 20927
rect 20821 20893 20855 20927
rect 23857 20893 23891 20927
rect 25973 20893 26007 20927
rect 26985 20893 27019 20927
rect 32505 20893 32539 20927
rect 33425 20893 33459 20927
rect 33609 20893 33643 20927
rect 34253 20893 34287 20927
rect 34713 20893 34747 20927
rect 34989 20893 35023 20927
rect 35081 20893 35115 20927
rect 35357 20893 35391 20927
rect 37565 20893 37599 20927
rect 39037 20893 39071 20927
rect 7389 20825 7423 20859
rect 10977 20825 11011 20859
rect 11193 20825 11227 20859
rect 18061 20825 18095 20859
rect 21557 20825 21591 20859
rect 24777 20825 24811 20859
rect 26433 20825 26467 20859
rect 27445 20825 27479 20859
rect 34897 20825 34931 20859
rect 38025 20825 38059 20859
rect 38853 20825 38887 20859
rect 39865 20825 39899 20859
rect 40877 20825 40911 20859
rect 3801 20757 3835 20791
rect 11345 20757 11379 20791
rect 17417 20757 17451 20791
rect 19993 20757 20027 20791
rect 20453 20757 20487 20791
rect 24409 20757 24443 20791
rect 25605 20757 25639 20791
rect 26065 20757 26099 20791
rect 31861 20757 31895 20791
rect 33701 20757 33735 20791
rect 36001 20757 36035 20791
rect 40969 20757 41003 20791
rect 5273 20553 5307 20587
rect 5457 20553 5491 20587
rect 5825 20553 5859 20587
rect 15025 20553 15059 20587
rect 17049 20553 17083 20587
rect 22293 20553 22327 20587
rect 24777 20553 24811 20587
rect 27445 20553 27479 20587
rect 29561 20553 29595 20587
rect 31953 20553 31987 20587
rect 34069 20553 34103 20587
rect 41521 20553 41555 20587
rect 10701 20485 10735 20519
rect 11774 20485 11808 20519
rect 15301 20485 15335 20519
rect 16129 20485 16163 20519
rect 20177 20485 20211 20519
rect 36746 20485 36780 20519
rect 37657 20485 37691 20519
rect 40325 20485 40359 20519
rect 3341 20417 3375 20451
rect 4905 20417 4939 20451
rect 5365 20417 5399 20451
rect 5549 20417 5583 20451
rect 5641 20417 5675 20451
rect 5825 20417 5859 20451
rect 8953 20417 8987 20451
rect 10241 20417 10275 20451
rect 11529 20417 11563 20451
rect 14197 20417 14231 20451
rect 14381 20417 14415 20451
rect 14565 20417 14599 20451
rect 14841 20417 14875 20451
rect 15117 20417 15151 20451
rect 16221 20417 16255 20451
rect 17949 20417 17983 20451
rect 19901 20417 19935 20451
rect 27353 20417 27387 20451
rect 27813 20417 27847 20451
rect 34428 20417 34462 20451
rect 40877 20417 40911 20451
rect 41275 20417 41309 20451
rect 41429 20417 41463 20451
rect 42073 20417 42107 20451
rect 2973 20349 3007 20383
rect 4997 20349 5031 20383
rect 9965 20349 9999 20383
rect 10333 20349 10367 20383
rect 11345 20349 11379 20383
rect 14105 20349 14139 20383
rect 17141 20349 17175 20383
rect 17325 20349 17359 20383
rect 17693 20349 17727 20383
rect 19809 20349 19843 20383
rect 21649 20349 21683 20383
rect 22385 20349 22419 20383
rect 22477 20349 22511 20383
rect 23029 20349 23063 20383
rect 23305 20349 23339 20383
rect 25053 20349 25087 20383
rect 25329 20349 25363 20383
rect 27537 20349 27571 20383
rect 28089 20349 28123 20383
rect 30205 20349 30239 20383
rect 30481 20349 30515 20383
rect 32321 20349 32355 20383
rect 32597 20349 32631 20383
rect 34161 20349 34195 20383
rect 37013 20349 37047 20383
rect 37749 20349 37783 20383
rect 37933 20349 37967 20383
rect 38117 20349 38151 20383
rect 39589 20349 39623 20383
rect 39865 20349 39899 20383
rect 4767 20281 4801 20315
rect 9321 20281 9355 20315
rect 21925 20281 21959 20315
rect 26985 20281 27019 20315
rect 35633 20281 35667 20315
rect 41061 20281 41095 20315
rect 5089 20213 5123 20247
rect 9137 20213 9171 20247
rect 10609 20213 10643 20247
rect 12909 20213 12943 20247
rect 14749 20213 14783 20247
rect 16313 20213 16347 20247
rect 16681 20213 16715 20247
rect 19073 20213 19107 20247
rect 19165 20213 19199 20247
rect 26801 20213 26835 20247
rect 35541 20213 35575 20247
rect 37289 20213 37323 20247
rect 10333 20009 10367 20043
rect 12173 20009 12207 20043
rect 16313 20009 16347 20043
rect 17785 20009 17819 20043
rect 18245 20009 18279 20043
rect 27077 20009 27111 20043
rect 27813 20009 27847 20043
rect 28457 20009 28491 20043
rect 31217 20009 31251 20043
rect 32781 20009 32815 20043
rect 34529 20009 34563 20043
rect 37841 20009 37875 20043
rect 38669 20009 38703 20043
rect 6009 19873 6043 19907
rect 6101 19873 6135 19907
rect 8125 19873 8159 19907
rect 13829 19873 13863 19907
rect 14933 19873 14967 19907
rect 25329 19873 25363 19907
rect 29009 19873 29043 19907
rect 31769 19873 31803 19907
rect 33241 19873 33275 19907
rect 33425 19873 33459 19907
rect 33885 19873 33919 19907
rect 35541 19873 35575 19907
rect 36093 19873 36127 19907
rect 39221 19873 39255 19907
rect 5825 19805 5859 19839
rect 5917 19805 5951 19839
rect 6653 19805 6687 19839
rect 8217 19805 8251 19839
rect 8953 19805 8987 19839
rect 10609 19805 10643 19839
rect 10865 19805 10899 19839
rect 12265 19805 12299 19839
rect 16405 19805 16439 19839
rect 17969 19805 18003 19839
rect 18061 19805 18095 19839
rect 18337 19805 18371 19839
rect 19073 19805 19107 19839
rect 19257 19805 19291 19839
rect 19524 19805 19558 19839
rect 27169 19805 27203 19839
rect 28825 19805 28859 19839
rect 31585 19805 31619 19839
rect 33149 19805 33183 19839
rect 34161 19805 34195 19839
rect 38117 19805 38151 19839
rect 38209 19805 38243 19839
rect 38485 19805 38519 19839
rect 39037 19805 39071 19839
rect 40049 19805 40083 19839
rect 40141 19805 40175 19839
rect 40417 19805 40451 19839
rect 41153 19805 41187 19839
rect 42165 19805 42199 19839
rect 3801 19737 3835 19771
rect 9198 19737 9232 19771
rect 13584 19737 13618 19771
rect 15200 19737 15234 19771
rect 25605 19737 25639 19771
rect 28917 19737 28951 19771
rect 36369 19737 36403 19771
rect 38301 19737 38335 19771
rect 39129 19737 39163 19771
rect 40233 19737 40267 19771
rect 6285 19669 6319 19703
rect 6469 19669 6503 19703
rect 8585 19669 8619 19703
rect 11989 19669 12023 19703
rect 12449 19669 12483 19703
rect 18429 19669 18463 19703
rect 20637 19669 20671 19703
rect 31677 19669 31711 19703
rect 34069 19669 34103 19703
rect 34897 19669 34931 19703
rect 37933 19669 37967 19703
rect 39865 19669 39899 19703
rect 40601 19669 40635 19703
rect 41521 19669 41555 19703
rect 5825 19465 5859 19499
rect 6009 19465 6043 19499
rect 8217 19465 8251 19499
rect 12081 19465 12115 19499
rect 16497 19465 16531 19499
rect 18429 19465 18463 19499
rect 23673 19465 23707 19499
rect 25605 19465 25639 19499
rect 25973 19465 26007 19499
rect 29285 19465 29319 19499
rect 33241 19465 33275 19499
rect 38485 19465 38519 19499
rect 40969 19465 41003 19499
rect 9444 19397 9478 19431
rect 10149 19397 10183 19431
rect 12173 19397 12207 19431
rect 13829 19397 13863 19431
rect 32689 19397 32723 19431
rect 39497 19397 39531 19431
rect 2421 19329 2455 19363
rect 2789 19329 2823 19363
rect 4353 19329 4387 19363
rect 5917 19329 5951 19363
rect 6377 19329 6411 19363
rect 6644 19329 6678 19363
rect 8033 19329 8067 19363
rect 8217 19329 8251 19363
rect 11161 19329 11195 19363
rect 11989 19329 12023 19363
rect 13461 19329 13495 19363
rect 13553 19329 13587 19363
rect 13921 19329 13955 19363
rect 14105 19329 14139 19363
rect 15117 19329 15151 19363
rect 15384 19329 15418 19363
rect 16681 19329 16715 19363
rect 19533 19329 19567 19363
rect 21833 19329 21867 19363
rect 27445 19329 27479 19363
rect 30205 19329 30239 19363
rect 32505 19329 32539 19363
rect 32781 19329 32815 19363
rect 32873 19329 32907 19363
rect 33241 19329 33275 19363
rect 33425 19329 33459 19363
rect 33977 19329 34011 19363
rect 34161 19329 34195 19363
rect 34253 19329 34287 19363
rect 34345 19329 34379 19363
rect 34621 19329 34655 19363
rect 34888 19329 34922 19363
rect 36737 19329 36771 19363
rect 36921 19329 36955 19363
rect 37105 19329 37139 19363
rect 37289 19329 37323 19363
rect 37473 19329 37507 19363
rect 37657 19329 37691 19363
rect 41797 19329 41831 19363
rect 4905 19261 4939 19295
rect 9689 19261 9723 19295
rect 10885 19261 10919 19295
rect 12817 19261 12851 19295
rect 13829 19261 13863 19295
rect 16957 19261 16991 19295
rect 19809 19261 19843 19295
rect 21281 19261 21315 19295
rect 22109 19261 22143 19295
rect 23581 19261 23615 19295
rect 24225 19261 24259 19295
rect 26065 19261 26099 19295
rect 26157 19261 26191 19295
rect 27721 19261 27755 19295
rect 29193 19261 29227 19295
rect 29837 19261 29871 19295
rect 30757 19261 30791 19295
rect 36093 19261 36127 19295
rect 39037 19261 39071 19295
rect 39221 19261 39255 19295
rect 41613 19261 41647 19295
rect 5641 19193 5675 19227
rect 8309 19193 8343 19227
rect 11805 19193 11839 19227
rect 13645 19193 13679 19227
rect 13921 19193 13955 19227
rect 41981 19193 42015 19227
rect 4215 19125 4249 19159
rect 6193 19125 6227 19159
rect 7757 19125 7791 19159
rect 11253 19125 11287 19159
rect 12357 19125 12391 19159
rect 32597 19125 32631 19159
rect 34529 19125 34563 19159
rect 36001 19125 36035 19159
rect 37013 19125 37047 19159
rect 37473 19125 37507 19159
rect 38209 19125 38243 19159
rect 41061 19125 41095 19159
rect 3203 18921 3237 18955
rect 4813 18921 4847 18955
rect 6561 18921 6595 18955
rect 6745 18921 6779 18955
rect 10333 18921 10367 18955
rect 11345 18921 11379 18955
rect 11713 18921 11747 18955
rect 11897 18921 11931 18955
rect 12173 18921 12207 18955
rect 12817 18921 12851 18955
rect 15393 18921 15427 18955
rect 17233 18921 17267 18955
rect 20269 18921 20303 18955
rect 28181 18921 28215 18955
rect 35449 18921 35483 18955
rect 37381 18921 37415 18955
rect 42165 18921 42199 18955
rect 5089 18853 5123 18887
rect 6193 18853 6227 18887
rect 32413 18853 32447 18887
rect 36645 18853 36679 18887
rect 40141 18853 40175 18887
rect 1409 18785 1443 18819
rect 3985 18785 4019 18819
rect 9229 18785 9263 18819
rect 9689 18785 9723 18819
rect 17785 18785 17819 18819
rect 20821 18785 20855 18819
rect 24133 18785 24167 18819
rect 24961 18785 24995 18819
rect 28825 18785 28859 18819
rect 30665 18785 30699 18819
rect 33057 18785 33091 18819
rect 34805 18785 34839 18819
rect 36185 18785 36219 18819
rect 36921 18785 36955 18819
rect 37473 18785 37507 18819
rect 38945 18785 38979 18819
rect 40325 18785 40359 18819
rect 40693 18785 40727 18819
rect 1777 18717 1811 18751
rect 4721 18717 4755 18751
rect 4997 18717 5031 18751
rect 5181 18717 5215 18751
rect 5273 18717 5307 18751
rect 5457 18717 5491 18751
rect 5549 18717 5583 18751
rect 5641 18717 5675 18751
rect 5825 18717 5859 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 9321 18717 9355 18751
rect 9505 18717 9539 18751
rect 10701 18717 10735 18751
rect 10885 18717 10919 18751
rect 11161 18717 11195 18751
rect 12633 18717 12667 18751
rect 14657 18717 14691 18751
rect 15577 18717 15611 18751
rect 15761 18717 15795 18751
rect 15853 18717 15887 18751
rect 17601 18717 17635 18751
rect 21281 18717 21315 18751
rect 22385 18717 22419 18751
rect 28365 18717 28399 18751
rect 28549 18717 28583 18751
rect 28687 18717 28721 18751
rect 29193 18717 29227 18751
rect 29377 18717 29411 18751
rect 29561 18717 29595 18751
rect 33977 18717 34011 18751
rect 36277 18717 36311 18751
rect 37013 18717 37047 18751
rect 37197 18717 37231 18751
rect 39221 18717 39255 18751
rect 40049 18717 40083 18751
rect 40417 18717 40451 18751
rect 6561 18649 6595 18683
rect 9781 18649 9815 18683
rect 11529 18649 11563 18683
rect 12141 18649 12175 18683
rect 12357 18649 12391 18683
rect 12449 18649 12483 18683
rect 20729 18649 20763 18683
rect 22109 18649 22143 18683
rect 22661 18649 22695 18683
rect 24409 18649 24443 18683
rect 28457 18649 28491 18683
rect 30941 18649 30975 18683
rect 6009 18581 6043 18615
rect 9965 18581 9999 18615
rect 10057 18581 10091 18615
rect 10149 18581 10183 18615
rect 10977 18581 11011 18615
rect 11729 18581 11763 18615
rect 11989 18581 12023 18615
rect 14105 18581 14139 18615
rect 17693 18581 17727 18615
rect 20637 18581 20671 18615
rect 29193 18581 29227 18615
rect 30205 18581 30239 18615
rect 32505 18581 32539 18615
rect 33425 18581 33459 18615
rect 40325 18581 40359 18615
rect 1593 18377 1627 18411
rect 4261 18377 4295 18411
rect 5273 18377 5307 18411
rect 9965 18377 9999 18411
rect 11805 18377 11839 18411
rect 11897 18377 11931 18411
rect 21833 18377 21867 18411
rect 22569 18377 22603 18411
rect 28457 18377 28491 18411
rect 28641 18377 28675 18411
rect 31217 18377 31251 18411
rect 32689 18377 32723 18411
rect 37381 18377 37415 18411
rect 38485 18377 38519 18411
rect 41061 18377 41095 18411
rect 41797 18377 41831 18411
rect 4445 18309 4479 18343
rect 4813 18309 4847 18343
rect 4905 18309 4939 18343
rect 11100 18309 11134 18343
rect 18613 18309 18647 18343
rect 19073 18309 19107 18343
rect 24593 18309 24627 18343
rect 30113 18309 30147 18343
rect 30481 18309 30515 18343
rect 30665 18309 30699 18343
rect 31493 18309 31527 18343
rect 31703 18309 31737 18343
rect 32321 18309 32355 18343
rect 33057 18309 33091 18343
rect 41337 18309 41371 18343
rect 41429 18309 41463 18343
rect 1409 18241 1443 18275
rect 4031 18241 4065 18275
rect 4169 18241 4203 18275
rect 4997 18241 5031 18275
rect 5641 18241 5675 18275
rect 7757 18241 7791 18275
rect 7849 18241 7883 18275
rect 7941 18241 7975 18275
rect 9321 18241 9355 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 13185 18241 13219 18275
rect 13645 18241 13679 18275
rect 13901 18241 13935 18275
rect 15117 18241 15151 18275
rect 15301 18241 15335 18275
rect 15393 18241 15427 18275
rect 18889 18241 18923 18275
rect 18981 18241 19015 18275
rect 19257 18241 19291 18275
rect 19625 18241 19659 18275
rect 19717 18241 19751 18275
rect 19901 18241 19935 18275
rect 21465 18241 21499 18275
rect 22017 18241 22051 18275
rect 22109 18241 22143 18275
rect 22201 18241 22235 18275
rect 22385 18241 22419 18275
rect 23489 18241 23523 18275
rect 23581 18241 23615 18275
rect 23673 18241 23707 18275
rect 23857 18241 23891 18275
rect 23949 18241 23983 18275
rect 24133 18241 24167 18275
rect 24317 18241 24351 18275
rect 26985 18241 27019 18275
rect 27169 18241 27203 18275
rect 27261 18241 27295 18275
rect 27445 18241 27479 18275
rect 28273 18241 28307 18275
rect 28457 18241 28491 18275
rect 28549 18241 28583 18275
rect 30389 18241 30423 18275
rect 31401 18241 31435 18275
rect 31585 18241 31619 18275
rect 32137 18241 32171 18275
rect 32413 18241 32447 18275
rect 32505 18241 32539 18275
rect 38025 18241 38059 18275
rect 39037 18241 39071 18275
rect 39865 18241 39899 18275
rect 41245 18241 41279 18275
rect 41613 18241 41647 18275
rect 41705 18241 41739 18275
rect 41889 18241 41923 18275
rect 41981 18241 42015 18275
rect 42165 18241 42199 18275
rect 2237 18173 2271 18207
rect 2605 18173 2639 18207
rect 5181 18173 5215 18207
rect 5457 18173 5491 18207
rect 5549 18173 5583 18207
rect 5733 18173 5767 18207
rect 11345 18173 11379 18207
rect 11529 18173 11563 18207
rect 12014 18173 12048 18207
rect 13093 18173 13127 18207
rect 13553 18173 13587 18207
rect 17325 18173 17359 18207
rect 18061 18173 18095 18207
rect 19349 18173 19383 18207
rect 19533 18173 19567 18207
rect 19809 18173 19843 18207
rect 23213 18173 23247 18207
rect 26065 18173 26099 18207
rect 26709 18173 26743 18207
rect 27353 18173 27387 18207
rect 31861 18173 31895 18207
rect 32781 18173 32815 18207
rect 35357 18173 35391 18207
rect 35633 18173 35667 18207
rect 39773 18173 39807 18207
rect 40233 18173 40267 18207
rect 8125 18105 8159 18139
rect 23305 18105 23339 18139
rect 23949 18105 23983 18139
rect 26157 18105 26191 18139
rect 37105 18105 37139 18139
rect 42073 18105 42107 18139
rect 7573 18037 7607 18071
rect 9137 18037 9171 18071
rect 9413 18037 9447 18071
rect 12173 18037 12207 18071
rect 15025 18037 15059 18071
rect 15117 18037 15151 18071
rect 16681 18037 16715 18071
rect 18705 18037 18739 18071
rect 19441 18037 19475 18071
rect 27077 18037 27111 18071
rect 30849 18037 30883 18071
rect 34529 18037 34563 18071
rect 3801 17833 3835 17867
rect 5365 17833 5399 17867
rect 5641 17833 5675 17867
rect 9137 17833 9171 17867
rect 10425 17833 10459 17867
rect 10609 17833 10643 17867
rect 13001 17833 13035 17867
rect 14197 17833 14231 17867
rect 17325 17833 17359 17867
rect 21557 17833 21591 17867
rect 22293 17833 22327 17867
rect 24869 17833 24903 17867
rect 28733 17833 28767 17867
rect 29561 17833 29595 17867
rect 30941 17833 30975 17867
rect 33241 17833 33275 17867
rect 33517 17833 33551 17867
rect 37289 17833 37323 17867
rect 37933 17833 37967 17867
rect 5825 17765 5859 17799
rect 7205 17765 7239 17799
rect 8769 17765 8803 17799
rect 10333 17765 10367 17799
rect 14657 17765 14691 17799
rect 21005 17765 21039 17799
rect 21649 17765 21683 17799
rect 30297 17765 30331 17799
rect 30849 17765 30883 17799
rect 31769 17765 31803 17799
rect 31861 17765 31895 17799
rect 38025 17765 38059 17799
rect 1409 17697 1443 17731
rect 4813 17697 4847 17731
rect 5733 17697 5767 17731
rect 6745 17697 6779 17731
rect 6837 17697 6871 17731
rect 12817 17697 12851 17731
rect 13921 17697 13955 17731
rect 15485 17697 15519 17731
rect 15761 17697 15795 17731
rect 18797 17697 18831 17731
rect 19073 17697 19107 17731
rect 21741 17697 21775 17731
rect 21925 17697 21959 17731
rect 23489 17697 23523 17731
rect 27353 17697 27387 17731
rect 31217 17697 31251 17731
rect 31953 17697 31987 17731
rect 38393 17697 38427 17731
rect 1777 17629 1811 17663
rect 3203 17629 3237 17663
rect 4353 17629 4387 17663
rect 5457 17629 5491 17663
rect 5549 17629 5583 17663
rect 5825 17629 5859 17663
rect 6009 17629 6043 17663
rect 6561 17629 6595 17663
rect 7389 17629 7423 17663
rect 9413 17629 9447 17663
rect 9505 17629 9539 17663
rect 9873 17629 9907 17663
rect 9965 17629 9999 17663
rect 10057 17629 10091 17663
rect 10149 17629 10183 17663
rect 10609 17629 10643 17663
rect 10701 17629 10735 17663
rect 12633 17629 12667 17663
rect 13277 17629 13311 17663
rect 14105 17629 14139 17663
rect 14473 17629 14507 17663
rect 14841 17629 14875 17663
rect 19257 17629 19291 17663
rect 19441 17629 19475 17663
rect 20913 17629 20947 17663
rect 21097 17629 21131 17663
rect 21189 17629 21223 17663
rect 21373 17629 21407 17663
rect 21465 17629 21499 17663
rect 22017 17629 22051 17663
rect 22477 17629 22511 17663
rect 22752 17629 22786 17663
rect 22845 17629 22879 17663
rect 23397 17629 23431 17663
rect 23581 17629 23615 17663
rect 24593 17629 24627 17663
rect 24777 17629 24811 17663
rect 25053 17629 25087 17663
rect 25237 17629 25271 17663
rect 25355 17629 25389 17663
rect 25513 17629 25547 17663
rect 27445 17629 27479 17663
rect 28273 17629 28307 17663
rect 28457 17629 28491 17663
rect 28917 17629 28951 17663
rect 29193 17629 29227 17663
rect 29745 17629 29779 17663
rect 29929 17629 29963 17663
rect 30113 17629 30147 17663
rect 30205 17629 30239 17663
rect 30665 17629 30699 17663
rect 31125 17629 31159 17663
rect 31309 17629 31343 17663
rect 31401 17629 31435 17663
rect 31585 17629 31619 17663
rect 31677 17629 31711 17663
rect 33517 17629 33551 17663
rect 33701 17629 33735 17663
rect 34713 17629 34747 17663
rect 37105 17629 37139 17663
rect 37473 17629 37507 17663
rect 37657 17629 37691 17663
rect 37841 17629 37875 17663
rect 41153 17629 41187 17663
rect 4905 17561 4939 17595
rect 7634 17561 7668 17595
rect 9045 17561 9079 17595
rect 10885 17561 10919 17595
rect 13093 17561 13127 17595
rect 20729 17561 20763 17595
rect 24685 17561 24719 17595
rect 25145 17561 25179 17595
rect 27077 17561 27111 17595
rect 29837 17561 29871 17595
rect 30481 17561 30515 17595
rect 32045 17561 32079 17595
rect 32781 17561 32815 17595
rect 34989 17561 35023 17595
rect 37565 17561 37599 17595
rect 41337 17561 41371 17595
rect 4997 17493 5031 17527
rect 6377 17493 6411 17527
rect 7297 17493 7331 17527
rect 9689 17493 9723 17527
rect 12449 17493 12483 17527
rect 15393 17493 15427 17527
rect 17233 17493 17267 17527
rect 19625 17493 19659 17527
rect 25605 17493 25639 17527
rect 27537 17493 27571 17527
rect 28365 17493 28399 17527
rect 29101 17493 29135 17527
rect 36461 17493 36495 17527
rect 36553 17493 36587 17527
rect 40969 17493 41003 17527
rect 1593 17289 1627 17323
rect 5089 17289 5123 17323
rect 5457 17289 5491 17323
rect 5825 17289 5859 17323
rect 7849 17289 7883 17323
rect 9689 17289 9723 17323
rect 13461 17289 13495 17323
rect 15485 17289 15519 17323
rect 17141 17289 17175 17323
rect 18705 17289 18739 17323
rect 20821 17289 20855 17323
rect 21925 17289 21959 17323
rect 23949 17289 23983 17323
rect 25605 17289 25639 17323
rect 27353 17289 27387 17323
rect 32137 17289 32171 17323
rect 32505 17289 32539 17323
rect 32781 17289 32815 17323
rect 34713 17289 34747 17323
rect 35081 17289 35115 17323
rect 38209 17289 38243 17323
rect 40049 17289 40083 17323
rect 6193 17221 6227 17255
rect 9229 17221 9263 17255
rect 9781 17221 9815 17255
rect 14596 17221 14630 17255
rect 14933 17221 14967 17255
rect 15133 17221 15167 17255
rect 18613 17221 18647 17255
rect 19717 17221 19751 17255
rect 19901 17221 19935 17255
rect 20637 17221 20671 17255
rect 21373 17221 21407 17255
rect 23489 17221 23523 17255
rect 23857 17221 23891 17255
rect 25237 17221 25271 17255
rect 25421 17221 25455 17255
rect 27169 17221 27203 17255
rect 28917 17221 28951 17255
rect 32965 17221 32999 17255
rect 35173 17221 35207 17255
rect 39313 17221 39347 17255
rect 39405 17221 39439 17255
rect 40141 17221 40175 17255
rect 40325 17221 40359 17255
rect 40785 17221 40819 17255
rect 1409 17153 1443 17187
rect 2605 17153 2639 17187
rect 4399 17153 4433 17187
rect 4537 17153 4571 17187
rect 4813 17153 4847 17187
rect 5181 17153 5215 17187
rect 5365 17153 5399 17187
rect 5641 17153 5675 17187
rect 6009 17153 6043 17187
rect 6633 17153 6667 17187
rect 8125 17153 8159 17187
rect 8493 17153 8527 17187
rect 8677 17153 8711 17187
rect 9505 17153 9539 17187
rect 12909 17153 12943 17187
rect 15393 17153 15427 17187
rect 15577 17153 15611 17187
rect 17049 17153 17083 17187
rect 17969 17153 18003 17187
rect 18889 17153 18923 17187
rect 18981 17153 19015 17187
rect 19073 17153 19107 17187
rect 19191 17153 19225 17187
rect 19497 17159 19531 17193
rect 19625 17153 19659 17187
rect 20177 17153 20211 17187
rect 20361 17153 20395 17187
rect 20453 17153 20487 17187
rect 21465 17153 21499 17187
rect 21649 17153 21683 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 23673 17153 23707 17187
rect 24133 17153 24167 17187
rect 24409 17153 24443 17187
rect 24593 17153 24627 17187
rect 24777 17153 24811 17187
rect 24961 17153 24995 17187
rect 25145 17153 25179 17187
rect 26433 17153 26467 17187
rect 26985 17153 27019 17187
rect 27721 17153 27755 17187
rect 27905 17153 27939 17187
rect 27997 17153 28031 17187
rect 28181 17153 28215 17187
rect 28457 17153 28491 17187
rect 28733 17153 28767 17187
rect 29469 17153 29503 17187
rect 30941 17153 30975 17187
rect 32321 17153 32355 17187
rect 32597 17153 32631 17187
rect 33149 17153 33183 17187
rect 39175 17153 39209 17187
rect 39497 17153 39531 17187
rect 40049 17153 40083 17187
rect 40601 17153 40635 17187
rect 40877 17153 40911 17187
rect 41797 17153 41831 17187
rect 41981 17153 42015 17187
rect 42165 17153 42199 17187
rect 2973 17085 3007 17119
rect 6377 17085 6411 17119
rect 8033 17085 8067 17119
rect 8217 17085 8251 17119
rect 8309 17085 8343 17119
rect 9321 17085 9355 17119
rect 9928 17085 9962 17119
rect 10149 17085 10183 17119
rect 12633 17085 12667 17119
rect 14841 17085 14875 17119
rect 17325 17085 17359 17119
rect 19349 17085 19383 17119
rect 24317 17085 24351 17119
rect 24685 17085 24719 17119
rect 27813 17085 27847 17119
rect 29193 17085 29227 17119
rect 30849 17085 30883 17119
rect 31401 17085 31435 17119
rect 31861 17085 31895 17119
rect 35357 17085 35391 17119
rect 38025 17085 38059 17119
rect 38117 17085 38151 17119
rect 39037 17085 39071 17119
rect 40417 17085 40451 17119
rect 42073 17085 42107 17119
rect 7757 17017 7791 17051
rect 10057 17017 10091 17051
rect 12357 17017 12391 17051
rect 19993 17017 20027 17051
rect 21097 17017 21131 17051
rect 21557 17017 21591 17051
rect 24225 17017 24259 17051
rect 28273 17017 28307 17051
rect 28365 17017 28399 17051
rect 29101 17017 29135 17051
rect 29377 17017 29411 17051
rect 31309 17017 31343 17051
rect 31585 17017 31619 17051
rect 4905 16949 4939 16983
rect 8585 16949 8619 16983
rect 9413 16949 9447 16983
rect 10425 16949 10459 16983
rect 12817 16949 12851 16983
rect 15117 16949 15151 16983
rect 15301 16949 15335 16983
rect 16681 16949 16715 16983
rect 19901 16949 19935 16983
rect 20177 16949 20211 16983
rect 20913 16949 20947 16983
rect 25789 16949 25823 16983
rect 28641 16949 28675 16983
rect 29285 16949 29319 16983
rect 38577 16949 38611 16983
rect 39681 16949 39715 16983
rect 41245 16949 41279 16983
rect 3801 16745 3835 16779
rect 5365 16745 5399 16779
rect 8769 16745 8803 16779
rect 9505 16745 9539 16779
rect 12817 16745 12851 16779
rect 14105 16745 14139 16779
rect 14565 16745 14599 16779
rect 17141 16745 17175 16779
rect 25145 16745 25179 16779
rect 26341 16745 26375 16779
rect 31861 16745 31895 16779
rect 33241 16745 33275 16779
rect 36921 16745 36955 16779
rect 38761 16745 38795 16779
rect 42165 16745 42199 16779
rect 24041 16677 24075 16711
rect 28641 16677 28675 16711
rect 28733 16677 28767 16711
rect 29653 16677 29687 16711
rect 4353 16609 4387 16643
rect 7021 16609 7055 16643
rect 9965 16609 9999 16643
rect 12449 16609 12483 16643
rect 13737 16609 13771 16643
rect 15301 16609 15335 16643
rect 15577 16609 15611 16643
rect 18521 16609 18555 16643
rect 20821 16609 20855 16643
rect 24685 16609 24719 16643
rect 28365 16609 28399 16643
rect 30021 16609 30055 16643
rect 32229 16609 32263 16643
rect 33149 16609 33183 16643
rect 35449 16609 35483 16643
rect 35725 16609 35759 16643
rect 38393 16609 38427 16643
rect 38669 16609 38703 16643
rect 39313 16609 39347 16643
rect 40417 16609 40451 16643
rect 5089 16541 5123 16575
rect 6929 16541 6963 16575
rect 7389 16541 7423 16575
rect 9505 16541 9539 16575
rect 9873 16541 9907 16575
rect 12541 16541 12575 16575
rect 12909 16541 12943 16575
rect 14249 16541 14283 16575
rect 14381 16541 14415 16575
rect 14565 16541 14599 16575
rect 17785 16541 17819 16575
rect 17877 16541 17911 16575
rect 18797 16541 18831 16575
rect 18981 16541 19015 16575
rect 20913 16541 20947 16575
rect 24593 16541 24627 16575
rect 25053 16541 25087 16575
rect 25237 16541 25271 16575
rect 25789 16541 25823 16575
rect 25973 16541 26007 16575
rect 26157 16541 26191 16575
rect 28273 16541 28307 16575
rect 28893 16541 28927 16575
rect 29101 16541 29135 16575
rect 29285 16541 29319 16575
rect 31309 16541 31343 16575
rect 31401 16541 31435 16575
rect 31677 16541 31711 16575
rect 31769 16541 31803 16575
rect 31953 16541 31987 16575
rect 33241 16541 33275 16575
rect 33425 16541 33459 16575
rect 35357 16541 35391 16575
rect 39865 16541 39899 16575
rect 40233 16541 40267 16575
rect 40325 16541 40359 16575
rect 5181 16473 5215 16507
rect 5365 16473 5399 16507
rect 7634 16473 7668 16507
rect 23765 16473 23799 16507
rect 26065 16473 26099 16507
rect 29009 16473 29043 16507
rect 31493 16473 31527 16507
rect 32965 16473 32999 16507
rect 40693 16473 40727 16507
rect 7297 16405 7331 16439
rect 9321 16405 9355 16439
rect 13093 16405 13127 16439
rect 13185 16405 13219 16439
rect 17049 16405 17083 16439
rect 18797 16405 18831 16439
rect 20545 16405 20579 16439
rect 24225 16405 24259 16439
rect 24961 16405 24995 16439
rect 29561 16405 29595 16439
rect 31125 16405 31159 16439
rect 32781 16405 32815 16439
rect 40141 16405 40175 16439
rect 4399 16201 4433 16235
rect 7941 16201 7975 16235
rect 11345 16201 11379 16235
rect 17049 16201 17083 16235
rect 24225 16201 24259 16235
rect 27353 16201 27387 16235
rect 27445 16201 27479 16235
rect 34529 16201 34563 16235
rect 36369 16201 36403 16235
rect 40049 16201 40083 16235
rect 40785 16201 40819 16235
rect 10977 16133 11011 16167
rect 11177 16133 11211 16167
rect 11774 16133 11808 16167
rect 13093 16133 13127 16167
rect 14412 16133 14446 16167
rect 14841 16133 14875 16167
rect 18731 16133 18765 16167
rect 20453 16133 20487 16167
rect 20545 16133 20579 16167
rect 20913 16133 20947 16167
rect 24685 16133 24719 16167
rect 24777 16133 24811 16167
rect 30481 16133 30515 16167
rect 37565 16133 37599 16167
rect 38577 16133 38611 16167
rect 40325 16133 40359 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 2605 16065 2639 16099
rect 4721 16065 4755 16099
rect 8585 16065 8619 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 14749 16065 14783 16099
rect 14933 16065 14967 16099
rect 17141 16065 17175 16099
rect 18153 16065 18187 16099
rect 18429 16065 18463 16099
rect 18521 16065 18555 16099
rect 18613 16065 18647 16099
rect 19441 16065 19475 16099
rect 19533 16065 19567 16099
rect 19625 16065 19659 16099
rect 19809 16065 19843 16099
rect 19901 16065 19935 16099
rect 20269 16065 20303 16099
rect 20637 16065 20671 16099
rect 24133 16065 24167 16099
rect 24317 16065 24351 16099
rect 24593 16065 24627 16099
rect 24961 16065 24995 16099
rect 28181 16065 28215 16099
rect 28365 16065 28399 16099
rect 30297 16065 30331 16099
rect 30573 16065 30607 16099
rect 30665 16065 30699 16099
rect 32229 16065 32263 16099
rect 34621 16065 34655 16099
rect 37013 16065 37047 16099
rect 37473 16065 37507 16099
rect 37657 16065 37691 16099
rect 37841 16065 37875 16099
rect 40141 16065 40175 16099
rect 40417 16065 40451 16099
rect 40509 16065 40543 16099
rect 41521 16065 41555 16099
rect 2973 15997 3007 16031
rect 4537 15997 4571 16031
rect 11529 15997 11563 16031
rect 14657 15997 14691 16031
rect 17233 15997 17267 16031
rect 17509 15997 17543 16031
rect 18889 15997 18923 16031
rect 21465 15997 21499 16031
rect 27537 15997 27571 16031
rect 27905 15997 27939 16031
rect 31125 15997 31159 16031
rect 32781 15997 32815 16031
rect 33057 15997 33091 16031
rect 34897 15997 34931 16031
rect 38301 15997 38335 16031
rect 41337 15997 41371 16031
rect 41613 15997 41647 16031
rect 13277 15929 13311 15963
rect 20085 15929 20119 15963
rect 24409 15929 24443 15963
rect 30849 15929 30883 15963
rect 40693 15929 40727 15963
rect 1593 15861 1627 15895
rect 1869 15861 1903 15895
rect 4905 15861 4939 15895
rect 11161 15861 11195 15895
rect 12909 15861 12943 15895
rect 16681 15861 16715 15895
rect 18245 15861 18279 15895
rect 19257 15861 19291 15895
rect 20821 15861 20855 15895
rect 26985 15861 27019 15895
rect 28628 15861 28662 15895
rect 30113 15861 30147 15895
rect 31769 15861 31803 15895
rect 36461 15861 36495 15895
rect 37289 15861 37323 15895
rect 41521 15861 41555 15895
rect 41889 15861 41923 15895
rect 3801 15657 3835 15691
rect 11345 15657 11379 15691
rect 11621 15657 11655 15691
rect 13093 15657 13127 15691
rect 17233 15657 17267 15691
rect 17325 15657 17359 15691
rect 19257 15657 19291 15691
rect 19809 15657 19843 15691
rect 27537 15657 27571 15691
rect 28549 15657 28583 15691
rect 32781 15657 32815 15691
rect 33609 15657 33643 15691
rect 35449 15657 35483 15691
rect 40233 15657 40267 15691
rect 12265 15589 12299 15623
rect 15209 15589 15243 15623
rect 28273 15589 28307 15623
rect 32689 15589 32723 15623
rect 1409 15521 1443 15555
rect 5733 15521 5767 15555
rect 6193 15521 6227 15555
rect 10793 15521 10827 15555
rect 11805 15521 11839 15555
rect 13369 15521 13403 15555
rect 13829 15521 13863 15555
rect 19073 15521 19107 15555
rect 20637 15521 20671 15555
rect 22385 15521 22419 15555
rect 23857 15521 23891 15555
rect 25789 15521 25823 15555
rect 27721 15521 27755 15555
rect 33333 15521 33367 15555
rect 34161 15521 34195 15555
rect 37197 15521 37231 15555
rect 40601 15521 40635 15555
rect 41521 15521 41555 15555
rect 42073 15521 42107 15555
rect 1777 15453 1811 15487
rect 3203 15453 3237 15487
rect 4353 15453 4387 15487
rect 5825 15453 5859 15487
rect 6653 15453 6687 15487
rect 6837 15453 6871 15487
rect 8953 15453 8987 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 9597 15453 9631 15487
rect 10977 15453 11011 15487
rect 11069 15453 11103 15487
rect 11897 15453 11931 15487
rect 11989 15453 12023 15487
rect 12081 15453 12115 15487
rect 12909 15453 12943 15487
rect 13001 15453 13035 15487
rect 13461 15453 13495 15487
rect 14105 15453 14139 15487
rect 14749 15453 14783 15487
rect 14841 15453 14875 15487
rect 15025 15453 15059 15487
rect 15485 15453 15519 15487
rect 19625 15453 19659 15487
rect 20361 15453 20395 15487
rect 23673 15453 23707 15487
rect 25421 15453 25455 15487
rect 29193 15453 29227 15487
rect 30205 15453 30239 15487
rect 30481 15453 30515 15487
rect 30665 15453 30699 15487
rect 30849 15453 30883 15487
rect 30941 15453 30975 15487
rect 33977 15453 34011 15487
rect 34805 15453 34839 15487
rect 37473 15453 37507 15487
rect 39037 15453 39071 15487
rect 40417 15453 40451 15487
rect 40785 15453 40819 15487
rect 40969 15453 41003 15487
rect 41153 15453 41187 15487
rect 11329 15385 11363 15419
rect 11529 15385 11563 15419
rect 15761 15385 15795 15419
rect 18797 15385 18831 15419
rect 19441 15385 19475 15419
rect 20913 15385 20947 15419
rect 23765 15385 23799 15419
rect 24869 15385 24903 15419
rect 26065 15385 26099 15419
rect 30573 15385 30607 15419
rect 31217 15385 31251 15419
rect 34069 15385 34103 15419
rect 38301 15385 38335 15419
rect 41061 15385 41095 15419
rect 6745 15317 6779 15351
rect 9505 15317 9539 15351
rect 10793 15317 10827 15351
rect 11161 15317 11195 15351
rect 23305 15317 23339 15351
rect 29561 15317 29595 15351
rect 30297 15317 30331 15351
rect 35725 15317 35759 15351
rect 41337 15317 41371 15351
rect 3203 15113 3237 15147
rect 6101 15113 6135 15147
rect 15025 15113 15059 15147
rect 18061 15113 18095 15147
rect 20637 15113 20671 15147
rect 11253 15045 11287 15079
rect 11774 15045 11808 15079
rect 19533 15045 19567 15079
rect 20269 15045 20303 15079
rect 21833 15045 21867 15079
rect 28825 15045 28859 15079
rect 32137 15045 32171 15079
rect 33885 15045 33919 15079
rect 34437 15045 34471 15079
rect 1409 14977 1443 15011
rect 1777 14977 1811 15011
rect 11161 14977 11195 15011
rect 11345 14977 11379 15011
rect 11529 14977 11563 15011
rect 13912 14977 13946 15011
rect 20085 14977 20119 15011
rect 20361 14977 20395 15011
rect 20453 14977 20487 15011
rect 22385 14977 22419 15011
rect 26709 14977 26743 15011
rect 29193 14977 29227 15011
rect 31401 14977 31435 15011
rect 31585 14977 31619 15011
rect 34253 14977 34287 15011
rect 34529 14977 34563 15011
rect 34621 14977 34655 15011
rect 35449 14977 35483 15011
rect 36001 14977 36035 15011
rect 39497 14977 39531 15011
rect 40509 14977 40543 15011
rect 40785 14977 40819 15011
rect 40969 14977 41003 15011
rect 41613 14977 41647 15011
rect 41797 14977 41831 15011
rect 41981 14977 42015 15011
rect 5549 14909 5583 14943
rect 6377 14909 6411 14943
rect 6653 14909 6687 14943
rect 9689 14909 9723 14943
rect 9965 14909 9999 14943
rect 13645 14909 13679 14943
rect 19809 14909 19843 14943
rect 21281 14909 21315 14943
rect 24593 14909 24627 14943
rect 24869 14909 24903 14943
rect 24961 14909 24995 14943
rect 26433 14909 26467 14943
rect 27353 14909 27387 14943
rect 29101 14909 29135 14943
rect 31125 14909 31159 14943
rect 34897 14909 34931 14943
rect 35909 14909 35943 14943
rect 36461 14909 36495 14943
rect 37105 14909 37139 14943
rect 37749 14909 37783 14943
rect 39221 14909 39255 14943
rect 39589 14909 39623 14943
rect 40141 14909 40175 14943
rect 29653 14841 29687 14875
rect 31861 14841 31895 14875
rect 34805 14841 34839 14875
rect 41797 14841 41831 14875
rect 8125 14773 8159 14807
rect 8217 14773 8251 14807
rect 12909 14773 12943 14807
rect 20729 14773 20763 14807
rect 23121 14773 23155 14807
rect 29377 14773 29411 14807
rect 36277 14773 36311 14807
rect 40325 14773 40359 14807
rect 41061 14773 41095 14807
rect 4997 14569 5031 14603
rect 9873 14569 9907 14603
rect 10333 14569 10367 14603
rect 11529 14569 11563 14603
rect 14933 14569 14967 14603
rect 24133 14569 24167 14603
rect 25053 14569 25087 14603
rect 32689 14569 32723 14603
rect 32781 14569 32815 14603
rect 38209 14569 38243 14603
rect 42165 14569 42199 14603
rect 22201 14501 22235 14535
rect 26249 14501 26283 14535
rect 26709 14501 26743 14535
rect 29561 14501 29595 14535
rect 39957 14501 39991 14535
rect 2237 14433 2271 14467
rect 8401 14433 8435 14467
rect 8677 14433 8711 14467
rect 11897 14433 11931 14467
rect 17233 14433 17267 14467
rect 17417 14433 17451 14467
rect 20729 14433 20763 14467
rect 22385 14433 22419 14467
rect 30941 14433 30975 14467
rect 33241 14433 33275 14467
rect 33425 14433 33459 14467
rect 34529 14433 34563 14467
rect 36185 14433 36219 14467
rect 36369 14433 36403 14467
rect 37105 14433 37139 14467
rect 37565 14433 37599 14467
rect 37749 14433 37783 14467
rect 40141 14433 40175 14467
rect 40693 14433 40727 14467
rect 2145 14365 2179 14399
rect 6745 14365 6779 14399
rect 7573 14365 7607 14399
rect 8585 14365 8619 14399
rect 8769 14365 8803 14399
rect 8953 14365 8987 14399
rect 9505 14365 9539 14399
rect 10149 14365 10183 14399
rect 10333 14365 10367 14399
rect 11713 14365 11747 14399
rect 13001 14365 13035 14399
rect 16681 14365 16715 14399
rect 18521 14365 18555 14399
rect 20453 14365 20487 14399
rect 24409 14365 24443 14399
rect 25697 14365 25731 14399
rect 25973 14365 26007 14399
rect 26433 14365 26467 14399
rect 26709 14365 26743 14399
rect 27169 14365 27203 14399
rect 28273 14365 28307 14399
rect 35265 14365 35299 14399
rect 36093 14365 36127 14399
rect 37013 14365 37047 14399
rect 38393 14365 38427 14399
rect 39865 14365 39899 14399
rect 40417 14365 40451 14399
rect 6469 14297 6503 14331
rect 6837 14297 6871 14331
rect 9715 14297 9749 14331
rect 16405 14297 16439 14331
rect 18153 14297 18187 14331
rect 18889 14297 18923 14331
rect 22661 14297 22695 14331
rect 29009 14297 29043 14331
rect 29745 14297 29779 14331
rect 31217 14297 31251 14331
rect 33149 14297 33183 14331
rect 34713 14297 34747 14331
rect 2513 14229 2547 14263
rect 7849 14229 7883 14263
rect 9889 14229 9923 14263
rect 10057 14229 10091 14263
rect 13645 14229 13679 14263
rect 16773 14229 16807 14263
rect 17141 14229 17175 14263
rect 18797 14229 18831 14263
rect 25145 14229 25179 14263
rect 26525 14229 26559 14263
rect 33885 14229 33919 14263
rect 35725 14229 35759 14263
rect 36553 14229 36587 14263
rect 36921 14229 36955 14263
rect 37841 14229 37875 14263
rect 40141 14229 40175 14263
rect 6738 14025 6772 14059
rect 7849 14025 7883 14059
rect 12626 14025 12660 14059
rect 18613 14025 18647 14059
rect 18981 14025 19015 14059
rect 21005 14025 21039 14059
rect 22293 14025 22327 14059
rect 24409 14025 24443 14059
rect 28733 14025 28767 14059
rect 30573 14025 30607 14059
rect 33425 14025 33459 14059
rect 33517 14025 33551 14059
rect 34253 14025 34287 14059
rect 34345 14025 34379 14059
rect 37013 14025 37047 14059
rect 39313 14025 39347 14059
rect 41429 14025 41463 14059
rect 2697 13957 2731 13991
rect 4445 13957 4479 13991
rect 6837 13957 6871 13991
rect 10333 13957 10367 13991
rect 20545 13957 20579 13991
rect 21281 13957 21315 13991
rect 24777 13957 24811 13991
rect 25605 13957 25639 13991
rect 27261 13957 27295 13991
rect 31125 13957 31159 13991
rect 31493 13957 31527 13991
rect 35541 13957 35575 13991
rect 5365 13889 5399 13923
rect 5549 13889 5583 13923
rect 6009 13889 6043 13923
rect 6561 13889 6595 13923
rect 6653 13889 6687 13923
rect 7573 13889 7607 13923
rect 7665 13889 7699 13923
rect 7941 13889 7975 13923
rect 10517 13889 10551 13923
rect 12449 13889 12483 13923
rect 12541 13889 12575 13923
rect 12725 13889 12759 13923
rect 12817 13889 12851 13923
rect 13553 13889 13587 13923
rect 13737 13889 13771 13923
rect 15301 13889 15335 13923
rect 15577 13889 15611 13923
rect 15761 13889 15795 13923
rect 18797 13889 18831 13923
rect 19349 13889 19383 13923
rect 19809 13889 19843 13923
rect 20821 13889 20855 13923
rect 21649 13889 21683 13923
rect 22201 13889 22235 13923
rect 22661 13889 22695 13923
rect 24593 13889 24627 13923
rect 24685 13889 24719 13923
rect 24961 13889 24995 13923
rect 25881 13889 25915 13923
rect 26157 13889 26191 13923
rect 26341 13889 26375 13923
rect 26433 13889 26467 13923
rect 26525 13889 26559 13923
rect 26985 13889 27019 13923
rect 28825 13889 28859 13923
rect 30757 13889 30791 13923
rect 31861 13889 31895 13923
rect 34713 13889 34747 13923
rect 34989 13889 35023 13923
rect 42073 13889 42107 13923
rect 2421 13821 2455 13855
rect 6929 13821 6963 13855
rect 10241 13821 10275 13855
rect 13369 13821 13403 13855
rect 15117 13821 15151 13855
rect 15853 13821 15887 13855
rect 16497 13821 16531 13855
rect 16681 13821 16715 13855
rect 16957 13821 16991 13855
rect 19441 13821 19475 13855
rect 19625 13821 19659 13855
rect 20361 13821 20395 13855
rect 20729 13821 20763 13855
rect 22477 13821 22511 13855
rect 23213 13821 23247 13855
rect 25697 13821 25731 13855
rect 32413 13821 32447 13855
rect 33701 13821 33735 13855
rect 34529 13821 34563 13855
rect 34805 13821 34839 13855
rect 35265 13821 35299 13855
rect 37565 13821 37599 13855
rect 37841 13821 37875 13855
rect 39681 13821 39715 13855
rect 39957 13821 39991 13855
rect 41521 13821 41555 13855
rect 5733 13753 5767 13787
rect 7665 13753 7699 13787
rect 33057 13753 33091 13787
rect 5365 13685 5399 13719
rect 9597 13685 9631 13719
rect 13737 13685 13771 13719
rect 18429 13685 18463 13719
rect 20637 13685 20671 13719
rect 21833 13685 21867 13719
rect 25697 13685 25731 13719
rect 26065 13685 26099 13719
rect 26709 13685 26743 13719
rect 29082 13685 29116 13719
rect 32965 13685 32999 13719
rect 33885 13685 33919 13719
rect 34897 13685 34931 13719
rect 35173 13685 35207 13719
rect 5549 13481 5583 13515
rect 5733 13481 5767 13515
rect 7113 13481 7147 13515
rect 7849 13481 7883 13515
rect 8769 13481 8803 13515
rect 9210 13481 9244 13515
rect 10701 13481 10735 13515
rect 17095 13481 17129 13515
rect 23029 13481 23063 13515
rect 26341 13481 26375 13515
rect 26525 13481 26559 13515
rect 28641 13481 28675 13515
rect 34713 13481 34747 13515
rect 34989 13481 35023 13515
rect 37197 13481 37231 13515
rect 38301 13481 38335 13515
rect 39865 13481 39899 13515
rect 26249 13413 26283 13447
rect 30205 13413 30239 13447
rect 34345 13413 34379 13447
rect 41981 13413 42015 13447
rect 3249 13345 3283 13379
rect 3525 13345 3559 13379
rect 3801 13345 3835 13379
rect 6193 13345 6227 13379
rect 7205 13345 7239 13379
rect 8493 13345 8527 13379
rect 11069 13345 11103 13379
rect 13921 13345 13955 13379
rect 15301 13345 15335 13379
rect 17969 13345 18003 13379
rect 18705 13345 18739 13379
rect 18889 13345 18923 13379
rect 21281 13345 21315 13379
rect 21557 13345 21591 13379
rect 26065 13345 26099 13379
rect 30757 13345 30791 13379
rect 32505 13345 32539 13379
rect 32873 13345 32907 13379
rect 35081 13345 35115 13379
rect 35357 13345 35391 13379
rect 35633 13345 35667 13379
rect 38853 13345 38887 13379
rect 3433 13277 3467 13311
rect 3617 13277 3651 13311
rect 6101 13277 6135 13311
rect 6929 13277 6963 13311
rect 7389 13277 7423 13311
rect 8401 13277 8435 13311
rect 8953 13277 8987 13311
rect 13654 13277 13688 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15669 13277 15703 13311
rect 19441 13277 19475 13311
rect 25053 13277 25087 13311
rect 26341 13277 26375 13311
rect 26433 13277 26467 13311
rect 28181 13277 28215 13311
rect 28825 13277 28859 13311
rect 29101 13277 29135 13311
rect 29653 13277 29687 13311
rect 30021 13277 30055 13311
rect 32597 13277 32631 13311
rect 34897 13277 34931 13311
rect 37749 13277 37783 13311
rect 38669 13277 38703 13311
rect 40049 13277 40083 13311
rect 40233 13277 40267 13311
rect 40351 13277 40385 13311
rect 40509 13277 40543 13311
rect 41797 13277 41831 13311
rect 2973 13209 3007 13243
rect 4077 13209 4111 13243
rect 7113 13209 7147 13243
rect 7817 13209 7851 13243
rect 8033 13209 8067 13243
rect 11336 13209 11370 13243
rect 17233 13209 17267 13243
rect 19717 13209 19751 13243
rect 30481 13209 30515 13243
rect 31033 13209 31067 13243
rect 35173 13209 35207 13243
rect 38761 13209 38795 13243
rect 40141 13209 40175 13243
rect 1501 13141 1535 13175
rect 7573 13141 7607 13175
rect 7665 13141 7699 13175
rect 12449 13141 12483 13175
rect 12541 13141 12575 13175
rect 14473 13141 14507 13175
rect 18245 13141 18279 13175
rect 18613 13141 18647 13175
rect 21189 13141 21223 13175
rect 24501 13141 24535 13175
rect 27629 13141 27663 13175
rect 29009 13141 29043 13175
rect 37105 13141 37139 13175
rect 2513 12937 2547 12971
rect 2789 12937 2823 12971
rect 3794 12937 3828 12971
rect 6193 12937 6227 12971
rect 6837 12937 6871 12971
rect 10977 12937 11011 12971
rect 11145 12937 11179 12971
rect 13185 12937 13219 12971
rect 14013 12937 14047 12971
rect 17049 12937 17083 12971
rect 17417 12937 17451 12971
rect 17785 12937 17819 12971
rect 20637 12937 20671 12971
rect 21097 12937 21131 12971
rect 22753 12937 22787 12971
rect 24041 12937 24075 12971
rect 24133 12937 24167 12971
rect 25053 12937 25087 12971
rect 32137 12937 32171 12971
rect 32505 12937 32539 12971
rect 35173 12937 35207 12971
rect 35357 12937 35391 12971
rect 2329 12869 2363 12903
rect 3893 12869 3927 12903
rect 4721 12869 4755 12903
rect 6545 12869 6579 12903
rect 6745 12869 6779 12903
rect 11345 12869 11379 12903
rect 14473 12869 14507 12903
rect 22661 12869 22695 12903
rect 27445 12869 27479 12903
rect 33333 12869 33367 12903
rect 35725 12869 35759 12903
rect 37933 12869 37967 12903
rect 38301 12869 38335 12903
rect 1685 12801 1719 12835
rect 2605 12801 2639 12835
rect 2697 12801 2731 12835
rect 2881 12801 2915 12835
rect 3617 12801 3651 12835
rect 3709 12801 3743 12835
rect 8125 12801 8159 12835
rect 9965 12801 9999 12835
rect 10149 12801 10183 12835
rect 11897 12801 11931 12835
rect 12265 12801 12299 12835
rect 13001 12801 13035 12835
rect 13185 12801 13219 12835
rect 13277 12801 13311 12835
rect 13829 12801 13863 12835
rect 14197 12801 14231 12835
rect 16865 12801 16899 12835
rect 17417 12801 17451 12835
rect 17601 12801 17635 12835
rect 18061 12801 18095 12835
rect 20085 12801 20119 12835
rect 20269 12801 20303 12835
rect 21005 12801 21039 12835
rect 21833 12801 21867 12835
rect 23581 12801 23615 12835
rect 24961 12801 24995 12835
rect 25605 12801 25639 12835
rect 27169 12801 27203 12835
rect 29469 12801 29503 12835
rect 30579 12801 30613 12835
rect 30757 12801 30791 12835
rect 32597 12801 32631 12835
rect 34989 12801 35023 12835
rect 35541 12801 35575 12835
rect 35817 12801 35851 12835
rect 37473 12801 37507 12835
rect 37565 12801 37599 12835
rect 37841 12801 37875 12835
rect 38485 12801 38519 12835
rect 4445 12733 4479 12767
rect 7389 12733 7423 12767
rect 8401 12733 8435 12767
rect 10057 12733 10091 12767
rect 10793 12733 10827 12767
rect 11529 12733 11563 12767
rect 11989 12733 12023 12767
rect 12817 12733 12851 12767
rect 14289 12733 14323 12767
rect 14565 12733 14599 12767
rect 16681 12733 16715 12767
rect 18245 12733 18279 12767
rect 18521 12733 18555 12767
rect 19993 12733 20027 12767
rect 21281 12733 21315 12767
rect 22477 12733 22511 12767
rect 24317 12733 24351 12767
rect 25237 12733 25271 12767
rect 26249 12733 26283 12767
rect 29653 12733 29687 12767
rect 29929 12733 29963 12767
rect 30849 12733 30883 12767
rect 32689 12733 32723 12767
rect 33057 12733 33091 12767
rect 36553 12733 36587 12767
rect 2329 12665 2363 12699
rect 6377 12665 6411 12699
rect 23397 12665 23431 12699
rect 34805 12665 34839 12699
rect 38669 12665 38703 12699
rect 1501 12597 1535 12631
rect 6561 12597 6595 12631
rect 9873 12597 9907 12631
rect 10241 12597 10275 12631
rect 11161 12597 11195 12631
rect 14197 12597 14231 12631
rect 15209 12597 15243 12631
rect 20085 12597 20119 12631
rect 23673 12597 23707 12631
rect 24593 12597 24627 12631
rect 28917 12597 28951 12631
rect 29377 12597 29411 12631
rect 30573 12597 30607 12631
rect 31493 12597 31527 12631
rect 37289 12597 37323 12631
rect 37749 12597 37783 12631
rect 1777 12393 1811 12427
rect 1961 12393 1995 12427
rect 4537 12393 4571 12427
rect 4721 12393 4755 12427
rect 7481 12393 7515 12427
rect 10241 12393 10275 12427
rect 11713 12393 11747 12427
rect 24672 12393 24706 12427
rect 26157 12393 26191 12427
rect 27721 12393 27755 12427
rect 31309 12393 31343 12427
rect 14105 12325 14139 12359
rect 39129 12325 39163 12359
rect 5733 12257 5767 12291
rect 6009 12257 6043 12291
rect 10609 12257 10643 12291
rect 10885 12257 10919 12291
rect 13921 12257 13955 12291
rect 19257 12257 19291 12291
rect 19809 12257 19843 12291
rect 20545 12257 20579 12291
rect 23397 12257 23431 12291
rect 26709 12257 26743 12291
rect 26801 12257 26835 12291
rect 28273 12257 28307 12291
rect 29561 12257 29595 12291
rect 29837 12257 29871 12291
rect 31953 12257 31987 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 9505 12189 9539 12223
rect 9965 12189 9999 12223
rect 10241 12189 10275 12223
rect 10517 12189 10551 12223
rect 13001 12189 13035 12223
rect 15485 12189 15519 12223
rect 17233 12189 17267 12223
rect 20637 12189 20671 12223
rect 21097 12189 21131 12223
rect 21373 12189 21407 12223
rect 21465 12189 21499 12223
rect 21925 12189 21959 12223
rect 22109 12189 22143 12223
rect 22201 12189 22235 12223
rect 23121 12189 23155 12223
rect 23305 12189 23339 12223
rect 23489 12189 23523 12223
rect 23673 12189 23707 12223
rect 24409 12189 24443 12223
rect 28181 12189 28215 12223
rect 29101 12189 29135 12223
rect 31769 12189 31803 12223
rect 31861 12189 31895 12223
rect 35449 12189 35483 12223
rect 36001 12189 36035 12223
rect 37289 12189 37323 12223
rect 39497 12189 39531 12223
rect 39681 12189 39715 12223
rect 2421 12121 2455 12155
rect 4905 12121 4939 12155
rect 9873 12121 9907 12155
rect 15218 12121 15252 12155
rect 17509 12121 17543 12155
rect 19993 12121 20027 12155
rect 20177 12121 20211 12155
rect 21281 12121 21315 12155
rect 28089 12121 28123 12155
rect 28549 12121 28583 12155
rect 37565 12121 37599 12155
rect 39313 12121 39347 12155
rect 39589 12121 39623 12155
rect 4705 12053 4739 12087
rect 9321 12053 9355 12087
rect 9597 12053 9631 12087
rect 9689 12053 9723 12087
rect 10057 12053 10091 12087
rect 13277 12053 13311 12087
rect 18981 12053 19015 12087
rect 20361 12053 20395 12087
rect 21649 12053 21683 12087
rect 21741 12053 21775 12087
rect 23857 12053 23891 12087
rect 26249 12053 26283 12087
rect 26617 12053 26651 12087
rect 31401 12053 31435 12087
rect 34897 12053 34931 12087
rect 39037 12053 39071 12087
rect 1777 11849 1811 11883
rect 3525 11849 3559 11883
rect 3985 11849 4019 11883
rect 5089 11849 5123 11883
rect 10517 11849 10551 11883
rect 12925 11849 12959 11883
rect 13093 11849 13127 11883
rect 13277 11849 13311 11883
rect 18889 11849 18923 11883
rect 20913 11849 20947 11883
rect 22477 11849 22511 11883
rect 26801 11849 26835 11883
rect 27997 11849 28031 11883
rect 28549 11849 28583 11883
rect 36277 11849 36311 11883
rect 5181 11781 5215 11815
rect 6653 11781 6687 11815
rect 9597 11781 9631 11815
rect 11529 11781 11563 11815
rect 12725 11781 12759 11815
rect 14390 11781 14424 11815
rect 19763 11781 19797 11815
rect 19993 11781 20027 11815
rect 20545 11781 20579 11815
rect 20761 11781 20795 11815
rect 22201 11781 22235 11815
rect 23305 11781 23339 11815
rect 25237 11781 25271 11815
rect 25789 11781 25823 11815
rect 25973 11781 26007 11815
rect 26433 11781 26467 11815
rect 27169 11781 27203 11815
rect 28917 11781 28951 11815
rect 31309 11781 31343 11815
rect 32413 11781 32447 11815
rect 34805 11781 34839 11815
rect 1685 11713 1719 11747
rect 1961 11713 1995 11747
rect 2329 11713 2363 11747
rect 2421 11713 2455 11747
rect 3157 11713 3191 11747
rect 3341 11713 3375 11747
rect 3801 11713 3835 11747
rect 4445 11713 4479 11747
rect 4629 11713 4663 11747
rect 4721 11713 4755 11747
rect 4905 11713 4939 11747
rect 5457 11713 5491 11747
rect 6929 11713 6963 11747
rect 7205 11713 7239 11747
rect 7389 11713 7423 11747
rect 9873 11713 9907 11747
rect 19533 11713 19567 11747
rect 19625 11713 19659 11747
rect 19901 11713 19935 11747
rect 20085 11713 20119 11747
rect 21833 11713 21867 11747
rect 21926 11713 21960 11747
rect 22109 11713 22143 11747
rect 22339 11713 22373 11747
rect 24869 11713 24903 11747
rect 24962 11713 24996 11747
rect 25145 11713 25179 11747
rect 25375 11713 25409 11747
rect 25605 11713 25639 11747
rect 26249 11713 26283 11747
rect 26525 11713 26559 11747
rect 26617 11713 26651 11747
rect 27905 11713 27939 11747
rect 28181 11713 28215 11747
rect 28733 11713 28767 11747
rect 28825 11713 28859 11747
rect 29101 11713 29135 11747
rect 32321 11713 32355 11747
rect 32505 11713 32539 11747
rect 32689 11713 32723 11747
rect 33977 11713 34011 11747
rect 34069 11713 34103 11747
rect 34253 11713 34287 11747
rect 36921 11713 36955 11747
rect 37841 11713 37875 11747
rect 40141 11713 40175 11747
rect 3617 11645 3651 11679
rect 4077 11645 4111 11679
rect 5365 11645 5399 11679
rect 6745 11645 6779 11679
rect 9689 11645 9723 11679
rect 11069 11645 11103 11679
rect 14657 11645 14691 11679
rect 21557 11645 21591 11679
rect 23029 11645 23063 11679
rect 24777 11645 24811 11679
rect 27721 11645 27755 11679
rect 31585 11645 31619 11679
rect 34529 11645 34563 11679
rect 37749 11645 37783 11679
rect 38117 11645 38151 11679
rect 38209 11645 38243 11679
rect 39865 11645 39899 11679
rect 40233 11645 40267 11679
rect 40785 11645 40819 11679
rect 4169 11577 4203 11611
rect 4813 11577 4847 11611
rect 20269 11577 20303 11611
rect 25513 11577 25547 11611
rect 37565 11577 37599 11611
rect 1501 11509 1535 11543
rect 2053 11509 2087 11543
rect 4261 11509 4295 11543
rect 4445 11509 4479 11543
rect 5181 11509 5215 11543
rect 5641 11509 5675 11543
rect 6929 11509 6963 11543
rect 7113 11509 7147 11543
rect 7205 11509 7239 11543
rect 9689 11509 9723 11543
rect 10057 11509 10091 11543
rect 12909 11509 12943 11543
rect 20729 11509 20763 11543
rect 21005 11509 21039 11543
rect 28365 11509 28399 11543
rect 29837 11509 29871 11543
rect 32137 11509 32171 11543
rect 34437 11509 34471 11543
rect 36369 11509 36403 11543
rect 38393 11509 38427 11543
rect 2329 11305 2363 11339
rect 5365 11305 5399 11339
rect 6377 11305 6411 11339
rect 10149 11305 10183 11339
rect 13185 11305 13219 11339
rect 18521 11305 18555 11339
rect 21373 11305 21407 11339
rect 21465 11305 21499 11339
rect 27537 11305 27571 11339
rect 28273 11305 28307 11339
rect 32413 11305 32447 11339
rect 34437 11305 34471 11339
rect 34989 11305 35023 11339
rect 36277 11305 36311 11339
rect 37841 11305 37875 11339
rect 38945 11305 38979 11339
rect 1777 11237 1811 11271
rect 2513 11237 2547 11271
rect 2973 11237 3007 11271
rect 4077 11237 4111 11271
rect 5549 11237 5583 11271
rect 7389 11237 7423 11271
rect 9505 11237 9539 11271
rect 9597 11237 9631 11271
rect 13921 11237 13955 11271
rect 33425 11237 33459 11271
rect 37749 11237 37783 11271
rect 2053 11169 2087 11203
rect 3157 11169 3191 11203
rect 6653 11169 6687 11203
rect 6837 11169 6871 11203
rect 7481 11169 7515 11203
rect 10517 11169 10551 11203
rect 12265 11169 12299 11203
rect 13461 11169 13495 11203
rect 18889 11169 18923 11203
rect 19625 11169 19659 11203
rect 22937 11169 22971 11203
rect 26065 11169 26099 11203
rect 27813 11169 27847 11203
rect 31401 11169 31435 11203
rect 33977 11169 34011 11203
rect 35449 11169 35483 11203
rect 35541 11169 35575 11203
rect 38117 11169 38151 11203
rect 39497 11169 39531 11203
rect 1685 11101 1719 11135
rect 1961 11101 1995 11135
rect 2421 11101 2455 11135
rect 2513 11101 2547 11135
rect 2789 11101 2823 11135
rect 3249 11101 3283 11135
rect 3893 11101 3927 11135
rect 6561 11101 6595 11135
rect 6745 11101 6779 11135
rect 7297 11101 7331 11135
rect 7573 11101 7607 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 9781 11101 9815 11135
rect 9873 11101 9907 11135
rect 12817 11101 12851 11135
rect 13553 11101 13587 11135
rect 18797 11101 18831 11135
rect 23213 11101 23247 11135
rect 24777 11101 24811 11135
rect 25789 11101 25823 11135
rect 27721 11101 27755 11135
rect 27997 11101 28031 11135
rect 28089 11101 28123 11135
rect 31309 11101 31343 11135
rect 31585 11101 31619 11135
rect 31677 11101 31711 11135
rect 31861 11101 31895 11135
rect 31953 11101 31987 11135
rect 32229 11101 32263 11135
rect 33241 11101 33275 11135
rect 33885 11101 33919 11135
rect 34161 11101 34195 11135
rect 34253 11101 34287 11135
rect 35357 11101 35391 11135
rect 36277 11101 36311 11135
rect 36553 11101 36587 11135
rect 36829 11101 36863 11135
rect 37105 11101 37139 11135
rect 37197 11101 37231 11135
rect 37473 11101 37507 11135
rect 37565 11101 37599 11135
rect 38209 11101 38243 11135
rect 3525 11033 3559 11067
rect 3617 11033 3651 11067
rect 5181 11033 5215 11067
rect 10117 11033 10151 11067
rect 10333 11033 10367 11067
rect 11989 11033 12023 11067
rect 13001 11033 13035 11067
rect 19901 11033 19935 11067
rect 32045 11033 32079 11067
rect 37381 11033 37415 11067
rect 1501 10965 1535 10999
rect 2697 10965 2731 10999
rect 5391 10965 5425 10999
rect 7757 10965 7791 10999
rect 7941 10965 7975 10999
rect 9965 10965 9999 10999
rect 3157 10761 3191 10795
rect 5825 10761 5859 10795
rect 6101 10761 6135 10795
rect 8493 10761 8527 10795
rect 18705 10761 18739 10795
rect 20637 10761 20671 10795
rect 20913 10761 20947 10795
rect 22569 10761 22603 10795
rect 23121 10761 23155 10795
rect 28089 10761 28123 10795
rect 29469 10761 29503 10795
rect 37473 10761 37507 10795
rect 38853 10761 38887 10795
rect 1685 10693 1719 10727
rect 5365 10693 5399 10727
rect 6745 10693 6779 10727
rect 6929 10693 6963 10727
rect 9965 10693 9999 10727
rect 10501 10693 10535 10727
rect 10701 10693 10735 10727
rect 20821 10693 20855 10727
rect 24869 10693 24903 10727
rect 25605 10693 25639 10727
rect 36001 10693 36035 10727
rect 36093 10693 36127 10727
rect 4169 10625 4203 10659
rect 7573 10625 7607 10659
rect 20453 10625 20487 10659
rect 20545 10625 20579 10659
rect 21097 10625 21131 10659
rect 21189 10625 21223 10659
rect 21281 10625 21315 10659
rect 21465 10625 21499 10659
rect 21833 10625 21867 10659
rect 22385 10625 22419 10659
rect 22753 10625 22787 10659
rect 22937 10625 22971 10659
rect 23029 10625 23063 10659
rect 23213 10625 23247 10659
rect 24225 10625 24259 10659
rect 24501 10625 24535 10659
rect 26341 10625 26375 10659
rect 27169 10625 27203 10659
rect 27261 10625 27295 10659
rect 27353 10625 27387 10659
rect 27537 10625 27571 10659
rect 28457 10625 28491 10659
rect 28917 10625 28951 10659
rect 29009 10625 29043 10659
rect 29101 10625 29135 10659
rect 29285 10625 29319 10659
rect 29653 10625 29687 10659
rect 30389 10625 30423 10659
rect 35725 10625 35759 10659
rect 35817 10625 35851 10659
rect 36185 10625 36219 10659
rect 37289 10625 37323 10659
rect 37473 10625 37507 10659
rect 37657 10625 37691 10659
rect 37841 10625 37875 10659
rect 37933 10625 37967 10659
rect 38025 10625 38059 10659
rect 38301 10625 38335 10659
rect 38485 10625 38519 10659
rect 38577 10625 38611 10659
rect 38669 10625 38703 10659
rect 39589 10625 39623 10659
rect 1409 10557 1443 10591
rect 5917 10557 5951 10591
rect 7481 10557 7515 10591
rect 7849 10557 7883 10591
rect 7941 10557 7975 10591
rect 10241 10557 10275 10591
rect 12909 10557 12943 10591
rect 13553 10557 13587 10591
rect 16865 10557 16899 10591
rect 17141 10557 17175 10591
rect 20177 10557 20211 10591
rect 24133 10557 24167 10591
rect 24593 10557 24627 10591
rect 25697 10557 25731 10591
rect 28365 10557 28399 10591
rect 29837 10557 29871 10591
rect 32137 10557 32171 10591
rect 32413 10557 32447 10591
rect 35449 10557 35483 10591
rect 5365 10489 5399 10523
rect 13001 10489 13035 10523
rect 38209 10489 38243 10523
rect 6561 10421 6595 10455
rect 7297 10421 7331 10455
rect 10333 10421 10367 10455
rect 10517 10421 10551 10455
rect 12265 10421 12299 10455
rect 18613 10421 18647 10455
rect 20821 10421 20855 10455
rect 22753 10421 22787 10455
rect 23949 10421 23983 10455
rect 26985 10421 27019 10455
rect 28733 10421 28767 10455
rect 33885 10421 33919 10455
rect 33977 10421 34011 10455
rect 36369 10421 36403 10455
rect 39497 10421 39531 10455
rect 3341 10217 3375 10251
rect 6009 10217 6043 10251
rect 6193 10217 6227 10251
rect 7665 10217 7699 10251
rect 9873 10217 9907 10251
rect 10425 10217 10459 10251
rect 10701 10217 10735 10251
rect 13369 10217 13403 10251
rect 18337 10217 18371 10251
rect 19993 10217 20027 10251
rect 22017 10217 22051 10251
rect 23305 10217 23339 10251
rect 24225 10217 24259 10251
rect 24869 10217 24903 10251
rect 26359 10217 26393 10251
rect 30665 10217 30699 10251
rect 32137 10217 32171 10251
rect 39865 10217 39899 10251
rect 9965 10149 9999 10183
rect 10885 10149 10919 10183
rect 29561 10149 29595 10183
rect 31217 10149 31251 10183
rect 34345 10149 34379 10183
rect 37197 10149 37231 10183
rect 6929 10081 6963 10115
rect 9229 10081 9263 10115
rect 9505 10081 9539 10115
rect 9597 10081 9631 10115
rect 9714 10081 9748 10115
rect 10333 10081 10367 10115
rect 11253 10081 11287 10115
rect 11529 10081 11563 10115
rect 11897 10081 11931 10115
rect 18521 10081 18555 10115
rect 19349 10081 19383 10115
rect 23121 10081 23155 10115
rect 23949 10081 23983 10115
rect 26617 10081 26651 10115
rect 27169 10081 27203 10115
rect 28917 10081 28951 10115
rect 30113 10081 30147 10115
rect 32321 10081 32355 10115
rect 33885 10081 33919 10115
rect 36921 10081 36955 10115
rect 37841 10081 37875 10115
rect 38485 10081 38519 10115
rect 40509 10081 40543 10115
rect 3249 10013 3283 10047
rect 4721 10013 4755 10047
rect 5549 10013 5583 10047
rect 6193 10013 6227 10047
rect 6377 10013 6411 10047
rect 7021 10013 7055 10047
rect 7941 10013 7975 10047
rect 8125 10013 8159 10047
rect 10149 10013 10183 10047
rect 10425 10013 10459 10047
rect 11161 10013 11195 10047
rect 11621 10013 11655 10047
rect 18613 10013 18647 10047
rect 18889 10013 18923 10047
rect 19901 10013 19935 10047
rect 20177 10013 20211 10047
rect 20269 10013 20303 10047
rect 20545 10013 20579 10047
rect 22201 10013 22235 10047
rect 22753 10013 22787 10047
rect 22937 10013 22971 10047
rect 23489 10013 23523 10047
rect 23857 10013 23891 10047
rect 29285 10013 29319 10047
rect 30941 10013 30975 10047
rect 31033 10013 31067 10047
rect 31585 10013 31619 10047
rect 31769 10013 31803 10047
rect 32413 10013 32447 10047
rect 32689 10013 32723 10047
rect 33333 10013 33367 10047
rect 34069 10013 34103 10047
rect 36829 10013 36863 10047
rect 37473 10013 37507 10047
rect 37565 10013 37599 10047
rect 39037 10013 39071 10047
rect 40601 10013 40635 10047
rect 3985 9945 4019 9979
rect 6653 9945 6687 9979
rect 7644 9945 7678 9979
rect 7849 9945 7883 9979
rect 10517 9945 10551 9979
rect 18981 9945 19015 9979
rect 20361 9945 20395 9979
rect 27445 9945 27479 9979
rect 30481 9945 30515 9979
rect 31217 9945 31251 9979
rect 32781 9945 32815 9979
rect 34345 9945 34379 9979
rect 37933 9945 37967 9979
rect 39313 9945 39347 9979
rect 4997 9877 5031 9911
rect 6745 9877 6779 9911
rect 7389 9877 7423 9911
rect 7481 9877 7515 9911
rect 8033 9877 8067 9911
rect 10717 9877 10751 9911
rect 29101 9877 29135 9911
rect 30681 9877 30715 9911
rect 30849 9877 30883 9911
rect 31677 9877 31711 9911
rect 34161 9877 34195 9911
rect 37289 9877 37323 9911
rect 39405 9877 39439 9911
rect 40785 9877 40819 9911
rect 4905 9673 4939 9707
rect 5825 9673 5859 9707
rect 7113 9673 7147 9707
rect 13277 9673 13311 9707
rect 25145 9673 25179 9707
rect 27169 9673 27203 9707
rect 27905 9673 27939 9707
rect 30389 9673 30423 9707
rect 34453 9673 34487 9707
rect 35909 9673 35943 9707
rect 36461 9673 36495 9707
rect 39037 9673 39071 9707
rect 40877 9673 40911 9707
rect 6009 9605 6043 9639
rect 7573 9605 7607 9639
rect 10701 9605 10735 9639
rect 23673 9605 23707 9639
rect 26985 9605 27019 9639
rect 27353 9605 27387 9639
rect 28457 9605 28491 9639
rect 28917 9605 28951 9639
rect 30665 9605 30699 9639
rect 31677 9605 31711 9639
rect 32137 9605 32171 9639
rect 32321 9605 32355 9639
rect 34253 9605 34287 9639
rect 34713 9605 34747 9639
rect 37565 9605 37599 9639
rect 39405 9605 39439 9639
rect 2881 9537 2915 9571
rect 4846 9537 4880 9571
rect 5273 9537 5307 9571
rect 5641 9537 5675 9571
rect 5733 9537 5767 9571
rect 6745 9537 6779 9571
rect 7481 9537 7515 9571
rect 7757 9537 7791 9571
rect 10057 9537 10091 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 10609 9537 10643 9571
rect 22753 9537 22787 9571
rect 26524 9537 26558 9571
rect 27261 9537 27295 9571
rect 28181 9537 28215 9571
rect 31401 9537 31435 9571
rect 31493 9537 31527 9571
rect 32965 9537 32999 9571
rect 33149 9537 33183 9571
rect 33241 9537 33275 9571
rect 33333 9537 33367 9571
rect 33977 9537 34011 9571
rect 34897 9537 34931 9571
rect 35541 9537 35575 9571
rect 36277 9537 36311 9571
rect 37289 9537 37323 9571
rect 3157 9469 3191 9503
rect 5365 9469 5399 9503
rect 5457 9469 5491 9503
rect 6561 9469 6595 9503
rect 6653 9469 6687 9503
rect 9965 9469 9999 9503
rect 11253 9469 11287 9503
rect 11529 9469 11563 9503
rect 11805 9469 11839 9503
rect 21833 9469 21867 9503
rect 22845 9469 22879 9503
rect 23397 9469 23431 9503
rect 26249 9469 26283 9503
rect 26340 9469 26374 9503
rect 26433 9469 26467 9503
rect 28089 9469 28123 9503
rect 28549 9469 28583 9503
rect 28641 9469 28675 9503
rect 31861 9469 31895 9503
rect 33885 9469 33919 9503
rect 35633 9469 35667 9503
rect 36093 9469 36127 9503
rect 39129 9469 39163 9503
rect 4721 9401 4755 9435
rect 10609 9401 10643 9435
rect 33517 9401 33551 9435
rect 34621 9401 34655 9435
rect 4629 9333 4663 9367
rect 7665 9333 7699 9367
rect 9689 9333 9723 9367
rect 22477 9333 22511 9367
rect 23029 9333 23063 9367
rect 26709 9333 26743 9367
rect 27537 9333 27571 9367
rect 32505 9333 32539 9367
rect 33701 9333 33735 9367
rect 34437 9333 34471 9367
rect 35081 9333 35115 9367
rect 5457 9129 5491 9163
rect 5641 9129 5675 9163
rect 6101 9129 6135 9163
rect 11161 9129 11195 9163
rect 11437 9129 11471 9163
rect 20913 9129 20947 9163
rect 22937 9129 22971 9163
rect 23581 9129 23615 9163
rect 24501 9129 24535 9163
rect 32505 9129 32539 9163
rect 33701 9129 33735 9163
rect 9413 8993 9447 9027
rect 22385 8993 22419 9027
rect 23949 8993 23983 9027
rect 30757 8993 30791 9027
rect 31033 8993 31067 9027
rect 32597 8993 32631 9027
rect 33333 8993 33367 9027
rect 36461 8993 36495 9027
rect 4353 8925 4387 8959
rect 4629 8925 4663 8959
rect 4721 8925 4755 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 11253 8925 11287 8959
rect 11437 8925 11471 8959
rect 19441 8925 19475 8959
rect 19809 8925 19843 8959
rect 22661 8925 22695 8959
rect 23857 8925 23891 8959
rect 24409 8925 24443 8959
rect 24593 8925 24627 8959
rect 26739 8925 26773 8959
rect 26893 8925 26927 8959
rect 27537 8925 27571 8959
rect 28365 8925 28399 8959
rect 28825 8925 28859 8959
rect 29009 8925 29043 8959
rect 29101 8925 29135 8959
rect 29193 8925 29227 8959
rect 30481 8925 30515 8959
rect 33149 8925 33183 8959
rect 33517 8925 33551 8959
rect 33977 8925 34011 8959
rect 34253 8925 34287 8959
rect 34345 8925 34379 8959
rect 35449 8925 35483 8959
rect 37105 8925 37139 8959
rect 37197 8925 37231 8959
rect 37565 8925 37599 8959
rect 5825 8857 5859 8891
rect 9689 8857 9723 8891
rect 19533 8857 19567 8891
rect 19625 8857 19659 8891
rect 22845 8857 22879 8891
rect 28733 8857 28767 8891
rect 34161 8857 34195 8891
rect 37381 8857 37415 8891
rect 37473 8857 37507 8891
rect 3801 8789 3835 8823
rect 4905 8789 4939 8823
rect 5625 8789 5659 8823
rect 19257 8789 19291 8823
rect 26525 8789 26559 8823
rect 28181 8789 28215 8823
rect 29377 8789 29411 8823
rect 34529 8789 34563 8823
rect 37749 8789 37783 8823
rect 3893 8585 3927 8619
rect 4445 8585 4479 8619
rect 5473 8585 5507 8619
rect 5641 8585 5675 8619
rect 5825 8585 5859 8619
rect 8861 8585 8895 8619
rect 18889 8585 18923 8619
rect 26801 8585 26835 8619
rect 32873 8585 32907 8619
rect 34253 8585 34287 8619
rect 36277 8585 36311 8619
rect 1685 8517 1719 8551
rect 4077 8517 4111 8551
rect 4277 8517 4311 8551
rect 5273 8517 5307 8551
rect 6561 8517 6595 8551
rect 8033 8517 8067 8551
rect 20361 8517 20395 8551
rect 20729 8517 20763 8551
rect 24041 8517 24075 8551
rect 26525 8517 26559 8551
rect 28273 8517 28307 8551
rect 28365 8517 28399 8551
rect 34069 8517 34103 8551
rect 36185 8517 36219 8551
rect 37841 8517 37875 8551
rect 3617 8449 3651 8483
rect 4537 8449 4571 8483
rect 4813 8449 4847 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 6469 8449 6503 8483
rect 6745 8449 6779 8483
rect 7297 8449 7331 8483
rect 8309 8449 8343 8483
rect 8953 8449 8987 8483
rect 9045 8449 9079 8483
rect 16957 8449 16991 8483
rect 21557 8449 21591 8483
rect 22661 8449 22695 8483
rect 23765 8449 23799 8483
rect 24409 8449 24443 8483
rect 24593 8449 24627 8483
rect 24685 8449 24719 8483
rect 24777 8449 24811 8483
rect 26249 8449 26283 8483
rect 26433 8449 26467 8483
rect 26617 8449 26651 8483
rect 27537 8449 27571 8483
rect 27997 8449 28031 8483
rect 28917 8449 28951 8483
rect 29469 8449 29503 8483
rect 30205 8449 30239 8483
rect 33057 8449 33091 8483
rect 33149 8449 33183 8483
rect 33241 8449 33275 8483
rect 33425 8449 33459 8483
rect 33686 8449 33720 8483
rect 33793 8449 33827 8483
rect 37565 8449 37599 8483
rect 37933 8449 37967 8483
rect 1409 8381 1443 8415
rect 3249 8381 3283 8415
rect 3709 8381 3743 8415
rect 4629 8381 4663 8415
rect 8217 8381 8251 8415
rect 8585 8381 8619 8415
rect 17233 8381 17267 8415
rect 20637 8381 20671 8415
rect 23673 8381 23707 8415
rect 24133 8381 24167 8415
rect 26985 8381 27019 8415
rect 27905 8381 27939 8415
rect 28825 8381 28859 8415
rect 29193 8381 29227 8415
rect 29285 8381 29319 8415
rect 30481 8381 30515 8415
rect 31953 8381 31987 8415
rect 32137 8381 32171 8415
rect 34161 8381 34195 8415
rect 34805 8381 34839 8415
rect 35449 8381 35483 8415
rect 36829 8381 36863 8415
rect 37473 8381 37507 8415
rect 3157 8313 3191 8347
rect 4997 8313 5031 8347
rect 7113 8313 7147 8347
rect 8493 8313 8527 8347
rect 18705 8313 18739 8347
rect 27721 8313 27755 8347
rect 37289 8313 37323 8347
rect 4261 8245 4295 8279
rect 4813 8245 4847 8279
rect 5457 8245 5491 8279
rect 6745 8245 6779 8279
rect 8217 8245 8251 8279
rect 23489 8245 23523 8279
rect 24961 8245 24995 8279
rect 28641 8245 28675 8279
rect 30113 8245 30147 8279
rect 32781 8245 32815 8279
rect 33517 8245 33551 8279
rect 3893 8041 3927 8075
rect 6469 8041 6503 8075
rect 7113 8041 7147 8075
rect 8125 8041 8159 8075
rect 8769 8041 8803 8075
rect 9505 8041 9539 8075
rect 19993 8041 20027 8075
rect 25237 8041 25271 8075
rect 27445 8041 27479 8075
rect 31401 8041 31435 8075
rect 34437 8041 34471 8075
rect 35436 8041 35470 8075
rect 37657 8041 37691 8075
rect 4537 7973 4571 8007
rect 7757 7973 7791 8007
rect 7849 7973 7883 8007
rect 31309 7973 31343 8007
rect 1409 7905 1443 7939
rect 1685 7905 1719 7939
rect 3157 7905 3191 7939
rect 3249 7905 3283 7939
rect 6653 7905 6687 7939
rect 8217 7905 8251 7939
rect 9045 7905 9079 7939
rect 9137 7905 9171 7939
rect 11437 7905 11471 7939
rect 19349 7905 19383 7939
rect 22385 7905 22419 7939
rect 22477 7905 22511 7939
rect 25697 7905 25731 7939
rect 25973 7905 26007 7939
rect 27537 7905 27571 7939
rect 29009 7905 29043 7939
rect 29285 7905 29319 7939
rect 29561 7905 29595 7939
rect 29837 7905 29871 7939
rect 31585 7905 31619 7939
rect 31953 7905 31987 7939
rect 32045 7905 32079 7939
rect 32689 7905 32723 7939
rect 35173 7905 35207 7939
rect 36921 7905 36955 7939
rect 37013 7905 37047 7939
rect 3433 7837 3467 7871
rect 4261 7837 4295 7871
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 5089 7837 5123 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 6429 7837 6463 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7849 7837 7883 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 8585 7837 8619 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 10701 7837 10735 7871
rect 24593 7837 24627 7871
rect 31677 7837 31711 7871
rect 32137 7837 32171 7871
rect 3617 7769 3651 7803
rect 4445 7769 4479 7803
rect 4813 7769 4847 7803
rect 7113 7769 7147 7803
rect 7297 7769 7331 7803
rect 7573 7769 7607 7803
rect 12265 7769 12299 7803
rect 22109 7769 22143 7803
rect 22753 7769 22787 7803
rect 32505 7769 32539 7803
rect 32965 7769 32999 7803
rect 4077 7701 4111 7735
rect 4169 7701 4203 7735
rect 5825 7701 5859 7735
rect 6285 7701 6319 7735
rect 7941 7701 7975 7735
rect 20637 7701 20671 7735
rect 24225 7701 24259 7735
rect 2697 7497 2731 7531
rect 3341 7497 3375 7531
rect 8125 7497 8159 7531
rect 8309 7497 8343 7531
rect 19257 7497 19291 7531
rect 21649 7497 21683 7531
rect 22569 7497 22603 7531
rect 23949 7497 23983 7531
rect 27353 7497 27387 7531
rect 29837 7497 29871 7531
rect 33241 7497 33275 7531
rect 35357 7497 35391 7531
rect 4629 7429 4663 7463
rect 9289 7429 9323 7463
rect 9505 7429 9539 7463
rect 11161 7429 11195 7463
rect 19809 7429 19843 7463
rect 19901 7429 19935 7463
rect 21281 7429 21315 7463
rect 21373 7429 21407 7463
rect 22477 7429 22511 7463
rect 23121 7429 23155 7463
rect 23213 7429 23247 7463
rect 25421 7429 25455 7463
rect 34713 7429 34747 7463
rect 2329 7361 2363 7395
rect 2421 7361 2455 7395
rect 2513 7361 2547 7395
rect 2973 7361 3007 7395
rect 3709 7361 3743 7395
rect 3801 7361 3835 7395
rect 3893 7361 3927 7395
rect 4077 7361 4111 7395
rect 4261 7361 4295 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 4721 7361 4755 7395
rect 5273 7361 5307 7395
rect 8217 7361 8251 7395
rect 8401 7361 8435 7395
rect 11713 7361 11747 7395
rect 12265 7361 12299 7395
rect 19441 7361 19475 7395
rect 19533 7361 19567 7395
rect 21097 7361 21131 7395
rect 21465 7361 21499 7395
rect 22845 7361 22879 7395
rect 25697 7361 25731 7395
rect 27445 7361 27479 7395
rect 27997 7361 28031 7395
rect 34989 7361 35023 7395
rect 37105 7361 37139 7395
rect 3065 7293 3099 7327
rect 3617 7293 3651 7327
rect 6377 7293 6411 7327
rect 6653 7293 6687 7327
rect 11897 7293 11931 7327
rect 11989 7293 12023 7327
rect 21833 7293 21867 7327
rect 22753 7293 22787 7327
rect 28273 7293 28307 7327
rect 29745 7293 29779 7327
rect 30389 7293 30423 7327
rect 36829 7293 36863 7327
rect 3433 7225 3467 7259
rect 11529 7225 11563 7259
rect 4169 7157 4203 7191
rect 4905 7157 4939 7191
rect 5089 7157 5123 7191
rect 9137 7157 9171 7191
rect 9321 7157 9355 7191
rect 11253 7157 11287 7191
rect 12173 7157 12207 7191
rect 4169 6953 4203 6987
rect 5653 6953 5687 6987
rect 9229 6953 9263 6987
rect 9413 6953 9447 6987
rect 12449 6953 12483 6987
rect 5917 6749 5951 6783
rect 6929 6749 6963 6783
rect 7021 6749 7055 6783
rect 7205 6749 7239 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9689 6749 9723 6783
rect 10701 6749 10735 6783
rect 12541 6749 12575 6783
rect 13001 6749 13035 6783
rect 6561 6681 6595 6715
rect 9597 6681 9631 6715
rect 10977 6681 11011 6715
rect 9045 6613 9079 6647
rect 9397 6613 9431 6647
rect 10333 6613 10367 6647
rect 12633 6613 12667 6647
rect 12725 6613 12759 6647
rect 9505 6409 9539 6443
rect 11161 6409 11195 6443
rect 9689 6273 9723 6307
rect 9781 6273 9815 6307
rect 9965 6273 9999 6307
rect 10149 6273 10183 6307
rect 10425 6273 10459 6307
rect 10609 6273 10643 6307
rect 10977 6273 11011 6307
rect 11253 6273 11287 6307
rect 11713 6273 11747 6307
rect 11897 6273 11931 6307
rect 11989 6273 12023 6307
rect 7665 6205 7699 6239
rect 7941 6205 7975 6239
rect 11529 6205 11563 6239
rect 11805 6205 11839 6239
rect 10241 6137 10275 6171
rect 10333 6137 10367 6171
rect 9413 6069 9447 6103
rect 9873 6069 9907 6103
rect 10793 6069 10827 6103
rect 4813 5865 4847 5899
rect 5089 5865 5123 5899
rect 5549 5865 5583 5899
rect 9229 5865 9263 5899
rect 9505 5865 9539 5899
rect 12357 5865 12391 5899
rect 2237 5729 2271 5763
rect 2513 5729 2547 5763
rect 7113 5729 7147 5763
rect 2145 5661 2179 5695
rect 2605 5661 2639 5695
rect 2697 5661 2731 5695
rect 2881 5661 2915 5695
rect 4261 5661 4295 5695
rect 4537 5661 4571 5695
rect 5089 5661 5123 5695
rect 5273 5661 5307 5695
rect 5365 5661 5399 5695
rect 6745 5661 6779 5695
rect 7021 5661 7055 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 8953 5661 8987 5695
rect 9045 5661 9079 5695
rect 9689 5661 9723 5695
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 10609 5661 10643 5695
rect 4445 5593 4479 5627
rect 4781 5593 4815 5627
rect 4997 5593 5031 5627
rect 9229 5593 9263 5627
rect 9873 5593 9907 5627
rect 10885 5593 10919 5627
rect 3065 5525 3099 5559
rect 4077 5525 4111 5559
rect 4629 5525 4663 5559
rect 6561 5525 6595 5559
rect 6929 5525 6963 5559
rect 2513 5321 2547 5355
rect 9321 5321 9355 5355
rect 10149 5321 10183 5355
rect 6009 5253 6043 5287
rect 6653 5253 6687 5287
rect 11897 5253 11931 5287
rect 2237 5185 2271 5219
rect 4261 5185 4295 5219
rect 9229 5185 9263 5219
rect 9413 5185 9447 5219
rect 9689 5185 9723 5219
rect 9873 5185 9907 5219
rect 9965 5185 9999 5219
rect 10241 5185 10275 5219
rect 10425 5185 10459 5219
rect 10517 5185 10551 5219
rect 2053 5117 2087 5151
rect 2421 5117 2455 5151
rect 3985 5117 4019 5151
rect 4353 5117 4387 5151
rect 5273 5117 5307 5151
rect 6377 5117 6411 5151
rect 9045 5049 9079 5083
rect 4997 4981 5031 5015
rect 8125 4981 8159 5015
rect 9597 4981 9631 5015
rect 9873 4981 9907 5015
rect 10241 4981 10275 5015
rect 11805 4981 11839 5015
rect 1409 4777 1443 4811
rect 4169 4777 4203 4811
rect 4997 4777 5031 4811
rect 7021 4777 7055 4811
rect 9137 4777 9171 4811
rect 9965 4777 9999 4811
rect 4445 4709 4479 4743
rect 7297 4709 7331 4743
rect 8677 4709 8711 4743
rect 3157 4641 3191 4675
rect 6745 4641 6779 4675
rect 10333 4641 10367 4675
rect 12081 4641 12115 4675
rect 3801 4573 3835 4607
rect 4629 4573 4663 4607
rect 4813 4573 4847 4607
rect 5549 4573 5583 4607
rect 6653 4573 6687 4607
rect 8401 4573 8435 4607
rect 8677 4573 8711 4607
rect 9781 4573 9815 4607
rect 9965 4573 9999 4607
rect 10057 4573 10091 4607
rect 10241 4573 10275 4607
rect 12541 4573 12575 4607
rect 2881 4505 2915 4539
rect 4169 4505 4203 4539
rect 4721 4505 4755 4539
rect 7481 4505 7515 4539
rect 8493 4505 8527 4539
rect 9105 4505 9139 4539
rect 9321 4505 9355 4539
rect 10149 4505 10183 4539
rect 11805 4505 11839 4539
rect 4353 4437 4387 4471
rect 8953 4437 8987 4471
rect 12265 4437 12299 4471
rect 4997 4233 5031 4267
rect 5365 4233 5399 4267
rect 5733 4165 5767 4199
rect 4261 4097 4295 4131
rect 5181 4097 5215 4131
rect 5457 4097 5491 4131
rect 5917 4097 5951 4131
rect 8217 4097 8251 4131
rect 8401 4097 8435 4131
rect 8677 4097 8711 4131
rect 8769 4097 8803 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 10057 4097 10091 4131
rect 10149 4097 10183 4131
rect 10425 4097 10459 4131
rect 4537 4029 4571 4063
rect 4629 4029 4663 4063
rect 4721 4029 4755 4063
rect 4813 4029 4847 4063
rect 9137 4029 9171 4063
rect 9689 4029 9723 4063
rect 4353 3961 4387 3995
rect 8493 3961 8527 3995
rect 9873 3961 9907 3995
rect 4169 3893 4203 3927
rect 5549 3893 5583 3927
rect 8401 3893 8435 3927
rect 11069 3893 11103 3927
rect 5641 3689 5675 3723
rect 10793 3689 10827 3723
rect 11253 3689 11287 3723
rect 3341 3621 3375 3655
rect 3433 3621 3467 3655
rect 10885 3621 10919 3655
rect 3893 3553 3927 3587
rect 6009 3553 6043 3587
rect 8125 3553 8159 3587
rect 8493 3553 8527 3587
rect 9413 3553 9447 3587
rect 11161 3553 11195 3587
rect 41889 3553 41923 3587
rect 3249 3485 3283 3519
rect 3525 3485 3559 3519
rect 5733 3485 5767 3519
rect 5825 3485 5859 3519
rect 6193 3485 6227 3519
rect 8585 3485 8619 3519
rect 10057 3485 10091 3519
rect 10241 3485 10275 3519
rect 10517 3485 10551 3519
rect 10609 3485 10643 3519
rect 11437 3485 11471 3519
rect 42165 3485 42199 3519
rect 4169 3417 4203 3451
rect 10425 3417 10459 3451
rect 3065 3349 3099 3383
rect 8769 3349 8803 3383
rect 4997 3145 5031 3179
rect 9413 3145 9447 3179
rect 3433 3077 3467 3111
rect 5273 3077 5307 3111
rect 5365 3077 5399 3111
rect 7941 3077 7975 3111
rect 9781 3077 9815 3111
rect 3157 3009 3191 3043
rect 5181 3009 5215 3043
rect 5549 3009 5583 3043
rect 7665 3009 7699 3043
rect 9505 3009 9539 3043
rect 4905 2941 4939 2975
rect 11253 2941 11287 2975
rect 11713 2397 11747 2431
rect 11897 2261 11931 2295
<< metal1 >>
rect 1104 43546 42504 43568
rect 1104 43494 4874 43546
rect 4926 43494 4938 43546
rect 4990 43494 5002 43546
rect 5054 43494 5066 43546
rect 5118 43494 5130 43546
rect 5182 43494 35594 43546
rect 35646 43494 35658 43546
rect 35710 43494 35722 43546
rect 35774 43494 35786 43546
rect 35838 43494 35850 43546
rect 35902 43494 42504 43546
rect 1104 43472 42504 43494
rect 17678 43392 17684 43444
rect 17736 43392 17742 43444
rect 19518 43392 19524 43444
rect 19576 43392 19582 43444
rect 20254 43392 20260 43444
rect 20312 43392 20318 43444
rect 20530 43392 20536 43444
rect 20588 43432 20594 43444
rect 20809 43435 20867 43441
rect 20809 43432 20821 43435
rect 20588 43404 20821 43432
rect 20588 43392 20594 43404
rect 20809 43401 20821 43404
rect 20855 43401 20867 43435
rect 20809 43395 20867 43401
rect 22830 43392 22836 43444
rect 22888 43392 22894 43444
rect 23382 43392 23388 43444
rect 23440 43392 23446 43444
rect 25314 43392 25320 43444
rect 25372 43392 25378 43444
rect 29178 43392 29184 43444
rect 29236 43392 29242 43444
rect 24394 43324 24400 43376
rect 24452 43364 24458 43376
rect 24673 43367 24731 43373
rect 24673 43364 24685 43367
rect 24452 43336 24685 43364
rect 24452 43324 24458 43336
rect 24673 43333 24685 43336
rect 24719 43333 24731 43367
rect 24673 43327 24731 43333
rect 28169 43367 28227 43373
rect 28169 43333 28181 43367
rect 28215 43364 28227 43367
rect 28442 43364 28448 43376
rect 28215 43336 28448 43364
rect 28215 43333 28227 43336
rect 28169 43327 28227 43333
rect 28442 43324 28448 43336
rect 28500 43324 28506 43376
rect 17494 43256 17500 43308
rect 17552 43256 17558 43308
rect 19705 43299 19763 43305
rect 19705 43265 19717 43299
rect 19751 43296 19763 43299
rect 19794 43296 19800 43308
rect 19751 43268 19800 43296
rect 19751 43265 19763 43268
rect 19705 43259 19763 43265
rect 19794 43256 19800 43268
rect 19852 43256 19858 43308
rect 20073 43299 20131 43305
rect 20073 43265 20085 43299
rect 20119 43265 20131 43299
rect 20073 43259 20131 43265
rect 19334 43188 19340 43240
rect 19392 43228 19398 43240
rect 20088 43228 20116 43259
rect 20990 43256 20996 43308
rect 21048 43256 21054 43308
rect 22649 43299 22707 43305
rect 22649 43265 22661 43299
rect 22695 43296 22707 43299
rect 22738 43296 22744 43308
rect 22695 43268 22744 43296
rect 22695 43265 22707 43268
rect 22649 43259 22707 43265
rect 22738 43256 22744 43268
rect 22796 43256 22802 43308
rect 23014 43256 23020 43308
rect 23072 43296 23078 43308
rect 23569 43299 23627 43305
rect 23569 43296 23581 43299
rect 23072 43268 23581 43296
rect 23072 43256 23078 43268
rect 23569 43265 23581 43268
rect 23615 43265 23627 43299
rect 23569 43259 23627 43265
rect 24578 43256 24584 43308
rect 24636 43256 24642 43308
rect 24765 43299 24823 43305
rect 24765 43265 24777 43299
rect 24811 43265 24823 43299
rect 24765 43259 24823 43265
rect 24949 43299 25007 43305
rect 24949 43265 24961 43299
rect 24995 43296 25007 43299
rect 25501 43299 25559 43305
rect 25501 43296 25513 43299
rect 24995 43268 25513 43296
rect 24995 43265 25007 43268
rect 24949 43259 25007 43265
rect 25501 43265 25513 43268
rect 25547 43296 25559 43299
rect 26142 43296 26148 43308
rect 25547 43268 26148 43296
rect 25547 43265 25559 43268
rect 25501 43259 25559 43265
rect 19392 43200 20116 43228
rect 19392 43188 19398 43200
rect 24670 43188 24676 43240
rect 24728 43228 24734 43240
rect 24780 43228 24808 43259
rect 26142 43256 26148 43268
rect 26200 43256 26206 43308
rect 28350 43256 28356 43308
rect 28408 43256 28414 43308
rect 29365 43299 29423 43305
rect 29365 43265 29377 43299
rect 29411 43296 29423 43299
rect 29546 43296 29552 43308
rect 29411 43268 29552 43296
rect 29411 43265 29423 43268
rect 29365 43259 29423 43265
rect 29546 43256 29552 43268
rect 29604 43256 29610 43308
rect 24728 43200 24808 43228
rect 24728 43188 24734 43200
rect 24026 43052 24032 43104
rect 24084 43092 24090 43104
rect 24397 43095 24455 43101
rect 24397 43092 24409 43095
rect 24084 43064 24409 43092
rect 24084 43052 24090 43064
rect 24397 43061 24409 43064
rect 24443 43061 24455 43095
rect 24397 43055 24455 43061
rect 28074 43052 28080 43104
rect 28132 43092 28138 43104
rect 28537 43095 28595 43101
rect 28537 43092 28549 43095
rect 28132 43064 28549 43092
rect 28132 43052 28138 43064
rect 28537 43061 28549 43064
rect 28583 43061 28595 43095
rect 28537 43055 28595 43061
rect 1104 43002 42504 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 42504 43002
rect 1104 42928 42504 42950
rect 17405 42891 17463 42897
rect 17405 42857 17417 42891
rect 17451 42888 17463 42891
rect 17494 42888 17500 42900
rect 17451 42860 17500 42888
rect 17451 42857 17463 42860
rect 17405 42851 17463 42857
rect 17494 42848 17500 42860
rect 17552 42848 17558 42900
rect 26142 42848 26148 42900
rect 26200 42848 26206 42900
rect 28350 42848 28356 42900
rect 28408 42888 28414 42900
rect 28445 42891 28503 42897
rect 28445 42888 28457 42891
rect 28408 42860 28457 42888
rect 28408 42848 28414 42860
rect 28445 42857 28457 42860
rect 28491 42857 28503 42891
rect 28445 42851 28503 42857
rect 24397 42755 24455 42761
rect 24397 42721 24409 42755
rect 24443 42752 24455 42755
rect 24762 42752 24768 42764
rect 24443 42724 24768 42752
rect 24443 42721 24455 42724
rect 24397 42715 24455 42721
rect 24762 42712 24768 42724
rect 24820 42752 24826 42764
rect 26329 42755 26387 42761
rect 26329 42752 26341 42755
rect 24820 42724 26341 42752
rect 24820 42712 24826 42724
rect 26329 42721 26341 42724
rect 26375 42752 26387 42755
rect 27614 42752 27620 42764
rect 26375 42724 27620 42752
rect 26375 42721 26387 42724
rect 26329 42715 26387 42721
rect 27614 42712 27620 42724
rect 27672 42712 27678 42764
rect 29638 42752 29644 42764
rect 27724 42724 29644 42752
rect 15654 42644 15660 42696
rect 15712 42644 15718 42696
rect 18325 42687 18383 42693
rect 18325 42653 18337 42687
rect 18371 42684 18383 42687
rect 19058 42684 19064 42696
rect 18371 42656 19064 42684
rect 18371 42653 18383 42656
rect 18325 42647 18383 42653
rect 19058 42644 19064 42656
rect 19116 42644 19122 42696
rect 19429 42687 19487 42693
rect 19429 42653 19441 42687
rect 19475 42684 19487 42687
rect 19475 42656 19748 42684
rect 19475 42653 19487 42656
rect 19429 42647 19487 42653
rect 15933 42619 15991 42625
rect 15933 42585 15945 42619
rect 15979 42616 15991 42619
rect 16206 42616 16212 42628
rect 15979 42588 16212 42616
rect 15979 42585 15991 42588
rect 15933 42579 15991 42585
rect 16206 42576 16212 42588
rect 16264 42576 16270 42628
rect 16390 42576 16396 42628
rect 16448 42576 16454 42628
rect 18509 42619 18567 42625
rect 18509 42585 18521 42619
rect 18555 42616 18567 42619
rect 18555 42588 19288 42616
rect 18555 42585 18567 42588
rect 18509 42579 18567 42585
rect 18138 42508 18144 42560
rect 18196 42548 18202 42560
rect 19260 42557 19288 42588
rect 19518 42576 19524 42628
rect 19576 42576 19582 42628
rect 19613 42619 19671 42625
rect 19613 42585 19625 42619
rect 19659 42585 19671 42619
rect 19720 42616 19748 42656
rect 19794 42644 19800 42696
rect 19852 42644 19858 42696
rect 19886 42644 19892 42696
rect 19944 42684 19950 42696
rect 20993 42687 21051 42693
rect 20993 42684 21005 42687
rect 19944 42656 21005 42684
rect 19944 42644 19950 42656
rect 20993 42653 21005 42656
rect 21039 42653 21051 42687
rect 20993 42647 21051 42653
rect 24026 42644 24032 42696
rect 24084 42644 24090 42696
rect 25682 42644 25688 42696
rect 25740 42684 25746 42696
rect 25740 42670 25806 42684
rect 27724 42670 27752 42724
rect 29638 42712 29644 42724
rect 29696 42712 29702 42764
rect 35161 42755 35219 42761
rect 35161 42721 35173 42755
rect 35207 42752 35219 42755
rect 37274 42752 37280 42764
rect 35207 42724 37280 42752
rect 35207 42721 35219 42724
rect 35161 42715 35219 42721
rect 37274 42712 37280 42724
rect 37332 42712 37338 42764
rect 25740 42656 25820 42670
rect 25740 42644 25746 42656
rect 20806 42616 20812 42628
rect 19720 42588 20812 42616
rect 19613 42579 19671 42585
rect 18693 42551 18751 42557
rect 18693 42548 18705 42551
rect 18196 42520 18705 42548
rect 18196 42508 18202 42520
rect 18693 42517 18705 42520
rect 18739 42517 18751 42551
rect 18693 42511 18751 42517
rect 19245 42551 19303 42557
rect 19245 42517 19257 42551
rect 19291 42517 19303 42551
rect 19245 42511 19303 42517
rect 19426 42508 19432 42560
rect 19484 42548 19490 42560
rect 19628 42548 19656 42579
rect 20806 42576 20812 42588
rect 20864 42576 20870 42628
rect 21269 42619 21327 42625
rect 21269 42585 21281 42619
rect 21315 42616 21327 42619
rect 21542 42616 21548 42628
rect 21315 42588 21548 42616
rect 21315 42585 21327 42588
rect 21269 42579 21327 42585
rect 21542 42576 21548 42588
rect 21600 42576 21606 42628
rect 22494 42588 23612 42616
rect 22186 42548 22192 42560
rect 19484 42520 22192 42548
rect 19484 42508 19490 42520
rect 22186 42508 22192 42520
rect 22244 42508 22250 42560
rect 22738 42508 22744 42560
rect 22796 42508 22802 42560
rect 23584 42548 23612 42588
rect 23658 42576 23664 42628
rect 23716 42616 23722 42628
rect 23845 42619 23903 42625
rect 23845 42616 23857 42619
rect 23716 42588 23857 42616
rect 23716 42576 23722 42588
rect 23845 42585 23857 42588
rect 23891 42585 23903 42619
rect 23845 42579 23903 42585
rect 24213 42619 24271 42625
rect 24213 42585 24225 42619
rect 24259 42616 24271 42619
rect 24673 42619 24731 42625
rect 24673 42616 24685 42619
rect 24259 42588 24685 42616
rect 24259 42585 24271 42588
rect 24213 42579 24271 42585
rect 24673 42585 24685 42588
rect 24719 42585 24731 42619
rect 24673 42579 24731 42585
rect 24026 42548 24032 42560
rect 23584 42520 24032 42548
rect 24026 42508 24032 42520
rect 24084 42508 24090 42560
rect 25792 42548 25820 42656
rect 27890 42644 27896 42696
rect 27948 42684 27954 42696
rect 28629 42687 28687 42693
rect 28629 42684 28641 42687
rect 27948 42656 28641 42684
rect 27948 42644 27954 42656
rect 28629 42653 28641 42656
rect 28675 42653 28687 42687
rect 28629 42647 28687 42653
rect 28997 42687 29055 42693
rect 28997 42653 29009 42687
rect 29043 42684 29055 42687
rect 29546 42684 29552 42696
rect 29043 42656 29552 42684
rect 29043 42653 29055 42656
rect 28997 42647 29055 42653
rect 29546 42644 29552 42656
rect 29604 42644 29610 42696
rect 26602 42576 26608 42628
rect 26660 42576 26666 42628
rect 28534 42616 28540 42628
rect 27908 42588 28540 42616
rect 27908 42548 27936 42588
rect 28534 42576 28540 42588
rect 28592 42576 28598 42628
rect 28721 42619 28779 42625
rect 28721 42585 28733 42619
rect 28767 42585 28779 42619
rect 28721 42579 28779 42585
rect 25792 42520 27936 42548
rect 28077 42551 28135 42557
rect 28077 42517 28089 42551
rect 28123 42548 28135 42551
rect 28258 42548 28264 42560
rect 28123 42520 28264 42548
rect 28123 42517 28135 42520
rect 28077 42511 28135 42517
rect 28258 42508 28264 42520
rect 28316 42548 28322 42560
rect 28736 42548 28764 42579
rect 28810 42576 28816 42628
rect 28868 42576 28874 42628
rect 35434 42576 35440 42628
rect 35492 42576 35498 42628
rect 36814 42616 36820 42628
rect 36662 42588 36820 42616
rect 36814 42576 36820 42588
rect 36872 42576 36878 42628
rect 28316 42520 28764 42548
rect 36909 42551 36967 42557
rect 28316 42508 28322 42520
rect 36909 42517 36921 42551
rect 36955 42548 36967 42551
rect 36998 42548 37004 42560
rect 36955 42520 37004 42548
rect 36955 42517 36967 42520
rect 36909 42511 36967 42517
rect 36998 42508 37004 42520
rect 37056 42508 37062 42560
rect 1104 42458 42504 42480
rect 1104 42406 4874 42458
rect 4926 42406 4938 42458
rect 4990 42406 5002 42458
rect 5054 42406 5066 42458
rect 5118 42406 5130 42458
rect 5182 42406 35594 42458
rect 35646 42406 35658 42458
rect 35710 42406 35722 42458
rect 35774 42406 35786 42458
rect 35838 42406 35850 42458
rect 35902 42406 42504 42458
rect 1104 42384 42504 42406
rect 16853 42347 16911 42353
rect 16853 42344 16865 42347
rect 16316 42316 16865 42344
rect 16316 42285 16344 42316
rect 16853 42313 16865 42316
rect 16899 42313 16911 42347
rect 18782 42344 18788 42356
rect 16853 42307 16911 42313
rect 17880 42316 18788 42344
rect 16301 42279 16359 42285
rect 16301 42245 16313 42279
rect 16347 42245 16359 42279
rect 16301 42239 16359 42245
rect 16574 42236 16580 42288
rect 16632 42276 16638 42288
rect 17129 42279 17187 42285
rect 17129 42276 17141 42279
rect 16632 42248 17141 42276
rect 16632 42236 16638 42248
rect 17129 42245 17141 42248
rect 17175 42245 17187 42279
rect 17129 42239 17187 42245
rect 15930 42168 15936 42220
rect 15988 42208 15994 42220
rect 16117 42211 16175 42217
rect 16117 42208 16129 42211
rect 15988 42180 16129 42208
rect 15988 42168 15994 42180
rect 16117 42177 16129 42180
rect 16163 42177 16175 42211
rect 16117 42171 16175 42177
rect 16206 42168 16212 42220
rect 16264 42208 16270 42220
rect 16485 42211 16543 42217
rect 16485 42208 16497 42211
rect 16264 42180 16497 42208
rect 16264 42168 16270 42180
rect 16485 42177 16497 42180
rect 16531 42177 16543 42211
rect 16485 42171 16543 42177
rect 17037 42211 17095 42217
rect 17037 42177 17049 42211
rect 17083 42208 17095 42211
rect 17221 42211 17279 42217
rect 17083 42180 17172 42208
rect 17083 42177 17095 42180
rect 17037 42171 17095 42177
rect 17144 42004 17172 42180
rect 17221 42177 17233 42211
rect 17267 42177 17279 42211
rect 17221 42171 17279 42177
rect 17405 42211 17463 42217
rect 17405 42177 17417 42211
rect 17451 42208 17463 42211
rect 17494 42208 17500 42220
rect 17451 42180 17500 42208
rect 17451 42177 17463 42180
rect 17405 42171 17463 42177
rect 17236 42140 17264 42171
rect 17494 42168 17500 42180
rect 17552 42168 17558 42220
rect 17880 42217 17908 42316
rect 18782 42304 18788 42316
rect 18840 42344 18846 42356
rect 19886 42344 19892 42356
rect 18840 42316 19892 42344
rect 18840 42304 18846 42316
rect 19886 42304 19892 42316
rect 19944 42304 19950 42356
rect 22002 42304 22008 42356
rect 22060 42344 22066 42356
rect 24578 42344 24584 42356
rect 22060 42316 24584 42344
rect 22060 42304 22066 42316
rect 24578 42304 24584 42316
rect 24636 42304 24642 42356
rect 24670 42304 24676 42356
rect 24728 42344 24734 42356
rect 24728 42316 25176 42344
rect 24728 42304 24734 42316
rect 18138 42236 18144 42288
rect 18196 42236 18202 42288
rect 19150 42236 19156 42288
rect 19208 42236 19214 42288
rect 20714 42236 20720 42288
rect 20772 42236 20778 42288
rect 25148 42276 25176 42316
rect 26602 42304 26608 42356
rect 26660 42344 26666 42356
rect 26973 42347 27031 42353
rect 26973 42344 26985 42347
rect 26660 42316 26985 42344
rect 26660 42304 26666 42316
rect 26973 42313 26985 42316
rect 27019 42313 27031 42347
rect 28258 42344 28264 42356
rect 26973 42307 27031 42313
rect 27632 42316 28264 42344
rect 27632 42285 27660 42316
rect 28258 42304 28264 42316
rect 28316 42304 28322 42356
rect 29546 42304 29552 42356
rect 29604 42304 29610 42356
rect 35345 42347 35403 42353
rect 35345 42313 35357 42347
rect 35391 42344 35403 42347
rect 35434 42344 35440 42356
rect 35391 42316 35440 42344
rect 35391 42313 35403 42316
rect 35345 42307 35403 42313
rect 35434 42304 35440 42316
rect 35492 42304 35498 42356
rect 39025 42347 39083 42353
rect 39025 42344 39037 42347
rect 36740 42316 39037 42344
rect 27617 42279 27675 42285
rect 25148 42248 27568 42276
rect 17865 42211 17923 42217
rect 17865 42177 17877 42211
rect 17911 42177 17923 42211
rect 17865 42171 17923 42177
rect 19886 42168 19892 42220
rect 19944 42168 19950 42220
rect 24026 42168 24032 42220
rect 24084 42208 24090 42220
rect 25590 42208 25596 42220
rect 24084 42180 25596 42208
rect 24084 42168 24090 42180
rect 25590 42168 25596 42180
rect 25648 42168 25654 42220
rect 27249 42211 27307 42217
rect 27249 42177 27261 42211
rect 27295 42208 27307 42211
rect 27430 42208 27436 42220
rect 27295 42180 27436 42208
rect 27295 42177 27307 42180
rect 27249 42171 27307 42177
rect 27430 42168 27436 42180
rect 27488 42168 27494 42220
rect 27540 42208 27568 42248
rect 27617 42245 27629 42279
rect 27663 42245 27675 42279
rect 27617 42239 27675 42245
rect 28074 42236 28080 42288
rect 28132 42236 28138 42288
rect 28534 42236 28540 42288
rect 28592 42236 28598 42288
rect 29638 42236 29644 42288
rect 29696 42276 29702 42288
rect 29696 42248 30958 42276
rect 34808 42248 35894 42276
rect 29696 42236 29702 42248
rect 34808 42220 34836 42248
rect 32401 42211 32459 42217
rect 27540 42180 27660 42208
rect 19426 42140 19432 42152
rect 17236 42112 19432 42140
rect 19426 42100 19432 42112
rect 19484 42100 19490 42152
rect 19613 42143 19671 42149
rect 19613 42109 19625 42143
rect 19659 42140 19671 42143
rect 19794 42140 19800 42152
rect 19659 42112 19800 42140
rect 19659 42109 19671 42112
rect 19613 42103 19671 42109
rect 19794 42100 19800 42112
rect 19852 42100 19858 42152
rect 20162 42100 20168 42152
rect 20220 42100 20226 42152
rect 22373 42143 22431 42149
rect 22373 42140 22385 42143
rect 21744 42112 22385 42140
rect 21744 42016 21772 42112
rect 22373 42109 22385 42112
rect 22419 42109 22431 42143
rect 22373 42103 22431 42109
rect 22646 42100 22652 42152
rect 22704 42100 22710 42152
rect 22925 42143 22983 42149
rect 22925 42109 22937 42143
rect 22971 42140 22983 42143
rect 23290 42140 23296 42152
rect 22971 42112 23296 42140
rect 22971 42109 22983 42112
rect 22925 42103 22983 42109
rect 23290 42100 23296 42112
rect 23348 42100 23354 42152
rect 27157 42143 27215 42149
rect 27157 42109 27169 42143
rect 27203 42140 27215 42143
rect 27338 42140 27344 42152
rect 27203 42112 27344 42140
rect 27203 42109 27215 42112
rect 27157 42103 27215 42109
rect 27338 42100 27344 42112
rect 27396 42100 27402 42152
rect 27525 42143 27583 42149
rect 27525 42109 27537 42143
rect 27571 42109 27583 42143
rect 27525 42103 27583 42109
rect 20806 42004 20812 42016
rect 17144 41976 20812 42004
rect 20806 41964 20812 41976
rect 20864 41964 20870 42016
rect 21637 42007 21695 42013
rect 21637 41973 21649 42007
rect 21683 42004 21695 42007
rect 21726 42004 21732 42016
rect 21683 41976 21732 42004
rect 21683 41973 21695 41976
rect 21637 41967 21695 41973
rect 21726 41964 21732 41976
rect 21784 41964 21790 42016
rect 21818 41964 21824 42016
rect 21876 41964 21882 42016
rect 24394 41964 24400 42016
rect 24452 42004 24458 42016
rect 25314 42004 25320 42016
rect 24452 41976 25320 42004
rect 24452 41964 24458 41976
rect 25314 41964 25320 41976
rect 25372 41964 25378 42016
rect 26878 41964 26884 42016
rect 26936 42004 26942 42016
rect 27540 42004 27568 42103
rect 27632 42072 27660 42180
rect 32401 42177 32413 42211
rect 32447 42208 32459 42211
rect 34790 42208 34796 42220
rect 32447 42180 34796 42208
rect 32447 42177 32459 42180
rect 32401 42171 32459 42177
rect 34790 42168 34796 42180
rect 34848 42168 34854 42220
rect 35618 42168 35624 42220
rect 35676 42168 35682 42220
rect 35866 42208 35894 42248
rect 36265 42211 36323 42217
rect 36265 42208 36277 42211
rect 35866 42180 36277 42208
rect 36265 42177 36277 42180
rect 36311 42177 36323 42211
rect 36265 42171 36323 42177
rect 36446 42168 36452 42220
rect 36504 42208 36510 42220
rect 36740 42217 36768 42316
rect 39025 42313 39037 42316
rect 39071 42313 39083 42347
rect 39025 42307 39083 42313
rect 36814 42236 36820 42288
rect 36872 42276 36878 42288
rect 36872 42248 38042 42276
rect 36872 42236 36878 42248
rect 36725 42211 36783 42217
rect 36725 42208 36737 42211
rect 36504 42180 36737 42208
rect 36504 42168 36510 42180
rect 36725 42177 36737 42180
rect 36771 42177 36783 42211
rect 36725 42171 36783 42177
rect 37274 42168 37280 42220
rect 37332 42168 37338 42220
rect 27706 42100 27712 42152
rect 27764 42140 27770 42152
rect 27801 42143 27859 42149
rect 27801 42140 27813 42143
rect 27764 42112 27813 42140
rect 27764 42100 27770 42112
rect 27801 42109 27813 42112
rect 27847 42109 27859 42143
rect 28718 42140 28724 42152
rect 27801 42103 27859 42109
rect 27908 42112 28724 42140
rect 27908 42072 27936 42112
rect 28718 42100 28724 42112
rect 28776 42100 28782 42152
rect 28810 42100 28816 42152
rect 28868 42140 28874 42152
rect 30193 42143 30251 42149
rect 30193 42140 30205 42143
rect 28868 42112 30205 42140
rect 28868 42100 28874 42112
rect 30193 42109 30205 42112
rect 30239 42109 30251 42143
rect 30193 42103 30251 42109
rect 30469 42143 30527 42149
rect 30469 42109 30481 42143
rect 30515 42140 30527 42143
rect 30834 42140 30840 42152
rect 30515 42112 30840 42140
rect 30515 42109 30527 42112
rect 30469 42103 30527 42109
rect 30834 42100 30840 42112
rect 30892 42100 30898 42152
rect 30926 42100 30932 42152
rect 30984 42140 30990 42152
rect 32030 42140 32036 42152
rect 30984 42112 32036 42140
rect 30984 42100 30990 42112
rect 27632 42044 27936 42072
rect 31570 42032 31576 42084
rect 31628 42072 31634 42084
rect 31726 42072 31754 42112
rect 32030 42100 32036 42112
rect 32088 42140 32094 42152
rect 32088 42112 32260 42140
rect 32088 42100 32094 42112
rect 32232 42081 32260 42112
rect 35342 42100 35348 42152
rect 35400 42140 35406 42152
rect 35529 42143 35587 42149
rect 35529 42140 35541 42143
rect 35400 42112 35541 42140
rect 35400 42100 35406 42112
rect 35529 42109 35541 42112
rect 35575 42109 35587 42143
rect 35529 42103 35587 42109
rect 35897 42143 35955 42149
rect 35897 42109 35909 42143
rect 35943 42109 35955 42143
rect 35897 42103 35955 42109
rect 35989 42143 36047 42149
rect 35989 42109 36001 42143
rect 36035 42109 36047 42143
rect 35989 42103 36047 42109
rect 31628 42044 31754 42072
rect 32217 42075 32275 42081
rect 31628 42032 31634 42044
rect 32217 42041 32229 42075
rect 32263 42041 32275 42075
rect 32217 42035 32275 42041
rect 30926 42004 30932 42016
rect 26936 41976 30932 42004
rect 26936 41964 26942 41976
rect 30926 41964 30932 41976
rect 30984 41964 30990 42016
rect 31202 41964 31208 42016
rect 31260 42004 31266 42016
rect 31941 42007 31999 42013
rect 31941 42004 31953 42007
rect 31260 41976 31953 42004
rect 31260 41964 31266 41976
rect 31941 41973 31953 41976
rect 31987 41973 31999 42007
rect 31941 41967 31999 41973
rect 32950 41964 32956 42016
rect 33008 42004 33014 42016
rect 35912 42004 35940 42103
rect 36004 42072 36032 42103
rect 36538 42100 36544 42152
rect 36596 42100 36602 42152
rect 36630 42100 36636 42152
rect 36688 42100 36694 42152
rect 37553 42143 37611 42149
rect 37553 42140 37565 42143
rect 37108 42112 37565 42140
rect 36998 42072 37004 42084
rect 36004 42044 37004 42072
rect 36998 42032 37004 42044
rect 37056 42032 37062 42084
rect 37108 42081 37136 42112
rect 37553 42109 37565 42112
rect 37599 42109 37611 42143
rect 37553 42103 37611 42109
rect 37093 42075 37151 42081
rect 37093 42041 37105 42075
rect 37139 42041 37151 42075
rect 37093 42035 37151 42041
rect 36078 42004 36084 42016
rect 33008 41976 36084 42004
rect 33008 41964 33014 41976
rect 36078 41964 36084 41976
rect 36136 41964 36142 42016
rect 1104 41914 42504 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 42504 41914
rect 1104 41840 42504 41862
rect 20162 41760 20168 41812
rect 20220 41800 20226 41812
rect 20441 41803 20499 41809
rect 20441 41800 20453 41803
rect 20220 41772 20453 41800
rect 20220 41760 20226 41772
rect 20441 41769 20453 41772
rect 20487 41769 20499 41803
rect 20441 41763 20499 41769
rect 21542 41760 21548 41812
rect 21600 41800 21606 41812
rect 21729 41803 21787 41809
rect 21729 41800 21741 41803
rect 21600 41772 21741 41800
rect 21600 41760 21606 41772
rect 21729 41769 21741 41772
rect 21775 41769 21787 41803
rect 21729 41763 21787 41769
rect 23290 41760 23296 41812
rect 23348 41760 23354 41812
rect 27338 41760 27344 41812
rect 27396 41760 27402 41812
rect 27430 41760 27436 41812
rect 27488 41800 27494 41812
rect 28445 41803 28503 41809
rect 28445 41800 28457 41803
rect 27488 41772 28457 41800
rect 27488 41760 27494 41772
rect 28445 41769 28457 41772
rect 28491 41769 28503 41803
rect 28445 41763 28503 41769
rect 28534 41760 28540 41812
rect 28592 41800 28598 41812
rect 28905 41803 28963 41809
rect 28905 41800 28917 41803
rect 28592 41772 28917 41800
rect 28592 41760 28598 41772
rect 28905 41769 28917 41772
rect 28951 41769 28963 41803
rect 28905 41763 28963 41769
rect 29012 41772 30696 41800
rect 28718 41732 28724 41744
rect 21100 41704 27292 41732
rect 21100 41676 21128 41704
rect 14829 41667 14887 41673
rect 14829 41633 14841 41667
rect 14875 41664 14887 41667
rect 15654 41664 15660 41676
rect 14875 41636 15660 41664
rect 14875 41633 14887 41636
rect 14829 41627 14887 41633
rect 15654 41624 15660 41636
rect 15712 41664 15718 41676
rect 17129 41667 17187 41673
rect 17129 41664 17141 41667
rect 15712 41636 17141 41664
rect 15712 41624 15718 41636
rect 17129 41633 17141 41636
rect 17175 41664 17187 41667
rect 18782 41664 18788 41676
rect 17175 41636 18788 41664
rect 17175 41633 17187 41636
rect 17129 41627 17187 41633
rect 18782 41624 18788 41636
rect 18840 41624 18846 41676
rect 20070 41624 20076 41676
rect 20128 41624 20134 41676
rect 21082 41624 21088 41676
rect 21140 41624 21146 41676
rect 21726 41624 21732 41676
rect 21784 41664 21790 41676
rect 23952 41673 23980 41704
rect 23937 41667 23995 41673
rect 21784 41636 22140 41664
rect 21784 41624 21790 41636
rect 16390 41596 16396 41608
rect 16238 41568 16396 41596
rect 16390 41556 16396 41568
rect 16448 41556 16454 41608
rect 19978 41556 19984 41608
rect 20036 41556 20042 41608
rect 20714 41596 20720 41608
rect 20088 41568 20720 41596
rect 15105 41531 15163 41537
rect 15105 41497 15117 41531
rect 15151 41528 15163 41531
rect 15378 41528 15384 41540
rect 15151 41500 15384 41528
rect 15151 41497 15163 41500
rect 15105 41491 15163 41497
rect 15378 41488 15384 41500
rect 15436 41488 15442 41540
rect 17402 41488 17408 41540
rect 17460 41488 17466 41540
rect 20088 41528 20116 41568
rect 20714 41556 20720 41568
rect 20772 41556 20778 41608
rect 20809 41599 20867 41605
rect 20809 41565 20821 41599
rect 20855 41596 20867 41599
rect 21818 41596 21824 41608
rect 20855 41568 21824 41596
rect 20855 41565 20867 41568
rect 20809 41559 20867 41565
rect 21818 41556 21824 41568
rect 21876 41556 21882 41608
rect 22002 41556 22008 41608
rect 22060 41556 22066 41608
rect 22112 41605 22140 41636
rect 23937 41633 23949 41667
rect 23983 41633 23995 41667
rect 23937 41627 23995 41633
rect 24026 41624 24032 41676
rect 24084 41664 24090 41676
rect 26145 41667 26203 41673
rect 24084 41636 26096 41664
rect 24084 41624 24090 41636
rect 26068 41608 26096 41636
rect 26145 41633 26157 41667
rect 26191 41664 26203 41667
rect 26878 41664 26884 41676
rect 26191 41636 26884 41664
rect 26191 41633 26203 41636
rect 26145 41627 26203 41633
rect 22097 41599 22155 41605
rect 22097 41565 22109 41599
rect 22143 41565 22155 41599
rect 22097 41559 22155 41565
rect 22373 41599 22431 41605
rect 22373 41565 22385 41599
rect 22419 41596 22431 41599
rect 22738 41596 22744 41608
rect 22419 41568 22744 41596
rect 22419 41565 22431 41568
rect 22373 41559 22431 41565
rect 22738 41556 22744 41568
rect 22796 41556 22802 41608
rect 23661 41599 23719 41605
rect 23661 41565 23673 41599
rect 23707 41596 23719 41599
rect 24394 41596 24400 41608
rect 23707 41568 24400 41596
rect 23707 41565 23719 41568
rect 23661 41559 23719 41565
rect 24394 41556 24400 41568
rect 24452 41556 24458 41608
rect 25866 41556 25872 41608
rect 25924 41556 25930 41608
rect 25958 41556 25964 41608
rect 26016 41556 26022 41608
rect 26050 41556 26056 41608
rect 26108 41556 26114 41608
rect 20901 41531 20959 41537
rect 20901 41528 20913 41531
rect 18630 41500 20116 41528
rect 20364 41500 20913 41528
rect 16574 41420 16580 41472
rect 16632 41420 16638 41472
rect 18322 41420 18328 41472
rect 18380 41460 18386 41472
rect 18877 41463 18935 41469
rect 18877 41460 18889 41463
rect 18380 41432 18889 41460
rect 18380 41420 18386 41432
rect 18877 41429 18889 41432
rect 18923 41460 18935 41463
rect 19426 41460 19432 41472
rect 18923 41432 19432 41460
rect 18923 41429 18935 41432
rect 18877 41423 18935 41429
rect 19426 41420 19432 41432
rect 19484 41420 19490 41472
rect 20364 41469 20392 41500
rect 20901 41497 20913 41500
rect 20947 41497 20959 41531
rect 20901 41491 20959 41497
rect 21358 41488 21364 41540
rect 21416 41488 21422 41540
rect 21545 41531 21603 41537
rect 21545 41497 21557 41531
rect 21591 41528 21603 41531
rect 21591 41500 21864 41528
rect 21591 41497 21603 41500
rect 21545 41491 21603 41497
rect 21836 41469 21864 41500
rect 22186 41488 22192 41540
rect 22244 41528 22250 41540
rect 22830 41528 22836 41540
rect 22244 41500 22836 41528
rect 22244 41488 22250 41500
rect 22830 41488 22836 41500
rect 22888 41528 22894 41540
rect 24670 41528 24676 41540
rect 22888 41500 24676 41528
rect 22888 41488 22894 41500
rect 24670 41488 24676 41500
rect 24728 41488 24734 41540
rect 25498 41488 25504 41540
rect 25556 41528 25562 41540
rect 26160 41528 26188 41627
rect 26878 41624 26884 41636
rect 26936 41624 26942 41676
rect 26973 41599 27031 41605
rect 26973 41565 26985 41599
rect 27019 41565 27031 41599
rect 26973 41559 27031 41565
rect 25556 41500 26188 41528
rect 25556 41488 25562 41500
rect 20349 41463 20407 41469
rect 20349 41429 20361 41463
rect 20395 41429 20407 41463
rect 20349 41423 20407 41429
rect 21821 41463 21879 41469
rect 21821 41429 21833 41463
rect 21867 41429 21879 41463
rect 21821 41423 21879 41429
rect 23750 41420 23756 41472
rect 23808 41420 23814 41472
rect 25682 41420 25688 41472
rect 25740 41420 25746 41472
rect 26988 41460 27016 41559
rect 27062 41556 27068 41608
rect 27120 41556 27126 41608
rect 27157 41599 27215 41605
rect 27157 41565 27169 41599
rect 27203 41565 27215 41599
rect 27264 41596 27292 41704
rect 27356 41704 28724 41732
rect 27356 41676 27384 41704
rect 28718 41692 28724 41704
rect 28776 41692 28782 41744
rect 29012 41732 29040 41772
rect 28828 41704 29040 41732
rect 29104 41704 30604 41732
rect 27338 41624 27344 41676
rect 27396 41624 27402 41676
rect 27614 41624 27620 41676
rect 27672 41624 27678 41676
rect 28828 41664 28856 41704
rect 29104 41673 29132 41704
rect 29089 41667 29147 41673
rect 29089 41664 29101 41667
rect 28644 41636 28856 41664
rect 28920 41636 29101 41664
rect 28166 41596 28172 41608
rect 27264 41568 28172 41596
rect 27157 41559 27215 41565
rect 27172 41528 27200 41559
rect 28166 41556 28172 41568
rect 28224 41556 28230 41608
rect 28353 41599 28411 41605
rect 28353 41565 28365 41599
rect 28399 41596 28411 41599
rect 28644 41596 28672 41636
rect 28399 41568 28672 41596
rect 28399 41565 28411 41568
rect 28353 41559 28411 41565
rect 28718 41556 28724 41608
rect 28776 41596 28782 41608
rect 28813 41599 28871 41605
rect 28813 41596 28825 41599
rect 28776 41568 28825 41596
rect 28776 41556 28782 41568
rect 28813 41565 28825 41568
rect 28859 41565 28871 41599
rect 28813 41559 28871 41565
rect 27798 41528 27804 41540
rect 27172 41500 27804 41528
rect 27798 41488 27804 41500
rect 27856 41528 27862 41540
rect 28445 41531 28503 41537
rect 28445 41528 28457 41531
rect 27856 41500 28457 41528
rect 27856 41488 27862 41500
rect 28445 41497 28457 41500
rect 28491 41528 28503 41531
rect 28534 41528 28540 41540
rect 28491 41500 28540 41528
rect 28491 41497 28503 41500
rect 28445 41491 28503 41497
rect 28534 41488 28540 41500
rect 28592 41488 28598 41540
rect 28629 41463 28687 41469
rect 28629 41460 28641 41463
rect 26988 41432 28641 41460
rect 28629 41429 28641 41432
rect 28675 41460 28687 41463
rect 28920 41460 28948 41636
rect 29089 41633 29101 41636
rect 29135 41633 29147 41667
rect 29089 41627 29147 41633
rect 30466 41556 30472 41608
rect 30524 41556 30530 41608
rect 30576 41605 30604 41704
rect 30668 41664 30696 41772
rect 30834 41760 30840 41812
rect 30892 41760 30898 41812
rect 30926 41760 30932 41812
rect 30984 41800 30990 41812
rect 32214 41800 32220 41812
rect 30984 41772 32220 41800
rect 30984 41760 30990 41772
rect 32214 41760 32220 41772
rect 32272 41800 32278 41812
rect 32858 41800 32864 41812
rect 32272 41772 32864 41800
rect 32272 41760 32278 41772
rect 32858 41760 32864 41772
rect 32916 41800 32922 41812
rect 33042 41800 33048 41812
rect 32916 41772 33048 41800
rect 32916 41760 32922 41772
rect 33042 41760 33048 41772
rect 33100 41760 33106 41812
rect 33137 41803 33195 41809
rect 33137 41769 33149 41803
rect 33183 41769 33195 41803
rect 33137 41763 33195 41769
rect 30745 41735 30803 41741
rect 30745 41701 30757 41735
rect 30791 41732 30803 41735
rect 31110 41732 31116 41744
rect 30791 41704 31116 41732
rect 30791 41701 30803 41704
rect 30745 41695 30803 41701
rect 31110 41692 31116 41704
rect 31168 41692 31174 41744
rect 33152 41732 33180 41763
rect 34790 41760 34796 41812
rect 34848 41760 34854 41812
rect 35342 41760 35348 41812
rect 35400 41760 35406 41812
rect 36354 41800 36360 41812
rect 35866 41772 36360 41800
rect 32232 41704 33180 41732
rect 35253 41735 35311 41741
rect 32122 41664 32128 41676
rect 30668 41636 32128 41664
rect 32122 41624 32128 41636
rect 32180 41624 32186 41676
rect 30561 41599 30619 41605
rect 30561 41565 30573 41599
rect 30607 41596 30619 41599
rect 30926 41596 30932 41608
rect 30607 41568 30932 41596
rect 30607 41565 30619 41568
rect 30561 41559 30619 41565
rect 30926 41556 30932 41568
rect 30984 41556 30990 41608
rect 31021 41599 31079 41605
rect 31021 41565 31033 41599
rect 31067 41565 31079 41599
rect 31021 41559 31079 41565
rect 30742 41488 30748 41540
rect 30800 41488 30806 41540
rect 28675 41432 28948 41460
rect 28675 41429 28687 41432
rect 28629 41423 28687 41429
rect 29086 41420 29092 41472
rect 29144 41420 29150 41472
rect 31036 41460 31064 41559
rect 31110 41556 31116 41608
rect 31168 41556 31174 41608
rect 31202 41556 31208 41608
rect 31260 41596 31266 41608
rect 31481 41599 31539 41605
rect 31481 41596 31493 41599
rect 31260 41568 31493 41596
rect 31260 41556 31266 41568
rect 31481 41565 31493 41568
rect 31527 41565 31539 41599
rect 31481 41559 31539 41565
rect 31570 41556 31576 41608
rect 31628 41556 31634 41608
rect 31757 41599 31815 41605
rect 31757 41565 31769 41599
rect 31803 41565 31815 41599
rect 31757 41559 31815 41565
rect 31389 41531 31447 41537
rect 31389 41497 31401 41531
rect 31435 41528 31447 41531
rect 31588 41528 31616 41556
rect 31435 41500 31616 41528
rect 31435 41497 31447 41500
rect 31389 41491 31447 41497
rect 31662 41488 31668 41540
rect 31720 41528 31726 41540
rect 31772 41528 31800 41559
rect 31846 41556 31852 41608
rect 31904 41556 31910 41608
rect 31938 41556 31944 41608
rect 31996 41556 32002 41608
rect 32030 41556 32036 41608
rect 32088 41556 32094 41608
rect 32232 41528 32260 41704
rect 35253 41701 35265 41735
rect 35299 41732 35311 41735
rect 35618 41732 35624 41744
rect 35299 41704 35624 41732
rect 35299 41701 35311 41704
rect 35253 41695 35311 41701
rect 35618 41692 35624 41704
rect 35676 41692 35682 41744
rect 35866 41664 35894 41772
rect 36354 41760 36360 41772
rect 36412 41760 36418 41812
rect 36449 41803 36507 41809
rect 36449 41769 36461 41803
rect 36495 41800 36507 41803
rect 36630 41800 36636 41812
rect 36495 41772 36636 41800
rect 36495 41769 36507 41772
rect 36449 41763 36507 41769
rect 36630 41760 36636 41772
rect 36688 41760 36694 41812
rect 32692 41636 33180 41664
rect 32398 41556 32404 41608
rect 32456 41596 32462 41608
rect 32692 41605 32720 41636
rect 32677 41599 32735 41605
rect 32677 41596 32689 41599
rect 32456 41568 32689 41596
rect 32456 41556 32462 41568
rect 32677 41565 32689 41568
rect 32723 41565 32735 41599
rect 32677 41559 32735 41565
rect 32766 41556 32772 41608
rect 32824 41556 32830 41608
rect 32858 41556 32864 41608
rect 32916 41556 32922 41608
rect 32950 41556 32956 41608
rect 33008 41556 33014 41608
rect 33152 41605 33180 41636
rect 34992 41636 35894 41664
rect 36096 41704 36676 41732
rect 33137 41599 33195 41605
rect 33137 41565 33149 41599
rect 33183 41565 33195 41599
rect 33137 41559 33195 41565
rect 33229 41599 33287 41605
rect 33229 41565 33241 41599
rect 33275 41565 33287 41599
rect 33229 41559 33287 41565
rect 33244 41528 33272 41559
rect 34514 41556 34520 41608
rect 34572 41596 34578 41608
rect 34992 41605 35020 41636
rect 35636 41605 35664 41636
rect 34701 41599 34759 41605
rect 34701 41596 34713 41599
rect 34572 41568 34713 41596
rect 34572 41556 34578 41568
rect 34701 41565 34713 41568
rect 34747 41565 34759 41599
rect 34701 41559 34759 41565
rect 34977 41599 35035 41605
rect 34977 41565 34989 41599
rect 35023 41565 35035 41599
rect 34977 41559 35035 41565
rect 35529 41599 35587 41605
rect 35529 41565 35541 41599
rect 35575 41565 35587 41599
rect 35529 41559 35587 41565
rect 35621 41599 35679 41605
rect 35621 41565 35633 41599
rect 35667 41565 35679 41599
rect 35621 41559 35679 41565
rect 34992 41528 35020 41559
rect 31720 41500 32260 41528
rect 32416 41500 33272 41528
rect 33520 41500 35020 41528
rect 35253 41531 35311 41537
rect 31720 41488 31726 41500
rect 31573 41463 31631 41469
rect 31573 41460 31585 41463
rect 31036 41432 31585 41460
rect 31573 41429 31585 41432
rect 31619 41429 31631 41463
rect 31573 41423 31631 41429
rect 31846 41420 31852 41472
rect 31904 41460 31910 41472
rect 32416 41460 32444 41500
rect 31904 41432 32444 41460
rect 32493 41463 32551 41469
rect 31904 41420 31910 41432
rect 32493 41429 32505 41463
rect 32539 41460 32551 41463
rect 32674 41460 32680 41472
rect 32539 41432 32680 41460
rect 32539 41429 32551 41432
rect 32493 41423 32551 41429
rect 32674 41420 32680 41432
rect 32732 41420 32738 41472
rect 33520 41469 33548 41500
rect 35253 41497 35265 41531
rect 35299 41528 35311 41531
rect 35544 41528 35572 41559
rect 35710 41556 35716 41608
rect 35768 41556 35774 41608
rect 35805 41599 35863 41605
rect 35805 41565 35817 41599
rect 35851 41596 35863 41599
rect 35894 41596 35900 41608
rect 35851 41568 35900 41596
rect 35851 41565 35863 41568
rect 35805 41559 35863 41565
rect 35894 41556 35900 41568
rect 35952 41556 35958 41608
rect 35299 41500 35572 41528
rect 35728 41528 35756 41556
rect 36096 41528 36124 41704
rect 36262 41624 36268 41676
rect 36320 41624 36326 41676
rect 36648 41673 36676 41704
rect 36633 41667 36691 41673
rect 36633 41633 36645 41667
rect 36679 41633 36691 41667
rect 36633 41627 36691 41633
rect 36173 41599 36231 41605
rect 36173 41565 36185 41599
rect 36219 41565 36231 41599
rect 36173 41559 36231 41565
rect 35728 41500 36124 41528
rect 36188 41528 36216 41559
rect 36814 41556 36820 41608
rect 36872 41556 36878 41608
rect 36906 41556 36912 41608
rect 36964 41556 36970 41608
rect 36633 41531 36691 41537
rect 36633 41528 36645 41531
rect 36188 41500 36645 41528
rect 35299 41497 35311 41500
rect 35253 41491 35311 41497
rect 33505 41463 33563 41469
rect 33505 41429 33517 41463
rect 33551 41429 33563 41463
rect 33505 41423 33563 41429
rect 35066 41420 35072 41472
rect 35124 41460 35130 41472
rect 35434 41460 35440 41472
rect 35124 41432 35440 41460
rect 35124 41420 35130 41432
rect 35434 41420 35440 41432
rect 35492 41420 35498 41472
rect 35544 41460 35572 41500
rect 36633 41497 36645 41500
rect 36679 41497 36691 41531
rect 36633 41491 36691 41497
rect 36814 41460 36820 41472
rect 35544 41432 36820 41460
rect 36814 41420 36820 41432
rect 36872 41420 36878 41472
rect 1104 41370 42504 41392
rect 1104 41318 4874 41370
rect 4926 41318 4938 41370
rect 4990 41318 5002 41370
rect 5054 41318 5066 41370
rect 5118 41318 5130 41370
rect 5182 41318 35594 41370
rect 35646 41318 35658 41370
rect 35710 41318 35722 41370
rect 35774 41318 35786 41370
rect 35838 41318 35850 41370
rect 35902 41318 42504 41370
rect 1104 41296 42504 41318
rect 15378 41216 15384 41268
rect 15436 41256 15442 41268
rect 15565 41259 15623 41265
rect 15565 41256 15577 41259
rect 15436 41228 15577 41256
rect 15436 41216 15442 41228
rect 15565 41225 15577 41228
rect 15611 41225 15623 41259
rect 15565 41219 15623 41225
rect 17420 41228 19288 41256
rect 16025 41191 16083 41197
rect 16025 41157 16037 41191
rect 16071 41188 16083 41191
rect 17034 41188 17040 41200
rect 16071 41160 17040 41188
rect 16071 41157 16083 41160
rect 16025 41151 16083 41157
rect 17034 41148 17040 41160
rect 17092 41188 17098 41200
rect 17420 41197 17448 41228
rect 17405 41191 17463 41197
rect 17405 41188 17417 41191
rect 17092 41160 17417 41188
rect 17092 41148 17098 41160
rect 17405 41157 17417 41160
rect 17451 41157 17463 41191
rect 17405 41151 17463 41157
rect 17586 41148 17592 41200
rect 17644 41197 17650 41200
rect 17644 41191 17663 41197
rect 17651 41157 17663 41191
rect 17644 41151 17663 41157
rect 17644 41148 17650 41151
rect 15933 41123 15991 41129
rect 15933 41089 15945 41123
rect 15979 41120 15991 41123
rect 16669 41123 16727 41129
rect 16669 41120 16681 41123
rect 15979 41092 16681 41120
rect 15979 41089 15991 41092
rect 15933 41083 15991 41089
rect 16669 41089 16681 41092
rect 16715 41089 16727 41123
rect 16669 41083 16727 41089
rect 17954 41080 17960 41132
rect 18012 41080 18018 41132
rect 19145 41123 19203 41129
rect 19145 41120 19157 41123
rect 19076 41110 19157 41120
rect 18892 41092 19157 41110
rect 18892 41082 19104 41092
rect 19145 41089 19157 41092
rect 19191 41089 19203 41123
rect 19260 41120 19288 41228
rect 19426 41216 19432 41268
rect 19484 41216 19490 41268
rect 19978 41216 19984 41268
rect 20036 41216 20042 41268
rect 23477 41259 23535 41265
rect 23477 41225 23489 41259
rect 23523 41256 23535 41259
rect 23750 41256 23756 41268
rect 23523 41228 23756 41256
rect 23523 41225 23535 41228
rect 23477 41219 23535 41225
rect 23750 41216 23756 41228
rect 23808 41216 23814 41268
rect 25866 41216 25872 41268
rect 25924 41256 25930 41268
rect 25924 41228 27016 41256
rect 25924 41216 25930 41228
rect 19318 41191 19376 41197
rect 19318 41157 19330 41191
rect 19364 41188 19376 41191
rect 19444 41188 19472 41216
rect 24026 41188 24032 41200
rect 19364 41160 19472 41188
rect 22940 41160 24032 41188
rect 19364 41157 19376 41160
rect 19318 41151 19376 41157
rect 22940 41132 22968 41160
rect 24026 41148 24032 41160
rect 24084 41148 24090 41200
rect 26988 41197 27016 41228
rect 27338 41216 27344 41268
rect 27396 41216 27402 41268
rect 28813 41259 28871 41265
rect 28813 41225 28825 41259
rect 28859 41256 28871 41259
rect 28859 41228 29224 41256
rect 28859 41225 28871 41228
rect 28813 41219 28871 41225
rect 26973 41191 27031 41197
rect 26973 41157 26985 41191
rect 27019 41157 27031 41191
rect 26973 41151 27031 41157
rect 27614 41148 27620 41200
rect 27672 41188 27678 41200
rect 28902 41188 28908 41200
rect 27672 41160 28908 41188
rect 27672 41148 27678 41160
rect 19429 41123 19487 41129
rect 19429 41120 19441 41123
rect 19260 41092 19441 41120
rect 19145 41083 19203 41089
rect 19429 41089 19441 41092
rect 19475 41089 19487 41123
rect 19429 41083 19487 41089
rect 19522 41123 19580 41129
rect 19522 41089 19534 41123
rect 19568 41089 19580 41123
rect 19889 41123 19947 41129
rect 19889 41120 19901 41123
rect 19522 41083 19580 41089
rect 19812 41092 19901 41120
rect 16209 41055 16267 41061
rect 16209 41021 16221 41055
rect 16255 41021 16267 41055
rect 16209 41015 16267 41021
rect 16224 40984 16252 41015
rect 16574 41012 16580 41064
rect 16632 41052 16638 41064
rect 17221 41055 17279 41061
rect 17221 41052 17233 41055
rect 16632 41024 17233 41052
rect 16632 41012 16638 41024
rect 17221 41021 17233 41024
rect 17267 41021 17279 41055
rect 17221 41015 17279 41021
rect 18138 41012 18144 41064
rect 18196 41052 18202 41064
rect 18693 41055 18751 41061
rect 18693 41052 18705 41055
rect 18196 41024 18705 41052
rect 18196 41012 18202 41024
rect 18693 41021 18705 41024
rect 18739 41052 18751 41055
rect 18782 41052 18788 41064
rect 18739 41024 18788 41052
rect 18739 41021 18751 41024
rect 18693 41015 18751 41021
rect 18782 41012 18788 41024
rect 18840 41012 18846 41064
rect 18046 40984 18052 40996
rect 16224 40956 18052 40984
rect 18046 40944 18052 40956
rect 18104 40984 18110 40996
rect 18892 40984 18920 41082
rect 19242 41012 19248 41064
rect 19300 41052 19306 41064
rect 19536 41052 19564 41083
rect 19300 41024 19564 41052
rect 19300 41012 19306 41024
rect 19812 40996 19840 41092
rect 19889 41089 19901 41092
rect 19935 41089 19947 41123
rect 19889 41083 19947 41089
rect 20073 41123 20131 41129
rect 20073 41089 20085 41123
rect 20119 41089 20131 41123
rect 20073 41083 20131 41089
rect 19978 41012 19984 41064
rect 20036 41052 20042 41064
rect 20088 41052 20116 41083
rect 20898 41080 20904 41132
rect 20956 41120 20962 41132
rect 22554 41120 22560 41132
rect 20956 41092 22560 41120
rect 20956 41080 20962 41092
rect 22554 41080 22560 41092
rect 22612 41120 22618 41132
rect 22649 41123 22707 41129
rect 22649 41120 22661 41123
rect 22612 41092 22661 41120
rect 22612 41080 22618 41092
rect 22649 41089 22661 41092
rect 22695 41089 22707 41123
rect 22649 41083 22707 41089
rect 22833 41123 22891 41129
rect 22833 41089 22845 41123
rect 22879 41120 22891 41123
rect 22922 41120 22928 41132
rect 22879 41092 22928 41120
rect 22879 41089 22891 41092
rect 22833 41083 22891 41089
rect 22922 41080 22928 41092
rect 22980 41080 22986 41132
rect 23109 41123 23167 41129
rect 23109 41089 23121 41123
rect 23155 41089 23167 41123
rect 23382 41120 23388 41132
rect 23109 41083 23167 41089
rect 23216 41092 23388 41120
rect 20990 41052 20996 41064
rect 20036 41024 20996 41052
rect 20036 41012 20042 41024
rect 20990 41012 20996 41024
rect 21048 41012 21054 41064
rect 22741 41055 22799 41061
rect 22741 41021 22753 41055
rect 22787 41052 22799 41055
rect 23124 41052 23152 41083
rect 23216 41061 23244 41092
rect 23382 41080 23388 41092
rect 23440 41120 23446 41132
rect 23569 41123 23627 41129
rect 23569 41120 23581 41123
rect 23440 41092 23581 41120
rect 23440 41080 23446 41092
rect 23569 41089 23581 41092
rect 23615 41089 23627 41123
rect 23569 41083 23627 41089
rect 23750 41080 23756 41132
rect 23808 41080 23814 41132
rect 24762 41080 24768 41132
rect 24820 41080 24826 41132
rect 27908 41129 27936 41160
rect 28902 41148 28908 41160
rect 28960 41148 28966 41200
rect 29196 41197 29224 41228
rect 30484 41228 34100 41256
rect 29181 41191 29239 41197
rect 29181 41157 29193 41191
rect 29227 41157 29239 41191
rect 29181 41151 29239 41157
rect 29638 41148 29644 41200
rect 29696 41148 29702 41200
rect 27157 41123 27215 41129
rect 26068 41092 26174 41120
rect 22787 41024 23152 41052
rect 23201 41055 23259 41061
rect 22787 41021 22799 41024
rect 22741 41015 22799 41021
rect 23201 41021 23213 41055
rect 23247 41021 23259 41055
rect 23201 41015 23259 41021
rect 25038 41012 25044 41064
rect 25096 41012 25102 41064
rect 25590 41012 25596 41064
rect 25648 41052 25654 41064
rect 25774 41052 25780 41064
rect 25648 41024 25780 41052
rect 25648 41012 25654 41024
rect 25774 41012 25780 41024
rect 25832 41052 25838 41064
rect 26068 41052 26096 41092
rect 27157 41089 27169 41123
rect 27203 41089 27215 41123
rect 27157 41083 27215 41089
rect 27893 41123 27951 41129
rect 27893 41089 27905 41123
rect 27939 41089 27951 41123
rect 28445 41123 28503 41129
rect 28445 41120 28457 41123
rect 27893 41083 27951 41089
rect 28092 41092 28457 41120
rect 27172 41052 27200 41083
rect 25832 41024 26096 41052
rect 26160 41024 27200 41052
rect 25832 41012 25838 41024
rect 18104 40956 19334 40984
rect 18104 40944 18110 40956
rect 17494 40876 17500 40928
rect 17552 40916 17558 40928
rect 17589 40919 17647 40925
rect 17589 40916 17601 40919
rect 17552 40888 17601 40916
rect 17552 40876 17558 40888
rect 17589 40885 17601 40888
rect 17635 40885 17647 40919
rect 17589 40879 17647 40885
rect 17770 40876 17776 40928
rect 17828 40876 17834 40928
rect 17862 40876 17868 40928
rect 17920 40916 17926 40928
rect 18969 40919 19027 40925
rect 18969 40916 18981 40919
rect 17920 40888 18981 40916
rect 17920 40876 17926 40888
rect 18969 40885 18981 40888
rect 19015 40885 19027 40919
rect 19306 40916 19334 40956
rect 19794 40944 19800 40996
rect 19852 40944 19858 40996
rect 26160 40928 26188 41024
rect 21082 40916 21088 40928
rect 19306 40888 21088 40916
rect 18969 40879 19027 40885
rect 21082 40876 21088 40888
rect 21140 40876 21146 40928
rect 23937 40919 23995 40925
rect 23937 40885 23949 40919
rect 23983 40916 23995 40919
rect 26142 40916 26148 40928
rect 23983 40888 26148 40916
rect 23983 40885 23995 40888
rect 23937 40879 23995 40885
rect 26142 40876 26148 40888
rect 26200 40876 26206 40928
rect 26234 40876 26240 40928
rect 26292 40916 26298 40928
rect 26513 40919 26571 40925
rect 26513 40916 26525 40919
rect 26292 40888 26525 40916
rect 26292 40876 26298 40888
rect 26513 40885 26525 40888
rect 26559 40885 26571 40919
rect 28092 40916 28120 41092
rect 28445 41089 28457 41092
rect 28491 41089 28503 41123
rect 28445 41083 28503 41089
rect 28166 41012 28172 41064
rect 28224 41052 28230 41064
rect 28261 41055 28319 41061
rect 28261 41052 28273 41055
rect 28224 41024 28273 41052
rect 28224 41012 28230 41024
rect 28261 41021 28273 41024
rect 28307 41021 28319 41055
rect 28261 41015 28319 41021
rect 28276 40984 28304 41015
rect 28350 41012 28356 41064
rect 28408 41012 28414 41064
rect 28902 41012 28908 41064
rect 28960 41012 28966 41064
rect 30484 41052 30512 41228
rect 31662 41188 31668 41200
rect 31588 41160 31668 41188
rect 30742 41080 30748 41132
rect 30800 41120 30806 41132
rect 31110 41120 31116 41132
rect 30800 41092 31116 41120
rect 30800 41080 30806 41092
rect 31110 41080 31116 41092
rect 31168 41120 31174 41132
rect 31588 41129 31616 41160
rect 31662 41148 31668 41160
rect 31720 41148 31726 41200
rect 31757 41191 31815 41197
rect 31757 41157 31769 41191
rect 31803 41188 31815 41191
rect 31846 41188 31852 41200
rect 31803 41160 31852 41188
rect 31803 41157 31815 41160
rect 31757 41151 31815 41157
rect 31573 41123 31631 41129
rect 31573 41120 31585 41123
rect 31168 41092 31585 41120
rect 31168 41080 31174 41092
rect 31573 41089 31585 41092
rect 31619 41089 31631 41123
rect 31573 41083 31631 41089
rect 29012 41024 30512 41052
rect 29012 40984 29040 41024
rect 30558 41012 30564 41064
rect 30616 41052 30622 41064
rect 31772 41052 31800 41151
rect 31846 41148 31852 41160
rect 31904 41148 31910 41200
rect 31941 41191 31999 41197
rect 31941 41157 31953 41191
rect 31987 41188 31999 41191
rect 32766 41188 32772 41200
rect 31987 41160 32772 41188
rect 31987 41157 31999 41160
rect 31941 41151 31999 41157
rect 32140 41129 32168 41160
rect 32766 41148 32772 41160
rect 32824 41148 32830 41200
rect 33226 41148 33232 41200
rect 33284 41148 33290 41200
rect 32125 41123 32183 41129
rect 32125 41089 32137 41123
rect 32171 41089 32183 41123
rect 32125 41083 32183 41089
rect 32214 41080 32220 41132
rect 32272 41080 32278 41132
rect 32398 41080 32404 41132
rect 32456 41080 32462 41132
rect 34072 41120 34100 41228
rect 34146 41148 34152 41200
rect 34204 41188 34210 41200
rect 36170 41188 36176 41200
rect 34204 41160 36176 41188
rect 34204 41148 34210 41160
rect 36170 41148 36176 41160
rect 36228 41188 36234 41200
rect 36722 41188 36728 41200
rect 36228 41160 36728 41188
rect 36228 41148 36234 41160
rect 36722 41148 36728 41160
rect 36780 41148 36786 41200
rect 36081 41123 36139 41129
rect 34072 41092 35894 41120
rect 30616 41024 31800 41052
rect 30616 41012 30622 41024
rect 32490 41012 32496 41064
rect 32548 41012 32554 41064
rect 32769 41055 32827 41061
rect 32769 41021 32781 41055
rect 32815 41052 32827 41055
rect 32858 41052 32864 41064
rect 32815 41024 32864 41052
rect 32815 41021 32827 41024
rect 32769 41015 32827 41021
rect 32858 41012 32864 41024
rect 32916 41012 32922 41064
rect 33134 41012 33140 41064
rect 33192 41052 33198 41064
rect 34698 41052 34704 41064
rect 33192 41024 34704 41052
rect 33192 41012 33198 41024
rect 34698 41012 34704 41024
rect 34756 41052 34762 41064
rect 35066 41052 35072 41064
rect 34756 41024 35072 41052
rect 34756 41012 34762 41024
rect 35066 41012 35072 41024
rect 35124 41012 35130 41064
rect 28276 40956 29040 40984
rect 35866 40984 35894 41092
rect 36081 41089 36093 41123
rect 36127 41120 36139 41123
rect 36262 41120 36268 41132
rect 36127 41092 36268 41120
rect 36127 41089 36139 41092
rect 36081 41083 36139 41089
rect 36262 41080 36268 41092
rect 36320 41120 36326 41132
rect 37182 41120 37188 41132
rect 36320 41092 37188 41120
rect 36320 41080 36326 41092
rect 37182 41080 37188 41092
rect 37240 41080 37246 41132
rect 37274 41080 37280 41132
rect 37332 41120 37338 41132
rect 38194 41120 38200 41132
rect 37332 41092 38200 41120
rect 37332 41080 37338 41092
rect 38194 41080 38200 41092
rect 38252 41080 38258 41132
rect 35989 41055 36047 41061
rect 35989 41021 36001 41055
rect 36035 41052 36047 41055
rect 36354 41052 36360 41064
rect 36035 41024 36360 41052
rect 36035 41021 36047 41024
rect 35989 41015 36047 41021
rect 36354 41012 36360 41024
rect 36412 41052 36418 41064
rect 36906 41052 36912 41064
rect 36412 41024 36912 41052
rect 36412 41012 36418 41024
rect 36906 41012 36912 41024
rect 36964 41012 36970 41064
rect 36538 40984 36544 40996
rect 35866 40956 36544 40984
rect 36538 40944 36544 40956
rect 36596 40984 36602 40996
rect 37366 40984 37372 40996
rect 36596 40956 37372 40984
rect 36596 40944 36602 40956
rect 37366 40944 37372 40956
rect 37424 40944 37430 40996
rect 30558 40916 30564 40928
rect 28092 40888 30564 40916
rect 26513 40879 26571 40885
rect 30558 40876 30564 40888
rect 30616 40916 30622 40928
rect 30653 40919 30711 40925
rect 30653 40916 30665 40919
rect 30616 40888 30665 40916
rect 30616 40876 30622 40888
rect 30653 40885 30665 40888
rect 30699 40885 30711 40919
rect 30653 40879 30711 40885
rect 32401 40919 32459 40925
rect 32401 40885 32413 40919
rect 32447 40916 32459 40919
rect 32766 40916 32772 40928
rect 32447 40888 32772 40916
rect 32447 40885 32459 40888
rect 32401 40879 32459 40885
rect 32766 40876 32772 40888
rect 32824 40876 32830 40928
rect 33318 40876 33324 40928
rect 33376 40916 33382 40928
rect 34241 40919 34299 40925
rect 34241 40916 34253 40919
rect 33376 40888 34253 40916
rect 33376 40876 33382 40888
rect 34241 40885 34253 40888
rect 34287 40885 34299 40919
rect 34241 40879 34299 40885
rect 35342 40876 35348 40928
rect 35400 40916 35406 40928
rect 35713 40919 35771 40925
rect 35713 40916 35725 40919
rect 35400 40888 35725 40916
rect 35400 40876 35406 40888
rect 35713 40885 35725 40888
rect 35759 40885 35771 40919
rect 35713 40879 35771 40885
rect 36081 40919 36139 40925
rect 36081 40885 36093 40919
rect 36127 40916 36139 40919
rect 36814 40916 36820 40928
rect 36127 40888 36820 40916
rect 36127 40885 36139 40888
rect 36081 40879 36139 40885
rect 36814 40876 36820 40888
rect 36872 40876 36878 40928
rect 1104 40826 42504 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 42504 40826
rect 1104 40752 42504 40774
rect 1302 40672 1308 40724
rect 1360 40712 1366 40724
rect 17126 40712 17132 40724
rect 1360 40684 17132 40712
rect 1360 40672 1366 40684
rect 17126 40672 17132 40684
rect 17184 40672 17190 40724
rect 17313 40715 17371 40721
rect 17313 40681 17325 40715
rect 17359 40712 17371 40715
rect 17402 40712 17408 40724
rect 17359 40684 17408 40712
rect 17359 40681 17371 40684
rect 17313 40675 17371 40681
rect 17402 40672 17408 40684
rect 17460 40672 17466 40724
rect 17494 40672 17500 40724
rect 17552 40712 17558 40724
rect 19978 40712 19984 40724
rect 17552 40684 19984 40712
rect 17552 40672 17558 40684
rect 19978 40672 19984 40684
rect 20036 40672 20042 40724
rect 20070 40672 20076 40724
rect 20128 40712 20134 40724
rect 20533 40715 20591 40721
rect 20533 40712 20545 40715
rect 20128 40684 20545 40712
rect 20128 40672 20134 40684
rect 20533 40681 20545 40684
rect 20579 40681 20591 40715
rect 20533 40675 20591 40681
rect 20898 40672 20904 40724
rect 20956 40672 20962 40724
rect 20993 40715 21051 40721
rect 20993 40681 21005 40715
rect 21039 40712 21051 40715
rect 21082 40712 21088 40724
rect 21039 40684 21088 40712
rect 21039 40681 21051 40684
rect 20993 40675 21051 40681
rect 21082 40672 21088 40684
rect 21140 40672 21146 40724
rect 25038 40672 25044 40724
rect 25096 40712 25102 40724
rect 25317 40715 25375 40721
rect 25317 40712 25329 40715
rect 25096 40684 25329 40712
rect 25096 40672 25102 40684
rect 25317 40681 25329 40684
rect 25363 40681 25375 40715
rect 25317 40675 25375 40681
rect 25866 40672 25872 40724
rect 25924 40712 25930 40724
rect 27433 40715 27491 40721
rect 27433 40712 27445 40715
rect 25924 40684 27445 40712
rect 25924 40672 25930 40684
rect 27433 40681 27445 40684
rect 27479 40681 27491 40715
rect 27433 40675 27491 40681
rect 28350 40672 28356 40724
rect 28408 40712 28414 40724
rect 28445 40715 28503 40721
rect 28445 40712 28457 40715
rect 28408 40684 28457 40712
rect 28408 40672 28414 40684
rect 28445 40681 28457 40684
rect 28491 40681 28503 40715
rect 28445 40675 28503 40681
rect 32493 40715 32551 40721
rect 32493 40681 32505 40715
rect 32539 40712 32551 40715
rect 32858 40712 32864 40724
rect 32539 40684 32864 40712
rect 32539 40681 32551 40684
rect 32493 40675 32551 40681
rect 32858 40672 32864 40684
rect 32916 40672 32922 40724
rect 33226 40672 33232 40724
rect 33284 40712 33290 40724
rect 34146 40712 34152 40724
rect 33284 40684 34152 40712
rect 33284 40672 33290 40684
rect 34146 40672 34152 40684
rect 34204 40672 34210 40724
rect 35529 40715 35587 40721
rect 35529 40712 35541 40715
rect 35176 40684 35541 40712
rect 17221 40647 17279 40653
rect 17221 40613 17233 40647
rect 17267 40644 17279 40647
rect 17681 40647 17739 40653
rect 17681 40644 17693 40647
rect 17267 40616 17693 40644
rect 17267 40613 17279 40616
rect 17221 40607 17279 40613
rect 17681 40613 17693 40616
rect 17727 40613 17739 40647
rect 17681 40607 17739 40613
rect 17770 40604 17776 40656
rect 17828 40604 17834 40656
rect 20441 40647 20499 40653
rect 20441 40613 20453 40647
rect 20487 40644 20499 40647
rect 20806 40644 20812 40656
rect 20487 40616 20812 40644
rect 20487 40613 20499 40616
rect 20441 40607 20499 40613
rect 20806 40604 20812 40616
rect 20864 40644 20870 40656
rect 26053 40647 26111 40653
rect 20864 40616 22048 40644
rect 20864 40604 20870 40616
rect 17402 40576 17408 40588
rect 16960 40548 17408 40576
rect 16960 40517 16988 40548
rect 17402 40536 17408 40548
rect 17460 40536 17466 40588
rect 17589 40579 17647 40585
rect 17589 40545 17601 40579
rect 17635 40576 17647 40579
rect 17788 40576 17816 40604
rect 17635 40548 17816 40576
rect 17635 40545 17647 40548
rect 17589 40539 17647 40545
rect 19794 40536 19800 40588
rect 19852 40576 19858 40588
rect 22020 40585 22048 40616
rect 26053 40613 26065 40647
rect 26099 40613 26111 40647
rect 26053 40607 26111 40613
rect 27893 40647 27951 40653
rect 27893 40613 27905 40647
rect 27939 40644 27951 40647
rect 30466 40644 30472 40656
rect 27939 40616 30472 40644
rect 27939 40613 27951 40616
rect 27893 40607 27951 40613
rect 20625 40579 20683 40585
rect 20625 40576 20637 40579
rect 19852 40548 20637 40576
rect 19852 40536 19858 40548
rect 16945 40511 17003 40517
rect 16945 40477 16957 40511
rect 16991 40477 17003 40511
rect 16945 40471 17003 40477
rect 17034 40468 17040 40520
rect 17092 40468 17098 40520
rect 17497 40511 17555 40517
rect 17497 40477 17509 40511
rect 17543 40508 17555 40511
rect 17773 40511 17831 40517
rect 17543 40480 17724 40508
rect 17543 40477 17555 40480
rect 17497 40471 17555 40477
rect 17221 40443 17279 40449
rect 17221 40409 17233 40443
rect 17267 40440 17279 40443
rect 17586 40440 17592 40452
rect 17267 40412 17592 40440
rect 17267 40409 17279 40412
rect 17221 40403 17279 40409
rect 17586 40400 17592 40412
rect 17644 40400 17650 40452
rect 17696 40440 17724 40480
rect 17773 40477 17785 40511
rect 17819 40508 17831 40511
rect 17862 40508 17868 40520
rect 17819 40480 17868 40508
rect 17819 40477 17831 40480
rect 17773 40471 17831 40477
rect 17862 40468 17868 40480
rect 17920 40468 17926 40520
rect 18138 40468 18144 40520
rect 18196 40468 18202 40520
rect 20272 40517 20300 40548
rect 20625 40545 20637 40548
rect 20671 40545 20683 40579
rect 20625 40539 20683 40545
rect 21177 40579 21235 40585
rect 21177 40545 21189 40579
rect 21223 40576 21235 40579
rect 21729 40579 21787 40585
rect 21729 40576 21741 40579
rect 21223 40548 21741 40576
rect 21223 40545 21235 40548
rect 21177 40539 21235 40545
rect 21729 40545 21741 40548
rect 21775 40545 21787 40579
rect 21729 40539 21787 40545
rect 22005 40579 22063 40585
rect 22005 40545 22017 40579
rect 22051 40545 22063 40579
rect 22005 40539 22063 40545
rect 22094 40536 22100 40588
rect 22152 40576 22158 40588
rect 22922 40576 22928 40588
rect 22152 40548 22928 40576
rect 22152 40536 22158 40548
rect 22922 40536 22928 40548
rect 22980 40536 22986 40588
rect 25501 40579 25559 40585
rect 25501 40545 25513 40579
rect 25547 40576 25559 40579
rect 25682 40576 25688 40588
rect 25547 40548 25688 40576
rect 25547 40545 25559 40548
rect 25501 40539 25559 40545
rect 25682 40536 25688 40548
rect 25740 40536 25746 40588
rect 25958 40536 25964 40588
rect 26016 40536 26022 40588
rect 20257 40511 20315 40517
rect 20257 40477 20269 40511
rect 20303 40477 20315 40511
rect 20257 40471 20315 40477
rect 20533 40511 20591 40517
rect 20533 40477 20545 40511
rect 20579 40477 20591 40511
rect 20533 40471 20591 40477
rect 18782 40440 18788 40452
rect 17696 40412 18788 40440
rect 18782 40400 18788 40412
rect 18840 40400 18846 40452
rect 20070 40400 20076 40452
rect 20128 40400 20134 40452
rect 20548 40440 20576 40471
rect 21266 40468 21272 40520
rect 21324 40468 21330 40520
rect 21913 40511 21971 40517
rect 21913 40508 21925 40511
rect 21376 40480 21925 40508
rect 20622 40440 20628 40452
rect 20548 40412 20628 40440
rect 20622 40400 20628 40412
rect 20680 40440 20686 40452
rect 21376 40440 21404 40480
rect 21913 40477 21925 40480
rect 21959 40477 21971 40511
rect 21913 40471 21971 40477
rect 22189 40511 22247 40517
rect 22189 40477 22201 40511
rect 22235 40508 22247 40511
rect 25593 40511 25651 40517
rect 22235 40480 25544 40508
rect 22235 40477 22247 40480
rect 22189 40471 22247 40477
rect 20680 40412 21404 40440
rect 21545 40443 21603 40449
rect 20680 40400 20686 40412
rect 21545 40409 21557 40443
rect 21591 40409 21603 40443
rect 21545 40403 21603 40409
rect 21637 40443 21695 40449
rect 21637 40409 21649 40443
rect 21683 40440 21695 40443
rect 21818 40440 21824 40452
rect 21683 40412 21824 40440
rect 21683 40409 21695 40412
rect 21637 40403 21695 40409
rect 18800 40372 18828 40400
rect 21560 40372 21588 40403
rect 21818 40400 21824 40412
rect 21876 40400 21882 40452
rect 22204 40372 22232 40471
rect 25516 40452 25544 40480
rect 25593 40477 25605 40511
rect 25639 40508 25651 40511
rect 26068 40508 26096 40607
rect 30466 40604 30472 40616
rect 30524 40604 30530 40656
rect 31110 40604 31116 40656
rect 31168 40604 31174 40656
rect 34790 40604 34796 40656
rect 34848 40644 34854 40656
rect 34977 40647 35035 40653
rect 34977 40644 34989 40647
rect 34848 40616 34989 40644
rect 34848 40604 34854 40616
rect 34977 40613 34989 40616
rect 35023 40613 35035 40647
rect 34977 40607 35035 40613
rect 27617 40579 27675 40585
rect 27617 40545 27629 40579
rect 27663 40576 27675 40579
rect 27798 40576 27804 40588
rect 27663 40548 27804 40576
rect 27663 40545 27675 40548
rect 27617 40539 27675 40545
rect 27798 40536 27804 40548
rect 27856 40536 27862 40588
rect 28261 40579 28319 40585
rect 28261 40545 28273 40579
rect 28307 40576 28319 40579
rect 29086 40576 29092 40588
rect 28307 40548 29092 40576
rect 28307 40545 28319 40548
rect 28261 40539 28319 40545
rect 29086 40536 29092 40548
rect 29144 40536 29150 40588
rect 30650 40536 30656 40588
rect 30708 40536 30714 40588
rect 32674 40536 32680 40588
rect 32732 40536 32738 40588
rect 32950 40536 32956 40588
rect 33008 40576 33014 40588
rect 33045 40579 33103 40585
rect 33045 40576 33057 40579
rect 33008 40548 33057 40576
rect 33008 40536 33014 40548
rect 33045 40545 33057 40548
rect 33091 40545 33103 40579
rect 33045 40539 33103 40545
rect 25639 40480 26096 40508
rect 25639 40477 25651 40480
rect 25593 40471 25651 40477
rect 26142 40468 26148 40520
rect 26200 40508 26206 40520
rect 26329 40511 26387 40517
rect 26329 40508 26341 40511
rect 26200 40480 26341 40508
rect 26200 40468 26206 40480
rect 26329 40477 26341 40480
rect 26375 40508 26387 40511
rect 27709 40511 27767 40517
rect 27709 40508 27721 40511
rect 26375 40480 27721 40508
rect 26375 40477 26387 40480
rect 26329 40471 26387 40477
rect 27709 40477 27721 40480
rect 27755 40477 27767 40511
rect 27709 40471 27767 40477
rect 28166 40468 28172 40520
rect 28224 40468 28230 40520
rect 30742 40468 30748 40520
rect 30800 40468 30806 40520
rect 32766 40468 32772 40520
rect 32824 40468 32830 40520
rect 34698 40468 34704 40520
rect 34756 40508 34762 40520
rect 35176 40517 35204 40684
rect 35529 40681 35541 40684
rect 35575 40681 35587 40715
rect 35529 40675 35587 40681
rect 35805 40647 35863 40653
rect 35805 40644 35817 40647
rect 35360 40616 35817 40644
rect 35360 40520 35388 40616
rect 35805 40613 35817 40616
rect 35851 40613 35863 40647
rect 35805 40607 35863 40613
rect 36814 40604 36820 40656
rect 36872 40644 36878 40656
rect 37461 40647 37519 40653
rect 37461 40644 37473 40647
rect 36872 40616 37473 40644
rect 36872 40604 36878 40616
rect 37461 40613 37473 40616
rect 37507 40613 37519 40647
rect 37461 40607 37519 40613
rect 37921 40579 37979 40585
rect 37921 40545 37933 40579
rect 37967 40545 37979 40579
rect 37921 40539 37979 40545
rect 35161 40511 35219 40517
rect 35161 40508 35173 40511
rect 34756 40480 35173 40508
rect 34756 40468 34762 40480
rect 35161 40477 35173 40480
rect 35207 40477 35219 40511
rect 35161 40471 35219 40477
rect 35250 40468 35256 40520
rect 35308 40468 35314 40520
rect 35342 40468 35348 40520
rect 35400 40468 35406 40520
rect 35989 40511 36047 40517
rect 35989 40477 36001 40511
rect 36035 40477 36047 40511
rect 35989 40471 36047 40477
rect 25498 40400 25504 40452
rect 25556 40440 25562 40452
rect 25869 40443 25927 40449
rect 25869 40440 25881 40443
rect 25556 40412 25881 40440
rect 25556 40400 25562 40412
rect 25869 40409 25881 40412
rect 25915 40409 25927 40443
rect 25869 40403 25927 40409
rect 26050 40400 26056 40452
rect 26108 40400 26114 40452
rect 27433 40443 27491 40449
rect 27433 40409 27445 40443
rect 27479 40440 27491 40443
rect 28184 40440 28212 40468
rect 27479 40412 28212 40440
rect 33137 40443 33195 40449
rect 27479 40409 27491 40412
rect 27433 40403 27491 40409
rect 33137 40409 33149 40443
rect 33183 40440 33195 40443
rect 33318 40440 33324 40452
rect 33183 40412 33324 40440
rect 33183 40409 33195 40412
rect 33137 40403 33195 40409
rect 33318 40400 33324 40412
rect 33376 40400 33382 40452
rect 34977 40443 35035 40449
rect 34977 40409 34989 40443
rect 35023 40440 35035 40443
rect 35434 40440 35440 40452
rect 35023 40412 35440 40440
rect 35023 40409 35035 40412
rect 34977 40403 35035 40409
rect 35434 40400 35440 40412
rect 35492 40400 35498 40452
rect 36004 40384 36032 40471
rect 37826 40468 37832 40520
rect 37884 40468 37890 40520
rect 37936 40508 37964 40539
rect 38194 40536 38200 40588
rect 38252 40576 38258 40588
rect 38841 40579 38899 40585
rect 38841 40576 38853 40579
rect 38252 40548 38853 40576
rect 38252 40536 38258 40548
rect 38841 40545 38853 40548
rect 38887 40545 38899 40579
rect 38841 40539 38899 40545
rect 39298 40508 39304 40520
rect 37936 40480 39304 40508
rect 39298 40468 39304 40480
rect 39356 40468 39362 40520
rect 42150 40468 42156 40520
rect 42208 40468 42214 40520
rect 38102 40400 38108 40452
rect 38160 40400 38166 40452
rect 18800 40344 22232 40372
rect 26234 40332 26240 40384
rect 26292 40332 26298 40384
rect 31938 40332 31944 40384
rect 31996 40372 32002 40384
rect 34422 40372 34428 40384
rect 31996 40344 34428 40372
rect 31996 40332 32002 40344
rect 34422 40332 34428 40344
rect 34480 40372 34486 40384
rect 35986 40372 35992 40384
rect 34480 40344 35992 40372
rect 34480 40332 34486 40344
rect 35986 40332 35992 40344
rect 36044 40332 36050 40384
rect 41046 40332 41052 40384
rect 41104 40372 41110 40384
rect 41509 40375 41567 40381
rect 41509 40372 41521 40375
rect 41104 40344 41521 40372
rect 41104 40332 41110 40344
rect 41509 40341 41521 40344
rect 41555 40341 41567 40375
rect 41509 40335 41567 40341
rect 1104 40282 42504 40304
rect 1104 40230 4874 40282
rect 4926 40230 4938 40282
rect 4990 40230 5002 40282
rect 5054 40230 5066 40282
rect 5118 40230 5130 40282
rect 5182 40230 35594 40282
rect 35646 40230 35658 40282
rect 35710 40230 35722 40282
rect 35774 40230 35786 40282
rect 35838 40230 35850 40282
rect 35902 40230 42504 40282
rect 1104 40208 42504 40230
rect 17497 40171 17555 40177
rect 17497 40137 17509 40171
rect 17543 40168 17555 40171
rect 17586 40168 17592 40180
rect 17543 40140 17592 40168
rect 17543 40137 17555 40140
rect 17497 40131 17555 40137
rect 17586 40128 17592 40140
rect 17644 40128 17650 40180
rect 19429 40171 19487 40177
rect 19429 40137 19441 40171
rect 19475 40168 19487 40171
rect 20070 40168 20076 40180
rect 19475 40140 20076 40168
rect 19475 40137 19487 40140
rect 19429 40131 19487 40137
rect 20070 40128 20076 40140
rect 20128 40128 20134 40180
rect 20622 40128 20628 40180
rect 20680 40168 20686 40180
rect 20986 40171 21044 40177
rect 20680 40140 20944 40168
rect 20680 40128 20686 40140
rect 15948 40072 16160 40100
rect 14550 39992 14556 40044
rect 14608 40032 14614 40044
rect 15948 40032 15976 40072
rect 14608 40004 15976 40032
rect 14608 39992 14614 40004
rect 16022 39992 16028 40044
rect 16080 39992 16086 40044
rect 16132 40032 16160 40072
rect 20806 40060 20812 40112
rect 20864 40060 20870 40112
rect 20916 40100 20944 40140
rect 20986 40137 20998 40171
rect 21032 40168 21044 40171
rect 21266 40168 21272 40180
rect 21032 40140 21272 40168
rect 21032 40137 21044 40140
rect 20986 40131 21044 40137
rect 21266 40128 21272 40140
rect 21324 40128 21330 40180
rect 23382 40128 23388 40180
rect 23440 40168 23446 40180
rect 23477 40171 23535 40177
rect 23477 40168 23489 40171
rect 23440 40140 23489 40168
rect 23440 40128 23446 40140
rect 23477 40137 23489 40140
rect 23523 40137 23535 40171
rect 23477 40131 23535 40137
rect 25409 40171 25467 40177
rect 25409 40137 25421 40171
rect 25455 40168 25467 40171
rect 26050 40168 26056 40180
rect 25455 40140 26056 40168
rect 25455 40137 25467 40140
rect 25409 40131 25467 40137
rect 26050 40128 26056 40140
rect 26108 40128 26114 40180
rect 30742 40128 30748 40180
rect 30800 40128 30806 40180
rect 32398 40128 32404 40180
rect 32456 40168 32462 40180
rect 32677 40171 32735 40177
rect 32677 40168 32689 40171
rect 32456 40140 32689 40168
rect 32456 40128 32462 40140
rect 32677 40137 32689 40140
rect 32723 40137 32735 40171
rect 35342 40168 35348 40180
rect 32677 40131 32735 40137
rect 34440 40140 35348 40168
rect 21085 40103 21143 40109
rect 21085 40100 21097 40103
rect 20916 40072 21097 40100
rect 21085 40069 21097 40072
rect 21131 40069 21143 40103
rect 21085 40063 21143 40069
rect 26234 40060 26240 40112
rect 26292 40100 26298 40112
rect 34440 40100 34468 40140
rect 35342 40128 35348 40140
rect 35400 40128 35406 40180
rect 37001 40171 37059 40177
rect 37001 40137 37013 40171
rect 37047 40168 37059 40171
rect 37826 40168 37832 40180
rect 37047 40140 37832 40168
rect 37047 40137 37059 40140
rect 37001 40131 37059 40137
rect 37826 40128 37832 40140
rect 37884 40128 37890 40180
rect 36170 40100 36176 40112
rect 26292 40072 34468 40100
rect 35282 40072 36176 40100
rect 26292 40060 26298 40072
rect 36170 40060 36176 40072
rect 36228 40060 36234 40112
rect 38194 40060 38200 40112
rect 38252 40100 38258 40112
rect 38252 40072 39804 40100
rect 38252 40060 38258 40072
rect 20812 40057 20870 40060
rect 16298 40032 16304 40044
rect 16132 40004 16304 40032
rect 16298 39992 16304 40004
rect 16356 39992 16362 40044
rect 17126 39992 17132 40044
rect 17184 39992 17190 40044
rect 18598 39992 18604 40044
rect 18656 40032 18662 40044
rect 19061 40035 19119 40041
rect 19061 40032 19073 40035
rect 18656 40004 19073 40032
rect 18656 39992 18662 40004
rect 19061 40001 19073 40004
rect 19107 40001 19119 40035
rect 20812 40023 20824 40057
rect 20858 40023 20870 40057
rect 20812 40017 20870 40023
rect 20901 40035 20959 40041
rect 19061 39995 19119 40001
rect 20901 40001 20913 40035
rect 20947 40032 20959 40035
rect 20990 40032 20996 40044
rect 20947 40004 20996 40032
rect 20947 40001 20959 40004
rect 20901 39995 20959 40001
rect 20990 39992 20996 40004
rect 21048 40032 21054 40044
rect 22094 40032 22100 40044
rect 21048 40004 22100 40032
rect 21048 39992 21054 40004
rect 22094 39992 22100 40004
rect 22152 39992 22158 40044
rect 23106 39992 23112 40044
rect 23164 39992 23170 40044
rect 25038 39992 25044 40044
rect 25096 39992 25102 40044
rect 26510 39992 26516 40044
rect 26568 40032 26574 40044
rect 27157 40035 27215 40041
rect 27157 40032 27169 40035
rect 26568 40004 27169 40032
rect 26568 39992 26574 40004
rect 27157 40001 27169 40004
rect 27203 40001 27215 40035
rect 27157 39995 27215 40001
rect 30282 39992 30288 40044
rect 30340 40032 30346 40044
rect 30653 40035 30711 40041
rect 30653 40032 30665 40035
rect 30340 40004 30665 40032
rect 30340 39992 30346 40004
rect 30653 40001 30665 40004
rect 30699 40001 30711 40035
rect 30653 39995 30711 40001
rect 30837 40035 30895 40041
rect 30837 40001 30849 40035
rect 30883 40032 30895 40035
rect 31386 40032 31392 40044
rect 30883 40004 31392 40032
rect 30883 40001 30895 40004
rect 30837 39995 30895 40001
rect 31386 39992 31392 40004
rect 31444 39992 31450 40044
rect 32030 39992 32036 40044
rect 32088 40032 32094 40044
rect 32309 40035 32367 40041
rect 32309 40032 32321 40035
rect 32088 40004 32321 40032
rect 32088 39992 32094 40004
rect 32309 40001 32321 40004
rect 32355 40001 32367 40035
rect 32309 39995 32367 40001
rect 35342 39992 35348 40044
rect 35400 40032 35406 40044
rect 35897 40035 35955 40041
rect 35897 40032 35909 40035
rect 35400 40004 35909 40032
rect 35400 39992 35406 40004
rect 35897 40001 35909 40004
rect 35943 40001 35955 40035
rect 35897 39995 35955 40001
rect 35986 39992 35992 40044
rect 36044 39992 36050 40044
rect 36909 40035 36967 40041
rect 36909 40001 36921 40035
rect 36955 40001 36967 40035
rect 36909 39995 36967 40001
rect 37093 40035 37151 40041
rect 37093 40001 37105 40035
rect 37139 40001 37151 40035
rect 37093 39995 37151 40001
rect 12894 39924 12900 39976
rect 12952 39964 12958 39976
rect 13265 39967 13323 39973
rect 13265 39964 13277 39967
rect 12952 39936 13277 39964
rect 12952 39924 12958 39936
rect 13265 39933 13277 39936
rect 13311 39933 13323 39967
rect 13265 39927 13323 39933
rect 13538 39924 13544 39976
rect 13596 39924 13602 39976
rect 15657 39967 15715 39973
rect 15657 39964 15669 39967
rect 15028 39936 15669 39964
rect 14826 39788 14832 39840
rect 14884 39828 14890 39840
rect 15028 39837 15056 39936
rect 15657 39933 15669 39936
rect 15703 39964 15715 39967
rect 15933 39967 15991 39973
rect 15933 39964 15945 39967
rect 15703 39936 15945 39964
rect 15703 39933 15715 39936
rect 15657 39927 15715 39933
rect 15933 39933 15945 39936
rect 15979 39933 15991 39967
rect 15933 39927 15991 39933
rect 16393 39967 16451 39973
rect 16393 39933 16405 39967
rect 16439 39964 16451 39967
rect 17034 39964 17040 39976
rect 16439 39936 17040 39964
rect 16439 39933 16451 39936
rect 16393 39927 16451 39933
rect 17034 39924 17040 39936
rect 17092 39924 17098 39976
rect 17221 39967 17279 39973
rect 17221 39933 17233 39967
rect 17267 39964 17279 39967
rect 17310 39964 17316 39976
rect 17267 39936 17316 39964
rect 17267 39933 17279 39936
rect 17221 39927 17279 39933
rect 17310 39924 17316 39936
rect 17368 39924 17374 39976
rect 18690 39924 18696 39976
rect 18748 39964 18754 39976
rect 18969 39967 19027 39973
rect 18969 39964 18981 39967
rect 18748 39936 18981 39964
rect 18748 39924 18754 39936
rect 18969 39933 18981 39936
rect 19015 39933 19027 39967
rect 18969 39927 19027 39933
rect 23198 39924 23204 39976
rect 23256 39924 23262 39976
rect 25130 39924 25136 39976
rect 25188 39924 25194 39976
rect 26786 39924 26792 39976
rect 26844 39964 26850 39976
rect 27065 39967 27123 39973
rect 27065 39964 27077 39967
rect 26844 39936 27077 39964
rect 26844 39924 26850 39936
rect 27065 39933 27077 39936
rect 27111 39933 27123 39967
rect 27065 39927 27123 39933
rect 32214 39924 32220 39976
rect 32272 39924 32278 39976
rect 32398 39924 32404 39976
rect 32456 39964 32462 39976
rect 33781 39967 33839 39973
rect 33781 39964 33793 39967
rect 32456 39936 33793 39964
rect 32456 39924 32462 39936
rect 33781 39933 33793 39936
rect 33827 39933 33839 39967
rect 33781 39927 33839 39933
rect 34057 39967 34115 39973
rect 34057 39933 34069 39967
rect 34103 39964 34115 39967
rect 34698 39964 34704 39976
rect 34103 39936 34704 39964
rect 34103 39933 34115 39936
rect 34057 39927 34115 39933
rect 34698 39924 34704 39936
rect 34756 39924 34762 39976
rect 35434 39924 35440 39976
rect 35492 39964 35498 39976
rect 35805 39967 35863 39973
rect 35805 39964 35817 39967
rect 35492 39936 35817 39964
rect 35492 39924 35498 39936
rect 35805 39933 35817 39936
rect 35851 39933 35863 39967
rect 35805 39927 35863 39933
rect 36078 39924 36084 39976
rect 36136 39924 36142 39976
rect 27525 39899 27583 39905
rect 27525 39865 27537 39899
rect 27571 39896 27583 39899
rect 27798 39896 27804 39908
rect 27571 39868 27804 39896
rect 27571 39865 27583 39868
rect 27525 39859 27583 39865
rect 27798 39856 27804 39868
rect 27856 39856 27862 39908
rect 35986 39856 35992 39908
rect 36044 39896 36050 39908
rect 36924 39896 36952 39995
rect 36998 39896 37004 39908
rect 36044 39868 37004 39896
rect 36044 39856 36050 39868
rect 36998 39856 37004 39868
rect 37056 39856 37062 39908
rect 15013 39831 15071 39837
rect 15013 39828 15025 39831
rect 14884 39800 15025 39828
rect 14884 39788 14890 39800
rect 15013 39797 15025 39800
rect 15059 39797 15071 39831
rect 15013 39791 15071 39797
rect 15102 39788 15108 39840
rect 15160 39788 15166 39840
rect 20714 39788 20720 39840
rect 20772 39828 20778 39840
rect 21542 39828 21548 39840
rect 20772 39800 21548 39828
rect 20772 39788 20778 39800
rect 21542 39788 21548 39800
rect 21600 39788 21606 39840
rect 35526 39788 35532 39840
rect 35584 39788 35590 39840
rect 35618 39788 35624 39840
rect 35676 39788 35682 39840
rect 35710 39788 35716 39840
rect 35768 39828 35774 39840
rect 37108 39828 37136 39995
rect 37182 39992 37188 40044
rect 37240 40032 37246 40044
rect 38381 40035 38439 40041
rect 37240 40004 38056 40032
rect 37240 39992 37246 40004
rect 37274 39924 37280 39976
rect 37332 39924 37338 39976
rect 38028 39905 38056 40004
rect 38381 40001 38393 40035
rect 38427 40032 38439 40035
rect 38657 40035 38715 40041
rect 38657 40032 38669 40035
rect 38427 40004 38669 40032
rect 38427 40001 38439 40004
rect 38381 39995 38439 40001
rect 38657 40001 38669 40004
rect 38703 40001 38715 40035
rect 38657 39995 38715 40001
rect 38853 40035 38911 40041
rect 38853 40001 38865 40035
rect 38899 40032 38911 40035
rect 39117 40035 39175 40041
rect 38899 40004 39068 40032
rect 38899 40001 38911 40004
rect 38853 39995 38911 40001
rect 38470 39924 38476 39976
rect 38528 39924 38534 39976
rect 39040 39964 39068 40004
rect 39117 40001 39129 40035
rect 39163 40032 39175 40035
rect 39574 40032 39580 40044
rect 39163 40004 39580 40032
rect 39163 40001 39175 40004
rect 39117 39995 39175 40001
rect 39574 39992 39580 40004
rect 39632 39992 39638 40044
rect 39666 39992 39672 40044
rect 39724 39992 39730 40044
rect 39776 40032 39804 40072
rect 40037 40035 40095 40041
rect 40037 40032 40049 40035
rect 39776 40004 40049 40032
rect 40037 40001 40049 40004
rect 40083 40001 40095 40035
rect 40037 39995 40095 40001
rect 41414 39992 41420 40044
rect 41472 39992 41478 40044
rect 39040 39936 39160 39964
rect 38013 39899 38071 39905
rect 38013 39865 38025 39899
rect 38059 39865 38071 39899
rect 38013 39859 38071 39865
rect 38930 39856 38936 39908
rect 38988 39856 38994 39908
rect 39022 39856 39028 39908
rect 39080 39856 39086 39908
rect 39132 39896 39160 39936
rect 39298 39924 39304 39976
rect 39356 39924 39362 39976
rect 40310 39924 40316 39976
rect 40368 39924 40374 39976
rect 39666 39896 39672 39908
rect 39132 39868 39672 39896
rect 39666 39856 39672 39868
rect 39724 39856 39730 39908
rect 37734 39828 37740 39840
rect 35768 39800 37740 39828
rect 35768 39788 35774 39800
rect 37734 39788 37740 39800
rect 37792 39788 37798 39840
rect 37918 39788 37924 39840
rect 37976 39788 37982 39840
rect 41782 39788 41788 39840
rect 41840 39788 41846 39840
rect 1104 39738 42504 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 42504 39738
rect 1104 39664 42504 39686
rect 13173 39627 13231 39633
rect 13173 39593 13185 39627
rect 13219 39624 13231 39627
rect 13538 39624 13544 39636
rect 13219 39596 13544 39624
rect 13219 39593 13231 39596
rect 13173 39587 13231 39593
rect 13538 39584 13544 39596
rect 13596 39584 13602 39636
rect 18138 39624 18144 39636
rect 15488 39596 18144 39624
rect 13725 39491 13783 39497
rect 13725 39457 13737 39491
rect 13771 39488 13783 39491
rect 14734 39488 14740 39500
rect 13771 39460 14740 39488
rect 13771 39457 13783 39460
rect 13725 39451 13783 39457
rect 14734 39448 14740 39460
rect 14792 39448 14798 39500
rect 14826 39448 14832 39500
rect 14884 39448 14890 39500
rect 15488 39497 15516 39596
rect 18138 39584 18144 39596
rect 18196 39624 18202 39636
rect 18196 39596 20852 39624
rect 18196 39584 18202 39596
rect 17310 39516 17316 39568
rect 17368 39516 17374 39568
rect 18233 39559 18291 39565
rect 17512 39528 18092 39556
rect 15473 39491 15531 39497
rect 15473 39457 15485 39491
rect 15519 39457 15531 39491
rect 15473 39451 15531 39457
rect 17126 39448 17132 39500
rect 17184 39488 17190 39500
rect 17512 39488 17540 39528
rect 17184 39460 17540 39488
rect 17184 39448 17190 39460
rect 17586 39448 17592 39500
rect 17644 39488 17650 39500
rect 17644 39460 18000 39488
rect 17644 39448 17650 39460
rect 13541 39423 13599 39429
rect 13541 39389 13553 39423
rect 13587 39420 13599 39423
rect 15102 39420 15108 39432
rect 13587 39392 15108 39420
rect 13587 39389 13599 39392
rect 13541 39383 13599 39389
rect 15102 39380 15108 39392
rect 15160 39380 15166 39432
rect 17972 39429 18000 39460
rect 17681 39423 17739 39429
rect 17681 39389 17693 39423
rect 17727 39389 17739 39423
rect 17681 39383 17739 39389
rect 17957 39423 18015 39429
rect 17957 39389 17969 39423
rect 18003 39389 18015 39423
rect 18064 39420 18092 39528
rect 18233 39525 18245 39559
rect 18279 39525 18291 39559
rect 18233 39519 18291 39525
rect 18248 39488 18276 39519
rect 18598 39516 18604 39568
rect 18656 39516 18662 39568
rect 18690 39516 18696 39568
rect 18748 39516 18754 39568
rect 20533 39559 20591 39565
rect 20533 39525 20545 39559
rect 20579 39556 20591 39559
rect 20622 39556 20628 39568
rect 20579 39528 20628 39556
rect 20579 39525 20591 39528
rect 20533 39519 20591 39525
rect 20622 39516 20628 39528
rect 20680 39516 20686 39568
rect 19242 39488 19248 39500
rect 18248 39460 19248 39488
rect 18233 39423 18291 39429
rect 18233 39420 18245 39423
rect 18064 39392 18245 39420
rect 17957 39383 18015 39389
rect 18233 39389 18245 39392
rect 18279 39389 18291 39423
rect 18233 39383 18291 39389
rect 14921 39355 14979 39361
rect 14921 39321 14933 39355
rect 14967 39352 14979 39355
rect 15194 39352 15200 39364
rect 14967 39324 15200 39352
rect 14967 39321 14979 39324
rect 14921 39315 14979 39321
rect 15194 39312 15200 39324
rect 15252 39312 15258 39364
rect 15746 39312 15752 39364
rect 15804 39312 15810 39364
rect 16298 39312 16304 39364
rect 16356 39312 16362 39364
rect 17494 39352 17500 39364
rect 17236 39324 17500 39352
rect 13633 39287 13691 39293
rect 13633 39253 13645 39287
rect 13679 39284 13691 39287
rect 13998 39284 14004 39296
rect 13679 39256 14004 39284
rect 13679 39253 13691 39256
rect 13633 39247 13691 39253
rect 13998 39244 14004 39256
rect 14056 39244 14062 39296
rect 15013 39287 15071 39293
rect 15013 39253 15025 39287
rect 15059 39284 15071 39287
rect 15102 39284 15108 39296
rect 15059 39256 15108 39284
rect 15059 39253 15071 39256
rect 15013 39247 15071 39253
rect 15102 39244 15108 39256
rect 15160 39244 15166 39296
rect 15381 39287 15439 39293
rect 15381 39253 15393 39287
rect 15427 39284 15439 39287
rect 17126 39284 17132 39296
rect 15427 39256 17132 39284
rect 15427 39253 15439 39256
rect 15381 39247 15439 39253
rect 17126 39244 17132 39256
rect 17184 39244 17190 39296
rect 17236 39293 17264 39324
rect 17494 39312 17500 39324
rect 17552 39352 17558 39364
rect 17696 39352 17724 39383
rect 18414 39380 18420 39432
rect 18472 39380 18478 39432
rect 18616 39429 18644 39460
rect 19242 39448 19248 39460
rect 19300 39488 19306 39500
rect 19613 39491 19671 39497
rect 19613 39488 19625 39491
rect 19300 39460 19625 39488
rect 19300 39448 19306 39460
rect 19613 39457 19625 39460
rect 19659 39457 19671 39491
rect 19613 39451 19671 39457
rect 20254 39448 20260 39500
rect 20312 39448 20318 39500
rect 20824 39497 20852 39596
rect 23106 39584 23112 39636
rect 23164 39584 23170 39636
rect 24213 39627 24271 39633
rect 23308 39596 23980 39624
rect 23198 39516 23204 39568
rect 23256 39516 23262 39568
rect 20809 39491 20867 39497
rect 20809 39457 20821 39491
rect 20855 39457 20867 39491
rect 20809 39451 20867 39457
rect 21082 39448 21088 39500
rect 21140 39448 21146 39500
rect 21818 39448 21824 39500
rect 21876 39488 21882 39500
rect 22557 39491 22615 39497
rect 22557 39488 22569 39491
rect 21876 39460 22569 39488
rect 21876 39448 21882 39460
rect 22557 39457 22569 39460
rect 22603 39457 22615 39491
rect 23308 39488 23336 39596
rect 23842 39556 23848 39568
rect 22557 39451 22615 39457
rect 22940 39460 23336 39488
rect 23400 39528 23848 39556
rect 22940 39432 22968 39460
rect 18601 39423 18659 39429
rect 18601 39389 18613 39423
rect 18647 39389 18659 39423
rect 18601 39383 18659 39389
rect 18968 39423 19026 39429
rect 18968 39389 18980 39423
rect 19014 39389 19026 39423
rect 18968 39383 19026 39389
rect 19061 39423 19119 39429
rect 19061 39389 19073 39423
rect 19107 39420 19119 39423
rect 19426 39420 19432 39432
rect 19107 39392 19432 39420
rect 19107 39389 19119 39392
rect 19061 39383 19119 39389
rect 18049 39355 18107 39361
rect 18049 39352 18061 39355
rect 17552 39324 18061 39352
rect 17552 39312 17558 39324
rect 18049 39321 18061 39324
rect 18095 39321 18107 39355
rect 18984 39352 19012 39383
rect 19426 39380 19432 39392
rect 19484 39380 19490 39432
rect 19518 39380 19524 39432
rect 19576 39380 19582 39432
rect 19702 39380 19708 39432
rect 19760 39380 19766 39432
rect 19889 39423 19947 39429
rect 19889 39389 19901 39423
rect 19935 39389 19947 39423
rect 19889 39383 19947 39389
rect 19720 39352 19748 39380
rect 18984 39324 19748 39352
rect 19904 39352 19932 39383
rect 20162 39380 20168 39432
rect 20220 39380 20226 39432
rect 22922 39380 22928 39432
rect 22980 39380 22986 39432
rect 23109 39423 23167 39429
rect 23109 39389 23121 39423
rect 23155 39420 23167 39423
rect 23400 39420 23428 39528
rect 23842 39516 23848 39528
rect 23900 39516 23906 39568
rect 23952 39497 23980 39596
rect 24213 39593 24225 39627
rect 24259 39624 24271 39627
rect 25038 39624 25044 39636
rect 24259 39596 25044 39624
rect 24259 39593 24271 39596
rect 24213 39587 24271 39593
rect 25038 39584 25044 39596
rect 25096 39584 25102 39636
rect 25130 39584 25136 39636
rect 25188 39584 25194 39636
rect 26510 39584 26516 39636
rect 26568 39584 26574 39636
rect 26786 39584 26792 39636
rect 26844 39584 26850 39636
rect 28166 39584 28172 39636
rect 28224 39584 28230 39636
rect 30561 39627 30619 39633
rect 30561 39593 30573 39627
rect 30607 39624 30619 39627
rect 30650 39624 30656 39636
rect 30607 39596 30656 39624
rect 30607 39593 30619 39596
rect 30561 39587 30619 39593
rect 30650 39584 30656 39596
rect 30708 39584 30714 39636
rect 31018 39584 31024 39636
rect 31076 39624 31082 39636
rect 31938 39624 31944 39636
rect 31076 39596 31944 39624
rect 31076 39584 31082 39596
rect 31938 39584 31944 39596
rect 31996 39584 32002 39636
rect 32030 39584 32036 39636
rect 32088 39624 32094 39636
rect 32125 39627 32183 39633
rect 32125 39624 32137 39627
rect 32088 39596 32137 39624
rect 32088 39584 32094 39596
rect 32125 39593 32137 39596
rect 32171 39593 32183 39627
rect 32125 39587 32183 39593
rect 32214 39584 32220 39636
rect 32272 39584 32278 39636
rect 34698 39584 34704 39636
rect 34756 39584 34762 39636
rect 35986 39624 35992 39636
rect 34808 39596 35992 39624
rect 24670 39516 24676 39568
rect 24728 39556 24734 39568
rect 24765 39559 24823 39565
rect 24765 39556 24777 39559
rect 24728 39528 24777 39556
rect 24728 39516 24734 39528
rect 24765 39525 24777 39528
rect 24811 39525 24823 39559
rect 24765 39519 24823 39525
rect 25222 39516 25228 39568
rect 25280 39516 25286 39568
rect 27246 39556 27252 39568
rect 26528 39528 27252 39556
rect 23937 39491 23995 39497
rect 23492 39460 23796 39488
rect 23492 39429 23520 39460
rect 23768 39432 23796 39460
rect 23937 39457 23949 39491
rect 23983 39488 23995 39491
rect 24302 39488 24308 39500
rect 23983 39460 24308 39488
rect 23983 39457 23995 39460
rect 23937 39451 23995 39457
rect 24302 39448 24308 39460
rect 24360 39448 24366 39500
rect 25240 39488 25268 39516
rect 26528 39488 26556 39528
rect 27246 39516 27252 39528
rect 27304 39516 27310 39568
rect 28534 39516 28540 39568
rect 28592 39516 28598 39568
rect 29178 39516 29184 39568
rect 29236 39556 29242 39568
rect 30282 39556 30288 39568
rect 29236 39528 30288 39556
rect 29236 39516 29242 39528
rect 30282 39516 30288 39528
rect 30340 39556 30346 39568
rect 31113 39559 31171 39565
rect 31113 39556 31125 39559
rect 30340 39528 31125 39556
rect 30340 39516 30346 39528
rect 31113 39525 31125 39528
rect 31159 39556 31171 39559
rect 31849 39559 31907 39565
rect 31849 39556 31861 39559
rect 31159 39528 31861 39556
rect 31159 39525 31171 39528
rect 31113 39519 31171 39525
rect 31849 39525 31861 39528
rect 31895 39525 31907 39559
rect 31849 39519 31907 39525
rect 32306 39516 32312 39568
rect 32364 39516 32370 39568
rect 34808 39556 34836 39596
rect 35986 39584 35992 39596
rect 36044 39584 36050 39636
rect 36078 39584 36084 39636
rect 36136 39584 36142 39636
rect 36998 39584 37004 39636
rect 37056 39624 37062 39636
rect 38930 39624 38936 39636
rect 37056 39596 38936 39624
rect 37056 39584 37062 39596
rect 36096 39556 36124 39584
rect 38580 39565 38608 39596
rect 38930 39584 38936 39596
rect 38988 39584 38994 39636
rect 39574 39584 39580 39636
rect 39632 39584 39638 39636
rect 42150 39624 42156 39636
rect 40512 39596 42156 39624
rect 38565 39559 38623 39565
rect 32692 39528 34836 39556
rect 35268 39528 36124 39556
rect 37936 39528 38332 39556
rect 27341 39491 27399 39497
rect 27341 39488 27353 39491
rect 24412 39460 25268 39488
rect 25884 39460 26556 39488
rect 23155 39392 23428 39420
rect 23476 39423 23534 39429
rect 23155 39389 23167 39392
rect 23109 39383 23167 39389
rect 23476 39389 23488 39423
rect 23522 39389 23534 39423
rect 23476 39383 23534 39389
rect 23569 39423 23627 39429
rect 23569 39389 23581 39423
rect 23615 39389 23627 39423
rect 23569 39383 23627 39389
rect 20990 39352 20996 39364
rect 19904 39324 20996 39352
rect 18049 39315 18107 39321
rect 20990 39312 20996 39324
rect 21048 39312 21054 39364
rect 21542 39312 21548 39364
rect 21600 39312 21606 39364
rect 17221 39287 17279 39293
rect 17221 39253 17233 39287
rect 17267 39253 17279 39287
rect 17221 39247 17279 39253
rect 19245 39287 19303 39293
rect 19245 39253 19257 39287
rect 19291 39284 19303 39287
rect 23124 39284 23152 39383
rect 23584 39296 23612 39383
rect 23750 39380 23756 39432
rect 23808 39380 23814 39432
rect 24026 39380 24032 39432
rect 24084 39380 24090 39432
rect 24412 39429 24440 39460
rect 24397 39423 24455 39429
rect 24397 39389 24409 39423
rect 24443 39389 24455 39423
rect 24397 39383 24455 39389
rect 24578 39380 24584 39432
rect 24636 39380 24642 39432
rect 24673 39423 24731 39429
rect 24673 39389 24685 39423
rect 24719 39389 24731 39423
rect 24673 39383 24731 39389
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39389 24915 39423
rect 24857 39383 24915 39389
rect 25041 39423 25099 39429
rect 25041 39389 25053 39423
rect 25087 39420 25099 39423
rect 25884 39420 25912 39460
rect 26528 39429 26556 39460
rect 26804 39460 27353 39488
rect 26329 39423 26387 39429
rect 26329 39420 26341 39423
rect 25087 39392 25912 39420
rect 25976 39392 26341 39420
rect 25087 39389 25099 39392
rect 25041 39383 25099 39389
rect 24118 39312 24124 39364
rect 24176 39352 24182 39364
rect 24688 39352 24716 39383
rect 24176 39324 24716 39352
rect 24176 39312 24182 39324
rect 19291 39256 23152 39284
rect 19291 39253 19303 39256
rect 19245 39247 19303 39253
rect 23566 39244 23572 39296
rect 23624 39284 23630 39296
rect 24026 39284 24032 39296
rect 23624 39256 24032 39284
rect 23624 39244 23630 39256
rect 24026 39244 24032 39256
rect 24084 39284 24090 39296
rect 24872 39284 24900 39383
rect 25976 39364 26004 39392
rect 26329 39389 26341 39392
rect 26375 39389 26387 39423
rect 26329 39383 26387 39389
rect 26513 39423 26571 39429
rect 26513 39389 26525 39423
rect 26559 39389 26571 39423
rect 26513 39383 26571 39389
rect 25593 39355 25651 39361
rect 25593 39321 25605 39355
rect 25639 39352 25651 39355
rect 25958 39352 25964 39364
rect 25639 39324 25964 39352
rect 25639 39321 25651 39324
rect 25593 39315 25651 39321
rect 25958 39312 25964 39324
rect 26016 39312 26022 39364
rect 26344 39352 26372 39383
rect 26804 39352 26832 39460
rect 27341 39457 27353 39460
rect 27387 39457 27399 39491
rect 27341 39451 27399 39457
rect 27985 39491 28043 39497
rect 27985 39457 27997 39491
rect 28031 39488 28043 39491
rect 28353 39491 28411 39497
rect 28353 39488 28365 39491
rect 28031 39460 28365 39488
rect 28031 39457 28043 39460
rect 27985 39451 28043 39457
rect 28353 39457 28365 39460
rect 28399 39457 28411 39491
rect 28353 39451 28411 39457
rect 30834 39448 30840 39500
rect 30892 39448 30898 39500
rect 31205 39491 31263 39497
rect 31205 39457 31217 39491
rect 31251 39488 31263 39491
rect 31386 39488 31392 39500
rect 31251 39460 31392 39488
rect 31251 39457 31263 39460
rect 31205 39451 31263 39457
rect 31386 39448 31392 39460
rect 31444 39448 31450 39500
rect 32324 39488 32352 39516
rect 31496 39460 32352 39488
rect 26880 39423 26938 39429
rect 26880 39389 26892 39423
rect 26926 39389 26938 39423
rect 26880 39383 26938 39389
rect 26973 39423 27031 39429
rect 26973 39389 26985 39423
rect 27019 39389 27031 39423
rect 26973 39383 27031 39389
rect 26344 39324 26832 39352
rect 24084 39256 24900 39284
rect 26896 39284 26924 39383
rect 26988 39352 27016 39383
rect 27154 39380 27160 39432
rect 27212 39380 27218 39432
rect 27433 39423 27491 39429
rect 27433 39389 27445 39423
rect 27479 39420 27491 39423
rect 27522 39420 27528 39432
rect 27479 39392 27528 39420
rect 27479 39389 27491 39392
rect 27433 39383 27491 39389
rect 27448 39352 27476 39383
rect 27522 39380 27528 39392
rect 27580 39380 27586 39432
rect 27617 39423 27675 39429
rect 27617 39389 27629 39423
rect 27663 39420 27675 39423
rect 27893 39423 27951 39429
rect 27893 39420 27905 39423
rect 27663 39392 27905 39420
rect 27663 39389 27675 39392
rect 27617 39383 27675 39389
rect 27893 39389 27905 39392
rect 27939 39389 27951 39423
rect 27893 39383 27951 39389
rect 30652 39423 30710 39429
rect 30652 39389 30664 39423
rect 30698 39389 30710 39423
rect 30652 39383 30710 39389
rect 30745 39423 30803 39429
rect 30745 39389 30757 39423
rect 30791 39420 30803 39423
rect 31018 39420 31024 39432
rect 30791 39392 31024 39420
rect 30791 39389 30803 39392
rect 30745 39383 30803 39389
rect 26988 39324 27476 39352
rect 28813 39355 28871 39361
rect 28813 39321 28825 39355
rect 28859 39352 28871 39355
rect 29178 39352 29184 39364
rect 28859 39324 29184 39352
rect 28859 39321 28871 39324
rect 28813 39315 28871 39321
rect 29178 39312 29184 39324
rect 29236 39312 29242 39364
rect 27154 39284 27160 39296
rect 26896 39256 27160 39284
rect 24084 39244 24090 39256
rect 27154 39244 27160 39256
rect 27212 39244 27218 39296
rect 30667 39284 30695 39383
rect 31018 39380 31024 39392
rect 31076 39380 31082 39432
rect 31496 39429 31524 39460
rect 32490 39448 32496 39500
rect 32548 39488 32554 39500
rect 32692 39497 32720 39528
rect 32677 39491 32735 39497
rect 32677 39488 32689 39491
rect 32548 39460 32689 39488
rect 32548 39448 32554 39460
rect 32677 39457 32689 39460
rect 32723 39457 32735 39491
rect 32677 39451 32735 39457
rect 34790 39448 34796 39500
rect 34848 39488 34854 39500
rect 35268 39497 35296 39528
rect 35253 39491 35311 39497
rect 34848 39460 35020 39488
rect 34848 39448 34854 39460
rect 31297 39423 31355 39429
rect 31297 39414 31309 39423
rect 31220 39389 31309 39414
rect 31343 39389 31355 39423
rect 31220 39386 31355 39389
rect 31220 39284 31248 39386
rect 31297 39383 31355 39386
rect 31481 39423 31539 39429
rect 31481 39389 31493 39423
rect 31527 39389 31539 39423
rect 31481 39383 31539 39389
rect 31662 39380 31668 39432
rect 31720 39380 31726 39432
rect 31754 39380 31760 39432
rect 31812 39380 31818 39432
rect 31938 39380 31944 39432
rect 31996 39380 32002 39432
rect 34992 39429 35020 39460
rect 35253 39457 35265 39491
rect 35299 39457 35311 39491
rect 35253 39451 35311 39457
rect 35713 39491 35771 39497
rect 35713 39457 35725 39491
rect 35759 39488 35771 39491
rect 36078 39488 36084 39500
rect 35759 39460 36084 39488
rect 35759 39457 35771 39460
rect 35713 39451 35771 39457
rect 36078 39448 36084 39460
rect 36136 39448 36142 39500
rect 37734 39448 37740 39500
rect 37792 39488 37798 39500
rect 37936 39488 37964 39528
rect 37792 39460 37964 39488
rect 38013 39491 38071 39497
rect 37792 39448 37798 39460
rect 38013 39457 38025 39491
rect 38059 39488 38071 39491
rect 38194 39488 38200 39500
rect 38059 39460 38200 39488
rect 38059 39457 38071 39460
rect 38013 39451 38071 39457
rect 38194 39448 38200 39460
rect 38252 39448 38258 39500
rect 38304 39488 38332 39528
rect 38565 39525 38577 39559
rect 38611 39525 38623 39559
rect 39022 39556 39028 39568
rect 38565 39519 38623 39525
rect 38672 39528 39028 39556
rect 38672 39497 38700 39528
rect 39022 39516 39028 39528
rect 39080 39516 39086 39568
rect 38657 39491 38715 39497
rect 38657 39488 38669 39491
rect 38304 39460 38669 39488
rect 38657 39457 38669 39460
rect 38703 39457 38715 39491
rect 39592 39488 39620 39584
rect 40512 39556 40540 39596
rect 42150 39584 42156 39596
rect 42208 39584 42214 39636
rect 38657 39451 38715 39457
rect 38764 39460 39620 39488
rect 40328 39528 40540 39556
rect 34885 39423 34943 39429
rect 34885 39389 34897 39423
rect 34931 39389 34943 39423
rect 34885 39383 34943 39389
rect 34977 39423 35035 39429
rect 34977 39389 34989 39423
rect 35023 39389 35035 39423
rect 35618 39420 35624 39432
rect 34977 39383 35035 39389
rect 35084 39392 35624 39420
rect 34900 39352 34928 39383
rect 35084 39352 35112 39392
rect 35618 39380 35624 39392
rect 35676 39380 35682 39432
rect 35805 39423 35863 39429
rect 35805 39389 35817 39423
rect 35851 39420 35863 39423
rect 35986 39420 35992 39432
rect 35851 39392 35992 39420
rect 35851 39389 35863 39392
rect 35805 39383 35863 39389
rect 35986 39380 35992 39392
rect 36044 39380 36050 39432
rect 36170 39380 36176 39432
rect 36228 39420 36234 39432
rect 38764 39429 38792 39460
rect 38473 39423 38531 39429
rect 36228 39392 36662 39420
rect 36228 39380 36234 39392
rect 38473 39389 38485 39423
rect 38519 39389 38531 39423
rect 38473 39383 38531 39389
rect 38749 39423 38807 39429
rect 38749 39389 38761 39423
rect 38795 39389 38807 39423
rect 38749 39383 38807 39389
rect 34900 39324 35112 39352
rect 35345 39355 35403 39361
rect 35345 39321 35357 39355
rect 35391 39352 35403 39355
rect 35526 39352 35532 39364
rect 35391 39324 35532 39352
rect 35391 39321 35403 39324
rect 35345 39315 35403 39321
rect 31662 39284 31668 39296
rect 30667 39256 31668 39284
rect 31662 39244 31668 39256
rect 31720 39284 31726 39296
rect 32766 39284 32772 39296
rect 31720 39256 32772 39284
rect 31720 39244 31726 39256
rect 32766 39244 32772 39256
rect 32824 39244 32830 39296
rect 34606 39244 34612 39296
rect 34664 39284 34670 39296
rect 35360 39284 35388 39315
rect 35526 39312 35532 39324
rect 35584 39312 35590 39364
rect 37458 39312 37464 39364
rect 37516 39352 37522 39364
rect 37737 39355 37795 39361
rect 37737 39352 37749 39355
rect 37516 39324 37749 39352
rect 37516 39312 37522 39324
rect 37737 39321 37749 39324
rect 37783 39321 37795 39355
rect 38488 39352 38516 39383
rect 38930 39380 38936 39432
rect 38988 39380 38994 39432
rect 39390 39380 39396 39432
rect 39448 39380 39454 39432
rect 39485 39423 39543 39429
rect 39485 39389 39497 39423
rect 39531 39420 39543 39423
rect 39942 39420 39948 39432
rect 39531 39392 39948 39420
rect 39531 39389 39543 39392
rect 39485 39383 39543 39389
rect 39942 39380 39948 39392
rect 40000 39380 40006 39432
rect 40218 39380 40224 39432
rect 40276 39420 40282 39432
rect 40328 39429 40356 39528
rect 40405 39491 40463 39497
rect 40405 39457 40417 39491
rect 40451 39488 40463 39491
rect 40770 39488 40776 39500
rect 40451 39460 40776 39488
rect 40451 39457 40463 39460
rect 40405 39451 40463 39457
rect 40770 39448 40776 39460
rect 40828 39448 40834 39500
rect 40313 39423 40371 39429
rect 40313 39420 40325 39423
rect 40276 39392 40325 39420
rect 40276 39380 40282 39392
rect 40313 39389 40325 39392
rect 40359 39389 40371 39423
rect 40313 39383 40371 39389
rect 39574 39352 39580 39364
rect 38488 39324 39580 39352
rect 37737 39315 37795 39321
rect 39574 39312 39580 39324
rect 39632 39312 39638 39364
rect 39669 39355 39727 39361
rect 39669 39321 39681 39355
rect 39715 39352 39727 39355
rect 40034 39352 40040 39364
rect 39715 39324 40040 39352
rect 39715 39321 39727 39324
rect 39669 39315 39727 39321
rect 40034 39312 40040 39324
rect 40092 39312 40098 39364
rect 40126 39312 40132 39364
rect 40184 39312 40190 39364
rect 40678 39312 40684 39364
rect 40736 39312 40742 39364
rect 41414 39312 41420 39364
rect 41472 39312 41478 39364
rect 34664 39256 35388 39284
rect 34664 39244 34670 39256
rect 36170 39244 36176 39296
rect 36228 39244 36234 39296
rect 36265 39287 36323 39293
rect 36265 39253 36277 39287
rect 36311 39284 36323 39287
rect 37090 39284 37096 39296
rect 36311 39256 37096 39284
rect 36311 39253 36323 39256
rect 36265 39247 36323 39253
rect 37090 39244 37096 39256
rect 37148 39244 37154 39296
rect 38286 39244 38292 39296
rect 38344 39244 38350 39296
rect 1104 39194 42504 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 42504 39194
rect 1104 39120 42504 39142
rect 15746 39040 15752 39092
rect 15804 39080 15810 39092
rect 16669 39083 16727 39089
rect 16669 39080 16681 39083
rect 15804 39052 16681 39080
rect 15804 39040 15810 39052
rect 16669 39049 16681 39052
rect 16715 39049 16727 39083
rect 16669 39043 16727 39049
rect 17589 39083 17647 39089
rect 17589 39049 17601 39083
rect 17635 39080 17647 39083
rect 18414 39080 18420 39092
rect 17635 39052 18420 39080
rect 17635 39049 17647 39052
rect 17589 39043 17647 39049
rect 18414 39040 18420 39052
rect 18472 39040 18478 39092
rect 19518 39080 19524 39092
rect 19352 39052 19524 39080
rect 18432 39012 18460 39040
rect 19352 39012 19380 39052
rect 19518 39040 19524 39052
rect 19576 39040 19582 39092
rect 19613 39083 19671 39089
rect 19613 39049 19625 39083
rect 19659 39080 19671 39083
rect 20162 39080 20168 39092
rect 19659 39052 20168 39080
rect 19659 39049 19671 39052
rect 19613 39043 19671 39049
rect 20162 39040 20168 39052
rect 20220 39040 20226 39092
rect 20254 39040 20260 39092
rect 20312 39080 20318 39092
rect 20809 39083 20867 39089
rect 20809 39080 20821 39083
rect 20312 39052 20821 39080
rect 20312 39040 20318 39052
rect 20809 39049 20821 39052
rect 20855 39049 20867 39083
rect 20809 39043 20867 39049
rect 23750 39040 23756 39092
rect 23808 39080 23814 39092
rect 24213 39083 24271 39089
rect 24213 39080 24225 39083
rect 23808 39052 24225 39080
rect 23808 39040 23814 39052
rect 24213 39049 24225 39052
rect 24259 39080 24271 39083
rect 24578 39080 24584 39092
rect 24259 39052 24584 39080
rect 24259 39049 24271 39052
rect 24213 39043 24271 39049
rect 24578 39040 24584 39052
rect 24636 39040 24642 39092
rect 25222 39040 25228 39092
rect 25280 39040 25286 39092
rect 31665 39083 31723 39089
rect 31665 39049 31677 39083
rect 31711 39080 31723 39083
rect 32306 39080 32312 39092
rect 31711 39052 32312 39080
rect 31711 39049 31723 39052
rect 31665 39043 31723 39049
rect 32306 39040 32312 39052
rect 32364 39040 32370 39092
rect 32490 39040 32496 39092
rect 32548 39040 32554 39092
rect 32766 39040 32772 39092
rect 32824 39040 32830 39092
rect 35342 39040 35348 39092
rect 35400 39040 35406 39092
rect 35802 39040 35808 39092
rect 35860 39040 35866 39092
rect 35897 39083 35955 39089
rect 35897 39049 35909 39083
rect 35943 39080 35955 39083
rect 35986 39080 35992 39092
rect 35943 39052 35992 39080
rect 35943 39049 35955 39052
rect 35897 39043 35955 39049
rect 35986 39040 35992 39052
rect 36044 39040 36050 39092
rect 36170 39040 36176 39092
rect 36228 39080 36234 39092
rect 37277 39083 37335 39089
rect 36228 39052 37044 39080
rect 36228 39040 36234 39052
rect 24121 39015 24179 39021
rect 24121 39012 24133 39015
rect 18432 38984 19380 39012
rect 3602 38904 3608 38956
rect 3660 38904 3666 38956
rect 14550 38904 14556 38956
rect 14608 38904 14614 38956
rect 15194 38944 15200 38956
rect 14936 38916 15200 38944
rect 12894 38836 12900 38888
rect 12952 38876 12958 38888
rect 13173 38879 13231 38885
rect 13173 38876 13185 38879
rect 12952 38848 13185 38876
rect 12952 38836 12958 38848
rect 13173 38845 13185 38848
rect 13219 38845 13231 38879
rect 13173 38839 13231 38845
rect 13449 38879 13507 38885
rect 13449 38845 13461 38879
rect 13495 38876 13507 38879
rect 14090 38876 14096 38888
rect 13495 38848 14096 38876
rect 13495 38845 13507 38848
rect 13449 38839 13507 38845
rect 14090 38836 14096 38848
rect 14148 38836 14154 38888
rect 14936 38885 14964 38916
rect 15194 38904 15200 38916
rect 15252 38944 15258 38956
rect 15657 38947 15715 38953
rect 15657 38944 15669 38947
rect 15252 38916 15669 38944
rect 15252 38904 15258 38916
rect 15657 38913 15669 38916
rect 15703 38944 15715 38947
rect 16022 38944 16028 38956
rect 15703 38916 16028 38944
rect 15703 38913 15715 38916
rect 15657 38907 15715 38913
rect 16022 38904 16028 38916
rect 16080 38904 16086 38956
rect 17037 38947 17095 38953
rect 17037 38913 17049 38947
rect 17083 38944 17095 38947
rect 17494 38944 17500 38956
rect 17083 38916 17500 38944
rect 17083 38913 17095 38916
rect 17037 38907 17095 38913
rect 17494 38904 17500 38916
rect 17552 38904 17558 38956
rect 17678 38904 17684 38956
rect 17736 38904 17742 38956
rect 19153 38947 19211 38953
rect 19153 38913 19165 38947
rect 19199 38913 19211 38947
rect 19153 38907 19211 38913
rect 14921 38879 14979 38885
rect 14921 38845 14933 38879
rect 14967 38845 14979 38879
rect 14921 38839 14979 38845
rect 17126 38836 17132 38888
rect 17184 38836 17190 38888
rect 17313 38879 17371 38885
rect 17313 38845 17325 38879
rect 17359 38845 17371 38879
rect 19168 38876 19196 38907
rect 19242 38904 19248 38956
rect 19300 38904 19306 38956
rect 19352 38953 19380 38984
rect 23768 38984 24133 39012
rect 23768 38956 23796 38984
rect 24121 38981 24133 38984
rect 24167 38981 24179 39015
rect 24121 38975 24179 38981
rect 27154 38972 27160 39024
rect 27212 39012 27218 39024
rect 30653 39015 30711 39021
rect 27212 38984 27660 39012
rect 27212 38972 27218 38984
rect 19337 38947 19395 38953
rect 19337 38913 19349 38947
rect 19383 38913 19395 38947
rect 19337 38907 19395 38913
rect 19429 38947 19487 38953
rect 19429 38913 19441 38947
rect 19475 38944 19487 38947
rect 19518 38944 19524 38956
rect 19475 38916 19524 38944
rect 19475 38913 19487 38916
rect 19429 38907 19487 38913
rect 19518 38904 19524 38916
rect 19576 38904 19582 38956
rect 20990 38904 20996 38956
rect 21048 38953 21054 38956
rect 21048 38947 21081 38953
rect 21069 38913 21081 38947
rect 21048 38907 21081 38913
rect 21177 38947 21235 38953
rect 21177 38913 21189 38947
rect 21223 38944 21235 38947
rect 22094 38944 22100 38956
rect 21223 38916 22100 38944
rect 21223 38913 21235 38916
rect 21177 38907 21235 38913
rect 21048 38904 21054 38907
rect 22094 38904 22100 38916
rect 22152 38944 22158 38956
rect 22922 38944 22928 38956
rect 22152 38916 22928 38944
rect 22152 38904 22158 38916
rect 22922 38904 22928 38916
rect 22980 38904 22986 38956
rect 23569 38947 23627 38953
rect 23569 38913 23581 38947
rect 23615 38913 23627 38947
rect 23569 38907 23627 38913
rect 19702 38876 19708 38888
rect 19168 38848 19708 38876
rect 17313 38839 17371 38845
rect 14734 38768 14740 38820
rect 14792 38808 14798 38820
rect 17328 38808 17356 38839
rect 19702 38836 19708 38848
rect 19760 38836 19766 38888
rect 23584 38876 23612 38907
rect 23750 38904 23756 38956
rect 23808 38904 23814 38956
rect 23845 38947 23903 38953
rect 23845 38913 23857 38947
rect 23891 38944 23903 38947
rect 23934 38944 23940 38956
rect 23891 38916 23940 38944
rect 23891 38913 23903 38916
rect 23845 38907 23903 38913
rect 23934 38904 23940 38916
rect 23992 38904 23998 38956
rect 24213 38947 24271 38953
rect 24213 38913 24225 38947
rect 24259 38913 24271 38947
rect 24213 38907 24271 38913
rect 24118 38876 24124 38888
rect 23584 38848 24124 38876
rect 24118 38836 24124 38848
rect 24176 38876 24182 38888
rect 24228 38876 24256 38907
rect 25130 38904 25136 38956
rect 25188 38904 25194 38956
rect 25222 38904 25228 38956
rect 25280 38904 25286 38956
rect 25409 38947 25467 38953
rect 25409 38913 25421 38947
rect 25455 38944 25467 38947
rect 25682 38944 25688 38956
rect 25455 38916 25688 38944
rect 25455 38913 25467 38916
rect 25409 38907 25467 38913
rect 25682 38904 25688 38916
rect 25740 38904 25746 38956
rect 27341 38947 27399 38953
rect 27341 38913 27353 38947
rect 27387 38944 27399 38947
rect 27522 38944 27528 38956
rect 27387 38916 27528 38944
rect 27387 38913 27399 38916
rect 27341 38907 27399 38913
rect 27522 38904 27528 38916
rect 27580 38904 27586 38956
rect 27632 38953 27660 38984
rect 30653 38981 30665 39015
rect 30699 39012 30711 39015
rect 30837 39015 30895 39021
rect 30837 39012 30849 39015
rect 30699 38984 30849 39012
rect 30699 38981 30711 38984
rect 30653 38975 30711 38981
rect 30837 38981 30849 38984
rect 30883 39012 30895 39015
rect 35360 39012 35388 39040
rect 37016 39012 37044 39052
rect 37277 39049 37289 39083
rect 37323 39080 37335 39083
rect 37458 39080 37464 39092
rect 37323 39052 37464 39080
rect 37323 39049 37335 39052
rect 37277 39043 37335 39049
rect 37458 39040 37464 39052
rect 37516 39040 37522 39092
rect 37645 39083 37703 39089
rect 37645 39049 37657 39083
rect 37691 39080 37703 39083
rect 37918 39080 37924 39092
rect 37691 39052 37924 39080
rect 37691 39049 37703 39052
rect 37645 39043 37703 39049
rect 37918 39040 37924 39052
rect 37976 39040 37982 39092
rect 38470 39040 38476 39092
rect 38528 39080 38534 39092
rect 38657 39083 38715 39089
rect 38657 39080 38669 39083
rect 38528 39052 38669 39080
rect 38528 39040 38534 39052
rect 38657 39049 38669 39052
rect 38703 39049 38715 39083
rect 38657 39043 38715 39049
rect 39942 39040 39948 39092
rect 40000 39040 40006 39092
rect 40034 39040 40040 39092
rect 40092 39080 40098 39092
rect 40129 39083 40187 39089
rect 40129 39080 40141 39083
rect 40092 39052 40141 39080
rect 40092 39040 40098 39052
rect 40129 39049 40141 39052
rect 40175 39049 40187 39083
rect 40129 39043 40187 39049
rect 40678 39040 40684 39092
rect 40736 39040 40742 39092
rect 41046 39040 41052 39092
rect 41104 39040 41110 39092
rect 37737 39015 37795 39021
rect 37737 39012 37749 39015
rect 30883 38984 32904 39012
rect 35360 38984 36216 39012
rect 37016 38984 37749 39012
rect 30883 38981 30895 38984
rect 30837 38975 30895 38981
rect 27617 38947 27675 38953
rect 27617 38913 27629 38947
rect 27663 38913 27675 38947
rect 27617 38907 27675 38913
rect 27801 38947 27859 38953
rect 27801 38913 27813 38947
rect 27847 38944 27859 38947
rect 28534 38944 28540 38956
rect 27847 38916 28540 38944
rect 27847 38913 27859 38916
rect 27801 38907 27859 38913
rect 24176 38848 24256 38876
rect 24176 38836 24182 38848
rect 25958 38836 25964 38888
rect 26016 38876 26022 38888
rect 27433 38879 27491 38885
rect 27433 38876 27445 38879
rect 26016 38848 27445 38876
rect 26016 38836 26022 38848
rect 27433 38845 27445 38848
rect 27479 38845 27491 38879
rect 27632 38876 27660 38907
rect 28534 38904 28540 38916
rect 28592 38904 28598 38956
rect 30190 38904 30196 38956
rect 30248 38944 30254 38956
rect 30285 38947 30343 38953
rect 30285 38944 30297 38947
rect 30248 38916 30297 38944
rect 30248 38904 30254 38916
rect 30285 38913 30297 38916
rect 30331 38913 30343 38947
rect 30285 38907 30343 38913
rect 30469 38947 30527 38953
rect 30469 38913 30481 38947
rect 30515 38944 30527 38947
rect 30558 38944 30564 38956
rect 30515 38916 30564 38944
rect 30515 38913 30527 38916
rect 30469 38907 30527 38913
rect 30558 38904 30564 38916
rect 30616 38904 30622 38956
rect 30742 38904 30748 38956
rect 30800 38904 30806 38956
rect 31018 38904 31024 38956
rect 31076 38904 31082 38956
rect 31389 38947 31447 38953
rect 31389 38913 31401 38947
rect 31435 38913 31447 38947
rect 31389 38907 31447 38913
rect 31573 38947 31631 38953
rect 31573 38913 31585 38947
rect 31619 38913 31631 38947
rect 31573 38907 31631 38913
rect 31665 38947 31723 38953
rect 31665 38913 31677 38947
rect 31711 38944 31723 38947
rect 31938 38944 31944 38956
rect 31711 38916 31944 38944
rect 31711 38913 31723 38916
rect 31665 38907 31723 38913
rect 27982 38876 27988 38888
rect 27632 38848 27988 38876
rect 27433 38839 27491 38845
rect 27982 38836 27988 38848
rect 28040 38836 28046 38888
rect 17494 38808 17500 38820
rect 14792 38780 17500 38808
rect 14792 38768 14798 38780
rect 17494 38768 17500 38780
rect 17552 38768 17558 38820
rect 23566 38768 23572 38820
rect 23624 38768 23630 38820
rect 27246 38768 27252 38820
rect 27304 38808 27310 38820
rect 27525 38811 27583 38817
rect 27525 38808 27537 38811
rect 27304 38780 27537 38808
rect 27304 38768 27310 38780
rect 27525 38777 27537 38780
rect 27571 38777 27583 38811
rect 27525 38771 27583 38777
rect 30926 38768 30932 38820
rect 30984 38808 30990 38820
rect 31021 38811 31079 38817
rect 31021 38808 31033 38811
rect 30984 38780 31033 38808
rect 30984 38768 30990 38780
rect 31021 38777 31033 38780
rect 31067 38777 31079 38811
rect 31404 38808 31432 38907
rect 31588 38876 31616 38907
rect 31938 38904 31944 38916
rect 31996 38944 32002 38956
rect 32125 38947 32183 38953
rect 32125 38944 32137 38947
rect 31996 38916 32137 38944
rect 31996 38904 32002 38916
rect 32125 38913 32137 38916
rect 32171 38913 32183 38947
rect 32125 38907 32183 38913
rect 32490 38904 32496 38956
rect 32548 38904 32554 38956
rect 32876 38953 32904 38984
rect 32861 38947 32919 38953
rect 32508 38876 32536 38904
rect 32766 38894 32772 38946
rect 32824 38894 32830 38946
rect 32861 38913 32873 38947
rect 32907 38913 32919 38947
rect 32861 38907 32919 38913
rect 33042 38904 33048 38956
rect 33100 38904 33106 38956
rect 34422 38904 34428 38956
rect 34480 38944 34486 38956
rect 35342 38944 35348 38956
rect 34480 38916 35348 38944
rect 34480 38904 34486 38916
rect 35342 38904 35348 38916
rect 35400 38904 35406 38956
rect 35636 38953 35664 38984
rect 35621 38947 35679 38953
rect 35621 38913 35633 38947
rect 35667 38913 35679 38947
rect 35986 38944 35992 38956
rect 35621 38907 35679 38913
rect 35728 38916 35992 38944
rect 31588 38848 32536 38876
rect 32674 38836 32680 38888
rect 32732 38836 32738 38888
rect 35437 38879 35495 38885
rect 35437 38845 35449 38879
rect 35483 38876 35495 38879
rect 35728 38876 35756 38916
rect 35986 38904 35992 38916
rect 36044 38904 36050 38956
rect 36188 38953 36216 38984
rect 37737 38981 37749 38984
rect 37783 38981 37795 39015
rect 37737 38975 37795 38981
rect 36173 38947 36231 38953
rect 36173 38913 36185 38947
rect 36219 38913 36231 38947
rect 36173 38907 36231 38913
rect 39390 38904 39396 38956
rect 39448 38944 39454 38956
rect 40052 38953 40080 39040
rect 39761 38947 39819 38953
rect 39761 38944 39773 38947
rect 39448 38916 39773 38944
rect 39448 38904 39454 38916
rect 39761 38913 39773 38916
rect 39807 38913 39819 38947
rect 39761 38907 39819 38913
rect 40037 38947 40095 38953
rect 40037 38913 40049 38947
rect 40083 38913 40095 38947
rect 40037 38907 40095 38913
rect 35483 38848 35756 38876
rect 35483 38845 35495 38848
rect 35437 38839 35495 38845
rect 35894 38836 35900 38888
rect 35952 38836 35958 38888
rect 37366 38836 37372 38888
rect 37424 38876 37430 38888
rect 37829 38879 37887 38885
rect 37829 38876 37841 38879
rect 37424 38848 37841 38876
rect 37424 38836 37430 38848
rect 37829 38845 37841 38848
rect 37875 38845 37887 38879
rect 37829 38839 37887 38845
rect 39114 38836 39120 38888
rect 39172 38836 39178 38888
rect 39776 38876 39804 38907
rect 40126 38904 40132 38956
rect 40184 38904 40190 38956
rect 40218 38904 40224 38956
rect 40276 38944 40282 38956
rect 40313 38947 40371 38953
rect 40313 38944 40325 38947
rect 40276 38916 40325 38944
rect 40276 38904 40282 38916
rect 40313 38913 40325 38916
rect 40359 38913 40371 38947
rect 41782 38944 41788 38956
rect 40313 38907 40371 38913
rect 40420 38916 41788 38944
rect 40420 38876 40448 38916
rect 41782 38904 41788 38916
rect 41840 38944 41846 38956
rect 42061 38947 42119 38953
rect 42061 38944 42073 38947
rect 41840 38916 42073 38944
rect 41840 38904 41846 38916
rect 42061 38913 42073 38916
rect 42107 38913 42119 38947
rect 42061 38907 42119 38913
rect 39776 38848 40448 38876
rect 41138 38836 41144 38888
rect 41196 38836 41202 38888
rect 41233 38879 41291 38885
rect 41233 38845 41245 38879
rect 41279 38845 41291 38879
rect 41233 38839 41291 38845
rect 31404 38780 31616 38808
rect 31021 38771 31079 38777
rect 3234 38700 3240 38752
rect 3292 38740 3298 38752
rect 3513 38743 3571 38749
rect 3513 38740 3525 38743
rect 3292 38712 3525 38740
rect 3292 38700 3298 38712
rect 3513 38709 3525 38712
rect 3559 38709 3571 38743
rect 3513 38703 3571 38709
rect 15010 38700 15016 38752
rect 15068 38700 15074 38752
rect 27157 38743 27215 38749
rect 27157 38709 27169 38743
rect 27203 38740 27215 38743
rect 31386 38740 31392 38752
rect 27203 38712 31392 38740
rect 27203 38709 27215 38712
rect 27157 38703 27215 38709
rect 31386 38700 31392 38712
rect 31444 38700 31450 38752
rect 31588 38740 31616 38780
rect 35526 38768 35532 38820
rect 35584 38768 35590 38820
rect 38841 38811 38899 38817
rect 38841 38777 38853 38811
rect 38887 38808 38899 38811
rect 38930 38808 38936 38820
rect 38887 38780 38936 38808
rect 38887 38777 38899 38780
rect 38841 38771 38899 38777
rect 32674 38740 32680 38752
rect 31588 38712 32680 38740
rect 32674 38700 32680 38712
rect 32732 38740 32738 38752
rect 32950 38740 32956 38752
rect 32732 38712 32956 38740
rect 32732 38700 32738 38712
rect 32950 38700 32956 38712
rect 33008 38700 33014 38752
rect 35342 38700 35348 38752
rect 35400 38740 35406 38752
rect 35894 38740 35900 38752
rect 35400 38712 35900 38740
rect 35400 38700 35406 38712
rect 35894 38700 35900 38712
rect 35952 38700 35958 38752
rect 36078 38700 36084 38752
rect 36136 38740 36142 38752
rect 37366 38740 37372 38752
rect 36136 38712 37372 38740
rect 36136 38700 36142 38712
rect 37366 38700 37372 38712
rect 37424 38700 37430 38752
rect 38856 38740 38884 38771
rect 38930 38768 38936 38780
rect 38988 38768 38994 38820
rect 39666 38768 39672 38820
rect 39724 38808 39730 38820
rect 39761 38811 39819 38817
rect 39761 38808 39773 38811
rect 39724 38780 39773 38808
rect 39724 38768 39730 38780
rect 39761 38777 39773 38780
rect 39807 38777 39819 38811
rect 39761 38771 39819 38777
rect 41046 38768 41052 38820
rect 41104 38808 41110 38820
rect 41248 38808 41276 38839
rect 41104 38780 41276 38808
rect 41104 38768 41110 38780
rect 40494 38740 40500 38752
rect 38856 38712 40500 38740
rect 40494 38700 40500 38712
rect 40552 38700 40558 38752
rect 40862 38700 40868 38752
rect 40920 38740 40926 38752
rect 41509 38743 41567 38749
rect 41509 38740 41521 38743
rect 40920 38712 41521 38740
rect 40920 38700 40926 38712
rect 41509 38709 41521 38712
rect 41555 38709 41567 38743
rect 41509 38703 41567 38709
rect 1104 38650 42504 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 42504 38650
rect 1104 38576 42504 38598
rect 7282 38536 7288 38548
rect 6288 38508 7288 38536
rect 1394 38360 1400 38412
rect 1452 38400 1458 38412
rect 1673 38403 1731 38409
rect 1673 38400 1685 38403
rect 1452 38372 1685 38400
rect 1452 38360 1458 38372
rect 1673 38369 1685 38372
rect 1719 38400 1731 38403
rect 3786 38400 3792 38412
rect 1719 38372 3792 38400
rect 1719 38369 1731 38372
rect 1673 38363 1731 38369
rect 3786 38360 3792 38372
rect 3844 38360 3850 38412
rect 5258 38400 5264 38412
rect 4724 38372 5264 38400
rect 3418 38292 3424 38344
rect 3476 38332 3482 38344
rect 4724 38341 4752 38372
rect 5258 38360 5264 38372
rect 5316 38360 5322 38412
rect 4341 38335 4399 38341
rect 4341 38332 4353 38335
rect 3476 38304 4353 38332
rect 3476 38292 3482 38304
rect 4341 38301 4353 38304
rect 4387 38332 4399 38335
rect 4709 38335 4767 38341
rect 4709 38332 4721 38335
rect 4387 38304 4721 38332
rect 4387 38301 4399 38304
rect 4341 38295 4399 38301
rect 4709 38301 4721 38304
rect 4755 38301 4767 38335
rect 4709 38295 4767 38301
rect 4985 38335 5043 38341
rect 4985 38301 4997 38335
rect 5031 38332 5043 38335
rect 5031 38304 5488 38332
rect 5031 38301 5043 38304
rect 4985 38295 5043 38301
rect 5460 38276 5488 38304
rect 6086 38292 6092 38344
rect 6144 38292 6150 38344
rect 6288 38341 6316 38508
rect 7282 38496 7288 38508
rect 7340 38496 7346 38548
rect 14090 38496 14096 38548
rect 14148 38496 14154 38548
rect 19518 38496 19524 38548
rect 19576 38496 19582 38548
rect 19702 38496 19708 38548
rect 19760 38496 19766 38548
rect 20990 38496 20996 38548
rect 21048 38536 21054 38548
rect 21177 38539 21235 38545
rect 21177 38536 21189 38539
rect 21048 38508 21189 38536
rect 21048 38496 21054 38508
rect 21177 38505 21189 38508
rect 21223 38505 21235 38539
rect 21177 38499 21235 38505
rect 21266 38496 21272 38548
rect 21324 38536 21330 38548
rect 21545 38539 21603 38545
rect 21545 38536 21557 38539
rect 21324 38508 21557 38536
rect 21324 38496 21330 38508
rect 21545 38505 21557 38508
rect 21591 38536 21603 38539
rect 22005 38539 22063 38545
rect 21591 38508 21956 38536
rect 21591 38505 21603 38508
rect 21545 38499 21603 38505
rect 13541 38471 13599 38477
rect 13541 38437 13553 38471
rect 13587 38468 13599 38471
rect 13814 38468 13820 38480
rect 13587 38440 13820 38468
rect 13587 38437 13599 38440
rect 13541 38431 13599 38437
rect 13814 38428 13820 38440
rect 13872 38468 13878 38480
rect 19610 38468 19616 38480
rect 13872 38440 19616 38468
rect 13872 38428 13878 38440
rect 19610 38428 19616 38440
rect 19668 38428 19674 38480
rect 6549 38403 6607 38409
rect 6549 38369 6561 38403
rect 6595 38400 6607 38403
rect 7098 38400 7104 38412
rect 6595 38372 7104 38400
rect 6595 38369 6607 38372
rect 6549 38363 6607 38369
rect 7098 38360 7104 38372
rect 7156 38360 7162 38412
rect 8294 38360 8300 38412
rect 8352 38400 8358 38412
rect 8573 38403 8631 38409
rect 8573 38400 8585 38403
rect 8352 38372 8585 38400
rect 8352 38360 8358 38372
rect 8573 38369 8585 38372
rect 8619 38400 8631 38403
rect 9493 38403 9551 38409
rect 9493 38400 9505 38403
rect 8619 38372 9505 38400
rect 8619 38369 8631 38372
rect 8573 38363 8631 38369
rect 9493 38369 9505 38372
rect 9539 38369 9551 38403
rect 9493 38363 9551 38369
rect 14734 38360 14740 38412
rect 14792 38360 14798 38412
rect 19518 38360 19524 38412
rect 19576 38400 19582 38412
rect 21928 38400 21956 38508
rect 22005 38505 22017 38539
rect 22051 38536 22063 38539
rect 22094 38536 22100 38548
rect 22051 38508 22100 38536
rect 22051 38505 22063 38508
rect 22005 38499 22063 38505
rect 22094 38496 22100 38508
rect 22152 38496 22158 38548
rect 23569 38539 23627 38545
rect 23569 38505 23581 38539
rect 23615 38536 23627 38539
rect 23750 38536 23756 38548
rect 23615 38508 23756 38536
rect 23615 38505 23627 38508
rect 23569 38499 23627 38505
rect 23750 38496 23756 38508
rect 23808 38496 23814 38548
rect 23934 38496 23940 38548
rect 23992 38536 23998 38548
rect 24121 38539 24179 38545
rect 24121 38536 24133 38539
rect 23992 38508 24133 38536
rect 23992 38496 23998 38508
rect 24121 38505 24133 38508
rect 24167 38505 24179 38539
rect 24121 38499 24179 38505
rect 25222 38496 25228 38548
rect 25280 38536 25286 38548
rect 25590 38536 25596 38548
rect 25280 38508 25596 38536
rect 25280 38496 25286 38508
rect 25590 38496 25596 38508
rect 25648 38496 25654 38548
rect 25682 38496 25688 38548
rect 25740 38536 25746 38548
rect 26145 38539 26203 38545
rect 26145 38536 26157 38539
rect 25740 38508 26157 38536
rect 25740 38496 25746 38508
rect 26145 38505 26157 38508
rect 26191 38505 26203 38539
rect 26145 38499 26203 38505
rect 28534 38496 28540 38548
rect 28592 38496 28598 38548
rect 29178 38496 29184 38548
rect 29236 38496 29242 38548
rect 31018 38496 31024 38548
rect 31076 38536 31082 38548
rect 31297 38539 31355 38545
rect 31297 38536 31309 38539
rect 31076 38508 31309 38536
rect 31076 38496 31082 38508
rect 31297 38505 31309 38508
rect 31343 38536 31355 38539
rect 31343 38508 31754 38536
rect 31343 38505 31355 38508
rect 31297 38499 31355 38505
rect 22278 38428 22284 38480
rect 22336 38468 22342 38480
rect 22465 38471 22523 38477
rect 22465 38468 22477 38471
rect 22336 38440 22477 38468
rect 22336 38428 22342 38440
rect 22465 38437 22477 38440
rect 22511 38437 22523 38471
rect 22465 38431 22523 38437
rect 25424 38440 25912 38468
rect 19576 38372 19932 38400
rect 19576 38360 19582 38372
rect 19904 38344 19932 38372
rect 21192 38372 21864 38400
rect 21928 38372 22232 38400
rect 6273 38335 6331 38341
rect 6273 38301 6285 38335
rect 6319 38301 6331 38335
rect 6273 38295 6331 38301
rect 6822 38292 6828 38344
rect 6880 38292 6886 38344
rect 11606 38292 11612 38344
rect 11664 38332 11670 38344
rect 11793 38335 11851 38341
rect 11793 38332 11805 38335
rect 11664 38304 11805 38332
rect 11664 38292 11670 38304
rect 11793 38301 11805 38304
rect 11839 38301 11851 38335
rect 11793 38295 11851 38301
rect 14461 38335 14519 38341
rect 14461 38301 14473 38335
rect 14507 38332 14519 38335
rect 15010 38332 15016 38344
rect 14507 38304 15016 38332
rect 14507 38301 14519 38304
rect 14461 38295 14519 38301
rect 15010 38292 15016 38304
rect 15068 38292 15074 38344
rect 19242 38292 19248 38344
rect 19300 38292 19306 38344
rect 19337 38335 19395 38341
rect 19337 38301 19349 38335
rect 19383 38332 19395 38335
rect 19426 38332 19432 38344
rect 19383 38304 19432 38332
rect 19383 38301 19395 38304
rect 19337 38295 19395 38301
rect 19426 38292 19432 38304
rect 19484 38332 19490 38344
rect 19797 38335 19855 38341
rect 19797 38332 19809 38335
rect 19484 38304 19809 38332
rect 19484 38292 19490 38304
rect 19797 38301 19809 38304
rect 19843 38301 19855 38335
rect 19797 38295 19855 38301
rect 19886 38292 19892 38344
rect 19944 38292 19950 38344
rect 20990 38292 20996 38344
rect 21048 38332 21054 38344
rect 21192 38341 21220 38372
rect 21177 38335 21235 38341
rect 21177 38332 21189 38335
rect 21048 38304 21189 38332
rect 21048 38292 21054 38304
rect 21177 38301 21189 38304
rect 21223 38301 21235 38335
rect 21177 38295 21235 38301
rect 21266 38292 21272 38344
rect 21324 38292 21330 38344
rect 21453 38335 21511 38341
rect 21453 38301 21465 38335
rect 21499 38332 21511 38335
rect 21634 38332 21640 38344
rect 21499 38304 21640 38332
rect 21499 38301 21511 38304
rect 21453 38295 21511 38301
rect 21634 38292 21640 38304
rect 21692 38292 21698 38344
rect 21836 38332 21864 38372
rect 22204 38341 22232 38372
rect 22388 38372 23796 38400
rect 22388 38344 22416 38372
rect 22005 38335 22063 38341
rect 22005 38334 22017 38335
rect 21928 38332 22017 38334
rect 21836 38306 22017 38332
rect 21836 38304 21956 38306
rect 22005 38301 22017 38306
rect 22051 38301 22063 38335
rect 22005 38295 22063 38301
rect 22189 38335 22247 38341
rect 22189 38301 22201 38335
rect 22235 38301 22247 38335
rect 22189 38295 22247 38301
rect 22278 38292 22284 38344
rect 22336 38292 22342 38344
rect 22370 38292 22376 38344
rect 22428 38292 22434 38344
rect 23768 38341 23796 38372
rect 25424 38344 25452 38440
rect 25590 38360 25596 38412
rect 25648 38400 25654 38412
rect 25884 38400 25912 38440
rect 25958 38428 25964 38480
rect 26016 38428 26022 38480
rect 28902 38428 28908 38480
rect 28960 38468 28966 38480
rect 28960 38440 29040 38468
rect 28960 38428 28966 38440
rect 29012 38400 29040 38440
rect 29549 38403 29607 38409
rect 29549 38400 29561 38403
rect 25648 38372 25820 38400
rect 25884 38372 26280 38400
rect 29012 38372 29561 38400
rect 25648 38360 25654 38372
rect 22557 38335 22615 38341
rect 22557 38301 22569 38335
rect 22603 38301 22615 38335
rect 22557 38295 22615 38301
rect 23753 38335 23811 38341
rect 23753 38301 23765 38335
rect 23799 38332 23811 38335
rect 24029 38335 24087 38341
rect 24029 38332 24041 38335
rect 23799 38304 24041 38332
rect 23799 38301 23811 38304
rect 23753 38295 23811 38301
rect 24029 38301 24041 38304
rect 24075 38301 24087 38335
rect 24029 38295 24087 38301
rect 24213 38335 24271 38341
rect 24213 38301 24225 38335
rect 24259 38301 24271 38335
rect 24213 38295 24271 38301
rect 1946 38224 1952 38276
rect 2004 38224 2010 38276
rect 2958 38224 2964 38276
rect 3016 38224 3022 38276
rect 4525 38267 4583 38273
rect 4525 38264 4537 38267
rect 3344 38236 4537 38264
rect 2590 38156 2596 38208
rect 2648 38196 2654 38208
rect 3344 38196 3372 38236
rect 4525 38233 4537 38236
rect 4571 38233 4583 38267
rect 5077 38267 5135 38273
rect 5077 38264 5089 38267
rect 4525 38227 4583 38233
rect 4724 38236 5089 38264
rect 4724 38208 4752 38236
rect 5077 38233 5089 38236
rect 5123 38233 5135 38267
rect 5077 38227 5135 38233
rect 5261 38267 5319 38273
rect 5261 38233 5273 38267
rect 5307 38233 5319 38267
rect 5261 38227 5319 38233
rect 2648 38168 3372 38196
rect 2648 38156 2654 38168
rect 3418 38156 3424 38208
rect 3476 38156 3482 38208
rect 3510 38156 3516 38208
rect 3568 38196 3574 38208
rect 3789 38199 3847 38205
rect 3789 38196 3801 38199
rect 3568 38168 3801 38196
rect 3568 38156 3574 38168
rect 3789 38165 3801 38168
rect 3835 38165 3847 38199
rect 3789 38159 3847 38165
rect 4706 38156 4712 38208
rect 4764 38156 4770 38208
rect 4798 38156 4804 38208
rect 4856 38196 4862 38208
rect 4893 38199 4951 38205
rect 4893 38196 4905 38199
rect 4856 38168 4905 38196
rect 4856 38156 4862 38168
rect 4893 38165 4905 38168
rect 4939 38196 4951 38199
rect 5276 38196 5304 38227
rect 5442 38224 5448 38276
rect 5500 38224 5506 38276
rect 6454 38273 6460 38276
rect 6181 38267 6239 38273
rect 6181 38233 6193 38267
rect 6227 38233 6239 38267
rect 6181 38227 6239 38233
rect 6411 38267 6460 38273
rect 6411 38233 6423 38267
rect 6457 38233 6460 38267
rect 6411 38227 6460 38233
rect 4939 38168 5304 38196
rect 4939 38165 4951 38168
rect 4893 38159 4951 38165
rect 5902 38156 5908 38208
rect 5960 38156 5966 38208
rect 6196 38196 6224 38227
rect 6454 38224 6460 38227
rect 6512 38224 6518 38276
rect 7006 38224 7012 38276
rect 7064 38264 7070 38276
rect 7101 38267 7159 38273
rect 7101 38264 7113 38267
rect 7064 38236 7113 38264
rect 7064 38224 7070 38236
rect 7101 38233 7113 38236
rect 7147 38233 7159 38267
rect 9674 38264 9680 38276
rect 8326 38236 9680 38264
rect 7101 38227 7159 38233
rect 9674 38224 9680 38236
rect 9732 38224 9738 38276
rect 12066 38224 12072 38276
rect 12124 38224 12130 38276
rect 14366 38264 14372 38276
rect 13294 38236 14372 38264
rect 14366 38224 14372 38236
rect 14424 38224 14430 38276
rect 19518 38224 19524 38276
rect 19576 38224 19582 38276
rect 19613 38267 19671 38273
rect 19613 38233 19625 38267
rect 19659 38233 19671 38267
rect 19613 38227 19671 38233
rect 7926 38196 7932 38208
rect 6196 38168 7932 38196
rect 7926 38156 7932 38168
rect 7984 38156 7990 38208
rect 8938 38156 8944 38208
rect 8996 38156 9002 38208
rect 14553 38199 14611 38205
rect 14553 38165 14565 38199
rect 14599 38196 14611 38199
rect 14642 38196 14648 38208
rect 14599 38168 14648 38196
rect 14599 38165 14611 38168
rect 14553 38159 14611 38165
rect 14642 38156 14648 38168
rect 14700 38156 14706 38208
rect 19242 38156 19248 38208
rect 19300 38196 19306 38208
rect 19628 38196 19656 38227
rect 21358 38224 21364 38276
rect 21416 38264 21422 38276
rect 21729 38267 21787 38273
rect 21729 38264 21741 38267
rect 21416 38236 21741 38264
rect 21416 38224 21422 38236
rect 21729 38233 21741 38236
rect 21775 38233 21787 38267
rect 21913 38267 21971 38273
rect 21913 38264 21925 38267
rect 21729 38227 21787 38233
rect 21836 38236 21925 38264
rect 21836 38208 21864 38236
rect 21913 38233 21925 38236
rect 21959 38233 21971 38267
rect 21913 38227 21971 38233
rect 22572 38208 22600 38295
rect 23934 38224 23940 38276
rect 23992 38264 23998 38276
rect 24228 38264 24256 38295
rect 25406 38292 25412 38344
rect 25464 38292 25470 38344
rect 25682 38292 25688 38344
rect 25740 38292 25746 38344
rect 25792 38341 25820 38372
rect 25777 38335 25835 38341
rect 25777 38301 25789 38335
rect 25823 38301 25835 38335
rect 26053 38335 26111 38341
rect 26053 38332 26065 38335
rect 25777 38295 25835 38301
rect 25884 38304 26065 38332
rect 23992 38236 24256 38264
rect 25593 38267 25651 38273
rect 23992 38224 23998 38236
rect 25593 38233 25605 38267
rect 25639 38264 25651 38267
rect 25884 38264 25912 38304
rect 26053 38301 26065 38304
rect 26099 38332 26111 38335
rect 26142 38332 26148 38344
rect 26099 38304 26148 38332
rect 26099 38301 26111 38304
rect 26053 38295 26111 38301
rect 26142 38292 26148 38304
rect 26200 38292 26206 38344
rect 26252 38341 26280 38372
rect 29549 38369 29561 38372
rect 29595 38369 29607 38403
rect 31726 38400 31754 38508
rect 36906 38496 36912 38548
rect 36964 38536 36970 38548
rect 37550 38536 37556 38548
rect 36964 38508 37556 38536
rect 36964 38496 36970 38508
rect 37550 38496 37556 38508
rect 37608 38496 37614 38548
rect 40310 38496 40316 38548
rect 40368 38536 40374 38548
rect 40497 38539 40555 38545
rect 40497 38536 40509 38539
rect 40368 38508 40509 38536
rect 40368 38496 40374 38508
rect 40497 38505 40509 38508
rect 40543 38505 40555 38539
rect 40497 38499 40555 38505
rect 38565 38471 38623 38477
rect 38565 38437 38577 38471
rect 38611 38437 38623 38471
rect 38565 38431 38623 38437
rect 32033 38403 32091 38409
rect 32033 38400 32045 38403
rect 31726 38372 32045 38400
rect 29549 38363 29607 38369
rect 32033 38369 32045 38372
rect 32079 38400 32091 38403
rect 32766 38400 32772 38412
rect 32079 38372 32772 38400
rect 32079 38369 32091 38372
rect 32033 38363 32091 38369
rect 32766 38360 32772 38372
rect 32824 38360 32830 38412
rect 34790 38360 34796 38412
rect 34848 38400 34854 38412
rect 35713 38403 35771 38409
rect 35713 38400 35725 38403
rect 34848 38372 35725 38400
rect 34848 38360 34854 38372
rect 35713 38369 35725 38372
rect 35759 38369 35771 38403
rect 35713 38363 35771 38369
rect 37366 38360 37372 38412
rect 37424 38360 37430 38412
rect 38580 38400 38608 38431
rect 38212 38372 38608 38400
rect 26237 38335 26295 38341
rect 26237 38301 26249 38335
rect 26283 38332 26295 38335
rect 28166 38332 28172 38344
rect 26283 38304 28172 38332
rect 26283 38301 26295 38304
rect 26237 38295 26295 38301
rect 28166 38292 28172 38304
rect 28224 38292 28230 38344
rect 28537 38335 28595 38341
rect 28537 38301 28549 38335
rect 28583 38332 28595 38335
rect 28813 38335 28871 38341
rect 28583 38304 28764 38332
rect 28583 38301 28595 38304
rect 28537 38295 28595 38301
rect 25639 38236 25912 38264
rect 25971 38267 26029 38273
rect 25639 38233 25651 38236
rect 25593 38227 25651 38233
rect 25971 38233 25983 38267
rect 26017 38264 26029 38267
rect 26017 38236 26096 38264
rect 26017 38233 26029 38236
rect 25971 38227 26029 38233
rect 26068 38208 26096 38236
rect 28626 38224 28632 38276
rect 28684 38224 28690 38276
rect 28736 38264 28764 38304
rect 28813 38301 28825 38335
rect 28859 38332 28871 38335
rect 28902 38332 28908 38344
rect 28859 38304 28908 38332
rect 28859 38301 28871 38304
rect 28813 38295 28871 38301
rect 28902 38292 28908 38304
rect 28960 38292 28966 38344
rect 32398 38292 32404 38344
rect 32456 38292 32462 38344
rect 35253 38335 35311 38341
rect 35253 38332 35265 38335
rect 34164 38304 35265 38332
rect 29178 38264 29184 38276
rect 28736 38236 29184 38264
rect 29178 38224 29184 38236
rect 29236 38224 29242 38276
rect 29546 38224 29552 38276
rect 29604 38264 29610 38276
rect 29825 38267 29883 38273
rect 29825 38264 29837 38267
rect 29604 38236 29837 38264
rect 29604 38224 29610 38236
rect 29825 38233 29837 38236
rect 29871 38233 29883 38267
rect 32306 38264 32312 38276
rect 31050 38236 32312 38264
rect 29825 38227 29883 38233
rect 32306 38224 32312 38236
rect 32364 38224 32370 38276
rect 32674 38224 32680 38276
rect 32732 38224 32738 38276
rect 33226 38224 33232 38276
rect 33284 38224 33290 38276
rect 19300 38168 19656 38196
rect 19300 38156 19306 38168
rect 21818 38156 21824 38208
rect 21876 38156 21882 38208
rect 22554 38156 22560 38208
rect 22612 38156 22618 38208
rect 25130 38156 25136 38208
rect 25188 38196 25194 38208
rect 26050 38196 26056 38208
rect 25188 38168 26056 38196
rect 25188 38156 25194 38168
rect 26050 38156 26056 38168
rect 26108 38156 26114 38208
rect 28644 38196 28672 38224
rect 28997 38199 29055 38205
rect 28997 38196 29009 38199
rect 28644 38168 29009 38196
rect 28997 38165 29009 38168
rect 29043 38165 29055 38199
rect 28997 38159 29055 38165
rect 31386 38156 31392 38208
rect 31444 38156 31450 38208
rect 33686 38156 33692 38208
rect 33744 38196 33750 38208
rect 34164 38205 34192 38304
rect 35253 38301 35265 38304
rect 35299 38301 35311 38335
rect 35253 38295 35311 38301
rect 35802 38292 35808 38344
rect 35860 38292 35866 38344
rect 37918 38292 37924 38344
rect 37976 38292 37982 38344
rect 38212 38341 38240 38372
rect 41046 38360 41052 38412
rect 41104 38360 41110 38412
rect 38197 38335 38255 38341
rect 38197 38301 38209 38335
rect 38243 38301 38255 38335
rect 38197 38295 38255 38301
rect 38286 38292 38292 38344
rect 38344 38332 38350 38344
rect 38565 38335 38623 38341
rect 38565 38332 38577 38335
rect 38344 38304 38577 38332
rect 38344 38292 38350 38304
rect 38565 38301 38577 38304
rect 38611 38301 38623 38335
rect 38565 38295 38623 38301
rect 38749 38335 38807 38341
rect 38749 38301 38761 38335
rect 38795 38332 38807 38335
rect 39114 38332 39120 38344
rect 38795 38304 39120 38332
rect 38795 38301 38807 38304
rect 38749 38295 38807 38301
rect 39114 38292 39120 38304
rect 39172 38332 39178 38344
rect 39390 38332 39396 38344
rect 39172 38304 39396 38332
rect 39172 38292 39178 38304
rect 39390 38292 39396 38304
rect 39448 38292 39454 38344
rect 40862 38292 40868 38344
rect 40920 38292 40926 38344
rect 41874 38292 41880 38344
rect 41932 38292 41938 38344
rect 40586 38224 40592 38276
rect 40644 38264 40650 38276
rect 41325 38267 41383 38273
rect 41325 38264 41337 38267
rect 40644 38236 41337 38264
rect 40644 38224 40650 38236
rect 41325 38233 41337 38236
rect 41371 38233 41383 38267
rect 41325 38227 41383 38233
rect 34149 38199 34207 38205
rect 34149 38196 34161 38199
rect 33744 38168 34161 38196
rect 33744 38156 33750 38168
rect 34149 38165 34161 38168
rect 34195 38165 34207 38199
rect 34149 38159 34207 38165
rect 34698 38156 34704 38208
rect 34756 38156 34762 38208
rect 35434 38156 35440 38208
rect 35492 38156 35498 38208
rect 40954 38156 40960 38208
rect 41012 38156 41018 38208
rect 1104 38106 42504 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 42504 38106
rect 1104 38032 42504 38054
rect 1946 37952 1952 38004
rect 2004 37992 2010 38004
rect 2317 37995 2375 38001
rect 2317 37992 2329 37995
rect 2004 37964 2329 37992
rect 2004 37952 2010 37964
rect 2317 37961 2329 37964
rect 2363 37961 2375 37995
rect 5810 37992 5816 38004
rect 2317 37955 2375 37961
rect 2838 37964 5816 37992
rect 2838 37933 2866 37964
rect 5810 37952 5816 37964
rect 5868 37992 5874 38004
rect 5868 37964 6040 37992
rect 5868 37952 5874 37964
rect 2823 37927 2881 37933
rect 2823 37893 2835 37927
rect 2869 37893 2881 37927
rect 6012 37924 6040 37964
rect 6086 37952 6092 38004
rect 6144 37992 6150 38004
rect 6365 37995 6423 38001
rect 6365 37992 6377 37995
rect 6144 37964 6377 37992
rect 6144 37952 6150 37964
rect 6365 37961 6377 37964
rect 6411 37961 6423 37995
rect 6365 37955 6423 37961
rect 7006 37952 7012 38004
rect 7064 37952 7070 38004
rect 7466 37992 7472 38004
rect 7116 37964 7472 37992
rect 6454 37924 6460 37936
rect 6012 37896 6460 37924
rect 2823 37887 2881 37893
rect 6454 37884 6460 37896
rect 6512 37924 6518 37936
rect 7116 37924 7144 37964
rect 7466 37952 7472 37964
rect 7524 37952 7530 38004
rect 15102 37952 15108 38004
rect 15160 37992 15166 38004
rect 15565 37995 15623 38001
rect 15565 37992 15577 37995
rect 15160 37964 15577 37992
rect 15160 37952 15166 37964
rect 15565 37961 15577 37964
rect 15611 37992 15623 37995
rect 18969 37995 19027 38001
rect 15611 37964 16988 37992
rect 15611 37961 15623 37964
rect 15565 37955 15623 37961
rect 7745 37927 7803 37933
rect 7745 37924 7757 37927
rect 6512 37896 7144 37924
rect 7208 37896 7757 37924
rect 6512 37884 6518 37896
rect 1765 37859 1823 37865
rect 1765 37825 1777 37859
rect 1811 37856 1823 37859
rect 1854 37856 1860 37868
rect 1811 37828 1860 37856
rect 1811 37825 1823 37828
rect 1765 37819 1823 37825
rect 1854 37816 1860 37828
rect 1912 37816 1918 37868
rect 2038 37816 2044 37868
rect 2096 37816 2102 37868
rect 2501 37859 2559 37865
rect 2501 37825 2513 37859
rect 2547 37825 2559 37859
rect 2501 37819 2559 37825
rect 1673 37791 1731 37797
rect 1673 37757 1685 37791
rect 1719 37788 1731 37791
rect 2516 37788 2544 37819
rect 2590 37816 2596 37868
rect 2648 37816 2654 37868
rect 2685 37859 2743 37865
rect 2685 37825 2697 37859
rect 2731 37825 2743 37859
rect 2685 37819 2743 37825
rect 2961 37859 3019 37865
rect 2961 37825 2973 37859
rect 3007 37856 3019 37859
rect 3510 37856 3516 37868
rect 3007 37828 3516 37856
rect 3007 37825 3019 37828
rect 2961 37819 3019 37825
rect 1719 37760 2544 37788
rect 2700 37788 2728 37819
rect 3510 37816 3516 37828
rect 3568 37816 3574 37868
rect 5534 37856 5540 37868
rect 5198 37828 5540 37856
rect 5534 37816 5540 37828
rect 5592 37816 5598 37868
rect 6733 37859 6791 37865
rect 6733 37825 6745 37859
rect 6779 37856 6791 37859
rect 6914 37856 6920 37868
rect 6779 37828 6920 37856
rect 6779 37825 6791 37828
rect 6733 37819 6791 37825
rect 6914 37816 6920 37828
rect 6972 37856 6978 37868
rect 7208 37865 7236 37896
rect 7745 37893 7757 37896
rect 7791 37893 7803 37927
rect 8938 37924 8944 37936
rect 7745 37887 7803 37893
rect 7852 37896 8944 37924
rect 7193 37859 7251 37865
rect 6972 37828 7144 37856
rect 6972 37816 6978 37828
rect 3326 37788 3332 37800
rect 2700 37760 3332 37788
rect 1719 37757 1731 37760
rect 1673 37751 1731 37757
rect 3326 37748 3332 37760
rect 3384 37748 3390 37800
rect 3694 37748 3700 37800
rect 3752 37748 3758 37800
rect 3786 37748 3792 37800
rect 3844 37748 3850 37800
rect 4065 37791 4123 37797
rect 4065 37757 4077 37791
rect 4111 37788 4123 37791
rect 4614 37788 4620 37800
rect 4111 37760 4620 37788
rect 4111 37757 4123 37760
rect 4065 37751 4123 37757
rect 4614 37748 4620 37760
rect 4672 37748 4678 37800
rect 6549 37791 6607 37797
rect 6549 37757 6561 37791
rect 6595 37757 6607 37791
rect 6549 37751 6607 37757
rect 5166 37680 5172 37732
rect 5224 37720 5230 37732
rect 5442 37720 5448 37732
rect 5224 37692 5448 37720
rect 5224 37680 5230 37692
rect 5442 37680 5448 37692
rect 5500 37720 5506 37732
rect 6564 37720 6592 37751
rect 6638 37748 6644 37800
rect 6696 37748 6702 37800
rect 6825 37791 6883 37797
rect 6825 37757 6837 37791
rect 6871 37788 6883 37791
rect 7006 37788 7012 37800
rect 6871 37760 7012 37788
rect 6871 37757 6883 37760
rect 6825 37751 6883 37757
rect 7006 37748 7012 37760
rect 7064 37748 7070 37800
rect 7116 37788 7144 37828
rect 7193 37825 7205 37859
rect 7239 37825 7251 37859
rect 7193 37819 7251 37825
rect 7282 37816 7288 37868
rect 7340 37816 7346 37868
rect 7374 37816 7380 37868
rect 7432 37816 7438 37868
rect 7466 37816 7472 37868
rect 7524 37865 7530 37868
rect 7524 37859 7553 37865
rect 7541 37825 7553 37859
rect 7524 37819 7553 37825
rect 7653 37859 7711 37865
rect 7653 37825 7665 37859
rect 7699 37856 7711 37859
rect 7852 37856 7880 37896
rect 8938 37884 8944 37896
rect 8996 37884 9002 37936
rect 7699 37828 7880 37856
rect 7929 37859 7987 37865
rect 7699 37825 7711 37828
rect 7653 37819 7711 37825
rect 7929 37825 7941 37859
rect 7975 37856 7987 37859
rect 8018 37856 8024 37868
rect 7975 37828 8024 37856
rect 7975 37825 7987 37828
rect 7929 37819 7987 37825
rect 7524 37816 7530 37819
rect 8018 37816 8024 37828
rect 8076 37816 8082 37868
rect 8113 37859 8171 37865
rect 8113 37825 8125 37859
rect 8159 37825 8171 37859
rect 8113 37819 8171 37825
rect 8205 37859 8263 37865
rect 8205 37825 8217 37859
rect 8251 37825 8263 37859
rect 8205 37819 8263 37825
rect 12805 37859 12863 37865
rect 12805 37825 12817 37859
rect 12851 37825 12863 37859
rect 12805 37819 12863 37825
rect 8128 37788 8156 37819
rect 7116 37760 8156 37788
rect 8018 37720 8024 37732
rect 5500 37692 5672 37720
rect 6564 37692 8024 37720
rect 5500 37680 5506 37692
rect 2225 37655 2283 37661
rect 2225 37621 2237 37655
rect 2271 37652 2283 37655
rect 2866 37652 2872 37664
rect 2271 37624 2872 37652
rect 2271 37621 2283 37624
rect 2225 37615 2283 37621
rect 2866 37612 2872 37624
rect 2924 37612 2930 37664
rect 3053 37655 3111 37661
rect 3053 37621 3065 37655
rect 3099 37652 3111 37655
rect 3142 37652 3148 37664
rect 3099 37624 3148 37652
rect 3099 37621 3111 37624
rect 3053 37615 3111 37621
rect 3142 37612 3148 37624
rect 3200 37612 3206 37664
rect 4798 37612 4804 37664
rect 4856 37652 4862 37664
rect 5537 37655 5595 37661
rect 5537 37652 5549 37655
rect 4856 37624 5549 37652
rect 4856 37612 4862 37624
rect 5537 37621 5549 37624
rect 5583 37621 5595 37655
rect 5644 37652 5672 37692
rect 8018 37680 8024 37692
rect 8076 37680 8082 37732
rect 8110 37680 8116 37732
rect 8168 37720 8174 37732
rect 8220 37720 8248 37819
rect 12820 37788 12848 37819
rect 14458 37816 14464 37868
rect 14516 37816 14522 37868
rect 15105 37859 15163 37865
rect 15105 37825 15117 37859
rect 15151 37825 15163 37859
rect 15105 37819 15163 37825
rect 15381 37859 15439 37865
rect 15381 37825 15393 37859
rect 15427 37825 15439 37859
rect 15381 37819 15439 37825
rect 12894 37788 12900 37800
rect 12820 37760 12900 37788
rect 12894 37748 12900 37760
rect 12952 37788 12958 37800
rect 13081 37791 13139 37797
rect 13081 37788 13093 37791
rect 12952 37760 13093 37788
rect 12952 37748 12958 37760
rect 13081 37757 13093 37760
rect 13127 37757 13139 37791
rect 13081 37751 13139 37757
rect 13357 37791 13415 37797
rect 13357 37757 13369 37791
rect 13403 37788 13415 37791
rect 14090 37788 14096 37800
rect 13403 37760 14096 37788
rect 13403 37757 13415 37760
rect 13357 37751 13415 37757
rect 14090 37748 14096 37760
rect 14148 37748 14154 37800
rect 14829 37791 14887 37797
rect 14829 37757 14841 37791
rect 14875 37788 14887 37791
rect 15120 37788 15148 37819
rect 14875 37760 15148 37788
rect 14875 37757 14887 37760
rect 14829 37751 14887 37757
rect 8570 37720 8576 37732
rect 8168 37692 8576 37720
rect 8168 37680 8174 37692
rect 8570 37680 8576 37692
rect 8628 37680 8634 37732
rect 15289 37723 15347 37729
rect 15289 37689 15301 37723
rect 15335 37720 15347 37723
rect 15396 37720 15424 37819
rect 16850 37816 16856 37868
rect 16908 37816 16914 37868
rect 16960 37856 16988 37964
rect 18969 37961 18981 37995
rect 19015 37992 19027 37995
rect 19242 37992 19248 38004
rect 19015 37964 19248 37992
rect 19015 37961 19027 37964
rect 18969 37955 19027 37961
rect 19242 37952 19248 37964
rect 19300 37952 19306 38004
rect 19426 37952 19432 38004
rect 19484 37992 19490 38004
rect 19521 37995 19579 38001
rect 19521 37992 19533 37995
rect 19484 37964 19533 37992
rect 19484 37952 19490 37964
rect 19521 37961 19533 37964
rect 19567 37961 19579 37995
rect 19521 37955 19579 37961
rect 19610 37952 19616 38004
rect 19668 37992 19674 38004
rect 19668 37964 27384 37992
rect 19668 37952 19674 37964
rect 19153 37927 19211 37933
rect 19153 37893 19165 37927
rect 19199 37924 19211 37927
rect 20070 37924 20076 37936
rect 19199 37896 20076 37924
rect 19199 37893 19211 37896
rect 19153 37887 19211 37893
rect 18417 37859 18475 37865
rect 18417 37856 18429 37859
rect 16960 37828 18429 37856
rect 16960 37797 16988 37828
rect 18417 37825 18429 37828
rect 18463 37856 18475 37859
rect 18877 37859 18935 37865
rect 18877 37856 18889 37859
rect 18463 37828 18889 37856
rect 18463 37825 18475 37828
rect 18417 37819 18475 37825
rect 18877 37825 18889 37828
rect 18923 37825 18935 37859
rect 18877 37819 18935 37825
rect 19061 37859 19119 37865
rect 19061 37825 19073 37859
rect 19107 37856 19119 37859
rect 19168 37856 19196 37887
rect 20070 37884 20076 37896
rect 20128 37884 20134 37936
rect 22281 37927 22339 37933
rect 22281 37893 22293 37927
rect 22327 37924 22339 37927
rect 22370 37924 22376 37936
rect 22327 37896 22376 37924
rect 22327 37893 22339 37896
rect 22281 37887 22339 37893
rect 22370 37884 22376 37896
rect 22428 37884 22434 37936
rect 19107 37828 19196 37856
rect 19337 37859 19395 37865
rect 19107 37825 19119 37828
rect 19061 37819 19119 37825
rect 19337 37825 19349 37859
rect 19383 37856 19395 37859
rect 21358 37856 21364 37868
rect 19383 37828 21364 37856
rect 19383 37825 19395 37828
rect 19337 37819 19395 37825
rect 16945 37791 17003 37797
rect 16945 37757 16957 37791
rect 16991 37757 17003 37791
rect 16945 37751 17003 37757
rect 17221 37791 17279 37797
rect 17221 37757 17233 37791
rect 17267 37788 17279 37791
rect 17678 37788 17684 37800
rect 17267 37760 17684 37788
rect 17267 37757 17279 37760
rect 17221 37751 17279 37757
rect 17678 37748 17684 37760
rect 17736 37748 17742 37800
rect 18892 37788 18920 37819
rect 19352 37788 19380 37819
rect 21358 37816 21364 37828
rect 21416 37816 21422 37868
rect 21637 37859 21695 37865
rect 21637 37825 21649 37859
rect 21683 37856 21695 37859
rect 22189 37859 22247 37865
rect 22189 37856 22201 37859
rect 21683 37828 22201 37856
rect 21683 37825 21695 37828
rect 21637 37819 21695 37825
rect 22189 37825 22201 37828
rect 22235 37825 22247 37859
rect 22189 37819 22247 37825
rect 22646 37816 22652 37868
rect 22704 37856 22710 37868
rect 23017 37859 23075 37865
rect 23017 37856 23029 37859
rect 22704 37828 23029 37856
rect 22704 37816 22710 37828
rect 23017 37825 23029 37828
rect 23063 37825 23075 37859
rect 23017 37819 23075 37825
rect 24118 37816 24124 37868
rect 24176 37816 24182 37868
rect 27062 37816 27068 37868
rect 27120 37816 27126 37868
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27249 37819 27307 37825
rect 18892 37760 19380 37788
rect 19886 37748 19892 37800
rect 19944 37788 19950 37800
rect 20349 37791 20407 37797
rect 20349 37788 20361 37791
rect 19944 37760 20361 37788
rect 19944 37748 19950 37760
rect 20349 37757 20361 37760
rect 20395 37757 20407 37791
rect 20349 37751 20407 37757
rect 20990 37748 20996 37800
rect 21048 37748 21054 37800
rect 22462 37748 22468 37800
rect 22520 37748 22526 37800
rect 25406 37720 25412 37732
rect 15335 37692 25412 37720
rect 15335 37689 15347 37692
rect 15289 37683 15347 37689
rect 25406 37680 25412 37692
rect 25464 37680 25470 37732
rect 8386 37652 8392 37664
rect 5644 37624 8392 37652
rect 5537 37615 5595 37621
rect 8386 37612 8392 37624
rect 8444 37612 8450 37664
rect 18509 37655 18567 37661
rect 18509 37621 18521 37655
rect 18555 37652 18567 37655
rect 18966 37652 18972 37664
rect 18555 37624 18972 37652
rect 18555 37621 18567 37624
rect 18509 37615 18567 37621
rect 18966 37612 18972 37624
rect 19024 37612 19030 37664
rect 19610 37612 19616 37664
rect 19668 37652 19674 37664
rect 19797 37655 19855 37661
rect 19797 37652 19809 37655
rect 19668 37624 19809 37652
rect 19668 37612 19674 37624
rect 19797 37621 19809 37624
rect 19843 37621 19855 37655
rect 19797 37615 19855 37621
rect 21821 37655 21879 37661
rect 21821 37621 21833 37655
rect 21867 37652 21879 37655
rect 22094 37652 22100 37664
rect 21867 37624 22100 37652
rect 21867 37621 21879 37624
rect 21821 37615 21879 37621
rect 22094 37612 22100 37624
rect 22152 37612 22158 37664
rect 23566 37612 23572 37664
rect 23624 37612 23630 37664
rect 27264 37652 27292 37819
rect 27356 37720 27384 37964
rect 27614 37952 27620 38004
rect 27672 38001 27678 38004
rect 27672 37955 27681 38001
rect 27672 37952 27678 37955
rect 27982 37952 27988 38004
rect 28040 37952 28046 38004
rect 28626 37952 28632 38004
rect 28684 37952 28690 38004
rect 28902 37952 28908 38004
rect 28960 37992 28966 38004
rect 29089 37995 29147 38001
rect 29089 37992 29101 37995
rect 28960 37964 29101 37992
rect 28960 37952 28966 37964
rect 29089 37961 29101 37964
rect 29135 37961 29147 37995
rect 29089 37955 29147 37961
rect 29546 37952 29552 38004
rect 29604 37952 29610 38004
rect 29917 37995 29975 38001
rect 29917 37961 29929 37995
rect 29963 37992 29975 37995
rect 31386 37992 31392 38004
rect 29963 37964 31392 37992
rect 29963 37961 29975 37964
rect 29917 37955 29975 37961
rect 31386 37952 31392 37964
rect 31444 37952 31450 38004
rect 32674 37952 32680 38004
rect 32732 37992 32738 38004
rect 33413 37995 33471 38001
rect 33413 37992 33425 37995
rect 32732 37964 33425 37992
rect 32732 37952 32738 37964
rect 33413 37961 33425 37964
rect 33459 37961 33471 37995
rect 33413 37955 33471 37961
rect 33781 37995 33839 38001
rect 33781 37961 33793 37995
rect 33827 37992 33839 37995
rect 34698 37992 34704 38004
rect 33827 37964 34704 37992
rect 33827 37961 33839 37964
rect 33781 37955 33839 37961
rect 34698 37952 34704 37964
rect 34756 37952 34762 38004
rect 34790 37952 34796 38004
rect 34848 37952 34854 38004
rect 35986 37952 35992 38004
rect 36044 37952 36050 38004
rect 37918 37952 37924 38004
rect 37976 37992 37982 38004
rect 38013 37995 38071 38001
rect 38013 37992 38025 37995
rect 37976 37964 38025 37992
rect 37976 37952 37982 37964
rect 38013 37961 38025 37964
rect 38059 37961 38071 37995
rect 38013 37955 38071 37961
rect 40494 37952 40500 38004
rect 40552 37952 40558 38004
rect 27433 37927 27491 37933
rect 27433 37893 27445 37927
rect 27479 37924 27491 37927
rect 27709 37927 27767 37933
rect 27709 37924 27721 37927
rect 27479 37896 27721 37924
rect 27479 37893 27491 37896
rect 27433 37887 27491 37893
rect 27709 37893 27721 37896
rect 27755 37924 27767 37927
rect 28077 37927 28135 37933
rect 28077 37924 28089 37927
rect 27755 37896 28089 37924
rect 27755 37893 27767 37896
rect 27709 37887 27767 37893
rect 28077 37893 28089 37896
rect 28123 37893 28135 37927
rect 28077 37887 28135 37893
rect 28997 37927 29055 37933
rect 28997 37893 29009 37927
rect 29043 37924 29055 37927
rect 30469 37927 30527 37933
rect 29043 37896 29316 37924
rect 29043 37893 29055 37896
rect 28997 37887 29055 37893
rect 29288 37868 29316 37896
rect 30469 37893 30481 37927
rect 30515 37924 30527 37927
rect 30742 37924 30748 37936
rect 30515 37896 30748 37924
rect 30515 37893 30527 37896
rect 30469 37887 30527 37893
rect 30742 37884 30748 37896
rect 30800 37884 30806 37936
rect 32398 37924 32404 37936
rect 31680 37896 32404 37924
rect 27525 37859 27583 37865
rect 27525 37825 27537 37859
rect 27571 37825 27583 37859
rect 27525 37819 27583 37825
rect 27801 37859 27859 37865
rect 27801 37825 27813 37859
rect 27847 37856 27859 37859
rect 27890 37856 27896 37868
rect 27847 37828 27896 37856
rect 27847 37825 27859 37828
rect 27801 37819 27859 37825
rect 27540 37788 27568 37819
rect 27890 37816 27896 37828
rect 27948 37816 27954 37868
rect 28169 37859 28227 37865
rect 28169 37825 28181 37859
rect 28215 37825 28227 37859
rect 28169 37819 28227 37825
rect 28813 37859 28871 37865
rect 28813 37825 28825 37859
rect 28859 37856 28871 37859
rect 28902 37856 28908 37868
rect 28859 37828 28908 37856
rect 28859 37825 28871 37828
rect 28813 37819 28871 37825
rect 27982 37788 27988 37800
rect 27540 37760 27988 37788
rect 27982 37748 27988 37760
rect 28040 37788 28046 37800
rect 28184 37788 28212 37819
rect 28902 37816 28908 37828
rect 28960 37856 28966 37868
rect 29089 37859 29147 37865
rect 29089 37856 29101 37859
rect 28960 37828 29101 37856
rect 28960 37816 28966 37828
rect 29089 37825 29101 37828
rect 29135 37825 29147 37859
rect 29089 37819 29147 37825
rect 29270 37816 29276 37868
rect 29328 37816 29334 37868
rect 30190 37816 30196 37868
rect 30248 37856 30254 37868
rect 30377 37859 30435 37865
rect 30377 37856 30389 37859
rect 30248 37828 30389 37856
rect 30248 37816 30254 37828
rect 30377 37825 30389 37828
rect 30423 37825 30435 37859
rect 30377 37819 30435 37825
rect 30558 37816 30564 37868
rect 30616 37816 30622 37868
rect 31294 37816 31300 37868
rect 31352 37856 31358 37868
rect 31680 37865 31708 37896
rect 32398 37884 32404 37896
rect 32456 37924 32462 37936
rect 32861 37927 32919 37933
rect 32861 37924 32873 37927
rect 32456 37896 32873 37924
rect 32456 37884 32462 37896
rect 32861 37893 32873 37896
rect 32907 37893 32919 37927
rect 32861 37887 32919 37893
rect 32950 37884 32956 37936
rect 33008 37924 33014 37936
rect 33229 37927 33287 37933
rect 33229 37924 33241 37927
rect 33008 37896 33241 37924
rect 33008 37884 33014 37896
rect 33229 37893 33241 37896
rect 33275 37893 33287 37927
rect 33229 37887 33287 37893
rect 33873 37927 33931 37933
rect 33873 37893 33885 37927
rect 33919 37924 33931 37927
rect 35434 37924 35440 37936
rect 33919 37896 35440 37924
rect 33919 37893 33931 37896
rect 33873 37887 33931 37893
rect 35434 37884 35440 37896
rect 35492 37884 35498 37936
rect 39850 37884 39856 37936
rect 39908 37924 39914 37936
rect 40405 37927 40463 37933
rect 40405 37924 40417 37927
rect 39908 37896 40417 37924
rect 39908 37884 39914 37896
rect 40405 37893 40417 37896
rect 40451 37893 40463 37927
rect 40405 37887 40463 37893
rect 31665 37859 31723 37865
rect 31665 37856 31677 37859
rect 31352 37828 31677 37856
rect 31352 37816 31358 37828
rect 31665 37825 31677 37828
rect 31711 37825 31723 37859
rect 31665 37819 31723 37825
rect 32122 37816 32128 37868
rect 32180 37816 32186 37868
rect 33134 37816 33140 37868
rect 33192 37816 33198 37868
rect 33321 37859 33379 37865
rect 33321 37825 33333 37859
rect 33367 37856 33379 37859
rect 33410 37856 33416 37868
rect 33367 37828 33416 37856
rect 33367 37825 33379 37828
rect 33321 37819 33379 37825
rect 28040 37760 28212 37788
rect 28040 37748 28046 37760
rect 30006 37748 30012 37800
rect 30064 37748 30070 37800
rect 30098 37748 30104 37800
rect 30156 37748 30162 37800
rect 30576 37788 30604 37816
rect 33336 37788 33364 37819
rect 33410 37816 33416 37828
rect 33468 37816 33474 37868
rect 34425 37859 34483 37865
rect 34425 37825 34437 37859
rect 34471 37825 34483 37859
rect 34425 37819 34483 37825
rect 36357 37859 36415 37865
rect 36357 37825 36369 37859
rect 36403 37856 36415 37859
rect 37369 37859 37427 37865
rect 37369 37856 37381 37859
rect 36403 37828 37381 37856
rect 36403 37825 36415 37828
rect 36357 37819 36415 37825
rect 37369 37825 37381 37828
rect 37415 37825 37427 37859
rect 37369 37819 37427 37825
rect 37553 37859 37611 37865
rect 37553 37825 37565 37859
rect 37599 37825 37611 37859
rect 37553 37819 37611 37825
rect 30576 37760 33364 37788
rect 33965 37791 34023 37797
rect 33965 37757 33977 37791
rect 34011 37757 34023 37791
rect 33965 37751 34023 37757
rect 33980 37720 34008 37751
rect 34238 37748 34244 37800
rect 34296 37788 34302 37800
rect 34333 37791 34391 37797
rect 34333 37788 34345 37791
rect 34296 37760 34345 37788
rect 34296 37748 34302 37760
rect 34333 37757 34345 37760
rect 34379 37757 34391 37791
rect 34440 37788 34468 37819
rect 35434 37788 35440 37800
rect 34440 37760 35440 37788
rect 34333 37751 34391 37757
rect 35434 37748 35440 37760
rect 35492 37748 35498 37800
rect 36446 37748 36452 37800
rect 36504 37748 36510 37800
rect 37568 37788 37596 37819
rect 37642 37816 37648 37868
rect 37700 37856 37706 37868
rect 37829 37859 37887 37865
rect 37829 37856 37841 37859
rect 37700 37828 37841 37856
rect 37700 37816 37706 37828
rect 37829 37825 37841 37828
rect 37875 37856 37887 37859
rect 38227 37859 38285 37865
rect 38227 37856 38239 37859
rect 37875 37828 38239 37856
rect 37875 37825 37887 37828
rect 37829 37819 37887 37825
rect 38227 37825 38239 37828
rect 38273 37825 38285 37859
rect 38227 37819 38285 37825
rect 38381 37859 38439 37865
rect 38381 37825 38393 37859
rect 38427 37856 38439 37859
rect 38470 37856 38476 37868
rect 38427 37828 38476 37856
rect 38427 37825 38439 37828
rect 38381 37819 38439 37825
rect 38396 37788 38424 37819
rect 38470 37816 38476 37828
rect 38528 37816 38534 37868
rect 39942 37816 39948 37868
rect 40000 37816 40006 37868
rect 40034 37816 40040 37868
rect 40092 37856 40098 37868
rect 40129 37859 40187 37865
rect 40129 37856 40141 37859
rect 40092 37828 40141 37856
rect 40092 37816 40098 37828
rect 40129 37825 40141 37828
rect 40175 37825 40187 37859
rect 40129 37819 40187 37825
rect 40310 37816 40316 37868
rect 40368 37856 40374 37868
rect 40589 37859 40647 37865
rect 40589 37856 40601 37859
rect 40368 37828 40601 37856
rect 40368 37816 40374 37828
rect 40589 37825 40601 37828
rect 40635 37825 40647 37859
rect 40589 37819 40647 37825
rect 40678 37816 40684 37868
rect 40736 37816 40742 37868
rect 40770 37816 40776 37868
rect 40828 37856 40834 37868
rect 40957 37859 41015 37865
rect 40957 37856 40969 37859
rect 40828 37828 40969 37856
rect 40828 37816 40834 37828
rect 40957 37825 40969 37828
rect 41003 37825 41015 37859
rect 40957 37819 41015 37825
rect 41690 37816 41696 37868
rect 41748 37856 41754 37868
rect 41877 37859 41935 37865
rect 41877 37856 41889 37859
rect 41748 37828 41889 37856
rect 41748 37816 41754 37828
rect 41877 37825 41889 37828
rect 41923 37825 41935 37859
rect 41877 37819 41935 37825
rect 37568 37760 38424 37788
rect 34514 37720 34520 37732
rect 27356 37692 31754 37720
rect 28902 37652 28908 37664
rect 27264 37624 28908 37652
rect 28902 37612 28908 37624
rect 28960 37612 28966 37664
rect 31726 37652 31754 37692
rect 33980 37692 34520 37720
rect 33980 37652 34008 37692
rect 34514 37680 34520 37692
rect 34572 37680 34578 37732
rect 37366 37680 37372 37732
rect 37424 37720 37430 37732
rect 37568 37720 37596 37760
rect 37424 37692 37596 37720
rect 37645 37723 37703 37729
rect 37424 37680 37430 37692
rect 37645 37689 37657 37723
rect 37691 37689 37703 37723
rect 37645 37683 37703 37689
rect 31726 37624 34008 37652
rect 37458 37612 37464 37664
rect 37516 37652 37522 37664
rect 37660 37652 37688 37683
rect 37734 37680 37740 37732
rect 37792 37720 37798 37732
rect 38286 37720 38292 37732
rect 37792 37692 38292 37720
rect 37792 37680 37798 37692
rect 38286 37680 38292 37692
rect 38344 37680 38350 37732
rect 41506 37680 41512 37732
rect 41564 37720 41570 37732
rect 41693 37723 41751 37729
rect 41693 37720 41705 37723
rect 41564 37692 41705 37720
rect 41564 37680 41570 37692
rect 41693 37689 41705 37692
rect 41739 37689 41751 37723
rect 41693 37683 41751 37689
rect 39390 37652 39396 37664
rect 37516 37624 39396 37652
rect 37516 37612 37522 37624
rect 39390 37612 39396 37624
rect 39448 37612 39454 37664
rect 40310 37612 40316 37664
rect 40368 37612 40374 37664
rect 1104 37562 42504 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 42504 37562
rect 1104 37488 42504 37510
rect 1854 37408 1860 37460
rect 1912 37448 1918 37460
rect 3237 37451 3295 37457
rect 3237 37448 3249 37451
rect 1912 37420 3249 37448
rect 1912 37408 1918 37420
rect 3237 37417 3249 37420
rect 3283 37417 3295 37451
rect 3237 37411 3295 37417
rect 3418 37408 3424 37460
rect 3476 37408 3482 37460
rect 5524 37451 5582 37457
rect 5524 37417 5536 37451
rect 5570 37448 5582 37451
rect 5902 37448 5908 37460
rect 5570 37420 5908 37448
rect 5570 37417 5582 37420
rect 5524 37411 5582 37417
rect 5902 37408 5908 37420
rect 5960 37408 5966 37460
rect 7006 37408 7012 37460
rect 7064 37408 7070 37460
rect 7282 37408 7288 37460
rect 7340 37448 7346 37460
rect 8481 37451 8539 37457
rect 8481 37448 8493 37451
rect 7340 37420 8493 37448
rect 7340 37408 7346 37420
rect 8481 37417 8493 37420
rect 8527 37417 8539 37451
rect 8481 37411 8539 37417
rect 12066 37408 12072 37460
rect 12124 37448 12130 37460
rect 12124 37420 12434 37448
rect 12124 37408 12130 37420
rect 3145 37383 3203 37389
rect 3145 37380 3157 37383
rect 2746 37352 3157 37380
rect 1394 37272 1400 37324
rect 1452 37272 1458 37324
rect 2038 37272 2044 37324
rect 2096 37312 2102 37324
rect 2746 37312 2774 37352
rect 3145 37349 3157 37352
rect 3191 37380 3203 37383
rect 3694 37380 3700 37392
rect 3191 37352 3700 37380
rect 3191 37349 3203 37352
rect 3145 37343 3203 37349
rect 3694 37340 3700 37352
rect 3752 37380 3758 37392
rect 4062 37380 4068 37392
rect 3752 37352 4068 37380
rect 3752 37340 3758 37352
rect 4062 37340 4068 37352
rect 4120 37340 4126 37392
rect 4154 37340 4160 37392
rect 4212 37380 4218 37392
rect 5166 37380 5172 37392
rect 4212 37352 5172 37380
rect 4212 37340 4218 37352
rect 5166 37340 5172 37352
rect 5224 37340 5230 37392
rect 2096 37284 2774 37312
rect 2096 37272 2102 37284
rect 3786 37272 3792 37324
rect 3844 37312 3850 37324
rect 6822 37312 6828 37324
rect 3844 37284 6828 37312
rect 3844 37272 3850 37284
rect 2774 37204 2780 37256
rect 2832 37244 2838 37256
rect 2958 37244 2964 37256
rect 2832 37216 2964 37244
rect 2832 37204 2838 37216
rect 2958 37204 2964 37216
rect 3016 37204 3022 37256
rect 4724 37253 4752 37284
rect 4709 37247 4767 37253
rect 4709 37213 4721 37247
rect 4755 37213 4767 37247
rect 4709 37207 4767 37213
rect 4985 37247 5043 37253
rect 4985 37213 4997 37247
rect 5031 37213 5043 37247
rect 4985 37207 5043 37213
rect 1670 37136 1676 37188
rect 1728 37136 1734 37188
rect 3605 37179 3663 37185
rect 3605 37145 3617 37179
rect 3651 37176 3663 37179
rect 4798 37176 4804 37188
rect 3651 37148 4804 37176
rect 3651 37145 3663 37148
rect 3605 37139 3663 37145
rect 4798 37136 4804 37148
rect 4856 37176 4862 37188
rect 5000 37176 5028 37207
rect 5166 37204 5172 37256
rect 5224 37204 5230 37256
rect 5276 37253 5304 37284
rect 6822 37272 6828 37284
rect 6880 37272 6886 37324
rect 7024 37312 7052 37408
rect 7926 37340 7932 37392
rect 7984 37380 7990 37392
rect 9033 37383 9091 37389
rect 9033 37380 9045 37383
rect 7984 37352 9045 37380
rect 7984 37340 7990 37352
rect 9033 37349 9045 37352
rect 9079 37349 9091 37383
rect 12406 37380 12434 37420
rect 14090 37408 14096 37460
rect 14148 37408 14154 37460
rect 14458 37408 14464 37460
rect 14516 37448 14522 37460
rect 15102 37448 15108 37460
rect 14516 37420 15108 37448
rect 14516 37408 14522 37420
rect 15102 37408 15108 37420
rect 15160 37448 15166 37460
rect 15565 37451 15623 37457
rect 15565 37448 15577 37451
rect 15160 37420 15577 37448
rect 15160 37408 15166 37420
rect 15565 37417 15577 37420
rect 15611 37417 15623 37451
rect 15565 37411 15623 37417
rect 20625 37451 20683 37457
rect 20625 37417 20637 37451
rect 20671 37448 20683 37451
rect 20990 37448 20996 37460
rect 20671 37420 20996 37448
rect 20671 37417 20683 37420
rect 20625 37411 20683 37417
rect 20990 37408 20996 37420
rect 21048 37408 21054 37460
rect 24118 37408 24124 37460
rect 24176 37448 24182 37460
rect 24213 37451 24271 37457
rect 24213 37448 24225 37451
rect 24176 37420 24225 37448
rect 24176 37408 24182 37420
rect 24213 37417 24225 37420
rect 24259 37417 24271 37451
rect 24213 37411 24271 37417
rect 26050 37408 26056 37460
rect 26108 37448 26114 37460
rect 26145 37451 26203 37457
rect 26145 37448 26157 37451
rect 26108 37420 26157 37448
rect 26108 37408 26114 37420
rect 26145 37417 26157 37420
rect 26191 37448 26203 37451
rect 26326 37448 26332 37460
rect 26191 37420 26332 37448
rect 26191 37417 26203 37420
rect 26145 37411 26203 37417
rect 26326 37408 26332 37420
rect 26384 37408 26390 37460
rect 27982 37408 27988 37460
rect 28040 37408 28046 37460
rect 34238 37408 34244 37460
rect 34296 37408 34302 37460
rect 36446 37408 36452 37460
rect 36504 37408 36510 37460
rect 39390 37408 39396 37460
rect 39448 37408 39454 37460
rect 39850 37408 39856 37460
rect 39908 37448 39914 37460
rect 39945 37451 40003 37457
rect 39945 37448 39957 37451
rect 39908 37420 39957 37448
rect 39908 37408 39914 37420
rect 39945 37417 39957 37420
rect 39991 37417 40003 37451
rect 39945 37411 40003 37417
rect 14550 37380 14556 37392
rect 12406 37352 14556 37380
rect 9033 37343 9091 37349
rect 14550 37340 14556 37352
rect 14608 37340 14614 37392
rect 14734 37340 14740 37392
rect 14792 37380 14798 37392
rect 14792 37352 16068 37380
rect 14792 37340 14798 37352
rect 7024 37284 7696 37312
rect 5261 37247 5319 37253
rect 5261 37213 5273 37247
rect 5307 37213 5319 37247
rect 5261 37207 5319 37213
rect 7098 37204 7104 37256
rect 7156 37204 7162 37256
rect 7668 37253 7696 37284
rect 8312 37284 8800 37312
rect 8312 37256 8340 37284
rect 7653 37247 7711 37253
rect 7653 37213 7665 37247
rect 7699 37244 7711 37247
rect 8113 37247 8171 37253
rect 8113 37244 8125 37247
rect 7699 37216 8125 37244
rect 7699 37213 7711 37216
rect 7653 37207 7711 37213
rect 8113 37213 8125 37216
rect 8159 37213 8171 37247
rect 8113 37207 8171 37213
rect 8205 37247 8263 37253
rect 8205 37213 8217 37247
rect 8251 37244 8263 37247
rect 8294 37244 8300 37256
rect 8251 37216 8300 37244
rect 8251 37213 8263 37216
rect 8205 37207 8263 37213
rect 8294 37204 8300 37216
rect 8352 37204 8358 37256
rect 8481 37247 8539 37253
rect 8481 37213 8493 37247
rect 8527 37213 8539 37247
rect 8481 37207 8539 37213
rect 4856 37148 5028 37176
rect 4856 37136 4862 37148
rect 3405 37111 3463 37117
rect 3405 37077 3417 37111
rect 3451 37108 3463 37111
rect 4154 37108 4160 37120
rect 3451 37080 4160 37108
rect 3451 37077 3463 37080
rect 3405 37071 3463 37077
rect 4154 37068 4160 37080
rect 4212 37068 4218 37120
rect 4430 37068 4436 37120
rect 4488 37108 4494 37120
rect 4985 37111 5043 37117
rect 4985 37108 4997 37111
rect 4488 37080 4997 37108
rect 4488 37068 4494 37080
rect 4985 37077 4997 37080
rect 5031 37077 5043 37111
rect 5184 37108 5212 37204
rect 6762 37148 6868 37176
rect 5350 37108 5356 37120
rect 5184 37080 5356 37108
rect 4985 37071 5043 37077
rect 5350 37068 5356 37080
rect 5408 37068 5414 37120
rect 5534 37068 5540 37120
rect 5592 37108 5598 37120
rect 6362 37108 6368 37120
rect 5592 37080 6368 37108
rect 5592 37068 5598 37080
rect 6362 37068 6368 37080
rect 6420 37108 6426 37120
rect 6840 37108 6868 37148
rect 6914 37136 6920 37188
rect 6972 37176 6978 37188
rect 7837 37179 7895 37185
rect 7837 37176 7849 37179
rect 6972 37148 7849 37176
rect 6972 37136 6978 37148
rect 7837 37145 7849 37148
rect 7883 37176 7895 37179
rect 8496 37176 8524 37207
rect 8570 37204 8576 37256
rect 8628 37204 8634 37256
rect 8772 37253 8800 37284
rect 9674 37272 9680 37324
rect 9732 37312 9738 37324
rect 13357 37315 13415 37321
rect 13357 37312 13369 37315
rect 9732 37284 13369 37312
rect 9732 37272 9738 37284
rect 13357 37281 13369 37284
rect 13403 37281 13415 37315
rect 15010 37312 15016 37324
rect 13357 37275 13415 37281
rect 14476 37284 15016 37312
rect 8757 37247 8815 37253
rect 8757 37213 8769 37247
rect 8803 37213 8815 37247
rect 8757 37207 8815 37213
rect 8941 37247 8999 37253
rect 8941 37213 8953 37247
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 7883 37148 8524 37176
rect 7883 37145 7895 37148
rect 7837 37139 7895 37145
rect 8128 37120 8156 37148
rect 7466 37108 7472 37120
rect 6420 37080 7472 37108
rect 6420 37068 6426 37080
rect 7466 37068 7472 37080
rect 7524 37068 7530 37120
rect 8018 37068 8024 37120
rect 8076 37068 8082 37120
rect 8110 37068 8116 37120
rect 8168 37068 8174 37120
rect 8386 37068 8392 37120
rect 8444 37108 8450 37120
rect 8956 37108 8984 37207
rect 12250 37204 12256 37256
rect 12308 37204 12314 37256
rect 12526 37204 12532 37256
rect 12584 37244 12590 37256
rect 13541 37247 13599 37253
rect 13541 37244 13553 37247
rect 12584 37216 13553 37244
rect 12584 37204 12590 37216
rect 13541 37213 13553 37216
rect 13587 37213 13599 37247
rect 13541 37207 13599 37213
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37244 14335 37247
rect 14366 37244 14372 37256
rect 14323 37216 14372 37244
rect 14323 37213 14335 37216
rect 14277 37207 14335 37213
rect 14366 37204 14372 37216
rect 14424 37204 14430 37256
rect 14476 37253 14504 37284
rect 15010 37272 15016 37284
rect 15068 37272 15074 37324
rect 16040 37321 16068 37352
rect 15289 37315 15347 37321
rect 15289 37281 15301 37315
rect 15335 37281 15347 37315
rect 15289 37275 15347 37281
rect 16025 37315 16083 37321
rect 16025 37281 16037 37315
rect 16071 37281 16083 37315
rect 16025 37275 16083 37281
rect 16301 37315 16359 37321
rect 16301 37281 16313 37315
rect 16347 37312 16359 37315
rect 17310 37312 17316 37324
rect 16347 37284 17316 37312
rect 16347 37281 16359 37284
rect 16301 37275 16359 37281
rect 14461 37247 14519 37253
rect 14461 37213 14473 37247
rect 14507 37213 14519 37247
rect 14461 37207 14519 37213
rect 14550 37204 14556 37256
rect 14608 37204 14614 37256
rect 12158 37136 12164 37188
rect 12216 37176 12222 37188
rect 12345 37179 12403 37185
rect 12345 37176 12357 37179
rect 12216 37148 12357 37176
rect 12216 37136 12222 37148
rect 12345 37145 12357 37148
rect 12391 37145 12403 37179
rect 12345 37139 12403 37145
rect 12894 37136 12900 37188
rect 12952 37176 12958 37188
rect 13081 37179 13139 37185
rect 13081 37176 13093 37179
rect 12952 37148 13093 37176
rect 12952 37136 12958 37148
rect 13081 37145 13093 37148
rect 13127 37145 13139 37179
rect 15304 37176 15332 37275
rect 17310 37272 17316 37284
rect 17368 37272 17374 37324
rect 17678 37272 17684 37324
rect 17736 37312 17742 37324
rect 18601 37315 18659 37321
rect 18601 37312 18613 37315
rect 17736 37284 18613 37312
rect 17736 37272 17742 37284
rect 18601 37281 18613 37284
rect 18647 37281 18659 37315
rect 18601 37275 18659 37281
rect 19702 37272 19708 37324
rect 19760 37312 19766 37324
rect 19797 37315 19855 37321
rect 19797 37312 19809 37315
rect 19760 37284 19809 37312
rect 19760 37272 19766 37284
rect 19797 37281 19809 37284
rect 19843 37281 19855 37315
rect 19797 37275 19855 37281
rect 22094 37272 22100 37324
rect 22152 37272 22158 37324
rect 24673 37315 24731 37321
rect 24673 37281 24685 37315
rect 24719 37312 24731 37315
rect 25038 37312 25044 37324
rect 24719 37284 25044 37312
rect 24719 37281 24731 37284
rect 24673 37275 24731 37281
rect 25038 37272 25044 37284
rect 25096 37272 25102 37324
rect 28000 37312 28028 37408
rect 28902 37340 28908 37392
rect 28960 37380 28966 37392
rect 29089 37383 29147 37389
rect 29089 37380 29101 37383
rect 28960 37352 29101 37380
rect 28960 37340 28966 37352
rect 29089 37349 29101 37352
rect 29135 37380 29147 37383
rect 30558 37380 30564 37392
rect 29135 37352 30564 37380
rect 29135 37349 29147 37352
rect 29089 37343 29147 37349
rect 30558 37340 30564 37352
rect 30616 37340 30622 37392
rect 34885 37383 34943 37389
rect 34885 37349 34897 37383
rect 34931 37380 34943 37383
rect 35342 37380 35348 37392
rect 34931 37352 35348 37380
rect 34931 37349 34943 37352
rect 34885 37343 34943 37349
rect 35342 37340 35348 37352
rect 35400 37380 35406 37392
rect 36357 37383 36415 37389
rect 35400 37352 35894 37380
rect 35400 37340 35406 37352
rect 28629 37315 28687 37321
rect 28629 37312 28641 37315
rect 28000 37284 28641 37312
rect 28629 37281 28641 37284
rect 28675 37281 28687 37315
rect 28629 37275 28687 37281
rect 30098 37272 30104 37324
rect 30156 37312 30162 37324
rect 31757 37315 31815 37321
rect 31757 37312 31769 37315
rect 30156 37284 31769 37312
rect 30156 37272 30162 37284
rect 31757 37281 31769 37284
rect 31803 37281 31815 37315
rect 31757 37275 31815 37281
rect 34057 37315 34115 37321
rect 34057 37281 34069 37315
rect 34103 37312 34115 37315
rect 34977 37315 35035 37321
rect 34103 37284 34836 37312
rect 34103 37281 34115 37284
rect 34057 37275 34115 37281
rect 17586 37244 17592 37256
rect 17434 37216 17592 37244
rect 17586 37204 17592 37216
rect 17644 37204 17650 37256
rect 17770 37204 17776 37256
rect 17828 37244 17834 37256
rect 18417 37247 18475 37253
rect 18417 37244 18429 37247
rect 17828 37216 18429 37244
rect 17828 37204 17834 37216
rect 18417 37213 18429 37216
rect 18463 37213 18475 37247
rect 18417 37207 18475 37213
rect 18782 37204 18788 37256
rect 18840 37204 18846 37256
rect 18966 37204 18972 37256
rect 19024 37204 19030 37256
rect 19061 37247 19119 37253
rect 19061 37213 19073 37247
rect 19107 37213 19119 37247
rect 19061 37207 19119 37213
rect 15841 37179 15899 37185
rect 15304 37148 15424 37176
rect 13081 37139 13139 37145
rect 15396 37120 15424 37148
rect 15841 37145 15853 37179
rect 15887 37176 15899 37179
rect 16206 37176 16212 37188
rect 15887 37148 16212 37176
rect 15887 37145 15899 37148
rect 15841 37139 15899 37145
rect 16206 37136 16212 37148
rect 16264 37136 16270 37188
rect 19076 37176 19104 37207
rect 19610 37204 19616 37256
rect 19668 37204 19674 37256
rect 22373 37247 22431 37253
rect 22373 37213 22385 37247
rect 22419 37244 22431 37247
rect 22465 37247 22523 37253
rect 22465 37244 22477 37247
rect 22419 37216 22477 37244
rect 22419 37213 22431 37216
rect 22373 37207 22431 37213
rect 22465 37213 22477 37216
rect 22511 37213 22523 37247
rect 22465 37207 22523 37213
rect 17604 37148 19104 37176
rect 8444 37080 8984 37108
rect 8444 37068 8450 37080
rect 14550 37068 14556 37120
rect 14608 37108 14614 37120
rect 14645 37111 14703 37117
rect 14645 37108 14657 37111
rect 14608 37080 14657 37108
rect 14608 37068 14614 37080
rect 14645 37077 14657 37080
rect 14691 37077 14703 37111
rect 14645 37071 14703 37077
rect 15378 37068 15384 37120
rect 15436 37108 15442 37120
rect 17604 37108 17632 37148
rect 21542 37136 21548 37188
rect 21600 37136 21606 37188
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 22480 37176 22508 37207
rect 24394 37204 24400 37256
rect 24452 37204 24458 37256
rect 25774 37204 25780 37256
rect 25832 37204 25838 37256
rect 26237 37247 26295 37253
rect 26237 37213 26249 37247
rect 26283 37213 26295 37247
rect 29454 37244 29460 37256
rect 27646 37216 29460 37244
rect 26237 37207 26295 37213
rect 22646 37176 22652 37188
rect 22244 37148 22652 37176
rect 22244 37136 22250 37148
rect 22646 37136 22652 37148
rect 22704 37136 22710 37188
rect 22738 37136 22744 37188
rect 22796 37136 22802 37188
rect 25130 37176 25136 37188
rect 23966 37148 25136 37176
rect 25130 37136 25136 37148
rect 25188 37136 25194 37188
rect 15436 37080 17632 37108
rect 15436 37068 15442 37080
rect 17770 37068 17776 37120
rect 17828 37068 17834 37120
rect 17862 37068 17868 37120
rect 17920 37068 17926 37120
rect 19242 37068 19248 37120
rect 19300 37068 19306 37120
rect 19705 37111 19763 37117
rect 19705 37077 19717 37111
rect 19751 37108 19763 37111
rect 19794 37108 19800 37120
rect 19751 37080 19800 37108
rect 19751 37077 19763 37080
rect 19705 37071 19763 37077
rect 19794 37068 19800 37080
rect 19852 37068 19858 37120
rect 24394 37068 24400 37120
rect 24452 37108 24458 37120
rect 26252 37108 26280 37207
rect 29454 37204 29460 37216
rect 29512 37204 29518 37256
rect 29546 37204 29552 37256
rect 29604 37244 29610 37256
rect 30190 37244 30196 37256
rect 29604 37216 30196 37244
rect 29604 37204 29610 37216
rect 30190 37204 30196 37216
rect 30248 37204 30254 37256
rect 31772 37244 31800 37275
rect 31846 37244 31852 37256
rect 31772 37216 31852 37244
rect 31846 37204 31852 37216
rect 31904 37204 31910 37256
rect 31938 37204 31944 37256
rect 31996 37244 32002 37256
rect 32585 37247 32643 37253
rect 32585 37244 32597 37247
rect 31996 37216 32597 37244
rect 31996 37204 32002 37216
rect 32585 37213 32597 37216
rect 32631 37213 32643 37247
rect 32585 37207 32643 37213
rect 32766 37204 32772 37256
rect 32824 37244 32830 37256
rect 33134 37244 33140 37256
rect 32824 37216 33140 37244
rect 32824 37204 32830 37216
rect 33134 37204 33140 37216
rect 33192 37204 33198 37256
rect 33962 37204 33968 37256
rect 34020 37204 34026 37256
rect 34146 37204 34152 37256
rect 34204 37244 34210 37256
rect 34808 37253 34836 37284
rect 34977 37281 34989 37315
rect 35023 37312 35035 37315
rect 35866 37312 35894 37352
rect 36357 37349 36369 37383
rect 36403 37380 36415 37383
rect 36906 37380 36912 37392
rect 36403 37352 36912 37380
rect 36403 37349 36415 37352
rect 36357 37343 36415 37349
rect 36906 37340 36912 37352
rect 36964 37340 36970 37392
rect 37458 37340 37464 37392
rect 37516 37340 37522 37392
rect 37553 37383 37611 37389
rect 37553 37349 37565 37383
rect 37599 37380 37611 37383
rect 37734 37380 37740 37392
rect 37599 37352 37740 37380
rect 37599 37349 37611 37352
rect 37553 37343 37611 37349
rect 37734 37340 37740 37352
rect 37792 37340 37798 37392
rect 37185 37315 37243 37321
rect 37185 37312 37197 37315
rect 35023 37284 35572 37312
rect 35866 37284 37197 37312
rect 35023 37281 35035 37284
rect 34977 37275 35035 37281
rect 34241 37247 34299 37253
rect 34241 37244 34253 37247
rect 34204 37216 34253 37244
rect 34204 37204 34210 37216
rect 34241 37213 34253 37216
rect 34287 37213 34299 37247
rect 34241 37207 34299 37213
rect 34425 37247 34483 37253
rect 34425 37213 34437 37247
rect 34471 37213 34483 37247
rect 34425 37207 34483 37213
rect 34793 37247 34851 37253
rect 34793 37213 34805 37247
rect 34839 37213 34851 37247
rect 34793 37207 34851 37213
rect 35069 37247 35127 37253
rect 35069 37213 35081 37247
rect 35115 37213 35127 37247
rect 35069 37207 35127 37213
rect 26510 37136 26516 37188
rect 26568 37136 26574 37188
rect 28166 37136 28172 37188
rect 28224 37176 28230 37188
rect 28905 37179 28963 37185
rect 28905 37176 28917 37179
rect 28224 37148 28917 37176
rect 28224 37136 28230 37148
rect 28905 37145 28917 37148
rect 28951 37176 28963 37179
rect 31386 37176 31392 37188
rect 28951 37148 31392 37176
rect 28951 37145 28963 37148
rect 28905 37139 28963 37145
rect 31386 37136 31392 37148
rect 31444 37136 31450 37188
rect 31573 37179 31631 37185
rect 31573 37145 31585 37179
rect 31619 37176 31631 37179
rect 32033 37179 32091 37185
rect 32033 37176 32045 37179
rect 31619 37148 32045 37176
rect 31619 37145 31631 37148
rect 31573 37139 31631 37145
rect 32033 37145 32045 37148
rect 32079 37145 32091 37179
rect 32033 37139 32091 37145
rect 32953 37179 33011 37185
rect 32953 37145 32965 37179
rect 32999 37145 33011 37179
rect 34440 37176 34468 37207
rect 34514 37176 34520 37188
rect 34440 37148 34520 37176
rect 32953 37139 33011 37145
rect 24452 37080 26280 37108
rect 24452 37068 24458 37080
rect 28074 37068 28080 37120
rect 28132 37068 28138 37120
rect 29638 37068 29644 37120
rect 29696 37068 29702 37120
rect 30466 37068 30472 37120
rect 30524 37108 30530 37120
rect 31205 37111 31263 37117
rect 31205 37108 31217 37111
rect 30524 37080 31217 37108
rect 30524 37068 30530 37080
rect 31205 37077 31217 37080
rect 31251 37077 31263 37111
rect 31205 37071 31263 37077
rect 31662 37068 31668 37120
rect 31720 37068 31726 37120
rect 32490 37068 32496 37120
rect 32548 37108 32554 37120
rect 32769 37111 32827 37117
rect 32769 37108 32781 37111
rect 32548 37080 32781 37108
rect 32548 37068 32554 37080
rect 32769 37077 32781 37080
rect 32815 37077 32827 37111
rect 32968 37108 32996 37139
rect 34514 37136 34520 37148
rect 34572 37176 34578 37188
rect 35084 37176 35112 37207
rect 35250 37204 35256 37256
rect 35308 37204 35314 37256
rect 35342 37204 35348 37256
rect 35400 37204 35406 37256
rect 35434 37204 35440 37256
rect 35492 37204 35498 37256
rect 35544 37253 35572 37284
rect 37185 37281 37197 37284
rect 37231 37281 37243 37315
rect 39868 37312 39896 37408
rect 37185 37275 37243 37281
rect 39684 37284 39896 37312
rect 40129 37315 40187 37321
rect 35529 37247 35587 37253
rect 35529 37213 35541 37247
rect 35575 37244 35587 37247
rect 35575 37216 35894 37244
rect 35575 37213 35587 37216
rect 35529 37207 35587 37213
rect 35866 37176 35894 37216
rect 37366 37204 37372 37256
rect 37424 37204 37430 37256
rect 37642 37204 37648 37256
rect 37700 37204 37706 37256
rect 39684 37253 39712 37284
rect 40129 37281 40141 37315
rect 40175 37312 40187 37315
rect 40770 37312 40776 37324
rect 40175 37284 40776 37312
rect 40175 37281 40187 37284
rect 40129 37275 40187 37281
rect 40770 37272 40776 37284
rect 40828 37272 40834 37324
rect 37829 37247 37887 37253
rect 37829 37213 37841 37247
rect 37875 37213 37887 37247
rect 37829 37207 37887 37213
rect 39669 37247 39727 37253
rect 39669 37213 39681 37247
rect 39715 37213 39727 37247
rect 39669 37207 39727 37213
rect 39853 37247 39911 37253
rect 39853 37213 39865 37247
rect 39899 37244 39911 37247
rect 39942 37244 39948 37256
rect 39899 37216 39948 37244
rect 39899 37213 39911 37216
rect 39853 37207 39911 37213
rect 35986 37176 35992 37188
rect 34572 37148 35112 37176
rect 35176 37148 35388 37176
rect 35866 37148 35992 37176
rect 34572 37136 34578 37148
rect 33410 37108 33416 37120
rect 32968 37080 33416 37108
rect 32769 37071 32827 37077
rect 33410 37068 33416 37080
rect 33468 37108 33474 37120
rect 35176 37108 35204 37148
rect 33468 37080 35204 37108
rect 35360 37108 35388 37148
rect 35986 37136 35992 37148
rect 36044 37136 36050 37188
rect 36906 37136 36912 37188
rect 36964 37176 36970 37188
rect 37844 37176 37872 37207
rect 39942 37204 39948 37216
rect 40000 37204 40006 37256
rect 40034 37204 40040 37256
rect 40092 37204 40098 37256
rect 36964 37148 37872 37176
rect 39393 37179 39451 37185
rect 36964 37136 36970 37148
rect 39393 37145 39405 37179
rect 39439 37145 39451 37179
rect 39393 37139 39451 37145
rect 39577 37179 39635 37185
rect 39577 37145 39589 37179
rect 39623 37176 39635 37179
rect 40310 37176 40316 37188
rect 39623 37148 40316 37176
rect 39623 37145 39635 37148
rect 39577 37139 39635 37145
rect 36262 37108 36268 37120
rect 35360 37080 36268 37108
rect 33468 37068 33474 37080
rect 36262 37068 36268 37080
rect 36320 37068 36326 37120
rect 39408 37108 39436 37139
rect 40310 37136 40316 37148
rect 40368 37136 40374 37188
rect 40402 37136 40408 37188
rect 40460 37136 40466 37188
rect 40494 37136 40500 37188
rect 40552 37176 40558 37188
rect 40552 37148 40894 37176
rect 40552 37136 40558 37148
rect 40678 37108 40684 37120
rect 39408 37080 40684 37108
rect 40678 37068 40684 37080
rect 40736 37108 40742 37120
rect 41874 37108 41880 37120
rect 40736 37080 41880 37108
rect 40736 37068 40742 37080
rect 41874 37068 41880 37080
rect 41932 37068 41938 37120
rect 1104 37018 42504 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 42504 37018
rect 1104 36944 42504 36966
rect 1670 36864 1676 36916
rect 1728 36904 1734 36916
rect 2501 36907 2559 36913
rect 2501 36904 2513 36907
rect 1728 36876 2513 36904
rect 1728 36864 1734 36876
rect 2501 36873 2513 36876
rect 2547 36873 2559 36907
rect 2866 36904 2872 36916
rect 2501 36867 2559 36873
rect 2792 36876 2872 36904
rect 2792 36845 2820 36876
rect 2866 36864 2872 36876
rect 2924 36864 2930 36916
rect 4249 36907 4307 36913
rect 4249 36873 4261 36907
rect 4295 36904 4307 36907
rect 4614 36904 4620 36916
rect 4295 36876 4620 36904
rect 4295 36873 4307 36876
rect 4249 36867 4307 36873
rect 4614 36864 4620 36876
rect 4672 36864 4678 36916
rect 5166 36864 5172 36916
rect 5224 36864 5230 36916
rect 5350 36864 5356 36916
rect 5408 36864 5414 36916
rect 6914 36864 6920 36916
rect 6972 36864 6978 36916
rect 8110 36864 8116 36916
rect 8168 36904 8174 36916
rect 8573 36907 8631 36913
rect 8573 36904 8585 36907
rect 8168 36876 8585 36904
rect 8168 36864 8174 36876
rect 8573 36873 8585 36876
rect 8619 36873 8631 36907
rect 12526 36904 12532 36916
rect 8573 36867 8631 36873
rect 9048 36876 12532 36904
rect 2777 36839 2835 36845
rect 2777 36805 2789 36839
rect 2823 36805 2835 36839
rect 2777 36799 2835 36805
rect 3007 36839 3065 36845
rect 3007 36805 3019 36839
rect 3053 36836 3065 36839
rect 3421 36839 3479 36845
rect 3053 36808 3372 36836
rect 3053 36805 3065 36808
rect 3007 36799 3065 36805
rect 2685 36771 2743 36777
rect 2685 36737 2697 36771
rect 2731 36737 2743 36771
rect 2685 36731 2743 36737
rect 2700 36700 2728 36731
rect 2866 36728 2872 36780
rect 2924 36728 2930 36780
rect 3142 36728 3148 36780
rect 3200 36728 3206 36780
rect 3344 36768 3372 36808
rect 3421 36805 3433 36839
rect 3467 36836 3479 36839
rect 3786 36836 3792 36848
rect 3467 36808 3792 36836
rect 3467 36805 3479 36808
rect 3421 36799 3479 36805
rect 3786 36796 3792 36808
rect 3844 36796 3850 36848
rect 4157 36839 4215 36845
rect 4157 36805 4169 36839
rect 4203 36836 4215 36839
rect 6638 36836 6644 36848
rect 4203 36808 6644 36836
rect 4203 36805 4215 36808
rect 4157 36799 4215 36805
rect 6638 36796 6644 36808
rect 6696 36796 6702 36848
rect 6932 36836 6960 36864
rect 9048 36845 9076 36876
rect 12526 36864 12532 36876
rect 12584 36864 12590 36916
rect 14182 36864 14188 36916
rect 14240 36904 14246 36916
rect 14645 36907 14703 36913
rect 14240 36876 14504 36904
rect 14240 36864 14246 36876
rect 8665 36839 8723 36845
rect 8665 36836 8677 36839
rect 6748 36808 6960 36836
rect 8326 36822 8677 36836
rect 8312 36808 8677 36822
rect 3510 36768 3516 36780
rect 3344 36740 3516 36768
rect 3510 36728 3516 36740
rect 3568 36728 3574 36780
rect 4430 36728 4436 36780
rect 4488 36728 4494 36780
rect 4522 36728 4528 36780
rect 4580 36728 4586 36780
rect 4617 36771 4675 36777
rect 4617 36737 4629 36771
rect 4663 36737 4675 36771
rect 4617 36731 4675 36737
rect 4755 36771 4813 36777
rect 4755 36737 4767 36771
rect 4801 36768 4813 36771
rect 4982 36768 4988 36780
rect 4801 36740 4988 36768
rect 4801 36737 4813 36740
rect 4755 36731 4813 36737
rect 3234 36700 3240 36712
rect 2700 36672 3240 36700
rect 3234 36660 3240 36672
rect 3292 36660 3298 36712
rect 3326 36660 3332 36712
rect 3384 36700 3390 36712
rect 4338 36700 4344 36712
rect 3384 36672 4344 36700
rect 3384 36660 3390 36672
rect 4338 36660 4344 36672
rect 4396 36700 4402 36712
rect 4632 36700 4660 36731
rect 4982 36728 4988 36740
rect 5040 36728 5046 36780
rect 5261 36771 5319 36777
rect 5092 36766 5212 36768
rect 5261 36766 5273 36771
rect 5092 36740 5273 36766
rect 4396 36672 4660 36700
rect 4893 36703 4951 36709
rect 4396 36660 4402 36672
rect 4893 36669 4905 36703
rect 4939 36700 4951 36703
rect 4939 36672 4973 36700
rect 4939 36669 4951 36672
rect 4893 36663 4951 36669
rect 4798 36592 4804 36644
rect 4856 36632 4862 36644
rect 4908 36632 4936 36663
rect 4985 36635 5043 36641
rect 4985 36632 4997 36635
rect 4856 36604 4997 36632
rect 4856 36592 4862 36604
rect 4985 36601 4997 36604
rect 5031 36601 5043 36635
rect 4985 36595 5043 36601
rect 4062 36524 4068 36576
rect 4120 36564 4126 36576
rect 5092 36564 5120 36740
rect 5184 36738 5273 36740
rect 5261 36737 5273 36738
rect 5307 36737 5319 36771
rect 5261 36731 5319 36737
rect 6546 36728 6552 36780
rect 6604 36728 6610 36780
rect 6748 36777 6776 36808
rect 6733 36771 6791 36777
rect 6733 36737 6745 36771
rect 6779 36737 6791 36771
rect 6733 36731 6791 36737
rect 6822 36660 6828 36712
rect 6880 36660 6886 36712
rect 7101 36703 7159 36709
rect 7101 36669 7113 36703
rect 7147 36700 7159 36703
rect 7190 36700 7196 36712
rect 7147 36672 7196 36700
rect 7147 36669 7159 36672
rect 7101 36663 7159 36669
rect 7190 36660 7196 36672
rect 7248 36660 7254 36712
rect 7466 36660 7472 36712
rect 7524 36700 7530 36712
rect 8312 36700 8340 36808
rect 8665 36805 8677 36808
rect 8711 36805 8723 36839
rect 8665 36799 8723 36805
rect 9033 36839 9091 36845
rect 9033 36805 9045 36839
rect 9079 36805 9091 36839
rect 9033 36799 9091 36805
rect 10336 36808 12664 36836
rect 10336 36777 10364 36808
rect 12636 36780 12664 36808
rect 13170 36796 13176 36848
rect 13228 36796 13234 36848
rect 14476 36836 14504 36876
rect 14645 36873 14657 36907
rect 14691 36904 14703 36907
rect 15378 36904 15384 36916
rect 14691 36876 15384 36904
rect 14691 36873 14703 36876
rect 14645 36867 14703 36873
rect 15378 36864 15384 36876
rect 15436 36864 15442 36916
rect 16485 36907 16543 36913
rect 16485 36873 16497 36907
rect 16531 36904 16543 36907
rect 16850 36904 16856 36916
rect 16531 36876 16856 36904
rect 16531 36873 16543 36876
rect 16485 36867 16543 36873
rect 16850 36864 16856 36876
rect 16908 36864 16914 36916
rect 17310 36864 17316 36916
rect 17368 36904 17374 36916
rect 17405 36907 17463 36913
rect 17405 36904 17417 36907
rect 17368 36876 17417 36904
rect 17368 36864 17374 36876
rect 17405 36873 17417 36876
rect 17451 36873 17463 36907
rect 17405 36867 17463 36873
rect 17586 36864 17592 36916
rect 17644 36904 17650 36916
rect 19242 36904 19248 36916
rect 17644 36876 18092 36904
rect 17644 36864 17650 36876
rect 15102 36836 15108 36848
rect 14398 36808 15108 36836
rect 15102 36796 15108 36808
rect 15160 36836 15166 36848
rect 15160 36808 15502 36836
rect 15160 36796 15166 36808
rect 10321 36771 10379 36777
rect 10321 36737 10333 36771
rect 10367 36737 10379 36771
rect 10321 36731 10379 36737
rect 10505 36771 10563 36777
rect 10505 36737 10517 36771
rect 10551 36737 10563 36771
rect 10505 36731 10563 36737
rect 10597 36771 10655 36777
rect 10597 36737 10609 36771
rect 10643 36737 10655 36771
rect 10597 36731 10655 36737
rect 7524 36672 8340 36700
rect 7524 36660 7530 36672
rect 10042 36660 10048 36712
rect 10100 36700 10106 36712
rect 10520 36700 10548 36731
rect 10100 36672 10548 36700
rect 10100 36660 10106 36672
rect 4120 36536 5120 36564
rect 5537 36567 5595 36573
rect 4120 36524 4126 36536
rect 5537 36533 5549 36567
rect 5583 36564 5595 36567
rect 5626 36564 5632 36576
rect 5583 36536 5632 36564
rect 5583 36533 5595 36536
rect 5537 36527 5595 36533
rect 5626 36524 5632 36536
rect 5684 36524 5690 36576
rect 6641 36567 6699 36573
rect 6641 36533 6653 36567
rect 6687 36564 6699 36567
rect 7098 36564 7104 36576
rect 6687 36536 7104 36564
rect 6687 36533 6699 36536
rect 6641 36527 6699 36533
rect 7098 36524 7104 36536
rect 7156 36524 7162 36576
rect 9858 36524 9864 36576
rect 9916 36564 9922 36576
rect 10137 36567 10195 36573
rect 10137 36564 10149 36567
rect 9916 36536 10149 36564
rect 9916 36524 9922 36536
rect 10137 36533 10149 36536
rect 10183 36533 10195 36567
rect 10137 36527 10195 36533
rect 10502 36524 10508 36576
rect 10560 36564 10566 36576
rect 10612 36564 10640 36731
rect 11974 36728 11980 36780
rect 12032 36768 12038 36780
rect 12437 36771 12495 36777
rect 12437 36768 12449 36771
rect 12032 36740 12449 36768
rect 12032 36728 12038 36740
rect 12437 36737 12449 36740
rect 12483 36737 12495 36771
rect 12437 36731 12495 36737
rect 12618 36728 12624 36780
rect 12676 36728 12682 36780
rect 16868 36768 16896 36864
rect 17221 36771 17279 36777
rect 17221 36768 17233 36771
rect 16868 36740 17233 36768
rect 17221 36737 17233 36740
rect 17267 36737 17279 36771
rect 17221 36731 17279 36737
rect 17402 36728 17408 36780
rect 17460 36768 17466 36780
rect 17589 36771 17647 36777
rect 17589 36768 17601 36771
rect 17460 36740 17601 36768
rect 17460 36728 17466 36740
rect 17589 36737 17601 36740
rect 17635 36737 17647 36771
rect 17589 36731 17647 36737
rect 17678 36728 17684 36780
rect 17736 36728 17742 36780
rect 17957 36771 18015 36777
rect 17957 36737 17969 36771
rect 18003 36737 18015 36771
rect 17957 36731 18015 36737
rect 11330 36660 11336 36712
rect 11388 36660 11394 36712
rect 12066 36660 12072 36712
rect 12124 36660 12130 36712
rect 12894 36660 12900 36712
rect 12952 36700 12958 36712
rect 14734 36700 14740 36712
rect 12952 36672 14740 36700
rect 12952 36660 12958 36672
rect 14734 36660 14740 36672
rect 14792 36660 14798 36712
rect 15013 36703 15071 36709
rect 15013 36669 15025 36703
rect 15059 36700 15071 36703
rect 15746 36700 15752 36712
rect 15059 36672 15752 36700
rect 15059 36669 15071 36672
rect 15013 36663 15071 36669
rect 15746 36660 15752 36672
rect 15804 36660 15810 36712
rect 16298 36660 16304 36712
rect 16356 36700 16362 36712
rect 16356 36672 16896 36700
rect 16356 36660 16362 36672
rect 11606 36592 11612 36644
rect 11664 36632 11670 36644
rect 12912 36632 12940 36660
rect 11664 36604 12940 36632
rect 11664 36592 11670 36604
rect 16206 36592 16212 36644
rect 16264 36632 16270 36644
rect 16868 36632 16896 36672
rect 17862 36660 17868 36712
rect 17920 36660 17926 36712
rect 17972 36632 18000 36731
rect 18064 36700 18092 36876
rect 18432 36876 19248 36904
rect 18432 36845 18460 36876
rect 19242 36864 19248 36876
rect 19300 36864 19306 36916
rect 19886 36864 19892 36916
rect 19944 36864 19950 36916
rect 22465 36907 22523 36913
rect 22465 36873 22477 36907
rect 22511 36904 22523 36907
rect 22738 36904 22744 36916
rect 22511 36876 22744 36904
rect 22511 36873 22523 36876
rect 22465 36867 22523 36873
rect 22738 36864 22744 36876
rect 22796 36864 22802 36916
rect 22833 36907 22891 36913
rect 22833 36873 22845 36907
rect 22879 36904 22891 36907
rect 23566 36904 23572 36916
rect 22879 36876 23572 36904
rect 22879 36873 22891 36876
rect 22833 36867 22891 36873
rect 23566 36864 23572 36876
rect 23624 36864 23630 36916
rect 24857 36907 24915 36913
rect 24857 36873 24869 36907
rect 24903 36904 24915 36907
rect 25038 36904 25044 36916
rect 24903 36876 25044 36904
rect 24903 36873 24915 36876
rect 24857 36867 24915 36873
rect 25038 36864 25044 36876
rect 25096 36864 25102 36916
rect 26510 36864 26516 36916
rect 26568 36904 26574 36916
rect 26973 36907 27031 36913
rect 26973 36904 26985 36907
rect 26568 36876 26985 36904
rect 26568 36864 26574 36876
rect 26973 36873 26985 36876
rect 27019 36873 27031 36907
rect 26973 36867 27031 36873
rect 27890 36864 27896 36916
rect 27948 36864 27954 36916
rect 31294 36904 31300 36916
rect 30208 36876 31300 36904
rect 18417 36839 18475 36845
rect 18417 36805 18429 36839
rect 18463 36805 18475 36839
rect 21542 36836 21548 36848
rect 19642 36822 21548 36836
rect 18417 36799 18475 36805
rect 19628 36808 21548 36822
rect 18138 36728 18144 36780
rect 18196 36728 18202 36780
rect 19628 36700 19656 36808
rect 21542 36796 21548 36808
rect 21600 36796 21606 36848
rect 22646 36796 22652 36848
rect 22704 36836 22710 36848
rect 23198 36836 23204 36848
rect 22704 36808 23204 36836
rect 22704 36796 22710 36808
rect 23198 36796 23204 36808
rect 23256 36836 23262 36848
rect 24029 36839 24087 36845
rect 24029 36836 24041 36839
rect 23256 36808 24041 36836
rect 23256 36796 23262 36808
rect 24029 36805 24041 36808
rect 24075 36836 24087 36839
rect 24394 36836 24400 36848
rect 24075 36808 24400 36836
rect 24075 36805 24087 36808
rect 24029 36799 24087 36805
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 25317 36839 25375 36845
rect 25317 36805 25329 36839
rect 25363 36836 25375 36839
rect 26050 36836 26056 36848
rect 25363 36808 26056 36836
rect 25363 36805 25375 36808
rect 25317 36799 25375 36805
rect 26050 36796 26056 36808
rect 26108 36796 26114 36848
rect 27341 36839 27399 36845
rect 27341 36805 27353 36839
rect 27387 36836 27399 36839
rect 28074 36836 28080 36848
rect 27387 36808 28080 36836
rect 27387 36805 27399 36808
rect 27341 36799 27399 36805
rect 28074 36796 28080 36808
rect 28132 36796 28138 36848
rect 21910 36728 21916 36780
rect 21968 36728 21974 36780
rect 22097 36771 22155 36777
rect 22097 36737 22109 36771
rect 22143 36768 22155 36771
rect 22462 36768 22468 36780
rect 22143 36740 22468 36768
rect 22143 36737 22155 36740
rect 22097 36731 22155 36737
rect 22462 36728 22468 36740
rect 22520 36768 22526 36780
rect 23293 36771 23351 36777
rect 22520 36740 23152 36768
rect 22520 36728 22526 36740
rect 23124 36712 23152 36740
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 24486 36768 24492 36780
rect 23339 36740 24492 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 24486 36728 24492 36740
rect 24544 36728 24550 36780
rect 25225 36771 25283 36777
rect 25225 36737 25237 36771
rect 25271 36768 25283 36771
rect 25777 36771 25835 36777
rect 25777 36768 25789 36771
rect 25271 36740 25789 36768
rect 25271 36737 25283 36740
rect 25225 36731 25283 36737
rect 25777 36737 25789 36740
rect 25823 36737 25835 36771
rect 25777 36731 25835 36737
rect 26326 36728 26332 36780
rect 26384 36728 26390 36780
rect 27433 36771 27491 36777
rect 27433 36737 27445 36771
rect 27479 36768 27491 36771
rect 27614 36768 27620 36780
rect 27479 36740 27620 36768
rect 27479 36737 27491 36740
rect 27433 36731 27491 36737
rect 27614 36728 27620 36740
rect 27672 36728 27678 36780
rect 27706 36728 27712 36780
rect 27764 36768 27770 36780
rect 27801 36771 27859 36777
rect 27801 36768 27813 36771
rect 27764 36740 27813 36768
rect 27764 36728 27770 36740
rect 27801 36737 27813 36740
rect 27847 36737 27859 36771
rect 27801 36731 27859 36737
rect 27985 36771 28043 36777
rect 27985 36737 27997 36771
rect 28031 36768 28043 36771
rect 28902 36768 28908 36780
rect 28031 36740 28908 36768
rect 28031 36737 28043 36740
rect 27985 36731 28043 36737
rect 28902 36728 28908 36740
rect 28960 36728 28966 36780
rect 29178 36728 29184 36780
rect 29236 36768 29242 36780
rect 30208 36777 30236 36876
rect 31294 36864 31300 36876
rect 31352 36864 31358 36916
rect 31386 36864 31392 36916
rect 31444 36904 31450 36916
rect 31444 36876 31800 36904
rect 31444 36864 31450 36876
rect 30466 36796 30472 36848
rect 30524 36796 30530 36848
rect 31772 36836 31800 36876
rect 31938 36864 31944 36916
rect 31996 36864 32002 36916
rect 32048 36876 34744 36904
rect 32048 36836 32076 36876
rect 31772 36808 32076 36836
rect 32306 36796 32312 36848
rect 32364 36836 32370 36848
rect 32490 36836 32496 36848
rect 32364 36808 32496 36836
rect 32364 36796 32370 36808
rect 32490 36796 32496 36808
rect 32548 36836 32554 36848
rect 34716 36845 34744 36876
rect 36906 36864 36912 36916
rect 36964 36864 36970 36916
rect 37642 36864 37648 36916
rect 37700 36904 37706 36916
rect 38013 36907 38071 36913
rect 38013 36904 38025 36907
rect 37700 36876 38025 36904
rect 37700 36864 37706 36876
rect 38013 36873 38025 36876
rect 38059 36873 38071 36907
rect 38013 36867 38071 36873
rect 38470 36864 38476 36916
rect 38528 36904 38534 36916
rect 38939 36907 38997 36913
rect 38939 36904 38951 36907
rect 38528 36876 38951 36904
rect 38528 36864 38534 36876
rect 38939 36873 38951 36876
rect 38985 36873 38997 36907
rect 38939 36867 38997 36873
rect 39942 36864 39948 36916
rect 40000 36904 40006 36916
rect 40129 36907 40187 36913
rect 40129 36904 40141 36907
rect 40000 36876 40141 36904
rect 40000 36864 40006 36876
rect 40129 36873 40141 36876
rect 40175 36873 40187 36907
rect 40129 36867 40187 36873
rect 40770 36864 40776 36916
rect 40828 36904 40834 36916
rect 41322 36904 41328 36916
rect 40828 36876 41328 36904
rect 40828 36864 40834 36876
rect 41322 36864 41328 36876
rect 41380 36904 41386 36916
rect 41380 36876 41828 36904
rect 41380 36864 41386 36876
rect 32861 36839 32919 36845
rect 32861 36836 32873 36839
rect 32548 36808 32873 36836
rect 32548 36796 32554 36808
rect 32861 36805 32873 36808
rect 32907 36805 32919 36839
rect 32861 36799 32919 36805
rect 33781 36839 33839 36845
rect 33781 36805 33793 36839
rect 33827 36805 33839 36839
rect 33781 36799 33839 36805
rect 33997 36839 34055 36845
rect 33997 36805 34009 36839
rect 34043 36836 34055 36839
rect 34701 36839 34759 36845
rect 34043 36808 34652 36836
rect 34043 36805 34055 36808
rect 33997 36799 34055 36805
rect 29641 36771 29699 36777
rect 29641 36768 29653 36771
rect 29236 36740 29653 36768
rect 29236 36728 29242 36740
rect 29641 36737 29653 36740
rect 29687 36737 29699 36771
rect 29641 36731 29699 36737
rect 30193 36771 30251 36777
rect 30193 36737 30205 36771
rect 30239 36737 30251 36771
rect 30193 36731 30251 36737
rect 31570 36728 31576 36780
rect 31628 36728 31634 36780
rect 32585 36771 32643 36777
rect 32585 36737 32597 36771
rect 32631 36737 32643 36771
rect 32585 36731 32643 36737
rect 18064 36672 19656 36700
rect 19536 36644 19564 36672
rect 20070 36660 20076 36712
rect 20128 36700 20134 36712
rect 20533 36703 20591 36709
rect 20533 36700 20545 36703
rect 20128 36672 20545 36700
rect 20128 36660 20134 36672
rect 20533 36669 20545 36672
rect 20579 36669 20591 36703
rect 20533 36663 20591 36669
rect 22925 36703 22983 36709
rect 22925 36669 22937 36703
rect 22971 36669 22983 36703
rect 22925 36663 22983 36669
rect 18046 36632 18052 36644
rect 16264 36604 16804 36632
rect 16868 36604 18052 36632
rect 16264 36592 16270 36604
rect 10689 36567 10747 36573
rect 10689 36564 10701 36567
rect 10560 36536 10701 36564
rect 10560 36524 10566 36536
rect 10689 36533 10701 36536
rect 10735 36533 10747 36567
rect 10689 36527 10747 36533
rect 11054 36524 11060 36576
rect 11112 36564 11118 36576
rect 11517 36567 11575 36573
rect 11517 36564 11529 36567
rect 11112 36536 11529 36564
rect 11112 36524 11118 36536
rect 11517 36533 11529 36536
rect 11563 36533 11575 36567
rect 11517 36527 11575 36533
rect 12250 36524 12256 36576
rect 12308 36524 12314 36576
rect 16666 36524 16672 36576
rect 16724 36524 16730 36576
rect 16776 36564 16804 36604
rect 18046 36592 18052 36604
rect 18104 36592 18110 36644
rect 19518 36592 19524 36644
rect 19576 36592 19582 36644
rect 22940 36632 22968 36663
rect 23106 36660 23112 36712
rect 23164 36700 23170 36712
rect 25501 36703 25559 36709
rect 25501 36700 25513 36703
rect 23164 36672 25513 36700
rect 23164 36660 23170 36672
rect 25501 36669 25513 36672
rect 25547 36700 25559 36703
rect 25590 36700 25596 36712
rect 25547 36672 25596 36700
rect 25547 36669 25559 36672
rect 25501 36663 25559 36669
rect 25590 36660 25596 36672
rect 25648 36660 25654 36712
rect 27338 36660 27344 36712
rect 27396 36700 27402 36712
rect 27525 36703 27583 36709
rect 27525 36700 27537 36703
rect 27396 36672 27537 36700
rect 27396 36660 27402 36672
rect 27525 36669 27537 36672
rect 27571 36669 27583 36703
rect 27525 36663 27583 36669
rect 29730 36660 29736 36712
rect 29788 36700 29794 36712
rect 31588 36700 31616 36728
rect 32600 36700 32628 36731
rect 33137 36703 33195 36709
rect 33137 36700 33149 36703
rect 29788 36672 31616 36700
rect 31726 36672 33149 36700
rect 29788 36660 29794 36672
rect 23474 36632 23480 36644
rect 22940 36604 23480 36632
rect 23474 36592 23480 36604
rect 23532 36592 23538 36644
rect 25774 36592 25780 36644
rect 25832 36632 25838 36644
rect 31726 36632 31754 36672
rect 33137 36669 33149 36672
rect 33183 36669 33195 36703
rect 33796 36700 33824 36799
rect 34256 36777 34284 36808
rect 34241 36771 34299 36777
rect 34241 36737 34253 36771
rect 34287 36737 34299 36771
rect 34241 36731 34299 36737
rect 34330 36728 34336 36780
rect 34388 36728 34394 36780
rect 34422 36728 34428 36780
rect 34480 36768 34486 36780
rect 34517 36771 34575 36777
rect 34517 36768 34529 36771
rect 34480 36740 34529 36768
rect 34480 36728 34486 36740
rect 34517 36737 34529 36740
rect 34563 36737 34575 36771
rect 34624 36768 34652 36808
rect 34701 36805 34713 36839
rect 34747 36805 34759 36839
rect 34701 36799 34759 36805
rect 35989 36839 36047 36845
rect 35989 36805 36001 36839
rect 36035 36836 36047 36839
rect 36633 36839 36691 36845
rect 36633 36836 36645 36839
rect 36035 36808 36645 36836
rect 36035 36805 36047 36808
rect 35989 36799 36047 36805
rect 36633 36805 36645 36808
rect 36679 36836 36691 36839
rect 37001 36839 37059 36845
rect 37001 36836 37013 36839
rect 36679 36808 37013 36836
rect 36679 36805 36691 36808
rect 36633 36799 36691 36805
rect 37001 36805 37013 36808
rect 37047 36805 37059 36839
rect 37001 36799 37059 36805
rect 38105 36839 38163 36845
rect 38105 36805 38117 36839
rect 38151 36836 38163 36839
rect 38381 36839 38439 36845
rect 38381 36836 38393 36839
rect 38151 36808 38393 36836
rect 38151 36805 38163 36808
rect 38105 36799 38163 36805
rect 38381 36805 38393 36808
rect 38427 36836 38439 36839
rect 39025 36839 39083 36845
rect 39025 36836 39037 36839
rect 38427 36808 39037 36836
rect 38427 36805 38439 36808
rect 38381 36799 38439 36805
rect 39025 36805 39037 36808
rect 39071 36805 39083 36839
rect 39025 36799 39083 36805
rect 35710 36768 35716 36780
rect 34624 36740 35716 36768
rect 34517 36731 34575 36737
rect 35710 36728 35716 36740
rect 35768 36728 35774 36780
rect 36173 36771 36231 36777
rect 36173 36737 36185 36771
rect 36219 36768 36231 36771
rect 36262 36768 36268 36780
rect 36219 36740 36268 36768
rect 36219 36737 36231 36740
rect 36173 36731 36231 36737
rect 36262 36728 36268 36740
rect 36320 36728 36326 36780
rect 36357 36771 36415 36777
rect 36357 36737 36369 36771
rect 36403 36737 36415 36771
rect 36357 36731 36415 36737
rect 36449 36771 36507 36777
rect 36449 36737 36461 36771
rect 36495 36768 36507 36771
rect 36538 36768 36544 36780
rect 36495 36740 36544 36768
rect 36495 36737 36507 36740
rect 36449 36731 36507 36737
rect 34440 36700 34468 36728
rect 33796 36672 34468 36700
rect 36372 36700 36400 36731
rect 36538 36728 36544 36740
rect 36596 36728 36602 36780
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36768 36783 36771
rect 36814 36768 36820 36780
rect 36771 36740 36820 36768
rect 36771 36737 36783 36740
rect 36725 36731 36783 36737
rect 36814 36728 36820 36740
rect 36872 36728 36878 36780
rect 37093 36771 37151 36777
rect 37093 36737 37105 36771
rect 37139 36737 37151 36771
rect 37093 36731 37151 36737
rect 38013 36771 38071 36777
rect 38013 36737 38025 36771
rect 38059 36768 38071 36771
rect 38194 36768 38200 36780
rect 38059 36740 38200 36768
rect 38059 36737 38071 36740
rect 38013 36731 38071 36737
rect 36906 36700 36912 36712
rect 36372 36672 36912 36700
rect 33137 36663 33195 36669
rect 36906 36660 36912 36672
rect 36964 36660 36970 36712
rect 36998 36660 37004 36712
rect 37056 36700 37062 36712
rect 37108 36700 37136 36731
rect 38194 36728 38200 36740
rect 38252 36728 38258 36780
rect 38286 36728 38292 36780
rect 38344 36728 38350 36780
rect 38565 36771 38623 36777
rect 38565 36737 38577 36771
rect 38611 36737 38623 36771
rect 38565 36731 38623 36737
rect 38749 36771 38807 36777
rect 38749 36737 38761 36771
rect 38795 36737 38807 36771
rect 38749 36731 38807 36737
rect 38841 36771 38899 36777
rect 38841 36737 38853 36771
rect 38887 36768 38899 36771
rect 38930 36768 38936 36780
rect 38887 36740 38936 36768
rect 38887 36737 38899 36740
rect 38841 36731 38899 36737
rect 38580 36700 38608 36731
rect 37056 36672 37136 36700
rect 38120 36672 38608 36700
rect 38764 36700 38792 36731
rect 38930 36728 38936 36740
rect 38988 36728 38994 36780
rect 39114 36728 39120 36780
rect 39172 36728 39178 36780
rect 39485 36771 39543 36777
rect 39485 36737 39497 36771
rect 39531 36768 39543 36771
rect 39960 36768 39988 36864
rect 41800 36836 41828 36876
rect 41800 36808 41920 36836
rect 39531 36740 39988 36768
rect 39531 36737 39543 36740
rect 39485 36731 39543 36737
rect 40494 36728 40500 36780
rect 40552 36728 40558 36780
rect 41892 36777 41920 36808
rect 41877 36771 41935 36777
rect 41877 36737 41889 36771
rect 41923 36737 41935 36771
rect 41877 36731 41935 36737
rect 39206 36700 39212 36712
rect 38764 36672 39212 36700
rect 37056 36660 37062 36672
rect 25832 36604 29224 36632
rect 25832 36592 25838 36604
rect 19150 36564 19156 36576
rect 16776 36536 19156 36564
rect 19150 36524 19156 36536
rect 19208 36564 19214 36576
rect 19610 36564 19616 36576
rect 19208 36536 19616 36564
rect 19208 36524 19214 36536
rect 19610 36524 19616 36536
rect 19668 36524 19674 36576
rect 19978 36524 19984 36576
rect 20036 36524 20042 36576
rect 29086 36524 29092 36576
rect 29144 36524 29150 36576
rect 29196 36564 29224 36604
rect 31496 36604 31754 36632
rect 31496 36564 31524 36604
rect 34146 36592 34152 36644
rect 34204 36592 34210 36644
rect 34514 36592 34520 36644
rect 34572 36592 34578 36644
rect 35986 36592 35992 36644
rect 36044 36632 36050 36644
rect 36449 36635 36507 36641
rect 36449 36632 36461 36635
rect 36044 36604 36461 36632
rect 36044 36592 36050 36604
rect 36449 36601 36461 36604
rect 36495 36601 36507 36635
rect 36449 36595 36507 36601
rect 36538 36592 36544 36644
rect 36596 36632 36602 36644
rect 37016 36632 37044 36660
rect 36596 36604 37044 36632
rect 36596 36592 36602 36604
rect 29196 36536 31524 36564
rect 31570 36524 31576 36576
rect 31628 36564 31634 36576
rect 32309 36567 32367 36573
rect 32309 36564 32321 36567
rect 31628 36536 32321 36564
rect 31628 36524 31634 36536
rect 32309 36533 32321 36536
rect 32355 36533 32367 36567
rect 32309 36527 32367 36533
rect 33965 36567 34023 36573
rect 33965 36533 33977 36567
rect 34011 36564 34023 36567
rect 34330 36564 34336 36576
rect 34011 36536 34336 36564
rect 34011 36533 34023 36536
rect 33965 36527 34023 36533
rect 34330 36524 34336 36536
rect 34388 36524 34394 36576
rect 34793 36567 34851 36573
rect 34793 36533 34805 36567
rect 34839 36564 34851 36567
rect 35618 36564 35624 36576
rect 34839 36536 35624 36564
rect 34839 36533 34851 36536
rect 34793 36527 34851 36533
rect 35618 36524 35624 36536
rect 35676 36564 35682 36576
rect 38120 36564 38148 36672
rect 38580 36632 38608 36672
rect 39206 36660 39212 36672
rect 39264 36660 39270 36712
rect 40512 36700 40540 36728
rect 41506 36700 41512 36712
rect 39960 36672 41512 36700
rect 39390 36632 39396 36644
rect 38580 36604 39396 36632
rect 39390 36592 39396 36604
rect 39448 36632 39454 36644
rect 39850 36632 39856 36644
rect 39448 36604 39856 36632
rect 39448 36592 39454 36604
rect 39850 36592 39856 36604
rect 39908 36592 39914 36644
rect 35676 36536 38148 36564
rect 35676 36524 35682 36536
rect 38194 36524 38200 36576
rect 38252 36564 38258 36576
rect 38930 36564 38936 36576
rect 38252 36536 38936 36564
rect 38252 36524 38258 36536
rect 38930 36524 38936 36536
rect 38988 36524 38994 36576
rect 39022 36524 39028 36576
rect 39080 36564 39086 36576
rect 39960 36564 39988 36672
rect 41506 36660 41512 36672
rect 41564 36660 41570 36712
rect 41598 36660 41604 36712
rect 41656 36660 41662 36712
rect 39080 36536 39988 36564
rect 39080 36524 39086 36536
rect 40034 36524 40040 36576
rect 40092 36524 40098 36576
rect 1104 36474 42504 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 42504 36474
rect 1104 36400 42504 36422
rect 4982 36320 4988 36372
rect 5040 36360 5046 36372
rect 5442 36360 5448 36372
rect 5040 36332 5448 36360
rect 5040 36320 5046 36332
rect 5442 36320 5448 36332
rect 5500 36320 5506 36372
rect 6917 36363 6975 36369
rect 6917 36329 6929 36363
rect 6963 36360 6975 36363
rect 7190 36360 7196 36372
rect 6963 36332 7196 36360
rect 6963 36329 6975 36332
rect 6917 36323 6975 36329
rect 7190 36320 7196 36332
rect 7248 36320 7254 36372
rect 11330 36320 11336 36372
rect 11388 36320 11394 36372
rect 13170 36320 13176 36372
rect 13228 36360 13234 36372
rect 14093 36363 14151 36369
rect 14093 36360 14105 36363
rect 13228 36332 14105 36360
rect 13228 36320 13234 36332
rect 14093 36329 14105 36332
rect 14139 36329 14151 36363
rect 14093 36323 14151 36329
rect 15746 36320 15752 36372
rect 15804 36320 15810 36372
rect 21910 36360 21916 36372
rect 16040 36332 16344 36360
rect 3068 36264 3924 36292
rect 2866 36116 2872 36168
rect 2924 36116 2930 36168
rect 2958 36116 2964 36168
rect 3016 36116 3022 36168
rect 3068 36165 3096 36264
rect 3421 36227 3479 36233
rect 3421 36193 3433 36227
rect 3467 36224 3479 36227
rect 3786 36224 3792 36236
rect 3467 36196 3792 36224
rect 3467 36193 3479 36196
rect 3421 36187 3479 36193
rect 3786 36184 3792 36196
rect 3844 36184 3850 36236
rect 3896 36224 3924 36264
rect 3970 36252 3976 36304
rect 4028 36292 4034 36304
rect 4065 36295 4123 36301
rect 4065 36292 4077 36295
rect 4028 36264 4077 36292
rect 4028 36252 4034 36264
rect 4065 36261 4077 36264
rect 4111 36261 4123 36295
rect 4065 36255 4123 36261
rect 6546 36252 6552 36304
rect 6604 36292 6610 36304
rect 7006 36292 7012 36304
rect 6604 36264 7012 36292
rect 6604 36252 6610 36264
rect 7006 36252 7012 36264
rect 7064 36292 7070 36304
rect 8018 36292 8024 36304
rect 7064 36264 8024 36292
rect 7064 36252 7070 36264
rect 8018 36252 8024 36264
rect 8076 36292 8082 36304
rect 8076 36264 8248 36292
rect 8076 36252 8082 36264
rect 6086 36224 6092 36236
rect 3896 36196 6092 36224
rect 6086 36184 6092 36196
rect 6144 36184 6150 36236
rect 7374 36224 7380 36236
rect 7300 36196 7380 36224
rect 3053 36159 3111 36165
rect 3053 36125 3065 36159
rect 3099 36125 3111 36159
rect 3053 36119 3111 36125
rect 3878 36116 3884 36168
rect 3936 36116 3942 36168
rect 3973 36159 4031 36165
rect 3973 36125 3985 36159
rect 4019 36156 4031 36159
rect 4062 36156 4068 36168
rect 4019 36128 4068 36156
rect 4019 36125 4031 36128
rect 3973 36119 4031 36125
rect 4062 36116 4068 36128
rect 4120 36116 4126 36168
rect 4157 36159 4215 36165
rect 4157 36125 4169 36159
rect 4203 36156 4215 36159
rect 5166 36156 5172 36168
rect 4203 36128 5172 36156
rect 4203 36125 4215 36128
rect 4157 36119 4215 36125
rect 5166 36116 5172 36128
rect 5224 36116 5230 36168
rect 7098 36116 7104 36168
rect 7156 36116 7162 36168
rect 7300 36165 7328 36196
rect 7374 36184 7380 36196
rect 7432 36184 7438 36236
rect 7561 36227 7619 36233
rect 7561 36193 7573 36227
rect 7607 36224 7619 36227
rect 8110 36224 8116 36236
rect 7607 36196 8116 36224
rect 7607 36193 7619 36196
rect 7561 36187 7619 36193
rect 7852 36165 7880 36196
rect 8110 36184 8116 36196
rect 8168 36184 8174 36236
rect 7285 36159 7343 36165
rect 7285 36125 7297 36159
rect 7331 36125 7343 36159
rect 7285 36119 7343 36125
rect 7837 36159 7895 36165
rect 7837 36125 7849 36159
rect 7883 36156 7895 36159
rect 8021 36159 8079 36165
rect 7883 36128 7917 36156
rect 7883 36125 7895 36128
rect 7837 36119 7895 36125
rect 8021 36125 8033 36159
rect 8067 36156 8079 36159
rect 8220 36156 8248 36264
rect 12342 36252 12348 36304
rect 12400 36292 12406 36304
rect 16040 36292 16068 36332
rect 12400 36264 16068 36292
rect 16316 36292 16344 36332
rect 18800 36332 21916 36360
rect 18800 36292 18828 36332
rect 21910 36320 21916 36332
rect 21968 36360 21974 36372
rect 21968 36332 26464 36360
rect 21968 36320 21974 36332
rect 25130 36292 25136 36304
rect 16316 36264 18828 36292
rect 23584 36264 25136 36292
rect 12400 36252 12406 36264
rect 9858 36184 9864 36236
rect 9916 36184 9922 36236
rect 10502 36184 10508 36236
rect 10560 36224 10566 36236
rect 10560 36196 12112 36224
rect 10560 36184 10566 36196
rect 8067 36128 8248 36156
rect 8067 36125 8079 36128
rect 8021 36119 8079 36125
rect 9582 36116 9588 36168
rect 9640 36116 9646 36168
rect 12084 36165 12112 36196
rect 12250 36184 12256 36236
rect 12308 36184 12314 36236
rect 14550 36184 14556 36236
rect 14608 36184 14614 36236
rect 14645 36227 14703 36233
rect 14645 36193 14657 36227
rect 14691 36193 14703 36227
rect 16298 36224 16304 36236
rect 14645 36187 14703 36193
rect 16040 36196 16304 36224
rect 12069 36159 12127 36165
rect 12069 36125 12081 36159
rect 12115 36125 12127 36159
rect 12069 36119 12127 36125
rect 12161 36159 12219 36165
rect 12161 36125 12173 36159
rect 12207 36156 12219 36159
rect 12805 36159 12863 36165
rect 12805 36156 12817 36159
rect 12207 36128 12817 36156
rect 12207 36125 12219 36128
rect 12161 36119 12219 36125
rect 12805 36125 12817 36128
rect 12851 36156 12863 36159
rect 13262 36156 13268 36168
rect 12851 36128 13268 36156
rect 12851 36125 12863 36128
rect 12805 36119 12863 36125
rect 13262 36116 13268 36128
rect 13320 36116 13326 36168
rect 13814 36116 13820 36168
rect 13872 36116 13878 36168
rect 14274 36116 14280 36168
rect 14332 36156 14338 36168
rect 14660 36156 14688 36187
rect 16040 36156 16068 36196
rect 16298 36184 16304 36196
rect 16356 36184 16362 36236
rect 16393 36227 16451 36233
rect 16393 36193 16405 36227
rect 16439 36224 16451 36227
rect 16439 36196 16804 36224
rect 16439 36193 16451 36196
rect 16393 36187 16451 36193
rect 14332 36128 14688 36156
rect 15488 36128 16068 36156
rect 16117 36159 16175 36165
rect 14332 36116 14338 36128
rect 2884 36088 2912 36116
rect 3145 36091 3203 36097
rect 3145 36088 3157 36091
rect 2884 36060 3157 36088
rect 3145 36057 3157 36060
rect 3191 36057 3203 36091
rect 3145 36051 3203 36057
rect 3283 36091 3341 36097
rect 3283 36057 3295 36091
rect 3329 36088 3341 36091
rect 3510 36088 3516 36100
rect 3329 36060 3516 36088
rect 3329 36057 3341 36060
rect 3283 36051 3341 36057
rect 2777 36023 2835 36029
rect 2777 35989 2789 36023
rect 2823 36020 2835 36023
rect 2866 36020 2872 36032
rect 2823 35992 2872 36020
rect 2823 35989 2835 35992
rect 2777 35983 2835 35989
rect 2866 35980 2872 35992
rect 2924 35980 2930 36032
rect 3160 36020 3188 36051
rect 3510 36048 3516 36060
rect 3568 36048 3574 36100
rect 3694 36048 3700 36100
rect 3752 36088 3758 36100
rect 6362 36088 6368 36100
rect 3752 36060 6368 36088
rect 3752 36048 3758 36060
rect 6362 36048 6368 36060
rect 6420 36048 6426 36100
rect 7193 36091 7251 36097
rect 7193 36057 7205 36091
rect 7239 36057 7251 36091
rect 7193 36051 7251 36057
rect 7423 36091 7481 36097
rect 7423 36057 7435 36091
rect 7469 36088 7481 36091
rect 7558 36088 7564 36100
rect 7469 36060 7564 36088
rect 7469 36057 7481 36060
rect 7423 36051 7481 36057
rect 4062 36020 4068 36032
rect 3160 35992 4068 36020
rect 4062 35980 4068 35992
rect 4120 35980 4126 36032
rect 4341 36023 4399 36029
rect 4341 35989 4353 36023
rect 4387 36020 4399 36023
rect 5350 36020 5356 36032
rect 4387 35992 5356 36020
rect 4387 35989 4399 35992
rect 4341 35983 4399 35989
rect 5350 35980 5356 35992
rect 5408 35980 5414 36032
rect 7208 36020 7236 36051
rect 7558 36048 7564 36060
rect 7616 36048 7622 36100
rect 9766 36048 9772 36100
rect 9824 36088 9830 36100
rect 9824 36060 10350 36088
rect 9824 36048 9830 36060
rect 12618 36048 12624 36100
rect 12676 36088 12682 36100
rect 15488 36088 15516 36128
rect 16117 36125 16129 36159
rect 16163 36156 16175 36159
rect 16666 36156 16672 36168
rect 16163 36128 16672 36156
rect 16163 36125 16175 36128
rect 16117 36119 16175 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 16776 36156 16804 36196
rect 16850 36184 16856 36236
rect 16908 36224 16914 36236
rect 17129 36227 17187 36233
rect 17129 36224 17141 36227
rect 16908 36196 17141 36224
rect 16908 36184 16914 36196
rect 17129 36193 17141 36196
rect 17175 36193 17187 36227
rect 17494 36224 17500 36236
rect 17129 36187 17187 36193
rect 17236 36196 17500 36224
rect 17236 36156 17264 36196
rect 17494 36184 17500 36196
rect 17552 36224 17558 36236
rect 19702 36224 19708 36236
rect 17552 36196 19708 36224
rect 17552 36184 17558 36196
rect 19702 36184 19708 36196
rect 19760 36224 19766 36236
rect 19797 36227 19855 36233
rect 19797 36224 19809 36227
rect 19760 36196 19809 36224
rect 19760 36184 19766 36196
rect 19797 36193 19809 36196
rect 19843 36193 19855 36227
rect 19797 36187 19855 36193
rect 19886 36184 19892 36236
rect 19944 36224 19950 36236
rect 20349 36227 20407 36233
rect 20349 36224 20361 36227
rect 19944 36196 20361 36224
rect 19944 36184 19950 36196
rect 20349 36193 20361 36196
rect 20395 36193 20407 36227
rect 20349 36187 20407 36193
rect 22186 36184 22192 36236
rect 22244 36184 22250 36236
rect 16776 36128 17264 36156
rect 19613 36159 19671 36165
rect 19613 36125 19625 36159
rect 19659 36156 19671 36159
rect 19978 36156 19984 36168
rect 19659 36128 19984 36156
rect 19659 36125 19671 36128
rect 19613 36119 19671 36125
rect 19978 36116 19984 36128
rect 20036 36116 20042 36168
rect 23584 36142 23612 36264
rect 25130 36252 25136 36264
rect 25188 36252 25194 36304
rect 23934 36184 23940 36236
rect 23992 36224 23998 36236
rect 25685 36227 25743 36233
rect 25685 36224 25697 36227
rect 23992 36196 25697 36224
rect 23992 36184 23998 36196
rect 25685 36193 25697 36196
rect 25731 36193 25743 36227
rect 25685 36187 25743 36193
rect 26436 36224 26464 36332
rect 29178 36320 29184 36372
rect 29236 36360 29242 36372
rect 29365 36363 29423 36369
rect 29365 36360 29377 36363
rect 29236 36332 29377 36360
rect 29236 36320 29242 36332
rect 29365 36329 29377 36332
rect 29411 36329 29423 36363
rect 29365 36323 29423 36329
rect 29546 36320 29552 36372
rect 29604 36320 29610 36372
rect 34330 36320 34336 36372
rect 34388 36360 34394 36372
rect 35437 36363 35495 36369
rect 35437 36360 35449 36363
rect 34388 36332 35449 36360
rect 34388 36320 34394 36332
rect 35437 36329 35449 36332
rect 35483 36329 35495 36363
rect 35437 36323 35495 36329
rect 35866 36332 36400 36360
rect 26697 36295 26755 36301
rect 26697 36261 26709 36295
rect 26743 36292 26755 36295
rect 27338 36292 27344 36304
rect 26743 36264 27344 36292
rect 26743 36261 26755 36264
rect 26697 36255 26755 36261
rect 27338 36252 27344 36264
rect 27396 36252 27402 36304
rect 35866 36292 35894 36332
rect 31220 36264 35894 36292
rect 31220 36224 31248 36264
rect 26436 36196 31248 36224
rect 26436 36165 26464 36196
rect 31294 36184 31300 36236
rect 31352 36184 31358 36236
rect 31478 36184 31484 36236
rect 31536 36224 31542 36236
rect 31849 36227 31907 36233
rect 31849 36224 31861 36227
rect 31536 36196 31861 36224
rect 31536 36184 31542 36196
rect 31849 36193 31861 36196
rect 31895 36193 31907 36227
rect 31849 36187 31907 36193
rect 31938 36184 31944 36236
rect 31996 36224 32002 36236
rect 33505 36227 33563 36233
rect 33505 36224 33517 36227
rect 31996 36196 33517 36224
rect 31996 36184 32002 36196
rect 33505 36193 33517 36196
rect 33551 36224 33563 36227
rect 34333 36227 34391 36233
rect 34333 36224 34345 36227
rect 33551 36196 34345 36224
rect 33551 36193 33563 36196
rect 33505 36187 33563 36193
rect 34333 36193 34345 36196
rect 34379 36193 34391 36227
rect 34333 36187 34391 36193
rect 35710 36184 35716 36236
rect 35768 36224 35774 36236
rect 35989 36227 36047 36233
rect 35989 36224 36001 36227
rect 35768 36196 36001 36224
rect 35768 36184 35774 36196
rect 35989 36193 36001 36196
rect 36035 36193 36047 36227
rect 35989 36187 36047 36193
rect 24949 36159 25007 36165
rect 24949 36125 24961 36159
rect 24995 36125 25007 36159
rect 24949 36119 25007 36125
rect 26421 36159 26479 36165
rect 26421 36125 26433 36159
rect 26467 36125 26479 36159
rect 26421 36119 26479 36125
rect 26973 36159 27031 36165
rect 26973 36125 26985 36159
rect 27019 36125 27031 36159
rect 26973 36119 27031 36125
rect 12676 36060 15516 36088
rect 15565 36091 15623 36097
rect 12676 36048 12682 36060
rect 7653 36023 7711 36029
rect 7653 36020 7665 36023
rect 7208 35992 7665 36020
rect 7653 35989 7665 35992
rect 7699 35989 7711 36023
rect 7653 35983 7711 35989
rect 11698 35980 11704 36032
rect 11756 35980 11762 36032
rect 13078 35980 13084 36032
rect 13136 36020 13142 36032
rect 13740 36029 13768 36060
rect 15565 36057 15577 36091
rect 15611 36088 15623 36091
rect 15654 36088 15660 36100
rect 15611 36060 15660 36088
rect 15611 36057 15623 36060
rect 15565 36051 15623 36057
rect 15654 36048 15660 36060
rect 15712 36048 15718 36100
rect 16850 36088 16856 36100
rect 16132 36060 16856 36088
rect 13357 36023 13415 36029
rect 13357 36020 13369 36023
rect 13136 35992 13369 36020
rect 13136 35980 13142 35992
rect 13357 35989 13369 35992
rect 13403 35989 13415 36023
rect 13357 35983 13415 35989
rect 13725 36023 13783 36029
rect 13725 35989 13737 36023
rect 13771 35989 13783 36023
rect 13725 35983 13783 35989
rect 14458 35980 14464 36032
rect 14516 35980 14522 36032
rect 15286 35980 15292 36032
rect 15344 36020 15350 36032
rect 15473 36023 15531 36029
rect 15473 36020 15485 36023
rect 15344 35992 15485 36020
rect 15344 35980 15350 35992
rect 15473 35989 15485 35992
rect 15519 36020 15531 36023
rect 16132 36020 16160 36060
rect 16850 36048 16856 36060
rect 16908 36048 16914 36100
rect 20625 36091 20683 36097
rect 20625 36057 20637 36091
rect 20671 36088 20683 36091
rect 20898 36088 20904 36100
rect 20671 36060 20904 36088
rect 20671 36057 20683 36060
rect 20625 36051 20683 36057
rect 20898 36048 20904 36060
rect 20956 36048 20962 36100
rect 21634 36048 21640 36100
rect 21692 36048 21698 36100
rect 22462 36048 22468 36100
rect 22520 36048 22526 36100
rect 24964 36088 24992 36119
rect 23768 36060 24992 36088
rect 26988 36088 27016 36119
rect 27430 36116 27436 36168
rect 27488 36156 27494 36168
rect 27617 36159 27675 36165
rect 27617 36156 27629 36159
rect 27488 36128 27629 36156
rect 27488 36116 27494 36128
rect 27617 36125 27629 36128
rect 27663 36125 27675 36159
rect 27617 36119 27675 36125
rect 32766 36116 32772 36168
rect 32824 36116 32830 36168
rect 35253 36159 35311 36165
rect 35253 36125 35265 36159
rect 35299 36125 35311 36159
rect 35253 36119 35311 36125
rect 27062 36088 27068 36100
rect 26988 36060 27068 36088
rect 15519 35992 16160 36020
rect 16209 36023 16267 36029
rect 15519 35989 15531 35992
rect 15473 35983 15531 35989
rect 16209 35989 16221 36023
rect 16255 36020 16267 36023
rect 16577 36023 16635 36029
rect 16577 36020 16589 36023
rect 16255 35992 16589 36020
rect 16255 35989 16267 35992
rect 16209 35983 16267 35989
rect 16577 35989 16589 35992
rect 16623 35989 16635 36023
rect 16577 35983 16635 35989
rect 16942 35980 16948 36032
rect 17000 35980 17006 36032
rect 17034 35980 17040 36032
rect 17092 35980 17098 36032
rect 18230 35980 18236 36032
rect 18288 36020 18294 36032
rect 19245 36023 19303 36029
rect 19245 36020 19257 36023
rect 18288 35992 19257 36020
rect 18288 35980 18294 35992
rect 19245 35989 19257 35992
rect 19291 35989 19303 36023
rect 19245 35983 19303 35989
rect 19702 35980 19708 36032
rect 19760 35980 19766 36032
rect 22097 36023 22155 36029
rect 22097 35989 22109 36023
rect 22143 36020 22155 36023
rect 22554 36020 22560 36032
rect 22143 35992 22560 36020
rect 22143 35989 22155 35992
rect 22097 35983 22155 35989
rect 22554 35980 22560 35992
rect 22612 36020 22618 36032
rect 23768 36020 23796 36060
rect 27062 36048 27068 36060
rect 27120 36088 27126 36100
rect 27120 36060 27752 36088
rect 27120 36048 27126 36060
rect 27724 36032 27752 36060
rect 27890 36048 27896 36100
rect 27948 36048 27954 36100
rect 29270 36088 29276 36100
rect 29118 36060 29276 36088
rect 29270 36048 29276 36060
rect 29328 36088 29334 36100
rect 29730 36088 29736 36100
rect 29328 36060 29736 36088
rect 29328 36048 29334 36060
rect 29730 36048 29736 36060
rect 29788 36088 29794 36100
rect 29788 36060 29854 36088
rect 29788 36048 29794 36060
rect 31018 36048 31024 36100
rect 31076 36048 31082 36100
rect 31757 36091 31815 36097
rect 31757 36057 31769 36091
rect 31803 36088 31815 36091
rect 32217 36091 32275 36097
rect 32217 36088 32229 36091
rect 31803 36060 32229 36088
rect 31803 36057 31815 36060
rect 31757 36051 31815 36057
rect 32217 36057 32229 36060
rect 32263 36057 32275 36091
rect 32217 36051 32275 36057
rect 33321 36091 33379 36097
rect 33321 36057 33333 36091
rect 33367 36088 33379 36091
rect 34054 36088 34060 36100
rect 33367 36060 34060 36088
rect 33367 36057 33379 36060
rect 33321 36051 33379 36057
rect 34054 36048 34060 36060
rect 34112 36048 34118 36100
rect 34149 36091 34207 36097
rect 34149 36057 34161 36091
rect 34195 36088 34207 36091
rect 34701 36091 34759 36097
rect 34701 36088 34713 36091
rect 34195 36060 34713 36088
rect 34195 36057 34207 36060
rect 34149 36051 34207 36057
rect 34701 36057 34713 36060
rect 34747 36057 34759 36091
rect 34701 36051 34759 36057
rect 22612 35992 23796 36020
rect 22612 35980 22618 35992
rect 24026 35980 24032 36032
rect 24084 36020 24090 36032
rect 24397 36023 24455 36029
rect 24397 36020 24409 36023
rect 24084 35992 24409 36020
rect 24084 35980 24090 35992
rect 24397 35989 24409 35992
rect 24443 35989 24455 36023
rect 24397 35983 24455 35989
rect 24578 35980 24584 36032
rect 24636 36020 24642 36032
rect 25133 36023 25191 36029
rect 25133 36020 25145 36023
rect 24636 35992 25145 36020
rect 24636 35980 24642 35992
rect 25133 35989 25145 35992
rect 25179 35989 25191 36023
rect 25133 35983 25191 35989
rect 27522 35980 27528 36032
rect 27580 35980 27586 36032
rect 27706 35980 27712 36032
rect 27764 35980 27770 36032
rect 30742 35980 30748 36032
rect 30800 36020 30806 36032
rect 31389 36023 31447 36029
rect 31389 36020 31401 36023
rect 30800 35992 31401 36020
rect 30800 35980 30806 35992
rect 31389 35989 31401 35992
rect 31435 35989 31447 36023
rect 31389 35983 31447 35989
rect 32674 35980 32680 36032
rect 32732 36020 32738 36032
rect 32953 36023 33011 36029
rect 32953 36020 32965 36023
rect 32732 35992 32965 36020
rect 32732 35980 32738 35992
rect 32953 35989 32965 35992
rect 32999 35989 33011 36023
rect 32953 35983 33011 35989
rect 33410 35980 33416 36032
rect 33468 35980 33474 36032
rect 33778 35980 33784 36032
rect 33836 35980 33842 36032
rect 34238 35980 34244 36032
rect 34296 35980 34302 36032
rect 34422 35980 34428 36032
rect 34480 36020 34486 36032
rect 35268 36020 35296 36119
rect 35434 36116 35440 36168
rect 35492 36156 35498 36168
rect 36372 36165 36400 36332
rect 36814 36320 36820 36372
rect 36872 36320 36878 36372
rect 38286 36320 38292 36372
rect 38344 36360 38350 36372
rect 39114 36360 39120 36372
rect 38344 36332 39120 36360
rect 38344 36320 38350 36332
rect 39114 36320 39120 36332
rect 39172 36360 39178 36372
rect 39301 36363 39359 36369
rect 39301 36360 39313 36363
rect 39172 36332 39313 36360
rect 39172 36320 39178 36332
rect 39301 36329 39313 36332
rect 39347 36329 39359 36363
rect 39301 36323 39359 36329
rect 40773 36363 40831 36369
rect 40773 36329 40785 36363
rect 40819 36360 40831 36363
rect 41598 36360 41604 36372
rect 40819 36332 41604 36360
rect 40819 36329 40831 36332
rect 40773 36323 40831 36329
rect 41598 36320 41604 36332
rect 41656 36320 41662 36372
rect 36446 36184 36452 36236
rect 36504 36224 36510 36236
rect 36504 36196 36768 36224
rect 36504 36184 36510 36196
rect 36740 36165 36768 36196
rect 38102 36184 38108 36236
rect 38160 36224 38166 36236
rect 38160 36196 39160 36224
rect 38160 36184 38166 36196
rect 35805 36159 35863 36165
rect 35805 36156 35817 36159
rect 35492 36128 35817 36156
rect 35492 36116 35498 36128
rect 35805 36125 35817 36128
rect 35851 36156 35863 36159
rect 35897 36159 35955 36165
rect 35897 36156 35909 36159
rect 35851 36128 35909 36156
rect 35851 36125 35863 36128
rect 35805 36119 35863 36125
rect 35897 36125 35909 36128
rect 35943 36125 35955 36159
rect 35897 36119 35955 36125
rect 36081 36159 36139 36165
rect 36081 36125 36093 36159
rect 36127 36125 36139 36159
rect 36081 36119 36139 36125
rect 36357 36159 36415 36165
rect 36357 36125 36369 36159
rect 36403 36125 36415 36159
rect 36357 36119 36415 36125
rect 36725 36159 36783 36165
rect 36725 36125 36737 36159
rect 36771 36125 36783 36159
rect 36725 36119 36783 36125
rect 35618 36048 35624 36100
rect 35676 36088 35682 36100
rect 36096 36088 36124 36119
rect 36906 36116 36912 36168
rect 36964 36116 36970 36168
rect 37366 36116 37372 36168
rect 37424 36116 37430 36168
rect 38746 36116 38752 36168
rect 38804 36156 38810 36168
rect 39022 36156 39028 36168
rect 38804 36128 39028 36156
rect 38804 36116 38810 36128
rect 39022 36116 39028 36128
rect 39080 36116 39086 36168
rect 35676 36060 36124 36088
rect 35676 36048 35682 36060
rect 36446 36048 36452 36100
rect 36504 36088 36510 36100
rect 36924 36088 36952 36116
rect 36504 36060 36952 36088
rect 36504 36048 36510 36060
rect 37642 36048 37648 36100
rect 37700 36048 37706 36100
rect 39132 36088 39160 36196
rect 40126 36184 40132 36236
rect 40184 36184 40190 36236
rect 41322 36184 41328 36236
rect 41380 36224 41386 36236
rect 41601 36227 41659 36233
rect 41601 36224 41613 36227
rect 41380 36196 41613 36224
rect 41380 36184 41386 36196
rect 41601 36193 41613 36196
rect 41647 36193 41659 36227
rect 41601 36187 41659 36193
rect 39206 36116 39212 36168
rect 39264 36116 39270 36168
rect 39390 36116 39396 36168
rect 39448 36116 39454 36168
rect 40865 36159 40923 36165
rect 40865 36156 40877 36159
rect 39500 36128 40877 36156
rect 39500 36088 39528 36128
rect 40865 36125 40877 36128
rect 40911 36125 40923 36159
rect 40865 36119 40923 36125
rect 39132 36060 39528 36088
rect 40034 36048 40040 36100
rect 40092 36088 40098 36100
rect 40405 36091 40463 36097
rect 40405 36088 40417 36091
rect 40092 36060 40417 36088
rect 40092 36048 40098 36060
rect 40405 36057 40417 36060
rect 40451 36057 40463 36091
rect 40405 36051 40463 36057
rect 34480 35992 35296 36020
rect 34480 35980 34486 35992
rect 36078 35980 36084 36032
rect 36136 36020 36142 36032
rect 36538 36020 36544 36032
rect 36136 35992 36544 36020
rect 36136 35980 36142 35992
rect 36538 35980 36544 35992
rect 36596 35980 36602 36032
rect 38930 35980 38936 36032
rect 38988 36020 38994 36032
rect 39117 36023 39175 36029
rect 39117 36020 39129 36023
rect 38988 35992 39129 36020
rect 38988 35980 38994 35992
rect 39117 35989 39129 35992
rect 39163 36020 39175 36023
rect 39298 36020 39304 36032
rect 39163 35992 39304 36020
rect 39163 35989 39175 35992
rect 39117 35983 39175 35989
rect 39298 35980 39304 35992
rect 39356 35980 39362 36032
rect 40313 36023 40371 36029
rect 40313 35989 40325 36023
rect 40359 36020 40371 36023
rect 41230 36020 41236 36032
rect 40359 35992 41236 36020
rect 40359 35989 40371 35992
rect 40313 35983 40371 35989
rect 41230 35980 41236 35992
rect 41288 35980 41294 36032
rect 1104 35930 42504 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 42504 35930
rect 1104 35856 42504 35878
rect 3602 35776 3608 35828
rect 3660 35816 3666 35828
rect 5626 35816 5632 35828
rect 3660 35788 5632 35816
rect 3660 35776 3666 35788
rect 5626 35776 5632 35788
rect 5684 35816 5690 35828
rect 5684 35788 5764 35816
rect 5684 35776 5690 35788
rect 5736 35757 5764 35788
rect 6086 35776 6092 35828
rect 6144 35776 6150 35828
rect 9674 35776 9680 35828
rect 9732 35816 9738 35828
rect 11011 35819 11069 35825
rect 9732 35788 9904 35816
rect 9732 35776 9738 35788
rect 5721 35751 5779 35757
rect 4556 35720 5488 35748
rect 2774 35640 2780 35692
rect 2832 35680 2838 35692
rect 3694 35680 3700 35692
rect 2832 35652 3700 35680
rect 2832 35640 2838 35652
rect 3694 35640 3700 35652
rect 3752 35640 3758 35692
rect 3878 35640 3884 35692
rect 3936 35680 3942 35692
rect 4249 35683 4307 35689
rect 4249 35680 4261 35683
rect 3936 35652 4261 35680
rect 3936 35640 3942 35652
rect 4249 35649 4261 35652
rect 4295 35649 4307 35683
rect 4249 35643 4307 35649
rect 1394 35572 1400 35624
rect 1452 35572 1458 35624
rect 1673 35615 1731 35621
rect 1673 35581 1685 35615
rect 1719 35612 1731 35615
rect 2866 35612 2872 35624
rect 1719 35584 2872 35612
rect 1719 35581 1731 35584
rect 1673 35575 1731 35581
rect 2866 35572 2872 35584
rect 2924 35572 2930 35624
rect 3329 35615 3387 35621
rect 3329 35581 3341 35615
rect 3375 35612 3387 35615
rect 3418 35612 3424 35624
rect 3375 35584 3424 35612
rect 3375 35581 3387 35584
rect 3329 35575 3387 35581
rect 3418 35572 3424 35584
rect 3476 35572 3482 35624
rect 3510 35572 3516 35624
rect 3568 35612 3574 35624
rect 3605 35615 3663 35621
rect 3605 35612 3617 35615
rect 3568 35584 3617 35612
rect 3568 35572 3574 35584
rect 3605 35581 3617 35584
rect 3651 35612 3663 35615
rect 4556 35612 4584 35720
rect 5460 35692 5488 35720
rect 5721 35717 5733 35751
rect 5767 35717 5779 35751
rect 9876 35748 9904 35788
rect 11011 35785 11023 35819
rect 11057 35816 11069 35819
rect 12066 35816 12072 35828
rect 11057 35788 12072 35816
rect 11057 35785 11069 35788
rect 11011 35779 11069 35785
rect 12066 35776 12072 35788
rect 12124 35776 12130 35828
rect 13541 35819 13599 35825
rect 13541 35785 13553 35819
rect 13587 35816 13599 35819
rect 14274 35816 14280 35828
rect 13587 35788 14280 35816
rect 13587 35785 13599 35788
rect 13541 35779 13599 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 14642 35776 14648 35828
rect 14700 35776 14706 35828
rect 16942 35776 16948 35828
rect 17000 35776 17006 35828
rect 17126 35776 17132 35828
rect 17184 35816 17190 35828
rect 17405 35819 17463 35825
rect 17405 35816 17417 35819
rect 17184 35788 17417 35816
rect 17184 35776 17190 35788
rect 17405 35785 17417 35788
rect 17451 35785 17463 35819
rect 17405 35779 17463 35785
rect 20898 35776 20904 35828
rect 20956 35816 20962 35828
rect 21821 35819 21879 35825
rect 21821 35816 21833 35819
rect 20956 35788 21833 35816
rect 20956 35776 20962 35788
rect 21821 35785 21833 35788
rect 21867 35785 21879 35819
rect 21821 35779 21879 35785
rect 22462 35776 22468 35828
rect 22520 35816 22526 35828
rect 22925 35819 22983 35825
rect 22925 35816 22937 35819
rect 22520 35788 22937 35816
rect 22520 35776 22526 35788
rect 22925 35785 22937 35788
rect 22971 35785 22983 35819
rect 22925 35779 22983 35785
rect 23293 35819 23351 35825
rect 23293 35785 23305 35819
rect 23339 35816 23351 35819
rect 24578 35816 24584 35828
rect 23339 35788 24584 35816
rect 23339 35785 23351 35788
rect 23293 35779 23351 35785
rect 24578 35776 24584 35788
rect 24636 35776 24642 35828
rect 27341 35819 27399 35825
rect 27341 35785 27353 35819
rect 27387 35816 27399 35819
rect 27522 35816 27528 35828
rect 27387 35788 27528 35816
rect 27387 35785 27399 35788
rect 27341 35779 27399 35785
rect 27522 35776 27528 35788
rect 27580 35776 27586 35828
rect 27890 35776 27896 35828
rect 27948 35816 27954 35828
rect 28261 35819 28319 35825
rect 28261 35816 28273 35819
rect 27948 35788 28273 35816
rect 27948 35776 27954 35788
rect 28261 35785 28273 35788
rect 28307 35785 28319 35819
rect 28261 35779 28319 35785
rect 28629 35819 28687 35825
rect 28629 35785 28641 35819
rect 28675 35816 28687 35819
rect 29086 35816 29092 35828
rect 28675 35788 29092 35816
rect 28675 35785 28687 35788
rect 28629 35779 28687 35785
rect 29086 35776 29092 35788
rect 29144 35776 29150 35828
rect 29638 35776 29644 35828
rect 29696 35816 29702 35828
rect 29733 35819 29791 35825
rect 29733 35816 29745 35819
rect 29696 35788 29745 35816
rect 29696 35776 29702 35788
rect 29733 35785 29745 35788
rect 29779 35785 29791 35819
rect 31202 35816 31208 35828
rect 29733 35779 29791 35785
rect 30300 35788 31208 35816
rect 9876 35720 9982 35748
rect 5721 35711 5779 35717
rect 11698 35708 11704 35760
rect 11756 35748 11762 35760
rect 11793 35751 11851 35757
rect 11793 35748 11805 35751
rect 11756 35720 11805 35748
rect 11756 35708 11762 35720
rect 11793 35717 11805 35720
rect 11839 35717 11851 35751
rect 14182 35748 14188 35760
rect 13018 35720 14188 35748
rect 11793 35711 11851 35717
rect 14182 35708 14188 35720
rect 14240 35708 14246 35760
rect 18230 35708 18236 35760
rect 18288 35708 18294 35760
rect 19518 35748 19524 35760
rect 19458 35720 19524 35748
rect 19518 35708 19524 35720
rect 19576 35708 19582 35760
rect 22830 35708 22836 35760
rect 22888 35748 22894 35760
rect 23198 35748 23204 35760
rect 22888 35720 23204 35748
rect 22888 35708 22894 35720
rect 23198 35708 23204 35720
rect 23256 35748 23262 35760
rect 25774 35748 25780 35760
rect 23256 35720 24164 35748
rect 25622 35720 25780 35748
rect 23256 35708 23262 35720
rect 4614 35640 4620 35692
rect 4672 35680 4678 35692
rect 5169 35683 5227 35689
rect 5169 35680 5181 35683
rect 4672 35652 5181 35680
rect 4672 35640 4678 35652
rect 5169 35649 5181 35652
rect 5215 35649 5227 35683
rect 5169 35643 5227 35649
rect 5258 35640 5264 35692
rect 5316 35640 5322 35692
rect 5353 35686 5411 35689
rect 5352 35683 5411 35686
rect 5352 35649 5365 35683
rect 5399 35649 5411 35683
rect 5352 35643 5411 35649
rect 3651 35584 4584 35612
rect 3651 35581 3663 35584
rect 3605 35575 3663 35581
rect 4890 35572 4896 35624
rect 4948 35572 4954 35624
rect 4985 35547 5043 35553
rect 4985 35544 4997 35547
rect 2700 35516 4997 35544
rect 2130 35436 2136 35488
rect 2188 35476 2194 35488
rect 2700 35476 2728 35516
rect 4985 35513 4997 35516
rect 5031 35513 5043 35547
rect 4985 35507 5043 35513
rect 5352 35544 5380 35643
rect 5442 35640 5448 35692
rect 5500 35689 5506 35692
rect 5500 35683 5549 35689
rect 5500 35649 5503 35683
rect 5537 35680 5549 35683
rect 5537 35652 5764 35680
rect 5537 35649 5549 35652
rect 5500 35643 5549 35649
rect 5500 35640 5506 35643
rect 5626 35572 5632 35624
rect 5684 35572 5690 35624
rect 5736 35612 5764 35652
rect 5902 35640 5908 35692
rect 5960 35640 5966 35692
rect 7561 35683 7619 35689
rect 7561 35649 7573 35683
rect 7607 35680 7619 35683
rect 7650 35680 7656 35692
rect 7607 35652 7656 35680
rect 7607 35649 7619 35652
rect 7561 35643 7619 35649
rect 7650 35640 7656 35652
rect 7708 35640 7714 35692
rect 7745 35683 7803 35689
rect 7745 35649 7757 35683
rect 7791 35680 7803 35683
rect 8202 35680 8208 35692
rect 7791 35652 8208 35680
rect 7791 35649 7803 35652
rect 7745 35643 7803 35649
rect 8202 35640 8208 35652
rect 8260 35640 8266 35692
rect 13816 35683 13874 35689
rect 13816 35649 13828 35683
rect 13862 35649 13874 35683
rect 13816 35643 13874 35649
rect 13909 35683 13967 35689
rect 13909 35649 13921 35683
rect 13955 35680 13967 35683
rect 14274 35680 14280 35692
rect 13955 35652 14280 35680
rect 13955 35649 13967 35652
rect 13909 35643 13967 35649
rect 6270 35612 6276 35624
rect 5736 35584 6276 35612
rect 6270 35572 6276 35584
rect 6328 35572 6334 35624
rect 9217 35615 9275 35621
rect 9217 35581 9229 35615
rect 9263 35612 9275 35615
rect 9490 35612 9496 35624
rect 9263 35584 9496 35612
rect 9263 35581 9275 35584
rect 9217 35575 9275 35581
rect 9490 35572 9496 35584
rect 9548 35572 9554 35624
rect 9585 35615 9643 35621
rect 9585 35581 9597 35615
rect 9631 35612 9643 35615
rect 9858 35612 9864 35624
rect 9631 35584 9864 35612
rect 9631 35581 9643 35584
rect 9585 35575 9643 35581
rect 9858 35572 9864 35584
rect 9916 35572 9922 35624
rect 11514 35572 11520 35624
rect 11572 35572 11578 35624
rect 13832 35612 13860 35643
rect 14274 35640 14280 35652
rect 14332 35640 14338 35692
rect 15013 35683 15071 35689
rect 15013 35649 15025 35683
rect 15059 35680 15071 35683
rect 15194 35680 15200 35692
rect 15059 35652 15200 35680
rect 15059 35649 15071 35652
rect 15013 35643 15071 35649
rect 15194 35640 15200 35652
rect 15252 35640 15258 35692
rect 15470 35640 15476 35692
rect 15528 35640 15534 35692
rect 17034 35680 17040 35692
rect 16592 35652 17040 35680
rect 16592 35624 16620 35652
rect 17034 35640 17040 35652
rect 17092 35640 17098 35692
rect 19886 35680 19892 35692
rect 19628 35652 19892 35680
rect 14366 35612 14372 35624
rect 13832 35584 14372 35612
rect 14366 35572 14372 35584
rect 14424 35572 14430 35624
rect 15102 35572 15108 35624
rect 15160 35572 15166 35624
rect 15286 35572 15292 35624
rect 15344 35572 15350 35624
rect 16485 35615 16543 35621
rect 16485 35581 16497 35615
rect 16531 35612 16543 35615
rect 16574 35612 16580 35624
rect 16531 35584 16580 35612
rect 16531 35581 16543 35584
rect 16485 35575 16543 35581
rect 16574 35572 16580 35584
rect 16632 35572 16638 35624
rect 16850 35572 16856 35624
rect 16908 35612 16914 35624
rect 16908 35584 17264 35612
rect 16908 35572 16914 35584
rect 5442 35544 5448 35556
rect 5352 35516 5448 35544
rect 2188 35448 2728 35476
rect 3145 35479 3203 35485
rect 2188 35436 2194 35448
rect 3145 35445 3157 35479
rect 3191 35476 3203 35479
rect 3970 35476 3976 35488
rect 3191 35448 3976 35476
rect 3191 35445 3203 35448
rect 3145 35439 3203 35445
rect 3970 35436 3976 35448
rect 4028 35436 4034 35488
rect 4062 35436 4068 35488
rect 4120 35476 4126 35488
rect 5352 35476 5380 35516
rect 5442 35504 5448 35516
rect 5500 35504 5506 35556
rect 4120 35448 5380 35476
rect 7745 35479 7803 35485
rect 4120 35436 4126 35448
rect 7745 35445 7757 35479
rect 7791 35476 7803 35479
rect 7834 35476 7840 35488
rect 7791 35448 7840 35476
rect 7791 35445 7803 35448
rect 7745 35439 7803 35445
rect 7834 35436 7840 35448
rect 7892 35436 7898 35488
rect 13262 35436 13268 35488
rect 13320 35436 13326 35488
rect 15654 35436 15660 35488
rect 15712 35436 15718 35488
rect 15841 35479 15899 35485
rect 15841 35445 15853 35479
rect 15887 35476 15899 35479
rect 16022 35476 16028 35488
rect 15887 35448 16028 35476
rect 15887 35445 15899 35448
rect 15841 35439 15899 35445
rect 16022 35436 16028 35448
rect 16080 35436 16086 35488
rect 17236 35476 17264 35584
rect 17310 35572 17316 35624
rect 17368 35612 17374 35624
rect 17957 35615 18015 35621
rect 17957 35612 17969 35615
rect 17368 35584 17969 35612
rect 17368 35572 17374 35584
rect 17957 35581 17969 35584
rect 18003 35612 18015 35615
rect 19628 35612 19656 35652
rect 19886 35640 19892 35652
rect 19944 35640 19950 35692
rect 20162 35640 20168 35692
rect 20220 35640 20226 35692
rect 20257 35683 20315 35689
rect 20257 35649 20269 35683
rect 20303 35680 20315 35683
rect 20530 35680 20536 35692
rect 20303 35652 20536 35680
rect 20303 35649 20315 35652
rect 20257 35643 20315 35649
rect 20530 35640 20536 35652
rect 20588 35640 20594 35692
rect 22189 35683 22247 35689
rect 22189 35649 22201 35683
rect 22235 35649 22247 35683
rect 22189 35643 22247 35649
rect 18003 35584 19656 35612
rect 19705 35615 19763 35621
rect 18003 35581 18015 35584
rect 17957 35575 18015 35581
rect 19705 35581 19717 35615
rect 19751 35612 19763 35615
rect 20070 35612 20076 35624
rect 19751 35584 20076 35612
rect 19751 35581 19763 35584
rect 19705 35575 19763 35581
rect 20070 35572 20076 35584
rect 20128 35572 20134 35624
rect 20438 35572 20444 35624
rect 20496 35572 20502 35624
rect 19794 35504 19800 35556
rect 19852 35504 19858 35556
rect 22204 35544 22232 35643
rect 23290 35640 23296 35692
rect 23348 35680 23354 35692
rect 24136 35689 24164 35720
rect 25774 35708 25780 35720
rect 25832 35708 25838 35760
rect 30300 35748 30328 35788
rect 31202 35776 31208 35788
rect 31260 35776 31266 35828
rect 31941 35819 31999 35825
rect 31941 35785 31953 35819
rect 31987 35816 31999 35819
rect 32766 35816 32772 35828
rect 31987 35788 32772 35816
rect 31987 35785 31999 35788
rect 31941 35779 31999 35785
rect 32766 35776 32772 35788
rect 32824 35776 32830 35828
rect 34241 35819 34299 35825
rect 34241 35785 34253 35819
rect 34287 35816 34299 35819
rect 34422 35816 34428 35828
rect 34287 35788 34428 35816
rect 34287 35785 34299 35788
rect 34241 35779 34299 35785
rect 34422 35776 34428 35788
rect 34480 35776 34486 35828
rect 37642 35776 37648 35828
rect 37700 35816 37706 35828
rect 37921 35819 37979 35825
rect 37921 35816 37933 35819
rect 37700 35788 37933 35816
rect 37700 35776 37706 35788
rect 37921 35785 37933 35788
rect 37967 35785 37979 35819
rect 40221 35819 40279 35825
rect 37921 35779 37979 35785
rect 38304 35788 40172 35816
rect 30208 35720 30328 35748
rect 30469 35751 30527 35757
rect 23385 35683 23443 35689
rect 23385 35680 23397 35683
rect 23348 35652 23397 35680
rect 23348 35640 23354 35652
rect 23385 35649 23397 35652
rect 23431 35649 23443 35683
rect 23385 35643 23443 35649
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35649 24179 35683
rect 30098 35680 30104 35692
rect 24121 35643 24179 35649
rect 29564 35652 30104 35680
rect 22278 35572 22284 35624
rect 22336 35572 22342 35624
rect 22465 35615 22523 35621
rect 22465 35581 22477 35615
rect 22511 35612 22523 35615
rect 23106 35612 23112 35624
rect 22511 35584 23112 35612
rect 22511 35581 22523 35584
rect 22465 35575 22523 35581
rect 23106 35572 23112 35584
rect 23164 35612 23170 35624
rect 23477 35615 23535 35621
rect 23477 35612 23489 35615
rect 23164 35584 23489 35612
rect 23164 35572 23170 35584
rect 23477 35581 23489 35584
rect 23523 35581 23535 35615
rect 23477 35575 23535 35581
rect 24397 35615 24455 35621
rect 24397 35581 24409 35615
rect 24443 35612 24455 35615
rect 24762 35612 24768 35624
rect 24443 35584 24768 35612
rect 24443 35581 24455 35584
rect 24397 35575 24455 35581
rect 24762 35572 24768 35584
rect 24820 35572 24826 35624
rect 25869 35615 25927 35621
rect 25869 35581 25881 35615
rect 25915 35612 25927 35615
rect 26142 35612 26148 35624
rect 25915 35584 26148 35612
rect 25915 35581 25927 35584
rect 25869 35575 25927 35581
rect 26142 35572 26148 35584
rect 26200 35612 26206 35624
rect 26513 35615 26571 35621
rect 26513 35612 26525 35615
rect 26200 35584 26525 35612
rect 26200 35572 26206 35584
rect 26513 35581 26525 35584
rect 26559 35581 26571 35615
rect 26513 35575 26571 35581
rect 26970 35572 26976 35624
rect 27028 35612 27034 35624
rect 27433 35615 27491 35621
rect 27433 35612 27445 35615
rect 27028 35584 27445 35612
rect 27028 35572 27034 35584
rect 27433 35581 27445 35584
rect 27479 35581 27491 35615
rect 27433 35575 27491 35581
rect 27617 35615 27675 35621
rect 27617 35581 27629 35615
rect 27663 35581 27675 35615
rect 27617 35575 27675 35581
rect 24026 35544 24032 35556
rect 22204 35516 24032 35544
rect 24026 35504 24032 35516
rect 24084 35504 24090 35556
rect 25406 35504 25412 35556
rect 25464 35544 25470 35556
rect 25961 35547 26019 35553
rect 25961 35544 25973 35547
rect 25464 35516 25973 35544
rect 25464 35504 25470 35516
rect 25961 35513 25973 35516
rect 26007 35513 26019 35547
rect 25961 35507 26019 35513
rect 27338 35504 27344 35556
rect 27396 35544 27402 35556
rect 27632 35544 27660 35575
rect 28718 35572 28724 35624
rect 28776 35572 28782 35624
rect 28905 35615 28963 35621
rect 28905 35581 28917 35615
rect 28951 35612 28963 35615
rect 28994 35612 29000 35624
rect 28951 35584 29000 35612
rect 28951 35581 28963 35584
rect 28905 35575 28963 35581
rect 28920 35544 28948 35575
rect 28994 35572 29000 35584
rect 29052 35612 29058 35624
rect 29564 35621 29592 35652
rect 30098 35640 30104 35652
rect 30156 35640 30162 35692
rect 30208 35689 30236 35720
rect 30469 35717 30481 35751
rect 30515 35748 30527 35751
rect 30742 35748 30748 35760
rect 30515 35720 30748 35748
rect 30515 35717 30527 35720
rect 30469 35711 30527 35717
rect 30742 35708 30748 35720
rect 30800 35708 30806 35760
rect 34054 35708 34060 35760
rect 34112 35748 34118 35760
rect 34333 35751 34391 35757
rect 34333 35748 34345 35751
rect 34112 35720 34345 35748
rect 34112 35708 34118 35720
rect 34333 35717 34345 35720
rect 34379 35717 34391 35751
rect 34333 35711 34391 35717
rect 37369 35751 37427 35757
rect 37369 35717 37381 35751
rect 37415 35748 37427 35751
rect 38304 35748 38332 35788
rect 37415 35720 38332 35748
rect 38381 35751 38439 35757
rect 37415 35717 37427 35720
rect 37369 35711 37427 35717
rect 38381 35717 38393 35751
rect 38427 35748 38439 35751
rect 39114 35748 39120 35760
rect 38427 35720 39120 35748
rect 38427 35717 38439 35720
rect 38381 35711 38439 35717
rect 39114 35708 39120 35720
rect 39172 35708 39178 35760
rect 40144 35748 40172 35788
rect 40221 35785 40233 35819
rect 40267 35816 40279 35819
rect 40402 35816 40408 35828
rect 40267 35788 40408 35816
rect 40267 35785 40279 35788
rect 40221 35779 40279 35785
rect 40402 35776 40408 35788
rect 40460 35776 40466 35828
rect 40586 35776 40592 35828
rect 40644 35776 40650 35828
rect 41049 35819 41107 35825
rect 41049 35785 41061 35819
rect 41095 35816 41107 35819
rect 41138 35816 41144 35828
rect 41095 35788 41144 35816
rect 41095 35785 41107 35788
rect 41049 35779 41107 35785
rect 41138 35776 41144 35788
rect 41196 35776 41202 35828
rect 41690 35748 41696 35760
rect 40144 35720 41696 35748
rect 41690 35708 41696 35720
rect 41748 35708 41754 35760
rect 30193 35683 30251 35689
rect 30193 35649 30205 35683
rect 30239 35649 30251 35683
rect 30193 35643 30251 35649
rect 31570 35640 31576 35692
rect 31628 35640 31634 35692
rect 33870 35640 33876 35692
rect 33928 35640 33934 35692
rect 35897 35683 35955 35689
rect 35897 35649 35909 35683
rect 35943 35680 35955 35683
rect 36357 35683 36415 35689
rect 36357 35680 36369 35683
rect 35943 35652 36369 35680
rect 35943 35649 35955 35652
rect 35897 35643 35955 35649
rect 36357 35649 36369 35652
rect 36403 35649 36415 35683
rect 36357 35643 36415 35649
rect 36906 35640 36912 35692
rect 36964 35640 36970 35692
rect 38289 35683 38347 35689
rect 38289 35649 38301 35683
rect 38335 35680 38347 35683
rect 38749 35683 38807 35689
rect 38749 35680 38761 35683
rect 38335 35652 38761 35680
rect 38335 35649 38347 35652
rect 38289 35643 38347 35649
rect 38749 35649 38761 35652
rect 38795 35649 38807 35683
rect 38749 35643 38807 35649
rect 39298 35640 39304 35692
rect 39356 35640 39362 35692
rect 41414 35640 41420 35692
rect 41472 35640 41478 35692
rect 29549 35615 29607 35621
rect 29549 35612 29561 35615
rect 29052 35584 29561 35612
rect 29052 35572 29058 35584
rect 29549 35581 29561 35584
rect 29595 35581 29607 35615
rect 29549 35575 29607 35581
rect 29641 35615 29699 35621
rect 29641 35581 29653 35615
rect 29687 35612 29699 35615
rect 30834 35612 30840 35624
rect 29687 35584 30840 35612
rect 29687 35581 29699 35584
rect 29641 35575 29699 35581
rect 30834 35572 30840 35584
rect 30892 35572 30898 35624
rect 31202 35572 31208 35624
rect 31260 35612 31266 35624
rect 32398 35612 32404 35624
rect 31260 35584 32404 35612
rect 31260 35572 31266 35584
rect 32398 35572 32404 35584
rect 32456 35612 32462 35624
rect 32493 35615 32551 35621
rect 32493 35612 32505 35615
rect 32456 35584 32505 35612
rect 32456 35572 32462 35584
rect 32493 35581 32505 35584
rect 32539 35581 32551 35615
rect 32493 35575 32551 35581
rect 32769 35615 32827 35621
rect 32769 35581 32781 35615
rect 32815 35612 32827 35615
rect 33778 35612 33784 35624
rect 32815 35584 33784 35612
rect 32815 35581 32827 35584
rect 32769 35575 32827 35581
rect 33778 35572 33784 35584
rect 33836 35572 33842 35624
rect 34698 35572 34704 35624
rect 34756 35612 34762 35624
rect 34885 35615 34943 35621
rect 34885 35612 34897 35615
rect 34756 35584 34897 35612
rect 34756 35572 34762 35584
rect 34885 35581 34897 35584
rect 34931 35612 34943 35615
rect 35434 35612 35440 35624
rect 34931 35584 35440 35612
rect 34931 35581 34943 35584
rect 34885 35575 34943 35581
rect 35434 35572 35440 35584
rect 35492 35572 35498 35624
rect 35986 35572 35992 35624
rect 36044 35572 36050 35624
rect 36078 35572 36084 35624
rect 36136 35572 36142 35624
rect 36538 35572 36544 35624
rect 36596 35612 36602 35624
rect 38470 35612 38476 35624
rect 36596 35584 38476 35612
rect 36596 35572 36602 35584
rect 38470 35572 38476 35584
rect 38528 35612 38534 35624
rect 40126 35612 40132 35624
rect 38528 35584 40132 35612
rect 38528 35572 38534 35584
rect 40126 35572 40132 35584
rect 40184 35572 40190 35624
rect 40402 35572 40408 35624
rect 40460 35612 40466 35624
rect 40681 35615 40739 35621
rect 40681 35612 40693 35615
rect 40460 35584 40693 35612
rect 40460 35572 40466 35584
rect 40681 35581 40693 35584
rect 40727 35581 40739 35615
rect 40681 35575 40739 35581
rect 40773 35615 40831 35621
rect 40773 35581 40785 35615
rect 40819 35612 40831 35615
rect 41046 35612 41052 35624
rect 40819 35584 41052 35612
rect 40819 35581 40831 35584
rect 40773 35575 40831 35581
rect 27396 35516 28948 35544
rect 40144 35544 40172 35572
rect 40788 35544 40816 35575
rect 41046 35572 41052 35584
rect 41104 35572 41110 35624
rect 41506 35572 41512 35624
rect 41564 35572 41570 35624
rect 41601 35615 41659 35621
rect 41601 35581 41613 35615
rect 41647 35581 41659 35615
rect 41601 35575 41659 35581
rect 40144 35516 40816 35544
rect 27396 35504 27402 35516
rect 41138 35504 41144 35556
rect 41196 35544 41202 35556
rect 41616 35544 41644 35575
rect 41196 35516 41644 35544
rect 41196 35504 41202 35516
rect 20438 35476 20444 35488
rect 17236 35448 20444 35476
rect 20438 35436 20444 35448
rect 20496 35436 20502 35488
rect 26142 35436 26148 35488
rect 26200 35476 26206 35488
rect 26973 35479 27031 35485
rect 26973 35476 26985 35479
rect 26200 35448 26985 35476
rect 26200 35436 26206 35448
rect 26973 35445 26985 35448
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 30101 35479 30159 35485
rect 30101 35445 30113 35479
rect 30147 35476 30159 35479
rect 31018 35476 31024 35488
rect 30147 35448 31024 35476
rect 30147 35445 30159 35448
rect 30101 35439 30159 35445
rect 31018 35436 31024 35448
rect 31076 35436 31082 35488
rect 33226 35436 33232 35488
rect 33284 35476 33290 35488
rect 33870 35476 33876 35488
rect 33284 35448 33876 35476
rect 33284 35436 33290 35448
rect 33870 35436 33876 35448
rect 33928 35436 33934 35488
rect 35526 35436 35532 35488
rect 35584 35436 35590 35488
rect 36354 35436 36360 35488
rect 36412 35476 36418 35488
rect 37461 35479 37519 35485
rect 37461 35476 37473 35479
rect 36412 35448 37473 35476
rect 36412 35436 36418 35448
rect 37461 35445 37473 35448
rect 37507 35445 37519 35479
rect 37461 35439 37519 35445
rect 1104 35386 42504 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 42504 35386
rect 1104 35312 42504 35334
rect 3605 35275 3663 35281
rect 3605 35241 3617 35275
rect 3651 35272 3663 35275
rect 3878 35272 3884 35284
rect 3651 35244 3884 35272
rect 3651 35241 3663 35244
rect 3605 35235 3663 35241
rect 3878 35232 3884 35244
rect 3936 35272 3942 35284
rect 4525 35275 4583 35281
rect 4525 35272 4537 35275
rect 3936 35244 4537 35272
rect 3936 35232 3942 35244
rect 4525 35241 4537 35244
rect 4571 35241 4583 35275
rect 5258 35272 5264 35284
rect 4525 35235 4583 35241
rect 4724 35244 5264 35272
rect 4249 35207 4307 35213
rect 4249 35173 4261 35207
rect 4295 35204 4307 35207
rect 4724 35204 4752 35244
rect 5258 35232 5264 35244
rect 5316 35232 5322 35284
rect 9858 35232 9864 35284
rect 9916 35232 9922 35284
rect 10704 35244 12020 35272
rect 4295 35176 4752 35204
rect 4295 35173 4307 35176
rect 4249 35167 4307 35173
rect 9674 35164 9680 35216
rect 9732 35204 9738 35216
rect 10704 35204 10732 35244
rect 9732 35176 10732 35204
rect 9732 35164 9738 35176
rect 1394 35096 1400 35148
rect 1452 35136 1458 35148
rect 1857 35139 1915 35145
rect 1857 35136 1869 35139
rect 1452 35108 1869 35136
rect 1452 35096 1458 35108
rect 1857 35105 1869 35108
rect 1903 35105 1915 35139
rect 1857 35099 1915 35105
rect 2130 35096 2136 35148
rect 2188 35096 2194 35148
rect 2682 35096 2688 35148
rect 2740 35136 2746 35148
rect 4801 35139 4859 35145
rect 4801 35136 4813 35139
rect 2740 35108 4813 35136
rect 2740 35096 2746 35108
rect 4801 35105 4813 35108
rect 4847 35136 4859 35139
rect 6822 35136 6828 35148
rect 4847 35108 6828 35136
rect 4847 35105 4859 35108
rect 4801 35099 4859 35105
rect 6822 35096 6828 35108
rect 6880 35136 6886 35148
rect 7009 35139 7067 35145
rect 7009 35136 7021 35139
rect 6880 35108 7021 35136
rect 6880 35096 6886 35108
rect 7009 35105 7021 35108
rect 7055 35136 7067 35139
rect 7282 35136 7288 35148
rect 7055 35108 7288 35136
rect 7055 35105 7067 35108
rect 7009 35099 7067 35105
rect 7282 35096 7288 35108
rect 7340 35096 7346 35148
rect 9582 35096 9588 35148
rect 9640 35136 9646 35148
rect 10597 35139 10655 35145
rect 10597 35136 10609 35139
rect 9640 35108 10609 35136
rect 9640 35096 9646 35108
rect 10597 35105 10609 35108
rect 10643 35136 10655 35139
rect 11514 35136 11520 35148
rect 10643 35108 11520 35136
rect 10643 35105 10655 35108
rect 10597 35099 10655 35105
rect 11514 35096 11520 35108
rect 11572 35096 11578 35148
rect 3602 35028 3608 35080
rect 3660 35068 3666 35080
rect 3789 35071 3847 35077
rect 3789 35068 3801 35071
rect 3660 35040 3801 35068
rect 3660 35028 3666 35040
rect 3789 35037 3801 35040
rect 3835 35037 3847 35071
rect 3789 35031 3847 35037
rect 3878 35028 3884 35080
rect 3936 35068 3942 35080
rect 4065 35071 4123 35077
rect 4065 35068 4077 35071
rect 3936 35040 4077 35068
rect 3936 35028 3942 35040
rect 4065 35037 4077 35040
rect 4111 35037 4123 35071
rect 4065 35031 4123 35037
rect 10042 35028 10048 35080
rect 10100 35028 10106 35080
rect 10321 35071 10379 35077
rect 10321 35037 10333 35071
rect 10367 35037 10379 35071
rect 10321 35031 10379 35037
rect 3694 35000 3700 35012
rect 3358 34972 3700 35000
rect 3694 34960 3700 34972
rect 3752 34960 3758 35012
rect 3970 35000 3976 35012
rect 3896 34972 3976 35000
rect 3896 34941 3924 34972
rect 3970 34960 3976 34972
rect 4028 35000 4034 35012
rect 4338 35000 4344 35012
rect 4028 34972 4344 35000
rect 4028 34960 4034 34972
rect 4338 34960 4344 34972
rect 4396 34960 4402 35012
rect 5084 35003 5142 35009
rect 5084 34969 5096 35003
rect 5130 35000 5142 35003
rect 6362 35000 6368 35012
rect 5130 34972 5212 35000
rect 6302 34972 6368 35000
rect 5130 34969 5142 34972
rect 5084 34963 5142 34969
rect 3881 34935 3939 34941
rect 3881 34901 3893 34935
rect 3927 34901 3939 34935
rect 3881 34895 3939 34901
rect 4062 34892 4068 34944
rect 4120 34932 4126 34944
rect 4541 34935 4599 34941
rect 4541 34932 4553 34935
rect 4120 34904 4553 34932
rect 4120 34892 4126 34904
rect 4541 34901 4553 34904
rect 4587 34901 4599 34935
rect 4541 34895 4599 34901
rect 4706 34892 4712 34944
rect 4764 34892 4770 34944
rect 5184 34932 5212 34972
rect 6362 34960 6368 34972
rect 6420 34960 6426 35012
rect 7285 35003 7343 35009
rect 7285 34969 7297 35003
rect 7331 35000 7343 35003
rect 7558 35000 7564 35012
rect 7331 34972 7564 35000
rect 7331 34969 7343 34972
rect 7285 34963 7343 34969
rect 7558 34960 7564 34972
rect 7616 34960 7622 35012
rect 9122 35000 9128 35012
rect 8510 34972 9128 35000
rect 9122 34960 9128 34972
rect 9180 35000 9186 35012
rect 9674 35000 9680 35012
rect 9180 34972 9680 35000
rect 9180 34960 9186 34972
rect 9674 34960 9680 34972
rect 9732 34960 9738 35012
rect 5258 34932 5264 34944
rect 5184 34904 5264 34932
rect 5258 34892 5264 34904
rect 5316 34892 5322 34944
rect 6454 34892 6460 34944
rect 6512 34932 6518 34944
rect 6549 34935 6607 34941
rect 6549 34932 6561 34935
rect 6512 34904 6561 34932
rect 6512 34892 6518 34904
rect 6549 34901 6561 34904
rect 6595 34901 6607 34935
rect 6549 34895 6607 34901
rect 8570 34892 8576 34944
rect 8628 34932 8634 34944
rect 8757 34935 8815 34941
rect 8757 34932 8769 34935
rect 8628 34904 8769 34932
rect 8628 34892 8634 34904
rect 8757 34901 8769 34904
rect 8803 34901 8815 34935
rect 10336 34932 10364 35031
rect 10502 35028 10508 35080
rect 10560 35028 10566 35080
rect 11992 35054 12020 35244
rect 12250 35232 12256 35284
rect 12308 35272 12314 35284
rect 12345 35275 12403 35281
rect 12345 35272 12357 35275
rect 12308 35244 12357 35272
rect 12308 35232 12314 35244
rect 12345 35241 12357 35244
rect 12391 35241 12403 35275
rect 12345 35235 12403 35241
rect 14185 35275 14243 35281
rect 14185 35241 14197 35275
rect 14231 35272 14243 35275
rect 15470 35272 15476 35284
rect 14231 35244 15476 35272
rect 14231 35241 14243 35244
rect 14185 35235 14243 35241
rect 15470 35232 15476 35244
rect 15528 35232 15534 35284
rect 15933 35275 15991 35281
rect 15933 35241 15945 35275
rect 15979 35272 15991 35275
rect 16574 35272 16580 35284
rect 15979 35244 16580 35272
rect 15979 35241 15991 35244
rect 15933 35235 15991 35241
rect 16574 35232 16580 35244
rect 16632 35232 16638 35284
rect 16942 35232 16948 35284
rect 17000 35272 17006 35284
rect 17862 35272 17868 35284
rect 17000 35244 17868 35272
rect 17000 35232 17006 35244
rect 17862 35232 17868 35244
rect 17920 35272 17926 35284
rect 19337 35275 19395 35281
rect 17920 35244 18460 35272
rect 17920 35232 17926 35244
rect 13998 35164 14004 35216
rect 14056 35204 14062 35216
rect 14645 35207 14703 35213
rect 14645 35204 14657 35207
rect 14056 35176 14657 35204
rect 14056 35164 14062 35176
rect 14645 35173 14657 35176
rect 14691 35173 14703 35207
rect 14645 35167 14703 35173
rect 13633 35139 13691 35145
rect 13633 35105 13645 35139
rect 13679 35136 13691 35139
rect 13679 35108 14044 35136
rect 13679 35105 13691 35108
rect 13633 35099 13691 35105
rect 14016 35080 14044 35108
rect 15286 35096 15292 35148
rect 15344 35096 15350 35148
rect 18432 35145 18460 35244
rect 19337 35241 19349 35275
rect 19383 35272 19395 35275
rect 19702 35272 19708 35284
rect 19383 35244 19708 35272
rect 19383 35241 19395 35244
rect 19337 35235 19395 35241
rect 19702 35232 19708 35244
rect 19760 35232 19766 35284
rect 22278 35232 22284 35284
rect 22336 35272 22342 35284
rect 22465 35275 22523 35281
rect 22465 35272 22477 35275
rect 22336 35244 22477 35272
rect 22336 35232 22342 35244
rect 22465 35241 22477 35244
rect 22511 35241 22523 35275
rect 22465 35235 22523 35241
rect 23290 35232 23296 35284
rect 23348 35272 23354 35284
rect 23477 35275 23535 35281
rect 23477 35272 23489 35275
rect 23348 35244 23489 35272
rect 23348 35232 23354 35244
rect 23477 35241 23489 35244
rect 23523 35241 23535 35275
rect 23477 35235 23535 35241
rect 24762 35232 24768 35284
rect 24820 35232 24826 35284
rect 27617 35275 27675 35281
rect 27617 35241 27629 35275
rect 27663 35272 27675 35275
rect 27706 35272 27712 35284
rect 27663 35244 27712 35272
rect 27663 35241 27675 35244
rect 27617 35235 27675 35241
rect 27706 35232 27712 35244
rect 27764 35232 27770 35284
rect 31389 35275 31447 35281
rect 31389 35241 31401 35275
rect 31435 35272 31447 35275
rect 31662 35272 31668 35284
rect 31435 35244 31668 35272
rect 31435 35241 31447 35244
rect 31389 35235 31447 35241
rect 31662 35232 31668 35244
rect 31720 35232 31726 35284
rect 36725 35275 36783 35281
rect 36725 35241 36737 35275
rect 36771 35272 36783 35275
rect 36906 35272 36912 35284
rect 36771 35244 36912 35272
rect 36771 35241 36783 35244
rect 36725 35235 36783 35241
rect 36906 35232 36912 35244
rect 36964 35232 36970 35284
rect 40402 35232 40408 35284
rect 40460 35232 40466 35284
rect 41230 35232 41236 35284
rect 41288 35232 41294 35284
rect 20438 35204 20444 35216
rect 19996 35176 20444 35204
rect 19996 35145 20024 35176
rect 20438 35164 20444 35176
rect 20496 35204 20502 35216
rect 20496 35176 21864 35204
rect 20496 35164 20502 35176
rect 18417 35139 18475 35145
rect 18417 35105 18429 35139
rect 18463 35105 18475 35139
rect 18417 35099 18475 35105
rect 19981 35139 20039 35145
rect 19981 35105 19993 35139
rect 20027 35105 20039 35139
rect 19981 35099 20039 35105
rect 20162 35096 20168 35148
rect 20220 35136 20226 35148
rect 21836 35145 21864 35176
rect 22370 35164 22376 35216
rect 22428 35164 22434 35216
rect 36446 35164 36452 35216
rect 36504 35204 36510 35216
rect 36504 35176 37412 35204
rect 36504 35164 36510 35176
rect 20349 35139 20407 35145
rect 20349 35136 20361 35139
rect 20220 35108 20361 35136
rect 20220 35096 20226 35108
rect 20349 35105 20361 35108
rect 20395 35105 20407 35139
rect 20349 35099 20407 35105
rect 21821 35139 21879 35145
rect 21821 35105 21833 35139
rect 21867 35136 21879 35139
rect 23017 35139 23075 35145
rect 23017 35136 23029 35139
rect 21867 35108 23029 35136
rect 21867 35105 21879 35108
rect 21821 35099 21879 35105
rect 23017 35105 23029 35108
rect 23063 35136 23075 35139
rect 23382 35136 23388 35148
rect 23063 35108 23388 35136
rect 23063 35105 23075 35108
rect 23017 35099 23075 35105
rect 23382 35096 23388 35108
rect 23440 35096 23446 35148
rect 24026 35136 24032 35148
rect 23952 35108 24032 35136
rect 13538 35028 13544 35080
rect 13596 35028 13602 35080
rect 13998 35028 14004 35080
rect 14056 35068 14062 35080
rect 14093 35071 14151 35077
rect 14093 35068 14105 35071
rect 14056 35040 14105 35068
rect 14056 35028 14062 35040
rect 14093 35037 14105 35040
rect 14139 35037 14151 35071
rect 14093 35031 14151 35037
rect 14274 35028 14280 35080
rect 14332 35028 14338 35080
rect 15013 35071 15071 35077
rect 15013 35037 15025 35071
rect 15059 35068 15071 35071
rect 15102 35068 15108 35080
rect 15059 35040 15108 35068
rect 15059 35037 15071 35040
rect 15013 35031 15071 35037
rect 15102 35028 15108 35040
rect 15160 35028 15166 35080
rect 15654 35028 15660 35080
rect 15712 35068 15718 35080
rect 15712 35040 17172 35068
rect 15712 35028 15718 35040
rect 10873 35003 10931 35009
rect 10873 34969 10885 35003
rect 10919 35000 10931 35003
rect 10962 35000 10968 35012
rect 10919 34972 10968 35000
rect 10919 34969 10931 34972
rect 10873 34963 10931 34969
rect 10962 34960 10968 34972
rect 11020 34960 11026 35012
rect 16482 34960 16488 35012
rect 16540 35000 16546 35012
rect 17046 35003 17104 35009
rect 17046 35000 17058 35003
rect 16540 34972 17058 35000
rect 16540 34960 16546 34972
rect 17046 34969 17058 34972
rect 17092 34969 17104 35003
rect 17144 35000 17172 35040
rect 17310 35028 17316 35080
rect 17368 35068 17374 35080
rect 17405 35071 17463 35077
rect 17405 35068 17417 35071
rect 17368 35040 17417 35068
rect 17368 35028 17374 35040
rect 17405 35037 17417 35040
rect 17451 35037 17463 35071
rect 17405 35031 17463 35037
rect 19797 35071 19855 35077
rect 19797 35037 19809 35071
rect 19843 35068 19855 35071
rect 20180 35068 20208 35096
rect 23952 35068 23980 35108
rect 24026 35096 24032 35108
rect 24084 35145 24090 35148
rect 24084 35139 24133 35145
rect 24084 35105 24087 35139
rect 24121 35105 24133 35139
rect 24084 35099 24133 35105
rect 25317 35139 25375 35145
rect 25317 35105 25329 35139
rect 25363 35136 25375 35139
rect 25590 35136 25596 35148
rect 25363 35108 25596 35136
rect 25363 35105 25375 35108
rect 25317 35099 25375 35105
rect 24084 35096 24090 35099
rect 25590 35096 25596 35108
rect 25648 35096 25654 35148
rect 25869 35139 25927 35145
rect 25869 35105 25881 35139
rect 25915 35136 25927 35139
rect 27430 35136 27436 35148
rect 25915 35108 27436 35136
rect 25915 35105 25927 35108
rect 25869 35099 25927 35105
rect 27430 35096 27436 35108
rect 27488 35096 27494 35148
rect 28813 35139 28871 35145
rect 28813 35105 28825 35139
rect 28859 35136 28871 35139
rect 28994 35136 29000 35148
rect 28859 35108 29000 35136
rect 28859 35105 28871 35108
rect 28813 35099 28871 35105
rect 28994 35096 29000 35108
rect 29052 35096 29058 35148
rect 29270 35136 29276 35148
rect 29104 35108 29276 35136
rect 19843 35040 20208 35068
rect 21928 35040 23980 35068
rect 25133 35071 25191 35077
rect 19843 35037 19855 35040
rect 19797 35031 19855 35037
rect 21928 35000 21956 35040
rect 25133 35037 25145 35071
rect 25179 35068 25191 35071
rect 25406 35068 25412 35080
rect 25179 35040 25412 35068
rect 25179 35037 25191 35040
rect 25133 35031 25191 35037
rect 25406 35028 25412 35040
rect 25464 35028 25470 35080
rect 29104 35068 29132 35108
rect 29270 35096 29276 35108
rect 29328 35096 29334 35148
rect 31938 35096 31944 35148
rect 31996 35096 32002 35148
rect 34790 35096 34796 35148
rect 34848 35136 34854 35148
rect 34977 35139 35035 35145
rect 34977 35136 34989 35139
rect 34848 35108 34989 35136
rect 34848 35096 34854 35108
rect 34977 35105 34989 35108
rect 35023 35136 35035 35139
rect 37274 35136 37280 35148
rect 35023 35108 37280 35136
rect 35023 35105 35035 35108
rect 34977 35099 35035 35105
rect 37274 35096 37280 35108
rect 37332 35096 37338 35148
rect 37384 35145 37412 35176
rect 37369 35139 37427 35145
rect 37369 35105 37381 35139
rect 37415 35105 37427 35139
rect 37369 35099 37427 35105
rect 38470 35096 38476 35148
rect 38528 35096 38534 35148
rect 39206 35096 39212 35148
rect 39264 35136 39270 35148
rect 39301 35139 39359 35145
rect 39301 35136 39313 35139
rect 39264 35108 39313 35136
rect 39264 35096 39270 35108
rect 39301 35105 39313 35108
rect 39347 35105 39359 35139
rect 39301 35099 39359 35105
rect 40034 35096 40040 35148
rect 40092 35136 40098 35148
rect 40957 35139 41015 35145
rect 40957 35136 40969 35139
rect 40092 35108 40969 35136
rect 40092 35096 40098 35108
rect 40957 35105 40969 35108
rect 41003 35136 41015 35139
rect 41138 35136 41144 35148
rect 41003 35108 41144 35136
rect 41003 35105 41015 35108
rect 40957 35099 41015 35105
rect 41138 35096 41144 35108
rect 41196 35136 41202 35148
rect 41785 35139 41843 35145
rect 41785 35136 41797 35139
rect 41196 35108 41797 35136
rect 41196 35096 41202 35108
rect 41785 35105 41797 35108
rect 41831 35105 41843 35139
rect 41785 35099 41843 35105
rect 27278 35040 29132 35068
rect 29178 35028 29184 35080
rect 29236 35068 29242 35080
rect 30101 35071 30159 35077
rect 30101 35068 30113 35071
rect 29236 35040 30113 35068
rect 29236 35028 29242 35040
rect 30101 35037 30113 35040
rect 30147 35037 30159 35071
rect 30101 35031 30159 35037
rect 36354 35028 36360 35080
rect 36412 35028 36418 35080
rect 17144 34972 21956 35000
rect 22005 35003 22063 35009
rect 17046 34963 17104 34969
rect 22005 34969 22017 35003
rect 22051 35000 22063 35003
rect 22278 35000 22284 35012
rect 22051 34972 22284 35000
rect 22051 34969 22063 34972
rect 22005 34963 22063 34969
rect 22278 34960 22284 34972
rect 22336 35000 22342 35012
rect 22925 35003 22983 35009
rect 22925 35000 22937 35003
rect 22336 34972 22937 35000
rect 22336 34960 22342 34972
rect 22925 34969 22937 34972
rect 22971 35000 22983 35003
rect 23198 35000 23204 35012
rect 22971 34972 23204 35000
rect 22971 34969 22983 34972
rect 22925 34963 22983 34969
rect 23198 34960 23204 34972
rect 23256 34960 23262 35012
rect 26142 34960 26148 35012
rect 26200 34960 26206 35012
rect 28537 35003 28595 35009
rect 28537 34969 28549 35003
rect 28583 35000 28595 35003
rect 29549 35003 29607 35009
rect 29549 35000 29561 35003
rect 28583 34972 29561 35000
rect 28583 34969 28595 34972
rect 28537 34963 28595 34969
rect 29549 34969 29561 34972
rect 29595 34969 29607 35003
rect 29549 34963 29607 34969
rect 32214 34960 32220 35012
rect 32272 34960 32278 35012
rect 35253 35003 35311 35009
rect 35253 34969 35265 35003
rect 35299 35000 35311 35003
rect 35526 35000 35532 35012
rect 35299 34972 35532 35000
rect 35299 34969 35311 34972
rect 35253 34963 35311 34969
rect 35526 34960 35532 34972
rect 35584 34960 35590 35012
rect 38102 35000 38108 35012
rect 36740 34972 38108 35000
rect 11054 34932 11060 34944
rect 10336 34904 11060 34932
rect 8757 34895 8815 34901
rect 11054 34892 11060 34904
rect 11112 34892 11118 34944
rect 13906 34892 13912 34944
rect 13964 34892 13970 34944
rect 15105 34935 15163 34941
rect 15105 34901 15117 34935
rect 15151 34932 15163 34935
rect 15194 34932 15200 34944
rect 15151 34904 15200 34932
rect 15151 34901 15163 34904
rect 15105 34895 15163 34901
rect 15194 34892 15200 34904
rect 15252 34932 15258 34944
rect 15654 34932 15660 34944
rect 15252 34904 15660 34932
rect 15252 34892 15258 34904
rect 15654 34892 15660 34904
rect 15712 34892 15718 34944
rect 17586 34892 17592 34944
rect 17644 34932 17650 34944
rect 17865 34935 17923 34941
rect 17865 34932 17877 34935
rect 17644 34904 17877 34932
rect 17644 34892 17650 34904
rect 17865 34901 17877 34904
rect 17911 34901 17923 34935
rect 17865 34895 17923 34901
rect 19705 34935 19763 34941
rect 19705 34901 19717 34935
rect 19751 34932 19763 34935
rect 20530 34932 20536 34944
rect 19751 34904 20536 34932
rect 19751 34901 19763 34904
rect 19705 34895 19763 34901
rect 20530 34892 20536 34904
rect 20588 34892 20594 34944
rect 20622 34892 20628 34944
rect 20680 34932 20686 34944
rect 20993 34935 21051 34941
rect 20993 34932 21005 34935
rect 20680 34904 21005 34932
rect 20680 34892 20686 34904
rect 20993 34901 21005 34904
rect 21039 34901 21051 34935
rect 20993 34895 21051 34901
rect 21913 34935 21971 34941
rect 21913 34901 21925 34935
rect 21959 34932 21971 34935
rect 22738 34932 22744 34944
rect 21959 34904 22744 34932
rect 21959 34901 21971 34904
rect 21913 34895 21971 34901
rect 22738 34892 22744 34904
rect 22796 34932 22802 34944
rect 22833 34935 22891 34941
rect 22833 34932 22845 34935
rect 22796 34904 22845 34932
rect 22796 34892 22802 34904
rect 22833 34901 22845 34904
rect 22879 34901 22891 34935
rect 22833 34895 22891 34901
rect 23842 34892 23848 34944
rect 23900 34892 23906 34944
rect 23934 34892 23940 34944
rect 23992 34892 23998 34944
rect 25222 34892 25228 34944
rect 25280 34892 25286 34944
rect 27706 34892 27712 34944
rect 27764 34932 27770 34944
rect 28169 34935 28227 34941
rect 28169 34932 28181 34935
rect 27764 34904 28181 34932
rect 27764 34892 27770 34904
rect 28169 34901 28181 34904
rect 28215 34901 28227 34935
rect 28169 34895 28227 34901
rect 28629 34935 28687 34941
rect 28629 34901 28641 34935
rect 28675 34932 28687 34935
rect 29454 34932 29460 34944
rect 28675 34904 29460 34932
rect 28675 34901 28687 34904
rect 28629 34895 28687 34901
rect 29454 34892 29460 34904
rect 29512 34892 29518 34944
rect 31754 34892 31760 34944
rect 31812 34892 31818 34944
rect 31849 34935 31907 34941
rect 31849 34901 31861 34935
rect 31895 34932 31907 34935
rect 32030 34932 32036 34944
rect 31895 34904 32036 34932
rect 31895 34901 31907 34904
rect 31849 34895 31907 34901
rect 32030 34892 32036 34904
rect 32088 34892 32094 34944
rect 32122 34892 32128 34944
rect 32180 34932 32186 34944
rect 33042 34932 33048 34944
rect 32180 34904 33048 34932
rect 32180 34892 32186 34904
rect 33042 34892 33048 34904
rect 33100 34932 33106 34944
rect 33505 34935 33563 34941
rect 33505 34932 33517 34935
rect 33100 34904 33517 34932
rect 33100 34892 33106 34904
rect 33505 34901 33517 34904
rect 33551 34932 33563 34935
rect 36740 34932 36768 34972
rect 38102 34960 38108 34972
rect 38160 34960 38166 35012
rect 38289 35003 38347 35009
rect 38289 34969 38301 35003
rect 38335 35000 38347 35003
rect 38749 35003 38807 35009
rect 38749 35000 38761 35003
rect 38335 34972 38761 35000
rect 38335 34969 38347 34972
rect 38289 34963 38347 34969
rect 38749 34969 38761 34972
rect 38795 34969 38807 35003
rect 38749 34963 38807 34969
rect 38930 34960 38936 35012
rect 38988 35000 38994 35012
rect 39945 35003 40003 35009
rect 39945 35000 39957 35003
rect 38988 34972 39957 35000
rect 38988 34960 38994 34972
rect 39945 34969 39957 34972
rect 39991 34969 40003 35003
rect 39945 34963 40003 34969
rect 40770 34960 40776 35012
rect 40828 35000 40834 35012
rect 41693 35003 41751 35009
rect 41693 35000 41705 35003
rect 40828 34972 41705 35000
rect 40828 34960 40834 34972
rect 41693 34969 41705 34972
rect 41739 34969 41751 35003
rect 41693 34963 41751 34969
rect 33551 34904 36768 34932
rect 33551 34901 33563 34904
rect 33505 34895 33563 34901
rect 36814 34892 36820 34944
rect 36872 34892 36878 34944
rect 37918 34892 37924 34944
rect 37976 34892 37982 34944
rect 38378 34892 38384 34944
rect 38436 34892 38442 34944
rect 40034 34892 40040 34944
rect 40092 34892 40098 34944
rect 40865 34935 40923 34941
rect 40865 34901 40877 34935
rect 40911 34932 40923 34935
rect 41230 34932 41236 34944
rect 40911 34904 41236 34932
rect 40911 34901 40923 34904
rect 40865 34895 40923 34901
rect 41230 34892 41236 34904
rect 41288 34932 41294 34944
rect 41601 34935 41659 34941
rect 41601 34932 41613 34935
rect 41288 34904 41613 34932
rect 41288 34892 41294 34904
rect 41601 34901 41613 34904
rect 41647 34901 41659 34935
rect 41601 34895 41659 34901
rect 1104 34842 42504 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 42504 34842
rect 1104 34768 42504 34790
rect 2958 34688 2964 34740
rect 3016 34728 3022 34740
rect 3421 34731 3479 34737
rect 3421 34728 3433 34731
rect 3016 34700 3433 34728
rect 3016 34688 3022 34700
rect 3421 34697 3433 34700
rect 3467 34697 3479 34731
rect 3421 34691 3479 34697
rect 4341 34731 4399 34737
rect 4341 34697 4353 34731
rect 4387 34728 4399 34731
rect 4614 34728 4620 34740
rect 4387 34700 4620 34728
rect 4387 34697 4399 34700
rect 4341 34691 4399 34697
rect 4614 34688 4620 34700
rect 4672 34688 4678 34740
rect 4801 34731 4859 34737
rect 4801 34697 4813 34731
rect 4847 34728 4859 34731
rect 5534 34728 5540 34740
rect 4847 34700 5540 34728
rect 4847 34697 4859 34700
rect 4801 34691 4859 34697
rect 5534 34688 5540 34700
rect 5592 34688 5598 34740
rect 6656 34700 11560 34728
rect 6656 34672 6684 34700
rect 3970 34660 3976 34672
rect 3436 34632 3976 34660
rect 3436 34601 3464 34632
rect 3970 34620 3976 34632
rect 4028 34620 4034 34672
rect 5626 34660 5632 34672
rect 5092 34632 5632 34660
rect 3421 34595 3479 34601
rect 3421 34561 3433 34595
rect 3467 34561 3479 34595
rect 3421 34555 3479 34561
rect 3602 34552 3608 34604
rect 3660 34592 3666 34604
rect 4062 34592 4068 34604
rect 3660 34564 4068 34592
rect 3660 34552 3666 34564
rect 4062 34552 4068 34564
rect 4120 34552 4126 34604
rect 4433 34595 4491 34601
rect 4433 34561 4445 34595
rect 4479 34592 4491 34595
rect 4706 34592 4712 34604
rect 4479 34564 4712 34592
rect 4479 34561 4491 34564
rect 4433 34555 4491 34561
rect 4706 34552 4712 34564
rect 4764 34592 4770 34604
rect 5092 34601 5120 34632
rect 5626 34620 5632 34632
rect 5684 34620 5690 34672
rect 6178 34620 6184 34672
rect 6236 34660 6242 34672
rect 6638 34660 6644 34672
rect 6236 34632 6644 34660
rect 6236 34620 6242 34632
rect 6638 34620 6644 34632
rect 6696 34620 6702 34672
rect 8202 34620 8208 34672
rect 8260 34660 8266 34672
rect 8541 34663 8599 34669
rect 8541 34660 8553 34663
rect 8260 34632 8553 34660
rect 8260 34620 8266 34632
rect 8541 34629 8553 34632
rect 8587 34629 8599 34663
rect 8541 34623 8599 34629
rect 8757 34663 8815 34669
rect 8757 34629 8769 34663
rect 8803 34660 8815 34663
rect 9398 34660 9404 34672
rect 8803 34632 9404 34660
rect 8803 34629 8815 34632
rect 8757 34623 8815 34629
rect 9398 34620 9404 34632
rect 9456 34620 9462 34672
rect 10962 34620 10968 34672
rect 11020 34620 11026 34672
rect 11532 34669 11560 34700
rect 11606 34688 11612 34740
rect 11664 34728 11670 34740
rect 12529 34731 12587 34737
rect 12529 34728 12541 34731
rect 11664 34700 12541 34728
rect 11664 34688 11670 34700
rect 12529 34697 12541 34700
rect 12575 34697 12587 34731
rect 12529 34691 12587 34697
rect 14001 34731 14059 34737
rect 14001 34697 14013 34731
rect 14047 34728 14059 34731
rect 14458 34728 14464 34740
rect 14047 34700 14464 34728
rect 14047 34697 14059 34700
rect 14001 34691 14059 34697
rect 14458 34688 14464 34700
rect 14516 34688 14522 34740
rect 16022 34688 16028 34740
rect 16080 34688 16086 34740
rect 16482 34688 16488 34740
rect 16540 34688 16546 34740
rect 16592 34700 17812 34728
rect 11517 34663 11575 34669
rect 11517 34629 11529 34663
rect 11563 34660 11575 34663
rect 12158 34660 12164 34672
rect 11563 34632 12164 34660
rect 11563 34629 11575 34632
rect 11517 34623 11575 34629
rect 12158 34620 12164 34632
rect 12216 34660 12222 34672
rect 12618 34660 12624 34672
rect 12216 34632 12624 34660
rect 12216 34620 12222 34632
rect 12618 34620 12624 34632
rect 12676 34620 12682 34672
rect 15562 34660 15568 34672
rect 14108 34632 15568 34660
rect 5077 34595 5135 34601
rect 5077 34592 5089 34595
rect 4764 34564 5089 34592
rect 4764 34552 4770 34564
rect 5077 34561 5089 34564
rect 5123 34561 5135 34595
rect 5077 34555 5135 34561
rect 5166 34552 5172 34604
rect 5224 34592 5230 34604
rect 5353 34595 5411 34601
rect 5353 34592 5365 34595
rect 5224 34564 5365 34592
rect 5224 34552 5230 34564
rect 5353 34561 5365 34564
rect 5399 34561 5411 34595
rect 5353 34555 5411 34561
rect 5445 34595 5503 34601
rect 5445 34561 5457 34595
rect 5491 34592 5503 34595
rect 6086 34592 6092 34604
rect 5491 34564 6092 34592
rect 5491 34561 5503 34564
rect 5445 34555 5503 34561
rect 6086 34552 6092 34564
rect 6144 34552 6150 34604
rect 6270 34552 6276 34604
rect 6328 34592 6334 34604
rect 6328 34564 7788 34592
rect 6328 34552 6334 34564
rect 4985 34527 5043 34533
rect 4985 34493 4997 34527
rect 5031 34524 5043 34527
rect 5537 34527 5595 34533
rect 5031 34496 5304 34524
rect 5031 34493 5043 34496
rect 4985 34487 5043 34493
rect 5276 34456 5304 34496
rect 5537 34493 5549 34527
rect 5583 34493 5595 34527
rect 5537 34487 5595 34493
rect 5552 34456 5580 34487
rect 7282 34484 7288 34536
rect 7340 34524 7346 34536
rect 7377 34527 7435 34533
rect 7377 34524 7389 34527
rect 7340 34496 7389 34524
rect 7340 34484 7346 34496
rect 7377 34493 7389 34496
rect 7423 34493 7435 34527
rect 7377 34487 7435 34493
rect 7558 34484 7564 34536
rect 7616 34524 7622 34536
rect 7760 34524 7788 34564
rect 7834 34552 7840 34604
rect 7892 34552 7898 34604
rect 7926 34552 7932 34604
rect 7984 34552 7990 34604
rect 10042 34552 10048 34604
rect 10100 34592 10106 34604
rect 10318 34592 10324 34604
rect 10100 34564 10324 34592
rect 10100 34552 10106 34564
rect 10318 34552 10324 34564
rect 10376 34592 10382 34604
rect 10597 34595 10655 34601
rect 10597 34592 10609 34595
rect 10376 34564 10609 34592
rect 10376 34552 10382 34564
rect 10597 34561 10609 34564
rect 10643 34561 10655 34595
rect 10597 34555 10655 34561
rect 10781 34595 10839 34601
rect 10781 34561 10793 34595
rect 10827 34592 10839 34595
rect 11054 34592 11060 34604
rect 10827 34564 11060 34592
rect 10827 34561 10839 34564
rect 10781 34555 10839 34561
rect 11054 34552 11060 34564
rect 11112 34552 11118 34604
rect 12894 34552 12900 34604
rect 12952 34552 12958 34604
rect 14108 34601 14136 34632
rect 15562 34620 15568 34632
rect 15620 34620 15626 34672
rect 16117 34663 16175 34669
rect 16117 34629 16129 34663
rect 16163 34660 16175 34663
rect 16592 34660 16620 34700
rect 17310 34660 17316 34672
rect 16163 34632 16620 34660
rect 16684 34632 17316 34660
rect 16163 34629 16175 34632
rect 16117 34623 16175 34629
rect 14093 34595 14151 34601
rect 14093 34561 14105 34595
rect 14139 34561 14151 34595
rect 14093 34555 14151 34561
rect 14360 34595 14418 34601
rect 14360 34561 14372 34595
rect 14406 34592 14418 34595
rect 14918 34592 14924 34604
rect 14406 34564 14924 34592
rect 14406 34561 14418 34564
rect 14360 34555 14418 34561
rect 14918 34552 14924 34564
rect 14976 34552 14982 34604
rect 15580 34592 15608 34620
rect 16684 34601 16712 34632
rect 17310 34620 17316 34632
rect 17368 34620 17374 34672
rect 17784 34660 17812 34700
rect 17862 34688 17868 34740
rect 17920 34728 17926 34740
rect 18049 34731 18107 34737
rect 18049 34728 18061 34731
rect 17920 34700 18061 34728
rect 17920 34688 17926 34700
rect 18049 34697 18061 34700
rect 18095 34697 18107 34731
rect 18049 34691 18107 34697
rect 20070 34688 20076 34740
rect 20128 34688 20134 34740
rect 20165 34731 20223 34737
rect 20165 34697 20177 34731
rect 20211 34697 20223 34731
rect 20165 34691 20223 34697
rect 18230 34660 18236 34672
rect 17784 34632 18236 34660
rect 18230 34620 18236 34632
rect 18288 34620 18294 34672
rect 18960 34663 19018 34669
rect 18960 34629 18972 34663
rect 19006 34660 19018 34663
rect 20180 34660 20208 34691
rect 20622 34688 20628 34740
rect 20680 34688 20686 34740
rect 23474 34688 23480 34740
rect 23532 34688 23538 34740
rect 23845 34731 23903 34737
rect 23845 34697 23857 34731
rect 23891 34728 23903 34731
rect 23934 34728 23940 34740
rect 23891 34700 23940 34728
rect 23891 34697 23903 34700
rect 23845 34691 23903 34697
rect 23934 34688 23940 34700
rect 23992 34688 23998 34740
rect 25222 34688 25228 34740
rect 25280 34688 25286 34740
rect 26050 34688 26056 34740
rect 26108 34688 26114 34740
rect 29178 34688 29184 34740
rect 29236 34688 29242 34740
rect 30006 34688 30012 34740
rect 30064 34688 30070 34740
rect 34149 34731 34207 34737
rect 30116 34700 34008 34728
rect 19006 34632 20208 34660
rect 22189 34663 22247 34669
rect 19006 34629 19018 34632
rect 18960 34623 19018 34629
rect 22189 34629 22201 34663
rect 22235 34660 22247 34663
rect 23290 34660 23296 34672
rect 22235 34632 23296 34660
rect 22235 34629 22247 34632
rect 22189 34623 22247 34629
rect 23290 34620 23296 34632
rect 23348 34620 23354 34672
rect 16942 34601 16948 34604
rect 16669 34595 16727 34601
rect 16669 34592 16681 34595
rect 15580 34564 16681 34592
rect 16669 34561 16681 34564
rect 16715 34561 16727 34595
rect 16669 34555 16727 34561
rect 16936 34555 16948 34601
rect 16942 34552 16948 34555
rect 17000 34552 17006 34604
rect 17328 34592 17356 34620
rect 18693 34595 18751 34601
rect 18693 34592 18705 34595
rect 17328 34564 18705 34592
rect 18693 34561 18705 34564
rect 18739 34561 18751 34595
rect 18693 34555 18751 34561
rect 20438 34552 20444 34604
rect 20496 34592 20502 34604
rect 20533 34595 20591 34601
rect 20533 34592 20545 34595
rect 20496 34564 20545 34592
rect 20496 34552 20502 34564
rect 20533 34561 20545 34564
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 22281 34595 22339 34601
rect 22281 34561 22293 34595
rect 22327 34592 22339 34595
rect 22649 34595 22707 34601
rect 22649 34592 22661 34595
rect 22327 34564 22661 34592
rect 22327 34561 22339 34564
rect 22281 34555 22339 34561
rect 22649 34561 22661 34564
rect 22695 34561 22707 34595
rect 22649 34555 22707 34561
rect 23198 34552 23204 34604
rect 23256 34552 23262 34604
rect 23952 34592 23980 34688
rect 25593 34663 25651 34669
rect 25593 34629 25605 34663
rect 25639 34660 25651 34663
rect 26142 34660 26148 34672
rect 25639 34632 26148 34660
rect 25639 34629 25651 34632
rect 25593 34623 25651 34629
rect 26142 34620 26148 34632
rect 26200 34660 26206 34672
rect 26513 34663 26571 34669
rect 26513 34660 26525 34663
rect 26200 34632 26525 34660
rect 26200 34620 26206 34632
rect 26513 34629 26525 34632
rect 26559 34629 26571 34663
rect 26513 34623 26571 34629
rect 27706 34620 27712 34672
rect 27764 34620 27770 34672
rect 29270 34660 29276 34672
rect 28934 34632 29276 34660
rect 29270 34620 29276 34632
rect 29328 34620 29334 34672
rect 30116 34660 30144 34700
rect 29380 34632 30144 34660
rect 30377 34663 30435 34669
rect 24857 34595 24915 34601
rect 24857 34592 24869 34595
rect 23952 34564 24869 34592
rect 24857 34561 24869 34564
rect 24903 34561 24915 34595
rect 26421 34595 26479 34601
rect 26421 34592 26433 34595
rect 24857 34555 24915 34561
rect 25700 34564 26433 34592
rect 25700 34536 25728 34564
rect 26421 34561 26433 34564
rect 26467 34561 26479 34595
rect 26421 34555 26479 34561
rect 29178 34552 29184 34604
rect 29236 34592 29242 34604
rect 29380 34601 29408 34632
rect 30377 34629 30389 34663
rect 30423 34660 30435 34663
rect 30926 34660 30932 34672
rect 30423 34632 30932 34660
rect 30423 34629 30435 34632
rect 30377 34623 30435 34629
rect 30926 34620 30932 34632
rect 30984 34660 30990 34672
rect 31297 34663 31355 34669
rect 31297 34660 31309 34663
rect 30984 34632 31309 34660
rect 30984 34620 30990 34632
rect 31297 34629 31309 34632
rect 31343 34629 31355 34663
rect 31297 34623 31355 34629
rect 32674 34620 32680 34672
rect 32732 34620 32738 34672
rect 33980 34660 34008 34700
rect 34149 34697 34161 34731
rect 34195 34728 34207 34731
rect 34698 34728 34704 34740
rect 34195 34700 34704 34728
rect 34195 34697 34207 34700
rect 34149 34691 34207 34697
rect 34698 34688 34704 34700
rect 34756 34688 34762 34740
rect 38930 34728 38936 34740
rect 34808 34700 38936 34728
rect 34808 34660 34836 34700
rect 38930 34688 38936 34700
rect 38988 34688 38994 34740
rect 39117 34731 39175 34737
rect 39117 34697 39129 34731
rect 39163 34728 39175 34731
rect 39206 34728 39212 34740
rect 39163 34700 39212 34728
rect 39163 34697 39175 34700
rect 39117 34691 39175 34697
rect 39206 34688 39212 34700
rect 39264 34688 39270 34740
rect 40770 34688 40776 34740
rect 40828 34688 40834 34740
rect 40954 34688 40960 34740
rect 41012 34688 41018 34740
rect 41322 34688 41328 34740
rect 41380 34688 41386 34740
rect 41414 34688 41420 34740
rect 41472 34688 41478 34740
rect 36354 34660 36360 34672
rect 33980 34632 34836 34660
rect 36294 34646 36360 34660
rect 36280 34632 36360 34646
rect 29365 34595 29423 34601
rect 29365 34592 29377 34595
rect 29236 34564 29377 34592
rect 29236 34552 29242 34564
rect 29365 34561 29377 34564
rect 29411 34561 29423 34595
rect 29365 34555 29423 34561
rect 30469 34595 30527 34601
rect 30469 34561 30481 34595
rect 30515 34592 30527 34595
rect 31205 34595 31263 34601
rect 31205 34592 31217 34595
rect 30515 34564 31217 34592
rect 30515 34561 30527 34564
rect 30469 34555 30527 34561
rect 31205 34561 31217 34564
rect 31251 34592 31263 34595
rect 31570 34592 31576 34604
rect 31251 34564 31576 34592
rect 31251 34561 31263 34564
rect 31205 34555 31263 34561
rect 31570 34552 31576 34564
rect 31628 34552 31634 34604
rect 32398 34552 32404 34604
rect 32456 34552 32462 34604
rect 8205 34527 8263 34533
rect 8205 34524 8217 34527
rect 7616 34496 7696 34524
rect 7760 34496 8217 34524
rect 7616 34484 7622 34496
rect 6454 34456 6460 34468
rect 5276 34428 6460 34456
rect 6454 34416 6460 34428
rect 6512 34416 6518 34468
rect 7668 34465 7696 34496
rect 8205 34493 8217 34496
rect 8251 34493 8263 34527
rect 8205 34487 8263 34493
rect 8297 34527 8355 34533
rect 8297 34493 8309 34527
rect 8343 34524 8355 34527
rect 8343 34496 8377 34524
rect 8343 34493 8355 34496
rect 8297 34487 8355 34493
rect 7653 34459 7711 34465
rect 7653 34425 7665 34459
rect 7699 34425 7711 34459
rect 7653 34419 7711 34425
rect 7742 34416 7748 34468
rect 7800 34456 7806 34468
rect 8312 34456 8340 34487
rect 12986 34484 12992 34536
rect 13044 34484 13050 34536
rect 13170 34484 13176 34536
rect 13228 34484 13234 34536
rect 13449 34527 13507 34533
rect 13449 34493 13461 34527
rect 13495 34524 13507 34527
rect 13998 34524 14004 34536
rect 13495 34496 14004 34524
rect 13495 34493 13507 34496
rect 13449 34487 13507 34493
rect 13998 34484 14004 34496
rect 14056 34484 14062 34536
rect 15470 34484 15476 34536
rect 15528 34524 15534 34536
rect 15841 34527 15899 34533
rect 15841 34524 15853 34527
rect 15528 34496 15853 34524
rect 15528 34484 15534 34496
rect 15841 34493 15853 34496
rect 15887 34493 15899 34527
rect 15841 34487 15899 34493
rect 20809 34527 20867 34533
rect 20809 34493 20821 34527
rect 20855 34524 20867 34527
rect 22370 34524 22376 34536
rect 20855 34496 22376 34524
rect 20855 34493 20867 34496
rect 20809 34487 20867 34493
rect 22370 34484 22376 34496
rect 22428 34484 22434 34536
rect 23842 34484 23848 34536
rect 23900 34524 23906 34536
rect 23937 34527 23995 34533
rect 23937 34524 23949 34527
rect 23900 34496 23949 34524
rect 23900 34484 23906 34496
rect 23937 34493 23949 34496
rect 23983 34493 23995 34527
rect 23937 34487 23995 34493
rect 24026 34484 24032 34536
rect 24084 34484 24090 34536
rect 25682 34484 25688 34536
rect 25740 34484 25746 34536
rect 25777 34527 25835 34533
rect 25777 34493 25789 34527
rect 25823 34493 25835 34527
rect 25777 34487 25835 34493
rect 26605 34527 26663 34533
rect 26605 34493 26617 34527
rect 26651 34493 26663 34527
rect 26605 34487 26663 34493
rect 7800 34428 8616 34456
rect 7800 34416 7806 34428
rect 8588 34400 8616 34428
rect 23382 34416 23388 34468
rect 23440 34456 23446 34468
rect 25792 34456 25820 34487
rect 26620 34456 26648 34487
rect 27430 34484 27436 34536
rect 27488 34484 27494 34536
rect 30653 34527 30711 34533
rect 30653 34493 30665 34527
rect 30699 34493 30711 34527
rect 30653 34487 30711 34493
rect 31481 34527 31539 34533
rect 31481 34493 31493 34527
rect 31527 34493 31539 34527
rect 33796 34524 33824 34578
rect 34790 34552 34796 34604
rect 34848 34552 34854 34604
rect 33870 34524 33876 34536
rect 33796 34496 33876 34524
rect 31481 34487 31539 34493
rect 23440 34428 26648 34456
rect 29641 34459 29699 34465
rect 23440 34416 23446 34428
rect 29641 34425 29653 34459
rect 29687 34456 29699 34459
rect 30190 34456 30196 34468
rect 29687 34428 30196 34456
rect 29687 34425 29699 34428
rect 29641 34419 29699 34425
rect 30190 34416 30196 34428
rect 30248 34456 30254 34468
rect 30668 34456 30696 34487
rect 31496 34456 31524 34487
rect 33870 34484 33876 34496
rect 33928 34524 33934 34536
rect 36280 34524 36308 34632
rect 36354 34620 36360 34632
rect 36412 34620 36418 34672
rect 37645 34663 37703 34669
rect 37645 34629 37657 34663
rect 37691 34660 37703 34663
rect 37918 34660 37924 34672
rect 37691 34632 37924 34660
rect 37691 34629 37703 34632
rect 37645 34623 37703 34629
rect 37918 34620 37924 34632
rect 37976 34620 37982 34672
rect 41340 34660 41368 34688
rect 39408 34632 41368 34660
rect 38746 34552 38752 34604
rect 38804 34552 38810 34604
rect 39408 34601 39436 34632
rect 41506 34620 41512 34672
rect 41564 34620 41570 34672
rect 39393 34595 39451 34601
rect 39393 34561 39405 34595
rect 39439 34561 39451 34595
rect 39393 34555 39451 34561
rect 39660 34595 39718 34601
rect 39660 34561 39672 34595
rect 39706 34592 39718 34595
rect 39942 34592 39948 34604
rect 39706 34564 39948 34592
rect 39706 34561 39718 34564
rect 39660 34555 39718 34561
rect 39942 34552 39948 34564
rect 40000 34552 40006 34604
rect 40402 34552 40408 34604
rect 40460 34592 40466 34604
rect 41325 34595 41383 34601
rect 41325 34592 41337 34595
rect 40460 34564 41337 34592
rect 40460 34552 40466 34564
rect 41325 34561 41337 34564
rect 41371 34592 41383 34595
rect 41524 34592 41552 34620
rect 41966 34592 41972 34604
rect 41371 34564 41972 34592
rect 41371 34561 41383 34564
rect 41325 34555 41383 34561
rect 41966 34552 41972 34564
rect 42024 34552 42030 34604
rect 33928 34496 36308 34524
rect 33928 34484 33934 34496
rect 36446 34484 36452 34536
rect 36504 34524 36510 34536
rect 36541 34527 36599 34533
rect 36541 34524 36553 34527
rect 36504 34496 36553 34524
rect 36504 34484 36510 34496
rect 36541 34493 36553 34496
rect 36587 34493 36599 34527
rect 36541 34487 36599 34493
rect 37366 34484 37372 34536
rect 37424 34484 37430 34536
rect 41138 34484 41144 34536
rect 41196 34524 41202 34536
rect 41509 34527 41567 34533
rect 41509 34524 41521 34527
rect 41196 34496 41521 34524
rect 41196 34484 41202 34496
rect 41509 34493 41521 34496
rect 41555 34493 41567 34527
rect 41509 34487 41567 34493
rect 31938 34456 31944 34468
rect 30248 34428 31944 34456
rect 30248 34416 30254 34428
rect 31938 34416 31944 34428
rect 31996 34456 32002 34468
rect 32122 34456 32128 34468
rect 31996 34428 32128 34456
rect 31996 34416 32002 34428
rect 32122 34416 32128 34428
rect 32180 34416 32186 34468
rect 5902 34348 5908 34400
rect 5960 34388 5966 34400
rect 6181 34391 6239 34397
rect 6181 34388 6193 34391
rect 5960 34360 6193 34388
rect 5960 34348 5966 34360
rect 6181 34357 6193 34360
rect 6227 34357 6239 34391
rect 6181 34351 6239 34357
rect 6362 34348 6368 34400
rect 6420 34388 6426 34400
rect 8110 34388 8116 34400
rect 6420 34360 8116 34388
rect 6420 34348 6426 34360
rect 8110 34348 8116 34360
rect 8168 34348 8174 34400
rect 8386 34348 8392 34400
rect 8444 34348 8450 34400
rect 8570 34348 8576 34400
rect 8628 34348 8634 34400
rect 15473 34391 15531 34397
rect 15473 34357 15485 34391
rect 15519 34388 15531 34391
rect 15654 34388 15660 34400
rect 15519 34360 15660 34388
rect 15519 34357 15531 34360
rect 15473 34351 15531 34357
rect 15654 34348 15660 34360
rect 15712 34388 15718 34400
rect 16022 34388 16028 34400
rect 15712 34360 16028 34388
rect 15712 34348 15718 34360
rect 16022 34348 16028 34360
rect 16080 34348 16086 34400
rect 21174 34348 21180 34400
rect 21232 34388 21238 34400
rect 21821 34391 21879 34397
rect 21821 34388 21833 34391
rect 21232 34360 21833 34388
rect 21232 34348 21238 34360
rect 21821 34357 21833 34360
rect 21867 34357 21879 34391
rect 21821 34351 21879 34357
rect 24302 34348 24308 34400
rect 24360 34348 24366 34400
rect 30834 34348 30840 34400
rect 30892 34348 30898 34400
rect 34790 34348 34796 34400
rect 34848 34388 34854 34400
rect 35050 34391 35108 34397
rect 35050 34388 35062 34391
rect 34848 34360 35062 34388
rect 34848 34348 34854 34360
rect 35050 34357 35062 34360
rect 35096 34357 35108 34391
rect 35050 34351 35108 34357
rect 1104 34298 42504 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 42504 34298
rect 1104 34224 42504 34246
rect 5258 34144 5264 34196
rect 5316 34144 5322 34196
rect 7926 34144 7932 34196
rect 7984 34184 7990 34196
rect 8021 34187 8079 34193
rect 8021 34184 8033 34187
rect 7984 34156 8033 34184
rect 7984 34144 7990 34156
rect 8021 34153 8033 34156
rect 8067 34153 8079 34187
rect 8021 34147 8079 34153
rect 8110 34144 8116 34196
rect 8168 34184 8174 34196
rect 9677 34187 9735 34193
rect 9677 34184 9689 34187
rect 8168 34156 9689 34184
rect 8168 34144 8174 34156
rect 9677 34153 9689 34156
rect 9723 34153 9735 34187
rect 9677 34147 9735 34153
rect 12986 34144 12992 34196
rect 13044 34184 13050 34196
rect 13173 34187 13231 34193
rect 13173 34184 13185 34187
rect 13044 34156 13185 34184
rect 13044 34144 13050 34156
rect 13173 34153 13185 34156
rect 13219 34153 13231 34187
rect 13173 34147 13231 34153
rect 14185 34187 14243 34193
rect 14185 34153 14197 34187
rect 14231 34184 14243 34187
rect 14274 34184 14280 34196
rect 14231 34156 14280 34184
rect 14231 34153 14243 34156
rect 14185 34147 14243 34153
rect 14274 34144 14280 34156
rect 14332 34144 14338 34196
rect 14918 34144 14924 34196
rect 14976 34144 14982 34196
rect 17862 34144 17868 34196
rect 17920 34184 17926 34196
rect 17920 34156 20944 34184
rect 17920 34144 17926 34156
rect 6638 34116 6644 34128
rect 6380 34088 6644 34116
rect 5445 34051 5503 34057
rect 5445 34017 5457 34051
rect 5491 34048 5503 34051
rect 5718 34048 5724 34060
rect 5491 34020 5724 34048
rect 5491 34017 5503 34020
rect 5445 34011 5503 34017
rect 5718 34008 5724 34020
rect 5776 34008 5782 34060
rect 5810 34008 5816 34060
rect 5868 34008 5874 34060
rect 5902 34008 5908 34060
rect 5960 34008 5966 34060
rect 5534 33940 5540 33992
rect 5592 33940 5598 33992
rect 5997 33983 6055 33989
rect 5997 33949 6009 33983
rect 6043 33949 6055 33983
rect 5997 33943 6055 33949
rect 6273 33983 6331 33989
rect 6273 33949 6285 33983
rect 6319 33980 6331 33983
rect 6380 33980 6408 34088
rect 6638 34076 6644 34088
rect 6696 34116 6702 34128
rect 17954 34116 17960 34128
rect 6696 34088 9996 34116
rect 6696 34076 6702 34088
rect 7650 34048 7656 34060
rect 7484 34020 7656 34048
rect 6319 33952 6408 33980
rect 6319 33949 6331 33952
rect 6273 33943 6331 33949
rect 6012 33912 6040 33943
rect 6454 33940 6460 33992
rect 6512 33940 6518 33992
rect 7282 33940 7288 33992
rect 7340 33940 7346 33992
rect 7374 33940 7380 33992
rect 7432 33980 7438 33992
rect 7484 33989 7512 34020
rect 7650 34008 7656 34020
rect 7708 34008 7714 34060
rect 7469 33983 7527 33989
rect 7469 33980 7481 33983
rect 7432 33952 7481 33980
rect 7432 33940 7438 33952
rect 7469 33949 7481 33952
rect 7515 33949 7527 33983
rect 7742 33980 7748 33992
rect 7469 33943 7527 33949
rect 7576 33952 7748 33980
rect 6362 33912 6368 33924
rect 6012 33884 6368 33912
rect 6362 33872 6368 33884
rect 6420 33872 6426 33924
rect 6914 33872 6920 33924
rect 6972 33912 6978 33924
rect 7576 33912 7604 33952
rect 7742 33940 7748 33952
rect 7800 33940 7806 33992
rect 7834 33940 7840 33992
rect 7892 33980 7898 33992
rect 8018 33980 8024 33992
rect 7892 33952 8024 33980
rect 7892 33940 7898 33952
rect 8018 33940 8024 33952
rect 8076 33940 8082 33992
rect 8389 33983 8447 33989
rect 8389 33949 8401 33983
rect 8435 33980 8447 33983
rect 8496 33980 8524 34088
rect 8435 33952 8524 33980
rect 8435 33949 8447 33952
rect 8389 33943 8447 33949
rect 8570 33940 8576 33992
rect 8628 33940 8634 33992
rect 9398 33940 9404 33992
rect 9456 33980 9462 33992
rect 9968 33989 9996 34088
rect 13096 34088 17960 34116
rect 10689 34051 10747 34057
rect 10689 34017 10701 34051
rect 10735 34048 10747 34051
rect 11606 34048 11612 34060
rect 10735 34020 11612 34048
rect 10735 34017 10747 34020
rect 10689 34011 10747 34017
rect 11606 34008 11612 34020
rect 11664 34008 11670 34060
rect 12618 34008 12624 34060
rect 12676 34048 12682 34060
rect 13096 34057 13124 34088
rect 17954 34076 17960 34088
rect 18012 34076 18018 34128
rect 13081 34051 13139 34057
rect 13081 34048 13093 34051
rect 12676 34020 13093 34048
rect 12676 34008 12682 34020
rect 13081 34017 13093 34020
rect 13127 34017 13139 34051
rect 13081 34011 13139 34017
rect 13906 34008 13912 34060
rect 13964 34048 13970 34060
rect 14369 34051 14427 34057
rect 14369 34048 14381 34051
rect 13964 34020 14381 34048
rect 13964 34008 13970 34020
rect 14369 34017 14381 34020
rect 14415 34017 14427 34051
rect 14369 34011 14427 34017
rect 15470 34008 15476 34060
rect 15528 34008 15534 34060
rect 19260 34057 19288 34156
rect 20916 34057 20944 34156
rect 22278 34144 22284 34196
rect 22336 34144 22342 34196
rect 23934 34144 23940 34196
rect 23992 34184 23998 34196
rect 24213 34187 24271 34193
rect 24213 34184 24225 34187
rect 23992 34156 24225 34184
rect 23992 34144 23998 34156
rect 24213 34153 24225 34156
rect 24259 34153 24271 34187
rect 27430 34184 27436 34196
rect 24213 34147 24271 34153
rect 24596 34156 27436 34184
rect 19245 34051 19303 34057
rect 15948 34020 19196 34048
rect 9493 33983 9551 33989
rect 9493 33980 9505 33983
rect 9456 33952 9505 33980
rect 9456 33940 9462 33952
rect 9493 33949 9505 33952
rect 9539 33949 9551 33983
rect 9493 33943 9551 33949
rect 9953 33983 10011 33989
rect 9953 33949 9965 33983
rect 9999 33949 10011 33983
rect 9953 33943 10011 33949
rect 10137 33983 10195 33989
rect 10137 33949 10149 33983
rect 10183 33949 10195 33983
rect 10137 33943 10195 33949
rect 6972 33884 7604 33912
rect 7653 33915 7711 33921
rect 6972 33872 6978 33884
rect 7653 33881 7665 33915
rect 7699 33881 7711 33915
rect 7653 33875 7711 33881
rect 6086 33804 6092 33856
rect 6144 33844 6150 33856
rect 6181 33847 6239 33853
rect 6181 33844 6193 33847
rect 6144 33816 6193 33844
rect 6144 33804 6150 33816
rect 6181 33813 6193 33816
rect 6227 33813 6239 33847
rect 7668 33844 7696 33875
rect 7926 33872 7932 33924
rect 7984 33912 7990 33924
rect 8941 33915 8999 33921
rect 8941 33912 8953 33915
rect 7984 33884 8953 33912
rect 7984 33872 7990 33884
rect 8941 33881 8953 33884
rect 8987 33881 8999 33915
rect 9508 33912 9536 33943
rect 10152 33912 10180 33943
rect 13814 33940 13820 33992
rect 13872 33980 13878 33992
rect 14461 33983 14519 33989
rect 14461 33980 14473 33983
rect 13872 33952 14473 33980
rect 13872 33940 13878 33952
rect 14461 33949 14473 33952
rect 14507 33949 14519 33983
rect 14461 33943 14519 33949
rect 15102 33940 15108 33992
rect 15160 33980 15166 33992
rect 15749 33983 15807 33989
rect 15749 33980 15761 33983
rect 15160 33952 15761 33980
rect 15160 33940 15166 33952
rect 15749 33949 15761 33952
rect 15795 33949 15807 33983
rect 15948 33980 15976 34020
rect 15749 33943 15807 33949
rect 15856 33952 15976 33980
rect 9508 33884 10180 33912
rect 11333 33915 11391 33921
rect 8941 33875 8999 33881
rect 11333 33881 11345 33915
rect 11379 33912 11391 33915
rect 15856 33912 15884 33952
rect 16022 33940 16028 33992
rect 16080 33980 16086 33992
rect 17037 33983 17095 33989
rect 17037 33980 17049 33983
rect 16080 33952 17049 33980
rect 16080 33940 16086 33952
rect 17037 33949 17049 33952
rect 17083 33949 17095 33983
rect 17037 33943 17095 33949
rect 17310 33940 17316 33992
rect 17368 33980 17374 33992
rect 17862 33980 17868 33992
rect 17368 33952 17868 33980
rect 17368 33940 17374 33952
rect 17862 33940 17868 33952
rect 17920 33980 17926 33992
rect 17957 33983 18015 33989
rect 17957 33980 17969 33983
rect 17920 33952 17969 33980
rect 17920 33940 17926 33952
rect 17957 33949 17969 33952
rect 18003 33949 18015 33983
rect 17957 33943 18015 33949
rect 18506 33940 18512 33992
rect 18564 33940 18570 33992
rect 19168 33980 19196 34020
rect 19245 34017 19257 34051
rect 19291 34017 19303 34051
rect 19245 34011 19303 34017
rect 20901 34051 20959 34057
rect 20901 34017 20913 34051
rect 20947 34017 20959 34051
rect 20901 34011 20959 34017
rect 22830 34008 22836 34060
rect 22888 34008 22894 34060
rect 24596 34057 24624 34156
rect 27430 34144 27436 34156
rect 27488 34144 27494 34196
rect 27614 34144 27620 34196
rect 27672 34184 27678 34196
rect 27801 34187 27859 34193
rect 27801 34184 27813 34187
rect 27672 34156 27813 34184
rect 27672 34144 27678 34156
rect 27801 34153 27813 34156
rect 27847 34153 27859 34187
rect 27801 34147 27859 34153
rect 28629 34187 28687 34193
rect 28629 34153 28641 34187
rect 28675 34184 28687 34187
rect 28718 34184 28724 34196
rect 28675 34156 28724 34184
rect 28675 34153 28687 34156
rect 28629 34147 28687 34153
rect 28718 34144 28724 34156
rect 28776 34144 28782 34196
rect 29454 34144 29460 34196
rect 29512 34184 29518 34196
rect 29549 34187 29607 34193
rect 29549 34184 29561 34187
rect 29512 34156 29561 34184
rect 29512 34144 29518 34156
rect 29549 34153 29561 34156
rect 29595 34153 29607 34187
rect 29549 34147 29607 34153
rect 31478 34144 31484 34196
rect 31536 34144 31542 34196
rect 34149 34187 34207 34193
rect 34149 34153 34161 34187
rect 34195 34184 34207 34187
rect 34238 34184 34244 34196
rect 34195 34156 34244 34184
rect 34195 34153 34207 34156
rect 34149 34147 34207 34153
rect 34238 34144 34244 34156
rect 34296 34144 34302 34196
rect 34790 34144 34796 34196
rect 34848 34184 34854 34196
rect 34977 34187 35035 34193
rect 34977 34184 34989 34187
rect 34848 34156 34989 34184
rect 34848 34144 34854 34156
rect 34977 34153 34989 34156
rect 35023 34153 35035 34187
rect 34977 34147 35035 34153
rect 35986 34144 35992 34196
rect 36044 34184 36050 34196
rect 36633 34187 36691 34193
rect 36633 34184 36645 34187
rect 36044 34156 36645 34184
rect 36044 34144 36050 34156
rect 36633 34153 36645 34156
rect 36679 34153 36691 34187
rect 36633 34147 36691 34153
rect 38197 34187 38255 34193
rect 38197 34153 38209 34187
rect 38243 34184 38255 34187
rect 38378 34184 38384 34196
rect 38243 34156 38384 34184
rect 38243 34153 38255 34156
rect 38197 34147 38255 34153
rect 38378 34144 38384 34156
rect 38436 34144 38442 34196
rect 40770 34184 40776 34196
rect 40512 34156 40776 34184
rect 25682 34076 25688 34128
rect 25740 34116 25746 34128
rect 25961 34119 26019 34125
rect 25961 34116 25973 34119
rect 25740 34088 25973 34116
rect 25740 34076 25746 34088
rect 25961 34085 25973 34088
rect 26007 34116 26019 34119
rect 26007 34088 26648 34116
rect 26007 34085 26019 34088
rect 25961 34079 26019 34085
rect 26620 34057 26648 34088
rect 26970 34076 26976 34128
rect 27028 34076 27034 34128
rect 36814 34116 36820 34128
rect 36356 34088 36820 34116
rect 24581 34051 24639 34057
rect 24581 34017 24593 34051
rect 24627 34017 24639 34051
rect 26605 34051 26663 34057
rect 24581 34011 24639 34017
rect 25608 34020 26004 34048
rect 21174 33989 21180 33992
rect 21168 33980 21180 33989
rect 19168 33952 20392 33980
rect 21135 33952 21180 33980
rect 16485 33915 16543 33921
rect 16485 33912 16497 33915
rect 11379 33884 15884 33912
rect 15948 33884 16497 33912
rect 11379 33881 11391 33884
rect 11333 33875 11391 33881
rect 8297 33847 8355 33853
rect 8297 33844 8309 33847
rect 7668 33816 8309 33844
rect 6181 33807 6239 33813
rect 8297 33813 8309 33816
rect 8343 33813 8355 33847
rect 8297 33807 8355 33813
rect 8478 33804 8484 33856
rect 8536 33844 8542 33856
rect 9861 33847 9919 33853
rect 9861 33844 9873 33847
rect 8536 33816 9873 33844
rect 8536 33804 8542 33816
rect 9861 33813 9873 33816
rect 9907 33813 9919 33847
rect 9861 33807 9919 33813
rect 11146 33804 11152 33856
rect 11204 33844 11210 33856
rect 11241 33847 11299 33853
rect 11241 33844 11253 33847
rect 11204 33816 11253 33844
rect 11204 33804 11210 33816
rect 11241 33813 11253 33816
rect 11287 33813 11299 33847
rect 11241 33807 11299 33813
rect 15286 33804 15292 33856
rect 15344 33804 15350 33856
rect 15381 33847 15439 33853
rect 15381 33813 15393 33847
rect 15427 33844 15439 33847
rect 15948 33844 15976 33884
rect 16485 33881 16497 33884
rect 16531 33881 16543 33915
rect 16485 33875 16543 33881
rect 17221 33915 17279 33921
rect 17221 33881 17233 33915
rect 17267 33881 17279 33915
rect 17221 33875 17279 33881
rect 19061 33915 19119 33921
rect 19061 33881 19073 33915
rect 19107 33912 19119 33915
rect 19490 33915 19548 33921
rect 19490 33912 19502 33915
rect 19107 33884 19502 33912
rect 19107 33881 19119 33884
rect 19061 33875 19119 33881
rect 19490 33881 19502 33884
rect 19536 33881 19548 33915
rect 20364 33912 20392 33952
rect 21168 33943 21180 33952
rect 21174 33940 21180 33943
rect 21232 33940 21238 33992
rect 25608 33980 25636 34020
rect 22066 33952 25636 33980
rect 22066 33912 22094 33952
rect 23216 33924 23244 33952
rect 23106 33921 23112 33924
rect 20364 33884 22094 33912
rect 19490 33875 19548 33881
rect 23100 33875 23112 33921
rect 15427 33816 15976 33844
rect 15427 33813 15439 33816
rect 15381 33807 15439 33813
rect 16114 33804 16120 33856
rect 16172 33844 16178 33856
rect 16393 33847 16451 33853
rect 16393 33844 16405 33847
rect 16172 33816 16405 33844
rect 16172 33804 16178 33816
rect 16393 33813 16405 33816
rect 16439 33813 16451 33847
rect 17236 33844 17264 33875
rect 23106 33872 23112 33875
rect 23164 33872 23170 33924
rect 23198 33872 23204 33924
rect 23256 33872 23262 33924
rect 24848 33915 24906 33921
rect 24848 33881 24860 33915
rect 24894 33912 24906 33915
rect 25038 33912 25044 33924
rect 24894 33884 25044 33912
rect 24894 33881 24906 33884
rect 24848 33875 24906 33881
rect 25038 33872 25044 33884
rect 25096 33872 25102 33924
rect 25976 33912 26004 34020
rect 26605 34017 26617 34051
rect 26651 34017 26663 34051
rect 26605 34011 26663 34017
rect 27522 34008 27528 34060
rect 27580 34048 27586 34060
rect 28353 34051 28411 34057
rect 28353 34048 28365 34051
rect 27580 34020 28365 34048
rect 27580 34008 27586 34020
rect 28353 34017 28365 34020
rect 28399 34048 28411 34051
rect 29178 34048 29184 34060
rect 28399 34020 29184 34048
rect 28399 34017 28411 34020
rect 28353 34011 28411 34017
rect 29178 34008 29184 34020
rect 29236 34008 29242 34060
rect 29273 34051 29331 34057
rect 29273 34017 29285 34051
rect 29319 34048 29331 34051
rect 30190 34048 30196 34060
rect 29319 34020 30196 34048
rect 29319 34017 29331 34020
rect 29273 34011 29331 34017
rect 30190 34008 30196 34020
rect 30248 34008 30254 34060
rect 31754 34008 31760 34060
rect 31812 34048 31818 34060
rect 31941 34051 31999 34057
rect 31941 34048 31953 34051
rect 31812 34020 31953 34048
rect 31812 34008 31818 34020
rect 31941 34017 31953 34020
rect 31987 34017 31999 34051
rect 31941 34011 31999 34017
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33980 27399 33983
rect 28626 33980 28632 33992
rect 27387 33952 28632 33980
rect 27387 33949 27399 33952
rect 27341 33943 27399 33949
rect 28626 33940 28632 33952
rect 28684 33940 28690 33992
rect 28997 33983 29055 33989
rect 28997 33949 29009 33983
rect 29043 33980 29055 33983
rect 30006 33980 30012 33992
rect 29043 33952 30012 33980
rect 29043 33949 29055 33952
rect 28997 33943 29055 33949
rect 30006 33940 30012 33952
rect 30064 33940 30070 33992
rect 31956 33980 31984 34011
rect 32122 34008 32128 34060
rect 32180 34048 32186 34060
rect 33597 34051 33655 34057
rect 33597 34048 33609 34051
rect 32180 34020 33609 34048
rect 32180 34008 32186 34020
rect 33597 34017 33609 34020
rect 33643 34017 33655 34051
rect 33597 34011 33655 34017
rect 35621 34051 35679 34057
rect 35621 34017 35633 34051
rect 35667 34048 35679 34051
rect 36078 34048 36084 34060
rect 35667 34020 36084 34048
rect 35667 34017 35679 34020
rect 35621 34011 35679 34017
rect 32306 33980 32312 33992
rect 31956 33952 32312 33980
rect 32306 33940 32312 33952
rect 32364 33980 32370 33992
rect 32401 33983 32459 33989
rect 32401 33980 32413 33983
rect 32364 33952 32413 33980
rect 32364 33940 32370 33952
rect 32401 33949 32413 33952
rect 32447 33949 32459 33983
rect 32401 33943 32459 33949
rect 32214 33912 32220 33924
rect 25976 33884 32220 33912
rect 32214 33872 32220 33884
rect 32272 33872 32278 33924
rect 33612 33912 33640 34011
rect 36078 34008 36084 34020
rect 36136 34008 36142 34060
rect 33689 33983 33747 33989
rect 33689 33949 33701 33983
rect 33735 33980 33747 33983
rect 33778 33980 33784 33992
rect 33735 33952 33784 33980
rect 33735 33949 33747 33952
rect 33689 33943 33747 33949
rect 33778 33940 33784 33952
rect 33836 33940 33842 33992
rect 35345 33983 35403 33989
rect 35345 33949 35357 33983
rect 35391 33980 35403 33983
rect 36356 33980 36384 34088
rect 36814 34076 36820 34088
rect 36872 34076 36878 34128
rect 36449 34051 36507 34057
rect 36449 34017 36461 34051
rect 36495 34048 36507 34051
rect 37185 34051 37243 34057
rect 37185 34048 37197 34051
rect 36495 34020 37197 34048
rect 36495 34017 36507 34020
rect 36449 34011 36507 34017
rect 37185 34017 37197 34020
rect 37231 34017 37243 34051
rect 37185 34011 37243 34017
rect 38841 34051 38899 34057
rect 38841 34017 38853 34051
rect 38887 34017 38899 34051
rect 38841 34011 38899 34017
rect 39117 34051 39175 34057
rect 39117 34017 39129 34051
rect 39163 34048 39175 34051
rect 40402 34048 40408 34060
rect 39163 34020 40408 34048
rect 39163 34017 39175 34020
rect 39117 34011 39175 34017
rect 35391 33952 36384 33980
rect 35391 33949 35403 33952
rect 35345 33943 35403 33949
rect 33962 33912 33968 33924
rect 33612 33884 33968 33912
rect 33962 33872 33968 33884
rect 34020 33912 34026 33924
rect 36464 33912 36492 34011
rect 38856 33980 38884 34011
rect 40402 34008 40408 34020
rect 40460 34008 40466 34060
rect 40512 34057 40540 34156
rect 40770 34144 40776 34156
rect 40828 34144 40834 34196
rect 41966 34144 41972 34196
rect 42024 34144 42030 34196
rect 40497 34051 40555 34057
rect 40497 34017 40509 34051
rect 40543 34017 40555 34051
rect 40497 34011 40555 34017
rect 40034 33980 40040 33992
rect 38856 33952 40040 33980
rect 40034 33940 40040 33952
rect 40092 33940 40098 33992
rect 40589 33983 40647 33989
rect 40589 33949 40601 33983
rect 40635 33980 40647 33983
rect 41322 33980 41328 33992
rect 40635 33952 41328 33980
rect 40635 33949 40647 33952
rect 40589 33943 40647 33949
rect 41322 33940 41328 33952
rect 41380 33940 41386 33992
rect 37001 33915 37059 33921
rect 37001 33912 37013 33915
rect 34020 33884 36492 33912
rect 36556 33884 37013 33912
rect 34020 33872 34026 33884
rect 17954 33844 17960 33856
rect 17236 33816 17960 33844
rect 16393 33807 16451 33813
rect 17954 33804 17960 33816
rect 18012 33844 18018 33856
rect 18138 33844 18144 33856
rect 18012 33816 18144 33844
rect 18012 33804 18018 33816
rect 18138 33804 18144 33816
rect 18196 33804 18202 33856
rect 20622 33804 20628 33856
rect 20680 33804 20686 33856
rect 22738 33804 22744 33856
rect 22796 33844 22802 33856
rect 23382 33844 23388 33856
rect 22796 33816 23388 33844
rect 22796 33804 22802 33816
rect 23382 33804 23388 33816
rect 23440 33804 23446 33856
rect 26050 33804 26056 33856
rect 26108 33804 26114 33856
rect 27433 33847 27491 33853
rect 27433 33813 27445 33847
rect 27479 33844 27491 33847
rect 28166 33844 28172 33856
rect 27479 33816 28172 33844
rect 27479 33813 27491 33816
rect 27433 33807 27491 33813
rect 28166 33804 28172 33816
rect 28224 33804 28230 33856
rect 28261 33847 28319 33853
rect 28261 33813 28273 33847
rect 28307 33844 28319 33847
rect 28626 33844 28632 33856
rect 28307 33816 28632 33844
rect 28307 33813 28319 33816
rect 28261 33807 28319 33813
rect 28626 33804 28632 33816
rect 28684 33804 28690 33856
rect 29089 33847 29147 33853
rect 29089 33813 29101 33847
rect 29135 33844 29147 33847
rect 29914 33844 29920 33856
rect 29135 33816 29920 33844
rect 29135 33813 29147 33816
rect 29089 33807 29147 33813
rect 29914 33804 29920 33816
rect 29972 33804 29978 33856
rect 30006 33804 30012 33856
rect 30064 33804 30070 33856
rect 31849 33847 31907 33853
rect 31849 33813 31861 33847
rect 31895 33844 31907 33847
rect 32030 33844 32036 33856
rect 31895 33816 32036 33844
rect 31895 33813 31907 33816
rect 31849 33807 31907 33813
rect 32030 33804 32036 33816
rect 32088 33804 32094 33856
rect 32582 33804 32588 33856
rect 32640 33844 32646 33856
rect 33045 33847 33103 33853
rect 33045 33844 33057 33847
rect 32640 33816 33057 33844
rect 32640 33804 32646 33816
rect 33045 33813 33057 33816
rect 33091 33813 33103 33847
rect 33045 33807 33103 33813
rect 33781 33847 33839 33853
rect 33781 33813 33793 33847
rect 33827 33844 33839 33847
rect 34054 33844 34060 33856
rect 33827 33816 34060 33844
rect 33827 33813 33839 33816
rect 33781 33807 33839 33813
rect 34054 33804 34060 33816
rect 34112 33804 34118 33856
rect 35437 33847 35495 33853
rect 35437 33813 35449 33847
rect 35483 33844 35495 33847
rect 35805 33847 35863 33853
rect 35805 33844 35817 33847
rect 35483 33816 35817 33844
rect 35483 33813 35495 33816
rect 35437 33807 35495 33813
rect 35805 33813 35817 33816
rect 35851 33813 35863 33847
rect 35805 33807 35863 33813
rect 36170 33804 36176 33856
rect 36228 33804 36234 33856
rect 36265 33847 36323 33853
rect 36265 33813 36277 33847
rect 36311 33844 36323 33847
rect 36446 33844 36452 33856
rect 36311 33816 36452 33844
rect 36311 33813 36323 33816
rect 36265 33807 36323 33813
rect 36446 33804 36452 33816
rect 36504 33844 36510 33856
rect 36556 33844 36584 33884
rect 37001 33881 37013 33884
rect 37047 33881 37059 33915
rect 37001 33875 37059 33881
rect 38565 33915 38623 33921
rect 38565 33881 38577 33915
rect 38611 33912 38623 33915
rect 38930 33912 38936 33924
rect 38611 33884 38936 33912
rect 38611 33881 38623 33884
rect 38565 33875 38623 33881
rect 38930 33872 38936 33884
rect 38988 33912 38994 33924
rect 39574 33912 39580 33924
rect 38988 33884 39580 33912
rect 38988 33872 38994 33884
rect 39574 33872 39580 33884
rect 39632 33872 39638 33924
rect 40862 33921 40868 33924
rect 40856 33875 40868 33921
rect 40862 33872 40868 33875
rect 40920 33872 40926 33924
rect 36504 33816 36584 33844
rect 36504 33804 36510 33816
rect 36814 33804 36820 33856
rect 36872 33844 36878 33856
rect 37093 33847 37151 33853
rect 37093 33844 37105 33847
rect 36872 33816 37105 33844
rect 36872 33804 36878 33816
rect 37093 33813 37105 33816
rect 37139 33813 37151 33847
rect 37093 33807 37151 33813
rect 38654 33804 38660 33856
rect 38712 33804 38718 33856
rect 39666 33804 39672 33856
rect 39724 33804 39730 33856
rect 39853 33847 39911 33853
rect 39853 33813 39865 33847
rect 39899 33844 39911 33847
rect 40402 33844 40408 33856
rect 39899 33816 40408 33844
rect 39899 33813 39911 33816
rect 39853 33807 39911 33813
rect 40402 33804 40408 33816
rect 40460 33804 40466 33856
rect 1104 33754 42504 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 42504 33754
rect 1104 33680 42504 33702
rect 1670 33640 1676 33652
rect 1504 33612 1676 33640
rect 1504 33572 1532 33612
rect 1670 33600 1676 33612
rect 1728 33640 1734 33652
rect 2682 33640 2688 33652
rect 1728 33612 2688 33640
rect 1728 33600 1734 33612
rect 2682 33600 2688 33612
rect 2740 33600 2746 33652
rect 3510 33600 3516 33652
rect 3568 33640 3574 33652
rect 4798 33640 4804 33652
rect 3568 33612 4804 33640
rect 3568 33600 3574 33612
rect 4798 33600 4804 33612
rect 4856 33640 4862 33652
rect 5261 33643 5319 33649
rect 5261 33640 5273 33643
rect 4856 33612 5273 33640
rect 4856 33600 4862 33612
rect 5261 33609 5273 33612
rect 5307 33609 5319 33643
rect 5261 33603 5319 33609
rect 5718 33600 5724 33652
rect 5776 33640 5782 33652
rect 6365 33643 6423 33649
rect 6365 33640 6377 33643
rect 5776 33612 6377 33640
rect 5776 33600 5782 33612
rect 6365 33609 6377 33612
rect 6411 33640 6423 33643
rect 6730 33640 6736 33652
rect 6411 33612 6736 33640
rect 6411 33609 6423 33612
rect 6365 33603 6423 33609
rect 6730 33600 6736 33612
rect 6788 33640 6794 33652
rect 6788 33612 7052 33640
rect 6788 33600 6794 33612
rect 1412 33544 1532 33572
rect 1412 33513 1440 33544
rect 3602 33532 3608 33584
rect 3660 33572 3666 33584
rect 3973 33575 4031 33581
rect 3973 33572 3985 33575
rect 3660 33544 3985 33572
rect 3660 33532 3666 33544
rect 3973 33541 3985 33544
rect 4019 33541 4031 33575
rect 3973 33535 4031 33541
rect 6454 33532 6460 33584
rect 6512 33572 6518 33584
rect 7024 33572 7052 33612
rect 7098 33600 7104 33652
rect 7156 33640 7162 33652
rect 9398 33640 9404 33652
rect 7156 33612 9404 33640
rect 7156 33600 7162 33612
rect 9398 33600 9404 33612
rect 9456 33640 9462 33652
rect 9861 33643 9919 33649
rect 9861 33640 9873 33643
rect 9456 33612 9873 33640
rect 9456 33600 9462 33612
rect 9861 33609 9873 33612
rect 9907 33609 9919 33643
rect 9861 33603 9919 33609
rect 13357 33643 13415 33649
rect 13357 33609 13369 33643
rect 13403 33640 13415 33643
rect 13538 33640 13544 33652
rect 13403 33612 13544 33640
rect 13403 33609 13415 33612
rect 13357 33603 13415 33609
rect 13538 33600 13544 33612
rect 13596 33600 13602 33652
rect 14185 33643 14243 33649
rect 14185 33609 14197 33643
rect 14231 33640 14243 33643
rect 15102 33640 15108 33652
rect 14231 33612 15108 33640
rect 14231 33609 14243 33612
rect 14185 33603 14243 33609
rect 15102 33600 15108 33612
rect 15160 33600 15166 33652
rect 15657 33643 15715 33649
rect 15657 33609 15669 33643
rect 15703 33609 15715 33643
rect 15657 33603 15715 33609
rect 7834 33572 7840 33584
rect 6512 33544 6684 33572
rect 7024 33544 7840 33572
rect 6512 33532 6518 33544
rect 1397 33507 1455 33513
rect 1397 33473 1409 33507
rect 1443 33473 1455 33507
rect 1397 33467 1455 33473
rect 2774 33464 2780 33516
rect 2832 33464 2838 33516
rect 3421 33507 3479 33513
rect 3421 33473 3433 33507
rect 3467 33504 3479 33507
rect 3881 33507 3939 33513
rect 3881 33504 3893 33507
rect 3467 33476 3893 33504
rect 3467 33473 3479 33476
rect 3421 33467 3479 33473
rect 3881 33473 3893 33476
rect 3927 33504 3939 33507
rect 4062 33504 4068 33516
rect 3927 33476 4068 33504
rect 3927 33473 3939 33476
rect 3881 33467 3939 33473
rect 4062 33464 4068 33476
rect 4120 33464 4126 33516
rect 4157 33507 4215 33513
rect 4157 33473 4169 33507
rect 4203 33504 4215 33507
rect 4798 33504 4804 33516
rect 4203 33476 4804 33504
rect 4203 33473 4215 33476
rect 4157 33467 4215 33473
rect 4798 33464 4804 33476
rect 4856 33464 4862 33516
rect 5077 33507 5135 33513
rect 5077 33473 5089 33507
rect 5123 33504 5135 33507
rect 5442 33504 5448 33516
rect 5123 33476 5448 33504
rect 5123 33473 5135 33476
rect 5077 33467 5135 33473
rect 5442 33464 5448 33476
rect 5500 33464 5506 33516
rect 5626 33464 5632 33516
rect 5684 33504 5690 33516
rect 6656 33513 6684 33544
rect 7834 33532 7840 33544
rect 7892 33532 7898 33584
rect 8021 33575 8079 33581
rect 8021 33541 8033 33575
rect 8067 33572 8079 33575
rect 8389 33575 8447 33581
rect 8389 33572 8401 33575
rect 8067 33544 8401 33572
rect 8067 33541 8079 33544
rect 8021 33535 8079 33541
rect 8389 33541 8401 33544
rect 8435 33541 8447 33575
rect 8389 33535 8447 33541
rect 9122 33532 9128 33584
rect 9180 33532 9186 33584
rect 6549 33507 6607 33513
rect 6549 33504 6561 33507
rect 5684 33476 6561 33504
rect 5684 33464 5690 33476
rect 6549 33473 6561 33476
rect 6595 33473 6607 33507
rect 6549 33467 6607 33473
rect 6641 33507 6699 33513
rect 6641 33473 6653 33507
rect 6687 33504 6699 33507
rect 7009 33507 7067 33513
rect 7009 33504 7021 33507
rect 6687 33476 7021 33504
rect 6687 33473 6699 33476
rect 6641 33467 6699 33473
rect 7009 33473 7021 33476
rect 7055 33473 7067 33507
rect 7009 33467 7067 33473
rect 7190 33464 7196 33516
rect 7248 33504 7254 33516
rect 7285 33507 7343 33513
rect 7285 33504 7297 33507
rect 7248 33476 7297 33504
rect 7248 33464 7254 33476
rect 7285 33473 7297 33476
rect 7331 33473 7343 33507
rect 7285 33467 7343 33473
rect 7745 33507 7803 33513
rect 7745 33473 7757 33507
rect 7791 33504 7803 33507
rect 7926 33504 7932 33516
rect 7791 33476 7932 33504
rect 7791 33473 7803 33476
rect 7745 33467 7803 33473
rect 7926 33464 7932 33476
rect 7984 33464 7990 33516
rect 10226 33513 10232 33516
rect 10220 33467 10232 33513
rect 10226 33464 10232 33467
rect 10284 33464 10290 33516
rect 11514 33464 11520 33516
rect 11572 33504 11578 33516
rect 11977 33507 12035 33513
rect 11977 33504 11989 33507
rect 11572 33476 11989 33504
rect 11572 33464 11578 33476
rect 11977 33473 11989 33476
rect 12023 33473 12035 33507
rect 11977 33467 12035 33473
rect 12244 33507 12302 33513
rect 12244 33473 12256 33507
rect 12290 33504 12302 33507
rect 12802 33504 12808 33516
rect 12290 33476 12808 33504
rect 12290 33473 12302 33476
rect 12244 33467 12302 33473
rect 12802 33464 12808 33476
rect 12860 33464 12866 33516
rect 13556 33504 13584 33600
rect 15320 33575 15378 33581
rect 15320 33541 15332 33575
rect 15366 33572 15378 33575
rect 15672 33572 15700 33603
rect 16114 33600 16120 33652
rect 16172 33600 16178 33652
rect 16942 33600 16948 33652
rect 17000 33640 17006 33652
rect 17129 33643 17187 33649
rect 17129 33640 17141 33643
rect 17000 33612 17141 33640
rect 17000 33600 17006 33612
rect 17129 33609 17141 33612
rect 17175 33609 17187 33643
rect 17129 33603 17187 33609
rect 17586 33600 17592 33652
rect 17644 33600 17650 33652
rect 18506 33600 18512 33652
rect 18564 33640 18570 33652
rect 19981 33643 20039 33649
rect 19981 33640 19993 33643
rect 18564 33612 19993 33640
rect 18564 33600 18570 33612
rect 19981 33609 19993 33612
rect 20027 33609 20039 33643
rect 19981 33603 20039 33609
rect 23106 33600 23112 33652
rect 23164 33640 23170 33652
rect 23385 33643 23443 33649
rect 23385 33640 23397 33643
rect 23164 33612 23397 33640
rect 23164 33600 23170 33612
rect 23385 33609 23397 33612
rect 23431 33609 23443 33643
rect 23385 33603 23443 33609
rect 23845 33643 23903 33649
rect 23845 33609 23857 33643
rect 23891 33640 23903 33643
rect 24302 33640 24308 33652
rect 23891 33612 24308 33640
rect 23891 33609 23903 33612
rect 23845 33603 23903 33609
rect 24302 33600 24308 33612
rect 24360 33600 24366 33652
rect 25038 33600 25044 33652
rect 25096 33600 25102 33652
rect 25501 33643 25559 33649
rect 25501 33609 25513 33643
rect 25547 33640 25559 33643
rect 26050 33640 26056 33652
rect 25547 33612 26056 33640
rect 25547 33609 25559 33612
rect 25501 33603 25559 33609
rect 26050 33600 26056 33612
rect 26108 33600 26114 33652
rect 30837 33643 30895 33649
rect 30837 33609 30849 33643
rect 30883 33640 30895 33643
rect 30926 33640 30932 33652
rect 30883 33612 30932 33640
rect 30883 33609 30895 33612
rect 30837 33603 30895 33609
rect 30926 33600 30932 33612
rect 30984 33600 30990 33652
rect 32582 33600 32588 33652
rect 32640 33600 32646 33652
rect 33410 33600 33416 33652
rect 33468 33600 33474 33652
rect 36170 33600 36176 33652
rect 36228 33640 36234 33652
rect 36814 33640 36820 33652
rect 36228 33612 36820 33640
rect 36228 33600 36234 33612
rect 36814 33600 36820 33612
rect 36872 33600 36878 33652
rect 38746 33600 38752 33652
rect 38804 33640 38810 33652
rect 39485 33643 39543 33649
rect 39485 33640 39497 33643
rect 38804 33612 39497 33640
rect 38804 33600 38810 33612
rect 39485 33609 39497 33612
rect 39531 33609 39543 33643
rect 39485 33603 39543 33609
rect 39574 33600 39580 33652
rect 39632 33600 39638 33652
rect 39942 33600 39948 33652
rect 40000 33600 40006 33652
rect 40402 33600 40408 33652
rect 40460 33600 40466 33652
rect 40773 33643 40831 33649
rect 40773 33609 40785 33643
rect 40819 33640 40831 33643
rect 40862 33640 40868 33652
rect 40819 33612 40868 33640
rect 40819 33609 40831 33612
rect 40773 33603 40831 33609
rect 40862 33600 40868 33612
rect 40920 33600 40926 33652
rect 15366 33544 15700 33572
rect 17497 33575 17555 33581
rect 15366 33541 15378 33544
rect 15320 33535 15378 33541
rect 17497 33541 17509 33575
rect 17543 33572 17555 33575
rect 18046 33572 18052 33584
rect 17543 33544 18052 33572
rect 17543 33541 17555 33544
rect 17497 33535 17555 33541
rect 18046 33532 18052 33544
rect 18104 33532 18110 33584
rect 20349 33575 20407 33581
rect 20349 33541 20361 33575
rect 20395 33572 20407 33575
rect 20530 33572 20536 33584
rect 20395 33544 20536 33572
rect 20395 33541 20407 33544
rect 20349 33535 20407 33541
rect 20530 33532 20536 33544
rect 20588 33532 20594 33584
rect 20622 33532 20628 33584
rect 20680 33572 20686 33584
rect 22830 33572 22836 33584
rect 20680 33544 21404 33572
rect 20680 33532 20686 33544
rect 14001 33507 14059 33513
rect 14001 33504 14013 33507
rect 13556 33476 14013 33504
rect 14001 33473 14013 33476
rect 14047 33473 14059 33507
rect 14001 33467 14059 33473
rect 15470 33464 15476 33516
rect 15528 33504 15534 33516
rect 16025 33507 16083 33513
rect 15528 33476 15700 33504
rect 15528 33464 15534 33476
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 2130 33436 2136 33448
rect 1719 33408 2136 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 2130 33396 2136 33408
rect 2188 33396 2194 33448
rect 3510 33396 3516 33448
rect 3568 33396 3574 33448
rect 3602 33396 3608 33448
rect 3660 33396 3666 33448
rect 3697 33439 3755 33445
rect 3697 33405 3709 33439
rect 3743 33405 3755 33439
rect 3697 33399 3755 33405
rect 3712 33368 3740 33399
rect 6914 33396 6920 33448
rect 6972 33436 6978 33448
rect 7101 33439 7159 33445
rect 7101 33436 7113 33439
rect 6972 33408 7113 33436
rect 6972 33396 6978 33408
rect 7101 33405 7113 33408
rect 7147 33405 7159 33439
rect 7101 33399 7159 33405
rect 7374 33396 7380 33448
rect 7432 33396 7438 33448
rect 7466 33396 7472 33448
rect 7524 33436 7530 33448
rect 7837 33439 7895 33445
rect 7837 33436 7849 33439
rect 7524 33408 7849 33436
rect 7524 33396 7530 33408
rect 7837 33405 7849 33408
rect 7883 33436 7895 33439
rect 8018 33436 8024 33448
rect 7883 33408 8024 33436
rect 7883 33405 7895 33408
rect 7837 33399 7895 33405
rect 8018 33396 8024 33408
rect 8076 33396 8082 33448
rect 8113 33439 8171 33445
rect 8113 33405 8125 33439
rect 8159 33405 8171 33439
rect 9950 33436 9956 33448
rect 8113 33399 8171 33405
rect 9416 33408 9956 33436
rect 3160 33340 3740 33368
rect 3160 33312 3188 33340
rect 7282 33328 7288 33380
rect 7340 33368 7346 33380
rect 8128 33368 8156 33399
rect 7340 33340 8156 33368
rect 7340 33328 7346 33340
rect 3142 33260 3148 33312
rect 3200 33260 3206 33312
rect 3234 33260 3240 33312
rect 3292 33260 3298 33312
rect 3786 33260 3792 33312
rect 3844 33300 3850 33312
rect 4157 33303 4215 33309
rect 4157 33300 4169 33303
rect 3844 33272 4169 33300
rect 3844 33260 3850 33272
rect 4157 33269 4169 33272
rect 4203 33269 4215 33303
rect 4157 33263 4215 33269
rect 6822 33260 6828 33312
rect 6880 33260 6886 33312
rect 7098 33260 7104 33312
rect 7156 33260 7162 33312
rect 8128 33300 8156 33340
rect 9416 33300 9444 33408
rect 9950 33396 9956 33408
rect 10008 33396 10014 33448
rect 15562 33396 15568 33448
rect 15620 33396 15626 33448
rect 15672 33436 15700 33476
rect 16025 33473 16037 33507
rect 16071 33504 16083 33507
rect 16482 33504 16488 33516
rect 16071 33476 16488 33504
rect 16071 33473 16083 33476
rect 16025 33467 16083 33473
rect 16482 33464 16488 33476
rect 16540 33464 16546 33516
rect 17862 33464 17868 33516
rect 17920 33504 17926 33516
rect 18141 33507 18199 33513
rect 18141 33504 18153 33507
rect 17920 33476 18153 33504
rect 17920 33464 17926 33476
rect 18141 33473 18153 33476
rect 18187 33473 18199 33507
rect 18141 33467 18199 33473
rect 19518 33464 19524 33516
rect 19576 33464 19582 33516
rect 21376 33513 21404 33544
rect 21836 33544 22836 33572
rect 21836 33513 21864 33544
rect 22830 33532 22836 33544
rect 22888 33532 22894 33584
rect 23753 33575 23811 33581
rect 23753 33541 23765 33575
rect 23799 33572 23811 33575
rect 23934 33572 23940 33584
rect 23799 33544 23940 33572
rect 23799 33541 23811 33544
rect 23753 33535 23811 33541
rect 23934 33532 23940 33544
rect 23992 33532 23998 33584
rect 22094 33513 22100 33516
rect 20441 33507 20499 33513
rect 20441 33473 20453 33507
rect 20487 33504 20499 33507
rect 20809 33507 20867 33513
rect 20809 33504 20821 33507
rect 20487 33476 20821 33504
rect 20487 33473 20499 33476
rect 20441 33467 20499 33473
rect 20809 33473 20821 33476
rect 20855 33473 20867 33507
rect 20809 33467 20867 33473
rect 21361 33507 21419 33513
rect 21361 33473 21373 33507
rect 21407 33473 21419 33507
rect 21361 33467 21419 33473
rect 21821 33507 21879 33513
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 22088 33467 22100 33513
rect 22094 33464 22100 33467
rect 22152 33464 22158 33516
rect 22370 33464 22376 33516
rect 22428 33504 22434 33516
rect 25409 33507 25467 33513
rect 22428 33476 24891 33504
rect 22428 33464 22434 33476
rect 16209 33439 16267 33445
rect 16209 33436 16221 33439
rect 15672 33408 16221 33436
rect 16209 33405 16221 33408
rect 16255 33436 16267 33439
rect 17681 33439 17739 33445
rect 17681 33436 17693 33439
rect 16255 33408 17693 33436
rect 16255 33405 16267 33408
rect 16209 33399 16267 33405
rect 17681 33405 17693 33408
rect 17727 33405 17739 33439
rect 17681 33399 17739 33405
rect 8128 33272 9444 33300
rect 11054 33260 11060 33312
rect 11112 33300 11118 33312
rect 11333 33303 11391 33309
rect 11333 33300 11345 33303
rect 11112 33272 11345 33300
rect 11112 33260 11118 33272
rect 11333 33269 11345 33272
rect 11379 33269 11391 33303
rect 11333 33263 11391 33269
rect 13446 33260 13452 33312
rect 13504 33260 13510 33312
rect 15286 33260 15292 33312
rect 15344 33300 15350 33312
rect 17034 33300 17040 33312
rect 15344 33272 17040 33300
rect 15344 33260 15350 33272
rect 17034 33260 17040 33272
rect 17092 33260 17098 33312
rect 17696 33300 17724 33399
rect 18414 33396 18420 33448
rect 18472 33396 18478 33448
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19889 33439 19947 33445
rect 19889 33436 19901 33439
rect 19484 33408 19901 33436
rect 19484 33396 19490 33408
rect 19889 33405 19901 33408
rect 19935 33436 19947 33439
rect 20070 33436 20076 33448
rect 19935 33408 20076 33436
rect 19935 33405 19947 33408
rect 19889 33399 19947 33405
rect 20070 33396 20076 33408
rect 20128 33396 20134 33448
rect 20622 33396 20628 33448
rect 20680 33396 20686 33448
rect 23937 33439 23995 33445
rect 23937 33436 23949 33439
rect 23124 33408 23949 33436
rect 23124 33300 23152 33408
rect 23937 33405 23949 33408
rect 23983 33436 23995 33439
rect 24026 33436 24032 33448
rect 23983 33408 24032 33436
rect 23983 33405 23995 33408
rect 23937 33399 23995 33405
rect 24026 33396 24032 33408
rect 24084 33396 24090 33448
rect 24765 33439 24823 33445
rect 24765 33405 24777 33439
rect 24811 33405 24823 33439
rect 24863 33436 24891 33476
rect 25409 33473 25421 33507
rect 25455 33504 25467 33507
rect 25866 33504 25872 33516
rect 25455 33476 25872 33504
rect 25455 33473 25467 33476
rect 25409 33467 25467 33473
rect 25866 33464 25872 33476
rect 25924 33464 25930 33516
rect 28350 33464 28356 33516
rect 28408 33504 28414 33516
rect 29730 33513 29736 33516
rect 28721 33507 28779 33513
rect 28721 33504 28733 33507
rect 28408 33476 28733 33504
rect 28408 33464 28414 33476
rect 28721 33473 28733 33476
rect 28767 33473 28779 33507
rect 28721 33467 28779 33473
rect 29724 33467 29736 33513
rect 29730 33464 29736 33467
rect 29788 33464 29794 33516
rect 30944 33504 30972 33600
rect 35805 33575 35863 33581
rect 35805 33541 35817 33575
rect 35851 33572 35863 33575
rect 36538 33572 36544 33584
rect 35851 33544 36544 33572
rect 35851 33541 35863 33544
rect 35805 33535 35863 33541
rect 36538 33532 36544 33544
rect 36596 33532 36602 33584
rect 38657 33575 38715 33581
rect 38657 33541 38669 33575
rect 38703 33572 38715 33575
rect 39298 33572 39304 33584
rect 38703 33544 39304 33572
rect 38703 33541 38715 33544
rect 38657 33535 38715 33541
rect 39298 33532 39304 33544
rect 39356 33532 39362 33584
rect 39666 33532 39672 33584
rect 39724 33572 39730 33584
rect 41233 33575 41291 33581
rect 41233 33572 41245 33575
rect 39724 33544 41245 33572
rect 39724 33532 39730 33544
rect 41233 33541 41245 33544
rect 41279 33541 41291 33575
rect 41233 33535 41291 33541
rect 31481 33507 31539 33513
rect 31481 33504 31493 33507
rect 30944 33476 31493 33504
rect 31481 33473 31493 33476
rect 31527 33473 31539 33507
rect 31481 33467 31539 33473
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33504 32551 33507
rect 32582 33504 32588 33516
rect 32539 33476 32588 33504
rect 32539 33473 32551 33476
rect 32493 33467 32551 33473
rect 32582 33464 32588 33476
rect 32640 33464 32646 33516
rect 33778 33464 33784 33516
rect 33836 33464 33842 33516
rect 33873 33507 33931 33513
rect 33873 33473 33885 33507
rect 33919 33504 33931 33507
rect 34054 33504 34060 33516
rect 33919 33476 34060 33504
rect 33919 33473 33931 33476
rect 33873 33467 33931 33473
rect 34054 33464 34060 33476
rect 34112 33464 34118 33516
rect 35897 33507 35955 33513
rect 35897 33473 35909 33507
rect 35943 33504 35955 33507
rect 36265 33507 36323 33513
rect 36265 33504 36277 33507
rect 35943 33476 36277 33504
rect 35943 33473 35955 33476
rect 35897 33467 35955 33473
rect 36265 33473 36277 33476
rect 36311 33473 36323 33507
rect 36265 33467 36323 33473
rect 37277 33507 37335 33513
rect 37277 33473 37289 33507
rect 37323 33504 37335 33507
rect 38102 33504 38108 33516
rect 37323 33476 38108 33504
rect 37323 33473 37335 33476
rect 37277 33467 37335 33473
rect 38102 33464 38108 33476
rect 38160 33504 38166 33516
rect 38562 33504 38568 33516
rect 38160 33476 38568 33504
rect 38160 33464 38166 33476
rect 38562 33464 38568 33476
rect 38620 33464 38626 33516
rect 38672 33476 40172 33504
rect 25685 33439 25743 33445
rect 25685 33436 25697 33439
rect 24863 33408 25697 33436
rect 24765 33399 24823 33405
rect 25685 33405 25697 33408
rect 25731 33436 25743 33439
rect 25774 33436 25780 33448
rect 25731 33408 25780 33436
rect 25731 33405 25743 33408
rect 25685 33399 25743 33405
rect 23201 33371 23259 33377
rect 23201 33337 23213 33371
rect 23247 33368 23259 33371
rect 23382 33368 23388 33380
rect 23247 33340 23388 33368
rect 23247 33337 23259 33340
rect 23201 33331 23259 33337
rect 23382 33328 23388 33340
rect 23440 33368 23446 33380
rect 24780 33368 24808 33399
rect 25774 33396 25780 33408
rect 25832 33396 25838 33448
rect 29454 33396 29460 33448
rect 29512 33396 29518 33448
rect 32769 33439 32827 33445
rect 32769 33405 32781 33439
rect 32815 33405 32827 33439
rect 32769 33399 32827 33405
rect 23440 33340 24808 33368
rect 23440 33328 23446 33340
rect 30558 33328 30564 33380
rect 30616 33368 30622 33380
rect 30929 33371 30987 33377
rect 30929 33368 30941 33371
rect 30616 33340 30941 33368
rect 30616 33328 30622 33340
rect 30929 33337 30941 33340
rect 30975 33337 30987 33371
rect 30929 33331 30987 33337
rect 32674 33328 32680 33380
rect 32732 33368 32738 33380
rect 32784 33368 32812 33399
rect 33962 33396 33968 33448
rect 34020 33396 34026 33448
rect 35802 33396 35808 33448
rect 35860 33436 35866 33448
rect 35989 33439 36047 33445
rect 35989 33436 36001 33439
rect 35860 33408 36001 33436
rect 35860 33396 35866 33408
rect 35989 33405 36001 33408
rect 36035 33405 36047 33439
rect 35989 33399 36047 33405
rect 36446 33396 36452 33448
rect 36504 33436 36510 33448
rect 36817 33439 36875 33445
rect 36817 33436 36829 33439
rect 36504 33408 36829 33436
rect 36504 33396 36510 33408
rect 36817 33405 36829 33408
rect 36863 33405 36875 33439
rect 36817 33399 36875 33405
rect 37366 33396 37372 33448
rect 37424 33436 37430 33448
rect 38013 33439 38071 33445
rect 38013 33436 38025 33439
rect 37424 33408 38025 33436
rect 37424 33396 37430 33408
rect 38013 33405 38025 33408
rect 38059 33405 38071 33439
rect 38013 33399 38071 33405
rect 38378 33396 38384 33448
rect 38436 33436 38442 33448
rect 38672 33436 38700 33476
rect 38436 33408 38700 33436
rect 38749 33439 38807 33445
rect 38436 33396 38442 33408
rect 38749 33405 38761 33439
rect 38795 33405 38807 33439
rect 38749 33399 38807 33405
rect 38933 33439 38991 33445
rect 38933 33405 38945 33439
rect 38979 33436 38991 33439
rect 39022 33436 39028 33448
rect 38979 33408 39028 33436
rect 38979 33405 38991 33408
rect 38933 33399 38991 33405
rect 35820 33368 35848 33396
rect 32732 33340 35848 33368
rect 32732 33328 32738 33340
rect 17696 33272 23152 33300
rect 23474 33260 23480 33312
rect 23532 33300 23538 33312
rect 24213 33303 24271 33309
rect 24213 33300 24225 33303
rect 23532 33272 24225 33300
rect 23532 33260 23538 33272
rect 24213 33269 24225 33272
rect 24259 33269 24271 33303
rect 24213 33263 24271 33269
rect 28629 33303 28687 33309
rect 28629 33269 28641 33303
rect 28675 33300 28687 33303
rect 30190 33300 30196 33312
rect 28675 33272 30196 33300
rect 28675 33269 28687 33272
rect 28629 33263 28687 33269
rect 30190 33260 30196 33272
rect 30248 33260 30254 33312
rect 32122 33260 32128 33312
rect 32180 33260 32186 33312
rect 35434 33260 35440 33312
rect 35492 33260 35498 33312
rect 37642 33260 37648 33312
rect 37700 33300 37706 33312
rect 38289 33303 38347 33309
rect 38289 33300 38301 33303
rect 37700 33272 38301 33300
rect 37700 33260 37706 33272
rect 38289 33269 38301 33272
rect 38335 33269 38347 33303
rect 38764 33300 38792 33399
rect 39022 33396 39028 33408
rect 39080 33436 39086 33448
rect 39761 33439 39819 33445
rect 39080 33408 39712 33436
rect 39080 33396 39086 33408
rect 39114 33328 39120 33380
rect 39172 33328 39178 33380
rect 39684 33368 39712 33408
rect 39761 33405 39773 33439
rect 39807 33436 39819 33439
rect 40034 33436 40040 33448
rect 39807 33408 40040 33436
rect 39807 33405 39819 33408
rect 39761 33399 39819 33405
rect 40034 33396 40040 33408
rect 40092 33396 40098 33448
rect 40144 33436 40172 33476
rect 40310 33464 40316 33516
rect 40368 33464 40374 33516
rect 41141 33507 41199 33513
rect 41141 33504 41153 33507
rect 40420 33476 41153 33504
rect 40420 33436 40448 33476
rect 41141 33473 41153 33476
rect 41187 33473 41199 33507
rect 41141 33467 41199 33473
rect 40144 33408 40448 33436
rect 40497 33439 40555 33445
rect 40497 33405 40509 33439
rect 40543 33436 40555 33439
rect 40954 33436 40960 33448
rect 40543 33408 40960 33436
rect 40543 33405 40555 33408
rect 40497 33399 40555 33405
rect 40512 33368 40540 33399
rect 40954 33396 40960 33408
rect 41012 33436 41018 33448
rect 41325 33439 41383 33445
rect 41325 33436 41337 33439
rect 41012 33408 41337 33436
rect 41012 33396 41018 33408
rect 41325 33405 41337 33408
rect 41371 33405 41383 33439
rect 41325 33399 41383 33405
rect 39684 33340 40540 33368
rect 38838 33300 38844 33312
rect 38764 33272 38844 33300
rect 38289 33263 38347 33269
rect 38838 33260 38844 33272
rect 38896 33260 38902 33312
rect 1104 33210 42504 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 42504 33210
rect 1104 33136 42504 33158
rect 5905 33099 5963 33105
rect 4724 33068 5488 33096
rect 4724 33037 4752 33068
rect 4709 33031 4767 33037
rect 4709 32997 4721 33031
rect 4755 32997 4767 33031
rect 4709 32991 4767 32997
rect 5350 32988 5356 33040
rect 5408 32988 5414 33040
rect 5460 33028 5488 33068
rect 5905 33065 5917 33099
rect 5951 33096 5963 33099
rect 6822 33096 6828 33108
rect 5951 33068 6828 33096
rect 5951 33065 5963 33068
rect 5905 33059 5963 33065
rect 6822 33056 6828 33068
rect 6880 33056 6886 33108
rect 7374 33056 7380 33108
rect 7432 33056 7438 33108
rect 10226 33056 10232 33108
rect 10284 33056 10290 33108
rect 10318 33056 10324 33108
rect 10376 33056 10382 33108
rect 10870 33056 10876 33108
rect 10928 33096 10934 33108
rect 10928 33068 12388 33096
rect 10928 33056 10934 33068
rect 6362 33028 6368 33040
rect 5460 33000 6368 33028
rect 6362 32988 6368 33000
rect 6420 32988 6426 33040
rect 7101 33031 7159 33037
rect 7101 32997 7113 33031
rect 7147 32997 7159 33031
rect 7101 32991 7159 32997
rect 1670 32920 1676 32972
rect 1728 32920 1734 32972
rect 3510 32920 3516 32972
rect 3568 32960 3574 32972
rect 4341 32963 4399 32969
rect 4341 32960 4353 32963
rect 3568 32932 4353 32960
rect 3568 32920 3574 32932
rect 4341 32929 4353 32932
rect 4387 32929 4399 32963
rect 5368 32960 5396 32988
rect 5997 32963 6055 32969
rect 5997 32960 6009 32963
rect 5368 32932 6009 32960
rect 4341 32923 4399 32929
rect 5997 32929 6009 32932
rect 6043 32929 6055 32963
rect 7116 32960 7144 32991
rect 9950 32988 9956 33040
rect 10008 33028 10014 33040
rect 10008 33000 11100 33028
rect 10008 32988 10014 33000
rect 10045 32963 10103 32969
rect 7116 32932 7880 32960
rect 5997 32923 6055 32929
rect 3602 32892 3608 32904
rect 3528 32864 3608 32892
rect 1949 32827 2007 32833
rect 1949 32793 1961 32827
rect 1995 32793 2007 32827
rect 1949 32787 2007 32793
rect 1964 32756 1992 32787
rect 2958 32784 2964 32836
rect 3016 32784 3022 32836
rect 3528 32768 3556 32864
rect 3602 32852 3608 32864
rect 3660 32892 3666 32904
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3660 32864 3985 32892
rect 3660 32852 3666 32864
rect 3973 32861 3985 32864
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 4062 32852 4068 32904
rect 4120 32892 4126 32904
rect 4249 32895 4307 32901
rect 4249 32892 4261 32895
rect 4120 32864 4261 32892
rect 4120 32852 4126 32864
rect 4249 32861 4261 32864
rect 4295 32861 4307 32895
rect 4249 32855 4307 32861
rect 4157 32827 4215 32833
rect 4157 32793 4169 32827
rect 4203 32824 4215 32827
rect 4356 32824 4384 32923
rect 5169 32895 5227 32901
rect 5169 32861 5181 32895
rect 5215 32861 5227 32895
rect 5169 32855 5227 32861
rect 4706 32824 4712 32836
rect 4203 32796 4712 32824
rect 4203 32793 4215 32796
rect 4157 32787 4215 32793
rect 4706 32784 4712 32796
rect 4764 32784 4770 32836
rect 5184 32824 5212 32855
rect 5350 32852 5356 32904
rect 5408 32852 5414 32904
rect 5445 32895 5503 32901
rect 5445 32861 5457 32895
rect 5491 32892 5503 32895
rect 5626 32892 5632 32904
rect 5491 32864 5632 32892
rect 5491 32861 5503 32864
rect 5445 32855 5503 32861
rect 5626 32852 5632 32864
rect 5684 32852 5690 32904
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32892 5779 32895
rect 5902 32892 5908 32904
rect 5767 32864 5908 32892
rect 5767 32861 5779 32864
rect 5721 32855 5779 32861
rect 5736 32824 5764 32855
rect 5902 32852 5908 32864
rect 5960 32852 5966 32904
rect 6730 32852 6736 32904
rect 6788 32892 6794 32904
rect 6825 32895 6883 32901
rect 6825 32892 6837 32895
rect 6788 32864 6837 32892
rect 6788 32852 6794 32864
rect 6825 32861 6837 32864
rect 6871 32861 6883 32895
rect 6825 32855 6883 32861
rect 6914 32852 6920 32904
rect 6972 32852 6978 32904
rect 7098 32852 7104 32904
rect 7156 32852 7162 32904
rect 7561 32895 7619 32901
rect 7561 32861 7573 32895
rect 7607 32861 7619 32895
rect 7561 32855 7619 32861
rect 5184 32796 5764 32824
rect 7576 32824 7604 32855
rect 7650 32852 7656 32904
rect 7708 32852 7714 32904
rect 7852 32901 7880 32932
rect 10045 32929 10057 32963
rect 10091 32960 10103 32963
rect 10318 32960 10324 32972
rect 10091 32932 10324 32960
rect 10091 32929 10103 32932
rect 10045 32923 10103 32929
rect 10318 32920 10324 32932
rect 10376 32920 10382 32972
rect 10962 32920 10968 32972
rect 11020 32920 11026 32972
rect 11072 32969 11100 33000
rect 11057 32963 11115 32969
rect 11057 32929 11069 32963
rect 11103 32929 11115 32963
rect 12360 32960 12388 33068
rect 12802 33056 12808 33108
rect 12860 33056 12866 33108
rect 13906 33056 13912 33108
rect 13964 33096 13970 33108
rect 13964 33068 16436 33096
rect 13964 33056 13970 33068
rect 12437 33031 12495 33037
rect 12437 32997 12449 33031
rect 12483 33028 12495 33031
rect 13814 33028 13820 33040
rect 12483 33000 13820 33028
rect 12483 32997 12495 33000
rect 12437 32991 12495 32997
rect 13814 32988 13820 33000
rect 13872 32988 13878 33040
rect 16408 33028 16436 33068
rect 16482 33056 16488 33108
rect 16540 33096 16546 33108
rect 16669 33099 16727 33105
rect 16669 33096 16681 33099
rect 16540 33068 16681 33096
rect 16540 33056 16546 33068
rect 16669 33065 16681 33068
rect 16715 33065 16727 33099
rect 16669 33059 16727 33065
rect 21729 33099 21787 33105
rect 21729 33065 21741 33099
rect 21775 33096 21787 33099
rect 22094 33096 22100 33108
rect 21775 33068 22100 33096
rect 21775 33065 21787 33068
rect 21729 33059 21787 33065
rect 22094 33056 22100 33068
rect 22152 33056 22158 33108
rect 22741 33099 22799 33105
rect 22741 33065 22753 33099
rect 22787 33096 22799 33099
rect 23842 33096 23848 33108
rect 22787 33068 23848 33096
rect 22787 33065 22799 33068
rect 22741 33059 22799 33065
rect 23842 33056 23848 33068
rect 23900 33096 23906 33108
rect 28353 33099 28411 33105
rect 28353 33096 28365 33099
rect 23900 33068 24992 33096
rect 23900 33056 23906 33068
rect 16408 33000 17172 33028
rect 13170 32960 13176 32972
rect 12360 32932 13176 32960
rect 11057 32923 11115 32929
rect 13170 32920 13176 32932
rect 13228 32960 13234 32972
rect 13357 32963 13415 32969
rect 13357 32960 13369 32963
rect 13228 32932 13369 32960
rect 13228 32920 13234 32932
rect 13357 32929 13369 32932
rect 13403 32960 13415 32963
rect 13538 32960 13544 32972
rect 13403 32932 13544 32960
rect 13403 32929 13415 32932
rect 13357 32923 13415 32929
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 15562 32960 15568 32972
rect 14936 32932 15568 32960
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32861 7895 32895
rect 7837 32855 7895 32861
rect 7929 32895 7987 32901
rect 7929 32861 7941 32895
rect 7975 32892 7987 32895
rect 8386 32892 8392 32904
rect 7975 32864 8392 32892
rect 7975 32861 7987 32864
rect 7929 32855 7987 32861
rect 8386 32852 8392 32864
rect 8444 32852 8450 32904
rect 9953 32895 10011 32901
rect 9953 32861 9965 32895
rect 9999 32892 10011 32895
rect 9999 32864 11100 32892
rect 9999 32861 10011 32864
rect 9953 32855 10011 32861
rect 8478 32824 8484 32836
rect 7576 32796 8484 32824
rect 8478 32784 8484 32796
rect 8536 32784 8542 32836
rect 9585 32827 9643 32833
rect 9585 32793 9597 32827
rect 9631 32824 9643 32827
rect 10870 32824 10876 32836
rect 9631 32796 10876 32824
rect 9631 32793 9643 32796
rect 9585 32787 9643 32793
rect 10870 32784 10876 32796
rect 10928 32784 10934 32836
rect 11072 32824 11100 32864
rect 11146 32852 11152 32904
rect 11204 32892 11210 32904
rect 11313 32895 11371 32901
rect 11313 32892 11325 32895
rect 11204 32864 11325 32892
rect 11204 32852 11210 32864
rect 11313 32861 11325 32864
rect 11359 32861 11371 32895
rect 11313 32855 11371 32861
rect 13265 32895 13323 32901
rect 13265 32861 13277 32895
rect 13311 32892 13323 32895
rect 13446 32892 13452 32904
rect 13311 32864 13452 32892
rect 13311 32861 13323 32864
rect 13265 32855 13323 32861
rect 13446 32852 13452 32864
rect 13504 32852 13510 32904
rect 13998 32852 14004 32904
rect 14056 32892 14062 32904
rect 14093 32895 14151 32901
rect 14093 32892 14105 32895
rect 14056 32864 14105 32892
rect 14056 32852 14062 32864
rect 14093 32861 14105 32864
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 14366 32852 14372 32904
rect 14424 32892 14430 32904
rect 14936 32901 14964 32932
rect 15562 32920 15568 32932
rect 15620 32960 15626 32972
rect 17037 32963 17095 32969
rect 17037 32960 17049 32963
rect 15620 32932 17049 32960
rect 15620 32920 15626 32932
rect 17037 32929 17049 32932
rect 17083 32929 17095 32963
rect 17144 32960 17172 33000
rect 17144 32932 18552 32960
rect 17037 32923 17095 32929
rect 14921 32895 14979 32901
rect 14921 32892 14933 32895
rect 14424 32864 14933 32892
rect 14424 32852 14430 32864
rect 14921 32861 14933 32864
rect 14967 32861 14979 32895
rect 18524 32892 18552 32932
rect 20070 32920 20076 32972
rect 20128 32920 20134 32972
rect 20622 32920 20628 32972
rect 20680 32960 20686 32972
rect 21085 32963 21143 32969
rect 21085 32960 21097 32963
rect 20680 32932 21097 32960
rect 20680 32920 20686 32932
rect 21085 32929 21097 32932
rect 21131 32960 21143 32963
rect 22370 32960 22376 32972
rect 21131 32932 22376 32960
rect 21131 32929 21143 32932
rect 21085 32923 21143 32929
rect 22370 32920 22376 32932
rect 22428 32920 22434 32972
rect 24964 32969 24992 33068
rect 26804 33068 28365 33096
rect 24949 32963 25007 32969
rect 24949 32929 24961 32963
rect 24995 32929 25007 32963
rect 24949 32923 25007 32929
rect 26142 32920 26148 32972
rect 26200 32960 26206 32972
rect 26329 32963 26387 32969
rect 26329 32960 26341 32963
rect 26200 32932 26341 32960
rect 26200 32920 26206 32932
rect 26329 32929 26341 32932
rect 26375 32929 26387 32963
rect 26329 32923 26387 32929
rect 26694 32920 26700 32972
rect 26752 32920 26758 32972
rect 26804 32969 26832 33068
rect 28353 33065 28365 33068
rect 28399 33065 28411 33099
rect 28353 33059 28411 33065
rect 29730 33056 29736 33108
rect 29788 33096 29794 33108
rect 29917 33099 29975 33105
rect 29917 33096 29929 33099
rect 29788 33068 29929 33096
rect 29788 33056 29794 33068
rect 29917 33065 29929 33068
rect 29963 33065 29975 33099
rect 29917 33059 29975 33065
rect 32217 33099 32275 33105
rect 32217 33065 32229 33099
rect 32263 33096 32275 33099
rect 32306 33096 32312 33108
rect 32263 33068 32312 33096
rect 32263 33065 32275 33068
rect 32217 33059 32275 33065
rect 32306 33056 32312 33068
rect 32364 33056 32370 33108
rect 38654 33056 38660 33108
rect 38712 33096 38718 33108
rect 38749 33099 38807 33105
rect 38749 33096 38761 33099
rect 38712 33068 38761 33096
rect 38712 33056 38718 33068
rect 38749 33065 38761 33068
rect 38795 33065 38807 33099
rect 38749 33059 38807 33065
rect 28092 33000 30880 33028
rect 26789 32963 26847 32969
rect 26789 32929 26801 32963
rect 26835 32929 26847 32963
rect 26789 32923 26847 32929
rect 20901 32895 20959 32901
rect 20901 32892 20913 32895
rect 18524 32864 20913 32892
rect 14921 32855 14979 32861
rect 20901 32861 20913 32864
rect 20947 32892 20959 32895
rect 21818 32892 21824 32904
rect 20947 32864 21824 32892
rect 20947 32861 20959 32864
rect 20901 32855 20959 32861
rect 21818 32852 21824 32864
rect 21876 32852 21882 32904
rect 22189 32895 22247 32901
rect 22189 32861 22201 32895
rect 22235 32892 22247 32895
rect 23474 32892 23480 32904
rect 22235 32864 23480 32892
rect 22235 32861 22247 32864
rect 22189 32855 22247 32861
rect 23474 32852 23480 32864
rect 23532 32852 23538 32904
rect 24118 32852 24124 32904
rect 24176 32852 24182 32904
rect 26881 32895 26939 32901
rect 26881 32861 26893 32895
rect 26927 32892 26939 32895
rect 27890 32892 27896 32904
rect 26927 32864 27896 32892
rect 26927 32861 26939 32864
rect 26881 32855 26939 32861
rect 27890 32852 27896 32864
rect 27948 32852 27954 32904
rect 12158 32824 12164 32836
rect 11072 32796 12164 32824
rect 12158 32784 12164 32796
rect 12216 32784 12222 32836
rect 15194 32784 15200 32836
rect 15252 32784 15258 32836
rect 15286 32784 15292 32836
rect 15344 32824 15350 32836
rect 15344 32796 15686 32824
rect 15344 32784 15350 32796
rect 17310 32784 17316 32836
rect 17368 32784 17374 32836
rect 19426 32824 19432 32836
rect 18538 32796 19432 32824
rect 19426 32784 19432 32796
rect 19484 32784 19490 32836
rect 23382 32784 23388 32836
rect 23440 32824 23446 32836
rect 23854 32827 23912 32833
rect 23854 32824 23866 32827
rect 23440 32796 23866 32824
rect 23440 32784 23446 32796
rect 23854 32793 23866 32796
rect 23900 32793 23912 32827
rect 23854 32787 23912 32793
rect 24486 32784 24492 32836
rect 24544 32824 24550 32836
rect 27341 32827 27399 32833
rect 27341 32824 27353 32827
rect 24544 32796 27353 32824
rect 24544 32784 24550 32796
rect 27341 32793 27353 32796
rect 27387 32824 27399 32827
rect 28092 32824 28120 33000
rect 28166 32920 28172 32972
rect 28224 32960 28230 32972
rect 28905 32963 28963 32969
rect 28905 32960 28917 32963
rect 28224 32932 28917 32960
rect 28224 32920 28230 32932
rect 28905 32929 28917 32932
rect 28951 32929 28963 32963
rect 28905 32923 28963 32929
rect 30190 32920 30196 32972
rect 30248 32960 30254 32972
rect 30469 32963 30527 32969
rect 30469 32960 30481 32963
rect 30248 32932 30481 32960
rect 30248 32920 30254 32932
rect 30469 32929 30481 32932
rect 30515 32929 30527 32963
rect 30852 32960 30880 33000
rect 38764 32960 38792 33059
rect 38838 33056 38844 33108
rect 38896 33056 38902 33108
rect 39393 32963 39451 32969
rect 39393 32960 39405 32963
rect 30852 32932 30972 32960
rect 38764 32932 39405 32960
rect 30469 32923 30527 32929
rect 30377 32895 30435 32901
rect 30377 32861 30389 32895
rect 30423 32892 30435 32895
rect 30558 32892 30564 32904
rect 30423 32864 30564 32892
rect 30423 32861 30435 32864
rect 30377 32855 30435 32861
rect 30558 32852 30564 32864
rect 30616 32852 30622 32904
rect 30837 32895 30895 32901
rect 30837 32861 30849 32895
rect 30883 32861 30895 32895
rect 30944 32892 30972 32932
rect 39393 32929 39405 32932
rect 39439 32929 39451 32963
rect 39393 32923 39451 32929
rect 40954 32920 40960 32972
rect 41012 32920 41018 32972
rect 41414 32920 41420 32972
rect 41472 32960 41478 32972
rect 41877 32963 41935 32969
rect 41877 32960 41889 32963
rect 41472 32932 41889 32960
rect 41472 32920 41478 32932
rect 41877 32929 41889 32932
rect 41923 32929 41935 32963
rect 41877 32923 41935 32929
rect 32122 32892 32128 32904
rect 30944 32864 31340 32892
rect 30837 32855 30895 32861
rect 27387 32796 28120 32824
rect 28169 32827 28227 32833
rect 27387 32793 27399 32796
rect 27341 32787 27399 32793
rect 28169 32793 28181 32827
rect 28215 32824 28227 32827
rect 29454 32824 29460 32836
rect 28215 32796 29460 32824
rect 28215 32793 28227 32796
rect 28169 32787 28227 32793
rect 29454 32784 29460 32796
rect 29512 32824 29518 32836
rect 30852 32824 30880 32855
rect 31312 32836 31340 32864
rect 31726 32864 32128 32892
rect 29512 32796 30880 32824
rect 31104 32827 31162 32833
rect 29512 32784 29518 32796
rect 31104 32793 31116 32827
rect 31150 32824 31162 32827
rect 31150 32796 31248 32824
rect 31150 32793 31162 32796
rect 31104 32787 31162 32793
rect 3326 32756 3332 32768
rect 1964 32728 3332 32756
rect 3326 32716 3332 32728
rect 3384 32716 3390 32768
rect 3421 32759 3479 32765
rect 3421 32725 3433 32759
rect 3467 32756 3479 32759
rect 3510 32756 3516 32768
rect 3467 32728 3516 32756
rect 3467 32725 3479 32728
rect 3421 32719 3479 32725
rect 3510 32716 3516 32728
rect 3568 32716 3574 32768
rect 3602 32716 3608 32768
rect 3660 32756 3666 32768
rect 3789 32759 3847 32765
rect 3789 32756 3801 32759
rect 3660 32728 3801 32756
rect 3660 32716 3666 32728
rect 3789 32725 3801 32728
rect 3835 32725 3847 32759
rect 3789 32719 3847 32725
rect 4798 32716 4804 32768
rect 4856 32716 4862 32768
rect 4985 32759 5043 32765
rect 4985 32725 4997 32759
rect 5031 32756 5043 32759
rect 5258 32756 5264 32768
rect 5031 32728 5264 32756
rect 5031 32725 5043 32728
rect 4985 32719 5043 32725
rect 5258 32716 5264 32728
rect 5316 32716 5322 32768
rect 5534 32716 5540 32768
rect 5592 32716 5598 32768
rect 13173 32759 13231 32765
rect 13173 32725 13185 32759
rect 13219 32756 13231 32759
rect 14274 32756 14280 32768
rect 13219 32728 14280 32756
rect 13219 32725 13231 32728
rect 13173 32719 13231 32725
rect 14274 32716 14280 32728
rect 14332 32716 14338 32768
rect 14550 32716 14556 32768
rect 14608 32756 14614 32768
rect 14737 32759 14795 32765
rect 14737 32756 14749 32759
rect 14608 32728 14749 32756
rect 14608 32716 14614 32728
rect 14737 32725 14749 32728
rect 14783 32725 14795 32759
rect 14737 32719 14795 32725
rect 18046 32716 18052 32768
rect 18104 32756 18110 32768
rect 18785 32759 18843 32765
rect 18785 32756 18797 32759
rect 18104 32728 18797 32756
rect 18104 32716 18110 32728
rect 18785 32725 18797 32728
rect 18831 32725 18843 32759
rect 18785 32719 18843 32725
rect 19150 32716 19156 32768
rect 19208 32756 19214 32768
rect 19521 32759 19579 32765
rect 19521 32756 19533 32759
rect 19208 32728 19533 32756
rect 19208 32716 19214 32728
rect 19521 32725 19533 32728
rect 19567 32725 19579 32759
rect 19521 32719 19579 32725
rect 22094 32716 22100 32768
rect 22152 32716 22158 32768
rect 24394 32716 24400 32768
rect 24452 32716 24458 32768
rect 25682 32716 25688 32768
rect 25740 32756 25746 32768
rect 25777 32759 25835 32765
rect 25777 32756 25789 32759
rect 25740 32728 25789 32756
rect 25740 32716 25746 32728
rect 25777 32725 25789 32728
rect 25823 32725 25835 32759
rect 25777 32719 25835 32725
rect 27246 32716 27252 32768
rect 27304 32716 27310 32768
rect 28350 32716 28356 32768
rect 28408 32756 28414 32768
rect 28810 32756 28816 32768
rect 28408 32728 28816 32756
rect 28408 32716 28414 32728
rect 28810 32716 28816 32728
rect 28868 32716 28874 32768
rect 30285 32759 30343 32765
rect 30285 32725 30297 32759
rect 30331 32756 30343 32759
rect 31018 32756 31024 32768
rect 30331 32728 31024 32756
rect 30331 32725 30343 32728
rect 30285 32719 30343 32725
rect 31018 32716 31024 32728
rect 31076 32716 31082 32768
rect 31220 32756 31248 32796
rect 31294 32784 31300 32836
rect 31352 32784 31358 32836
rect 31726 32756 31754 32864
rect 32122 32852 32128 32864
rect 32180 32852 32186 32904
rect 32585 32895 32643 32901
rect 32585 32861 32597 32895
rect 32631 32892 32643 32895
rect 35066 32892 35072 32904
rect 32631 32864 35072 32892
rect 32631 32861 32643 32864
rect 32585 32855 32643 32861
rect 35066 32852 35072 32864
rect 35124 32892 35130 32904
rect 36909 32895 36967 32901
rect 36909 32892 36921 32895
rect 35124 32864 36921 32892
rect 35124 32852 35130 32864
rect 36909 32861 36921 32864
rect 36955 32892 36967 32895
rect 37366 32892 37372 32904
rect 36955 32864 37372 32892
rect 36955 32861 36967 32864
rect 36909 32855 36967 32861
rect 37366 32852 37372 32864
rect 37424 32852 37430 32904
rect 37642 32901 37648 32904
rect 37636 32892 37648 32901
rect 37603 32864 37648 32892
rect 37636 32855 37648 32864
rect 37642 32852 37648 32855
rect 37700 32852 37706 32904
rect 32852 32827 32910 32833
rect 32852 32793 32864 32827
rect 32898 32824 32910 32827
rect 33134 32824 33140 32836
rect 32898 32796 33140 32824
rect 32898 32793 32910 32796
rect 32852 32787 32910 32793
rect 33134 32784 33140 32796
rect 33192 32784 33198 32836
rect 35342 32833 35348 32836
rect 35336 32787 35348 32833
rect 35342 32784 35348 32787
rect 35400 32784 35406 32836
rect 38838 32784 38844 32836
rect 38896 32824 38902 32836
rect 40773 32827 40831 32833
rect 40773 32824 40785 32827
rect 38896 32796 40785 32824
rect 38896 32784 38902 32796
rect 40773 32793 40785 32796
rect 40819 32793 40831 32827
rect 40773 32787 40831 32793
rect 31220 32728 31754 32756
rect 33965 32759 34023 32765
rect 33965 32725 33977 32759
rect 34011 32756 34023 32759
rect 34054 32756 34060 32768
rect 34011 32728 34060 32756
rect 34011 32725 34023 32728
rect 33965 32719 34023 32725
rect 34054 32716 34060 32728
rect 34112 32716 34118 32768
rect 36449 32759 36507 32765
rect 36449 32725 36461 32759
rect 36495 32756 36507 32759
rect 36814 32756 36820 32768
rect 36495 32728 36820 32756
rect 36495 32725 36507 32728
rect 36449 32719 36507 32725
rect 36814 32716 36820 32728
rect 36872 32716 36878 32768
rect 40405 32759 40463 32765
rect 40405 32725 40417 32759
rect 40451 32756 40463 32759
rect 40586 32756 40592 32768
rect 40451 32728 40592 32756
rect 40451 32725 40463 32728
rect 40405 32719 40463 32725
rect 40586 32716 40592 32728
rect 40644 32716 40650 32768
rect 40865 32759 40923 32765
rect 40865 32725 40877 32759
rect 40911 32756 40923 32759
rect 41325 32759 41383 32765
rect 41325 32756 41337 32759
rect 40911 32728 41337 32756
rect 40911 32725 40923 32728
rect 40865 32719 40923 32725
rect 41325 32725 41337 32728
rect 41371 32725 41383 32759
rect 41325 32719 41383 32725
rect 1104 32666 42504 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 42504 32666
rect 1104 32592 42504 32614
rect 2130 32512 2136 32564
rect 2188 32512 2194 32564
rect 2777 32555 2835 32561
rect 2777 32521 2789 32555
rect 2823 32521 2835 32555
rect 2777 32515 2835 32521
rect 2590 32484 2596 32496
rect 2332 32456 2596 32484
rect 2332 32425 2360 32456
rect 2590 32444 2596 32456
rect 2648 32484 2654 32496
rect 2792 32484 2820 32515
rect 3326 32512 3332 32564
rect 3384 32552 3390 32564
rect 3421 32555 3479 32561
rect 3421 32552 3433 32555
rect 3384 32524 3433 32552
rect 3384 32512 3390 32524
rect 3421 32521 3433 32524
rect 3467 32521 3479 32555
rect 5810 32552 5816 32564
rect 3421 32515 3479 32521
rect 3896 32524 5816 32552
rect 2648 32456 2820 32484
rect 2648 32444 2654 32456
rect 2317 32419 2375 32425
rect 2317 32385 2329 32419
rect 2363 32385 2375 32419
rect 2317 32379 2375 32385
rect 2501 32419 2559 32425
rect 2501 32385 2513 32419
rect 2547 32416 2559 32419
rect 3234 32416 3240 32428
rect 2547 32388 3240 32416
rect 2547 32385 2559 32388
rect 2501 32379 2559 32385
rect 3234 32376 3240 32388
rect 3292 32376 3298 32428
rect 3326 32376 3332 32428
rect 3384 32376 3390 32428
rect 3602 32376 3608 32428
rect 3660 32376 3666 32428
rect 3786 32376 3792 32428
rect 3844 32376 3850 32428
rect 3896 32425 3924 32524
rect 5810 32512 5816 32524
rect 5868 32512 5874 32564
rect 12621 32555 12679 32561
rect 12621 32521 12633 32555
rect 12667 32552 12679 32555
rect 13998 32552 14004 32564
rect 12667 32524 14004 32552
rect 12667 32521 12679 32524
rect 12621 32515 12679 32521
rect 13998 32512 14004 32524
rect 14056 32512 14062 32564
rect 14093 32555 14151 32561
rect 14093 32521 14105 32555
rect 14139 32521 14151 32555
rect 14093 32515 14151 32521
rect 6270 32484 6276 32496
rect 5750 32456 6276 32484
rect 6270 32444 6276 32456
rect 6328 32444 6334 32496
rect 7650 32444 7656 32496
rect 7708 32484 7714 32496
rect 8113 32487 8171 32493
rect 8113 32484 8125 32487
rect 7708 32456 8125 32484
rect 7708 32444 7714 32456
rect 8113 32453 8125 32456
rect 8159 32453 8171 32487
rect 8113 32447 8171 32453
rect 13538 32444 13544 32496
rect 13596 32444 13602 32496
rect 13756 32487 13814 32493
rect 13756 32453 13768 32487
rect 13802 32484 13814 32487
rect 14108 32484 14136 32515
rect 14550 32512 14556 32564
rect 14608 32512 14614 32564
rect 17310 32512 17316 32564
rect 17368 32552 17374 32564
rect 17773 32555 17831 32561
rect 17773 32552 17785 32555
rect 17368 32524 17785 32552
rect 17368 32512 17374 32524
rect 17773 32521 17785 32524
rect 17819 32521 17831 32555
rect 17773 32515 17831 32521
rect 18046 32512 18052 32564
rect 18104 32552 18110 32564
rect 18141 32555 18199 32561
rect 18141 32552 18153 32555
rect 18104 32524 18153 32552
rect 18104 32512 18110 32524
rect 18141 32521 18153 32524
rect 18187 32521 18199 32555
rect 18141 32515 18199 32521
rect 18414 32512 18420 32564
rect 18472 32552 18478 32564
rect 18601 32555 18659 32561
rect 18601 32552 18613 32555
rect 18472 32524 18613 32552
rect 18472 32512 18478 32524
rect 18601 32521 18613 32524
rect 18647 32521 18659 32555
rect 22646 32552 22652 32564
rect 18601 32515 18659 32521
rect 18984 32524 22652 32552
rect 18984 32493 19012 32524
rect 22646 32512 22652 32524
rect 22704 32552 22710 32564
rect 23198 32552 23204 32564
rect 22704 32524 23204 32552
rect 22704 32512 22710 32524
rect 23198 32512 23204 32524
rect 23256 32512 23262 32564
rect 23382 32512 23388 32564
rect 23440 32512 23446 32564
rect 23845 32555 23903 32561
rect 23845 32521 23857 32555
rect 23891 32552 23903 32555
rect 24394 32552 24400 32564
rect 23891 32524 24400 32552
rect 23891 32521 23903 32524
rect 23845 32515 23903 32521
rect 24394 32512 24400 32524
rect 24452 32512 24458 32564
rect 26142 32512 26148 32564
rect 26200 32512 26206 32564
rect 28166 32512 28172 32564
rect 28224 32552 28230 32564
rect 28353 32555 28411 32561
rect 28353 32552 28365 32555
rect 28224 32524 28365 32552
rect 28224 32512 28230 32524
rect 28353 32521 28365 32524
rect 28399 32521 28411 32555
rect 28353 32515 28411 32521
rect 33134 32512 33140 32564
rect 33192 32512 33198 32564
rect 36446 32512 36452 32564
rect 36504 32512 36510 32564
rect 38749 32555 38807 32561
rect 38749 32521 38761 32555
rect 38795 32552 38807 32555
rect 38930 32552 38936 32564
rect 38795 32524 38936 32552
rect 38795 32521 38807 32524
rect 38749 32515 38807 32521
rect 38930 32512 38936 32524
rect 38988 32512 38994 32564
rect 41414 32512 41420 32564
rect 41472 32552 41478 32564
rect 41693 32555 41751 32561
rect 41693 32552 41705 32555
rect 41472 32524 41705 32552
rect 41472 32512 41478 32524
rect 41693 32521 41705 32524
rect 41739 32521 41751 32555
rect 41693 32515 41751 32521
rect 13802 32456 14136 32484
rect 18969 32487 19027 32493
rect 13802 32453 13814 32456
rect 13756 32447 13814 32453
rect 18969 32453 18981 32487
rect 19015 32453 19027 32487
rect 18969 32447 19027 32453
rect 19337 32487 19395 32493
rect 19337 32453 19349 32487
rect 19383 32484 19395 32487
rect 19426 32484 19432 32496
rect 19383 32456 19432 32484
rect 19383 32453 19395 32456
rect 19337 32447 19395 32453
rect 19426 32444 19432 32456
rect 19484 32444 19490 32496
rect 19610 32444 19616 32496
rect 19668 32484 19674 32496
rect 19705 32487 19763 32493
rect 19705 32484 19717 32487
rect 19668 32456 19717 32484
rect 19668 32444 19674 32456
rect 19705 32453 19717 32456
rect 19751 32453 19763 32487
rect 19705 32447 19763 32453
rect 20070 32444 20076 32496
rect 20128 32484 20134 32496
rect 20128 32456 20654 32484
rect 20128 32444 20134 32456
rect 24118 32444 24124 32496
rect 24176 32484 24182 32496
rect 27430 32484 27436 32496
rect 24176 32456 27436 32484
rect 24176 32444 24182 32456
rect 3881 32419 3939 32425
rect 3881 32385 3893 32419
rect 3927 32385 3939 32419
rect 3881 32379 3939 32385
rect 3050 32308 3056 32360
rect 3108 32348 3114 32360
rect 3896 32348 3924 32379
rect 6914 32376 6920 32428
rect 6972 32416 6978 32428
rect 7190 32416 7196 32428
rect 6972 32388 7196 32416
rect 6972 32376 6978 32388
rect 7190 32376 7196 32388
rect 7248 32416 7254 32428
rect 7285 32419 7343 32425
rect 7285 32416 7297 32419
rect 7248 32388 7297 32416
rect 7248 32376 7254 32388
rect 7285 32385 7297 32388
rect 7331 32416 7343 32419
rect 7331 32388 8248 32416
rect 7331 32385 7343 32388
rect 7285 32379 7343 32385
rect 8220 32360 8248 32388
rect 8386 32376 8392 32428
rect 8444 32416 8450 32428
rect 8941 32419 8999 32425
rect 8941 32416 8953 32419
rect 8444 32388 8953 32416
rect 8444 32376 8450 32388
rect 8941 32385 8953 32388
rect 8987 32385 8999 32419
rect 13556 32416 13584 32444
rect 14001 32419 14059 32425
rect 13556 32388 13952 32416
rect 8941 32379 8999 32385
rect 3108 32320 3924 32348
rect 4249 32351 4307 32357
rect 3108 32308 3114 32320
rect 4249 32317 4261 32351
rect 4295 32317 4307 32351
rect 4249 32311 4307 32317
rect 4525 32351 4583 32357
rect 4525 32317 4537 32351
rect 4571 32348 4583 32351
rect 4614 32348 4620 32360
rect 4571 32320 4620 32348
rect 4571 32317 4583 32320
rect 4525 32311 4583 32317
rect 3237 32215 3295 32221
rect 3237 32181 3249 32215
rect 3283 32212 3295 32215
rect 3786 32212 3792 32224
rect 3283 32184 3792 32212
rect 3283 32181 3295 32184
rect 3237 32175 3295 32181
rect 3786 32172 3792 32184
rect 3844 32172 3850 32224
rect 4264 32212 4292 32311
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 7374 32308 7380 32360
rect 7432 32348 7438 32360
rect 8021 32351 8079 32357
rect 8021 32348 8033 32351
rect 7432 32320 8033 32348
rect 7432 32308 7438 32320
rect 8021 32317 8033 32320
rect 8067 32317 8079 32351
rect 8021 32311 8079 32317
rect 8202 32308 8208 32360
rect 8260 32348 8266 32360
rect 8481 32351 8539 32357
rect 8481 32348 8493 32351
rect 8260 32320 8493 32348
rect 8260 32308 8266 32320
rect 8481 32317 8493 32320
rect 8527 32348 8539 32351
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 8527 32320 9137 32348
rect 8527 32317 8539 32320
rect 8481 32311 8539 32317
rect 9125 32317 9137 32320
rect 9171 32317 9183 32351
rect 9125 32311 9183 32317
rect 9306 32308 9312 32360
rect 9364 32348 9370 32360
rect 10045 32351 10103 32357
rect 10045 32348 10057 32351
rect 9364 32320 10057 32348
rect 9364 32308 9370 32320
rect 10045 32317 10057 32320
rect 10091 32348 10103 32351
rect 12066 32348 12072 32360
rect 10091 32320 12072 32348
rect 10091 32317 10103 32320
rect 10045 32311 10103 32317
rect 12066 32308 12072 32320
rect 12124 32308 12130 32360
rect 13924 32348 13952 32388
rect 14001 32385 14013 32419
rect 14047 32416 14059 32419
rect 14366 32416 14372 32428
rect 14047 32388 14372 32416
rect 14047 32385 14059 32388
rect 14001 32379 14059 32385
rect 14366 32376 14372 32388
rect 14424 32376 14430 32428
rect 14458 32376 14464 32428
rect 14516 32376 14522 32428
rect 18414 32376 18420 32428
rect 18472 32416 18478 32428
rect 18739 32419 18797 32425
rect 18739 32416 18751 32419
rect 18472 32388 18751 32416
rect 18472 32376 18478 32388
rect 18739 32385 18751 32388
rect 18785 32385 18797 32419
rect 18739 32379 18797 32385
rect 18877 32419 18935 32425
rect 18877 32385 18889 32419
rect 18923 32385 18935 32419
rect 19150 32416 19156 32428
rect 19111 32388 19156 32416
rect 18877 32379 18935 32385
rect 14645 32351 14703 32357
rect 14645 32348 14657 32351
rect 13924 32320 14657 32348
rect 14645 32317 14657 32320
rect 14691 32348 14703 32351
rect 15470 32348 15476 32360
rect 14691 32320 15476 32348
rect 14691 32317 14703 32320
rect 14645 32311 14703 32317
rect 15470 32308 15476 32320
rect 15528 32308 15534 32360
rect 18046 32308 18052 32360
rect 18104 32348 18110 32360
rect 18233 32351 18291 32357
rect 18233 32348 18245 32351
rect 18104 32320 18245 32348
rect 18104 32308 18110 32320
rect 18233 32317 18245 32320
rect 18279 32317 18291 32351
rect 18233 32311 18291 32317
rect 18325 32351 18383 32357
rect 18325 32317 18337 32351
rect 18371 32317 18383 32351
rect 18325 32311 18383 32317
rect 7742 32240 7748 32292
rect 7800 32280 7806 32292
rect 8757 32283 8815 32289
rect 8757 32280 8769 32283
rect 7800 32252 8769 32280
rect 7800 32240 7806 32252
rect 8757 32249 8769 32252
rect 8803 32249 8815 32283
rect 8757 32243 8815 32249
rect 16022 32240 16028 32292
rect 16080 32280 16086 32292
rect 18340 32280 18368 32311
rect 18782 32280 18788 32292
rect 16080 32252 18788 32280
rect 16080 32240 16086 32252
rect 18782 32240 18788 32252
rect 18840 32240 18846 32292
rect 4614 32212 4620 32224
rect 4264 32184 4620 32212
rect 4614 32172 4620 32184
rect 4672 32172 4678 32224
rect 5074 32172 5080 32224
rect 5132 32212 5138 32224
rect 5626 32212 5632 32224
rect 5132 32184 5632 32212
rect 5132 32172 5138 32184
rect 5626 32172 5632 32184
rect 5684 32172 5690 32224
rect 5902 32172 5908 32224
rect 5960 32212 5966 32224
rect 5997 32215 6055 32221
rect 5997 32212 6009 32215
rect 5960 32184 6009 32212
rect 5960 32172 5966 32184
rect 5997 32181 6009 32184
rect 6043 32181 6055 32215
rect 5997 32175 6055 32181
rect 7926 32172 7932 32224
rect 7984 32172 7990 32224
rect 8662 32172 8668 32224
rect 8720 32172 8726 32224
rect 10502 32172 10508 32224
rect 10560 32212 10566 32224
rect 10597 32215 10655 32221
rect 10597 32212 10609 32215
rect 10560 32184 10609 32212
rect 10560 32172 10566 32184
rect 10597 32181 10609 32184
rect 10643 32181 10655 32215
rect 10597 32175 10655 32181
rect 17494 32172 17500 32224
rect 17552 32212 17558 32224
rect 17770 32212 17776 32224
rect 17552 32184 17776 32212
rect 17552 32172 17558 32184
rect 17770 32172 17776 32184
rect 17828 32212 17834 32224
rect 18892 32212 18920 32379
rect 19150 32376 19156 32388
rect 19208 32376 19214 32428
rect 19242 32376 19248 32428
rect 19300 32376 19306 32428
rect 24780 32425 24808 32456
rect 26988 32428 27016 32456
rect 27430 32444 27436 32456
rect 27488 32484 27494 32496
rect 27488 32456 28488 32484
rect 27488 32444 27494 32456
rect 25038 32425 25044 32428
rect 23753 32419 23811 32425
rect 23753 32385 23765 32419
rect 23799 32416 23811 32419
rect 24765 32419 24823 32425
rect 23799 32388 24164 32416
rect 23799 32385 23811 32388
rect 23753 32379 23811 32385
rect 24136 32360 24164 32388
rect 24765 32385 24777 32419
rect 24811 32385 24823 32419
rect 24765 32379 24823 32385
rect 25032 32379 25044 32425
rect 25038 32376 25044 32379
rect 25096 32376 25102 32428
rect 26970 32376 26976 32428
rect 27028 32376 27034 32428
rect 27246 32425 27252 32428
rect 27240 32416 27252 32425
rect 27207 32388 27252 32416
rect 27240 32379 27252 32388
rect 27246 32376 27252 32379
rect 27304 32376 27310 32428
rect 19889 32351 19947 32357
rect 19889 32348 19901 32351
rect 18984 32320 19901 32348
rect 18984 32292 19012 32320
rect 19889 32317 19901 32320
rect 19935 32317 19947 32351
rect 19889 32311 19947 32317
rect 20162 32308 20168 32360
rect 20220 32308 20226 32360
rect 20530 32308 20536 32360
rect 20588 32348 20594 32360
rect 21637 32351 21695 32357
rect 21637 32348 21649 32351
rect 20588 32320 21649 32348
rect 20588 32308 20594 32320
rect 21637 32317 21649 32320
rect 21683 32348 21695 32351
rect 21910 32348 21916 32360
rect 21683 32320 21916 32348
rect 21683 32317 21695 32320
rect 21637 32311 21695 32317
rect 21910 32308 21916 32320
rect 21968 32308 21974 32360
rect 24026 32308 24032 32360
rect 24084 32308 24090 32360
rect 24118 32308 24124 32360
rect 24176 32308 24182 32360
rect 28460 32357 28488 32456
rect 28810 32444 28816 32496
rect 28868 32484 28874 32496
rect 33410 32484 33416 32496
rect 28868 32456 33416 32484
rect 28868 32444 28874 32456
rect 33410 32444 33416 32456
rect 33468 32444 33474 32496
rect 35336 32487 35394 32493
rect 35336 32453 35348 32487
rect 35382 32484 35394 32487
rect 35434 32484 35440 32496
rect 35382 32456 35440 32484
rect 35382 32453 35394 32456
rect 35336 32447 35394 32453
rect 35434 32444 35440 32456
rect 35492 32444 35498 32496
rect 28534 32376 28540 32428
rect 28592 32416 28598 32428
rect 28701 32419 28759 32425
rect 28701 32416 28713 32419
rect 28592 32388 28713 32416
rect 28592 32376 28598 32388
rect 28701 32385 28713 32388
rect 28747 32385 28759 32419
rect 28701 32379 28759 32385
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 29914 32416 29920 32428
rect 29696 32388 29920 32416
rect 29696 32376 29702 32388
rect 29914 32376 29920 32388
rect 29972 32376 29978 32428
rect 33502 32376 33508 32428
rect 33560 32376 33566 32428
rect 33597 32419 33655 32425
rect 33597 32385 33609 32419
rect 33643 32416 33655 32419
rect 33965 32419 34023 32425
rect 33965 32416 33977 32419
rect 33643 32388 33977 32416
rect 33643 32385 33655 32388
rect 33597 32379 33655 32385
rect 33965 32385 33977 32388
rect 34011 32385 34023 32419
rect 33965 32379 34023 32385
rect 34054 32376 34060 32428
rect 34112 32416 34118 32428
rect 34517 32419 34575 32425
rect 34517 32416 34529 32419
rect 34112 32388 34529 32416
rect 34112 32376 34118 32388
rect 34517 32385 34529 32388
rect 34563 32385 34575 32419
rect 34517 32379 34575 32385
rect 34698 32376 34704 32428
rect 34756 32416 34762 32428
rect 35066 32416 35072 32428
rect 34756 32388 35072 32416
rect 34756 32376 34762 32388
rect 35066 32376 35072 32388
rect 35124 32376 35130 32428
rect 37642 32425 37648 32428
rect 37636 32379 37648 32425
rect 37642 32376 37648 32379
rect 37700 32376 37706 32428
rect 38948 32416 38976 32512
rect 40586 32493 40592 32496
rect 40580 32484 40592 32493
rect 40547 32456 40592 32484
rect 40580 32447 40592 32456
rect 40586 32444 40592 32447
rect 40644 32444 40650 32496
rect 39393 32419 39451 32425
rect 39393 32416 39405 32419
rect 38948 32388 39405 32416
rect 39393 32385 39405 32388
rect 39439 32385 39451 32419
rect 39393 32379 39451 32385
rect 40313 32419 40371 32425
rect 40313 32385 40325 32419
rect 40359 32416 40371 32419
rect 40402 32416 40408 32428
rect 40359 32388 40408 32416
rect 40359 32385 40371 32388
rect 40313 32379 40371 32385
rect 40402 32376 40408 32388
rect 40460 32376 40466 32428
rect 41877 32419 41935 32425
rect 41877 32385 41889 32419
rect 41923 32416 41935 32419
rect 41966 32416 41972 32428
rect 41923 32388 41972 32416
rect 41923 32385 41935 32388
rect 41877 32379 41935 32385
rect 41966 32376 41972 32388
rect 42024 32376 42030 32428
rect 28445 32351 28503 32357
rect 28445 32317 28457 32351
rect 28491 32317 28503 32351
rect 30006 32348 30012 32360
rect 28445 32311 28503 32317
rect 29840 32320 30012 32348
rect 18966 32240 18972 32292
rect 19024 32240 19030 32292
rect 19076 32252 19334 32280
rect 19076 32212 19104 32252
rect 17828 32184 19104 32212
rect 19306 32212 19334 32252
rect 20898 32212 20904 32224
rect 19306 32184 20904 32212
rect 17828 32172 17834 32184
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21818 32172 21824 32224
rect 21876 32212 21882 32224
rect 28350 32212 28356 32224
rect 21876 32184 28356 32212
rect 21876 32172 21882 32184
rect 28350 32172 28356 32184
rect 28408 32172 28414 32224
rect 28460 32212 28488 32311
rect 29840 32289 29868 32320
rect 30006 32308 30012 32320
rect 30064 32348 30070 32360
rect 31205 32351 31263 32357
rect 31205 32348 31217 32351
rect 30064 32320 31217 32348
rect 30064 32308 30070 32320
rect 31205 32317 31217 32320
rect 31251 32317 31263 32351
rect 31205 32311 31263 32317
rect 32122 32308 32128 32360
rect 32180 32308 32186 32360
rect 33781 32351 33839 32357
rect 33781 32317 33793 32351
rect 33827 32348 33839 32351
rect 34238 32348 34244 32360
rect 33827 32320 34244 32348
rect 33827 32317 33839 32320
rect 33781 32311 33839 32317
rect 34238 32308 34244 32320
rect 34296 32308 34302 32360
rect 37366 32308 37372 32360
rect 37424 32308 37430 32360
rect 29825 32283 29883 32289
rect 29825 32249 29837 32283
rect 29871 32249 29883 32283
rect 29825 32243 29883 32249
rect 31294 32240 31300 32292
rect 31352 32280 31358 32292
rect 33042 32280 33048 32292
rect 31352 32252 33048 32280
rect 31352 32240 31358 32252
rect 33042 32240 33048 32252
rect 33100 32240 33106 32292
rect 29454 32212 29460 32224
rect 28460 32184 29460 32212
rect 29454 32172 29460 32184
rect 29512 32172 29518 32224
rect 30558 32172 30564 32224
rect 30616 32172 30622 32224
rect 30650 32172 30656 32224
rect 30708 32172 30714 32224
rect 31018 32172 31024 32224
rect 31076 32212 31082 32224
rect 31386 32212 31392 32224
rect 31076 32184 31392 32212
rect 31076 32172 31082 32184
rect 31386 32172 31392 32184
rect 31444 32172 31450 32224
rect 32766 32172 32772 32224
rect 32824 32172 32830 32224
rect 38286 32172 38292 32224
rect 38344 32212 38350 32224
rect 38841 32215 38899 32221
rect 38841 32212 38853 32215
rect 38344 32184 38853 32212
rect 38344 32172 38350 32184
rect 38841 32181 38853 32184
rect 38887 32181 38899 32215
rect 38841 32175 38899 32181
rect 42058 32172 42064 32224
rect 42116 32172 42122 32224
rect 1104 32122 42504 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 42504 32122
rect 1104 32048 42504 32070
rect 3050 31968 3056 32020
rect 3108 32008 3114 32020
rect 3145 32011 3203 32017
rect 3145 32008 3157 32011
rect 3108 31980 3157 32008
rect 3108 31968 3114 31980
rect 3145 31977 3157 31980
rect 3191 31977 3203 32011
rect 3145 31971 3203 31977
rect 4706 31968 4712 32020
rect 4764 31968 4770 32020
rect 5350 31968 5356 32020
rect 5408 32008 5414 32020
rect 5629 32011 5687 32017
rect 5629 32008 5641 32011
rect 5408 31980 5641 32008
rect 5408 31968 5414 31980
rect 5629 31977 5641 31980
rect 5675 31977 5687 32011
rect 5629 31971 5687 31977
rect 5718 31968 5724 32020
rect 5776 32008 5782 32020
rect 6362 32008 6368 32020
rect 5776 31980 6368 32008
rect 5776 31968 5782 31980
rect 6362 31968 6368 31980
rect 6420 31968 6426 32020
rect 6641 32011 6699 32017
rect 6641 31977 6653 32011
rect 6687 32008 6699 32011
rect 7374 32008 7380 32020
rect 6687 31980 7380 32008
rect 6687 31977 6699 31980
rect 6641 31971 6699 31977
rect 7374 31968 7380 31980
rect 7432 31968 7438 32020
rect 8202 31968 8208 32020
rect 8260 32008 8266 32020
rect 8665 32011 8723 32017
rect 8665 32008 8677 32011
rect 8260 31980 8677 32008
rect 8260 31968 8266 31980
rect 8665 31977 8677 31980
rect 8711 31977 8723 32011
rect 8665 31971 8723 31977
rect 9306 31968 9312 32020
rect 9364 31968 9370 32020
rect 12345 32011 12403 32017
rect 12345 31977 12357 32011
rect 12391 32008 12403 32011
rect 12894 32008 12900 32020
rect 12391 31980 12900 32008
rect 12391 31977 12403 31980
rect 12345 31971 12403 31977
rect 12894 31968 12900 31980
rect 12952 31968 12958 32020
rect 13538 31968 13544 32020
rect 13596 31968 13602 32020
rect 15194 31968 15200 32020
rect 15252 32008 15258 32020
rect 15657 32011 15715 32017
rect 15657 32008 15669 32011
rect 15252 31980 15669 32008
rect 15252 31968 15258 31980
rect 15657 31977 15669 31980
rect 15703 31977 15715 32011
rect 15657 31971 15715 31977
rect 16022 31968 16028 32020
rect 16080 32008 16086 32020
rect 16117 32011 16175 32017
rect 16117 32008 16129 32011
rect 16080 31980 16129 32008
rect 16080 31968 16086 31980
rect 16117 31977 16129 31980
rect 16163 31977 16175 32011
rect 16117 31971 16175 31977
rect 16758 31968 16764 32020
rect 16816 32008 16822 32020
rect 16816 31980 18000 32008
rect 16816 31968 16822 31980
rect 5902 31940 5908 31952
rect 5552 31912 5908 31940
rect 4798 31832 4804 31884
rect 4856 31872 4862 31884
rect 4985 31875 5043 31881
rect 4985 31872 4997 31875
rect 4856 31844 4997 31872
rect 4856 31832 4862 31844
rect 4985 31841 4997 31844
rect 5031 31841 5043 31875
rect 4985 31835 5043 31841
rect 5077 31875 5135 31881
rect 5077 31841 5089 31875
rect 5123 31872 5135 31875
rect 5445 31875 5503 31881
rect 5445 31872 5457 31875
rect 5123 31844 5457 31872
rect 5123 31841 5135 31844
rect 5077 31835 5135 31841
rect 5445 31841 5457 31844
rect 5491 31841 5503 31875
rect 5445 31835 5503 31841
rect 3329 31807 3387 31813
rect 3329 31773 3341 31807
rect 3375 31804 3387 31807
rect 3418 31804 3424 31816
rect 3375 31776 3424 31804
rect 3375 31773 3387 31776
rect 3329 31767 3387 31773
rect 3418 31764 3424 31776
rect 3476 31764 3482 31816
rect 4893 31807 4951 31813
rect 4893 31804 4905 31807
rect 4871 31776 4905 31804
rect 4893 31773 4905 31776
rect 4939 31773 4951 31807
rect 4893 31767 4951 31773
rect 5169 31807 5227 31813
rect 5169 31773 5181 31807
rect 5215 31804 5227 31807
rect 5258 31804 5264 31816
rect 5215 31776 5264 31804
rect 5215 31773 5227 31776
rect 5169 31767 5227 31773
rect 4908 31736 4936 31767
rect 5258 31764 5264 31776
rect 5316 31764 5322 31816
rect 5552 31813 5580 31912
rect 5902 31900 5908 31912
rect 5960 31900 5966 31952
rect 16301 31943 16359 31949
rect 16301 31940 16313 31943
rect 16040 31912 16313 31940
rect 6362 31832 6368 31884
rect 6420 31872 6426 31884
rect 7742 31872 7748 31884
rect 6420 31844 7748 31872
rect 6420 31832 6426 31844
rect 7742 31832 7748 31844
rect 7800 31832 7806 31884
rect 10410 31832 10416 31884
rect 10468 31872 10474 31884
rect 11149 31875 11207 31881
rect 11149 31872 11161 31875
rect 10468 31844 11161 31872
rect 10468 31832 10474 31844
rect 11149 31841 11161 31844
rect 11195 31841 11207 31875
rect 11149 31835 11207 31841
rect 11716 31844 12388 31872
rect 5537 31807 5595 31813
rect 5537 31773 5549 31807
rect 5583 31773 5595 31807
rect 5537 31767 5595 31773
rect 5626 31764 5632 31816
rect 5684 31764 5690 31816
rect 5813 31807 5871 31813
rect 5813 31804 5825 31807
rect 5791 31776 5825 31804
rect 5813 31773 5825 31776
rect 5859 31806 5871 31807
rect 5859 31804 5948 31806
rect 6380 31804 6408 31832
rect 6638 31804 6644 31816
rect 5859 31778 6408 31804
rect 5859 31773 5871 31778
rect 5920 31776 6408 31778
rect 6619 31776 6644 31804
rect 5813 31767 5871 31773
rect 5350 31736 5356 31748
rect 4908 31708 5356 31736
rect 5350 31696 5356 31708
rect 5408 31736 5414 31748
rect 5828 31736 5856 31767
rect 6638 31764 6644 31776
rect 6696 31764 6702 31816
rect 6822 31764 6828 31816
rect 6880 31764 6886 31816
rect 6914 31764 6920 31816
rect 6972 31764 6978 31816
rect 11057 31807 11115 31813
rect 11057 31773 11069 31807
rect 11103 31773 11115 31807
rect 11057 31767 11115 31773
rect 5408 31708 5856 31736
rect 5408 31696 5414 31708
rect 5994 31696 6000 31748
rect 6052 31736 6058 31748
rect 6656 31736 6684 31764
rect 6052 31708 6684 31736
rect 6052 31696 6058 31708
rect 7190 31696 7196 31748
rect 7248 31696 7254 31748
rect 8418 31708 8524 31736
rect 10350 31708 10456 31736
rect 3970 31628 3976 31680
rect 4028 31668 4034 31680
rect 6012 31668 6040 31696
rect 4028 31640 6040 31668
rect 4028 31628 4034 31640
rect 8202 31628 8208 31680
rect 8260 31668 8266 31680
rect 8496 31668 8524 31708
rect 10428 31668 10456 31708
rect 10778 31696 10784 31748
rect 10836 31696 10842 31748
rect 10870 31696 10876 31748
rect 10928 31736 10934 31748
rect 11072 31736 11100 31767
rect 11514 31764 11520 31816
rect 11572 31804 11578 31816
rect 11716 31813 11744 31844
rect 11701 31807 11759 31813
rect 11701 31804 11713 31807
rect 11572 31776 11713 31804
rect 11572 31764 11578 31776
rect 11701 31773 11713 31776
rect 11747 31773 11759 31807
rect 11701 31767 11759 31773
rect 12158 31764 12164 31816
rect 12216 31764 12222 31816
rect 12360 31813 12388 31844
rect 12345 31807 12403 31813
rect 12345 31773 12357 31807
rect 12391 31773 12403 31807
rect 12345 31767 12403 31773
rect 13814 31764 13820 31816
rect 13872 31764 13878 31816
rect 15838 31764 15844 31816
rect 15896 31764 15902 31816
rect 15933 31807 15991 31813
rect 15933 31773 15945 31807
rect 15979 31804 15991 31807
rect 16040 31804 16068 31912
rect 16301 31909 16313 31912
rect 16347 31909 16359 31943
rect 16301 31903 16359 31909
rect 16942 31900 16948 31952
rect 17000 31940 17006 31952
rect 17037 31943 17095 31949
rect 17037 31940 17049 31943
rect 17000 31912 17049 31940
rect 17000 31900 17006 31912
rect 17037 31909 17049 31912
rect 17083 31909 17095 31943
rect 17037 31903 17095 31909
rect 17972 31872 18000 31980
rect 18046 31968 18052 32020
rect 18104 31968 18110 32020
rect 18782 31968 18788 32020
rect 18840 32008 18846 32020
rect 21174 32008 21180 32020
rect 18840 31980 21180 32008
rect 18840 31968 18846 31980
rect 21174 31968 21180 31980
rect 21232 32008 21238 32020
rect 21821 32011 21879 32017
rect 21821 32008 21833 32011
rect 21232 31980 21833 32008
rect 21232 31968 21238 31980
rect 21821 31977 21833 31980
rect 21867 32008 21879 32011
rect 21867 31980 22094 32008
rect 21867 31977 21879 31980
rect 21821 31971 21879 31977
rect 20162 31900 20168 31952
rect 20220 31940 20226 31952
rect 21269 31943 21327 31949
rect 20220 31912 21220 31940
rect 20220 31900 20226 31912
rect 18877 31875 18935 31881
rect 18877 31872 18889 31875
rect 16500 31844 17080 31872
rect 17972 31844 18460 31872
rect 15979 31776 16068 31804
rect 16209 31807 16267 31813
rect 15979 31773 15991 31776
rect 15933 31767 15991 31773
rect 16209 31773 16221 31807
rect 16255 31804 16267 31807
rect 16390 31804 16396 31816
rect 16255 31776 16396 31804
rect 16255 31773 16267 31776
rect 16209 31767 16267 31773
rect 16390 31764 16396 31776
rect 16448 31764 16454 31816
rect 16500 31813 16528 31844
rect 16485 31807 16543 31813
rect 16485 31773 16497 31807
rect 16531 31773 16543 31807
rect 16485 31767 16543 31773
rect 16574 31764 16580 31816
rect 16632 31764 16638 31816
rect 16669 31807 16727 31813
rect 16669 31773 16681 31807
rect 16715 31804 16727 31807
rect 16758 31804 16764 31816
rect 16715 31776 16764 31804
rect 16715 31773 16727 31776
rect 16669 31767 16727 31773
rect 16758 31764 16764 31776
rect 16816 31764 16822 31816
rect 16850 31764 16856 31816
rect 16908 31764 16914 31816
rect 10928 31708 11100 31736
rect 11885 31739 11943 31745
rect 10928 31696 10934 31708
rect 11885 31705 11897 31739
rect 11931 31736 11943 31739
rect 12066 31736 12072 31748
rect 11931 31708 12072 31736
rect 11931 31705 11943 31708
rect 11885 31699 11943 31705
rect 12066 31696 12072 31708
rect 12124 31696 12130 31748
rect 16408 31736 16436 31764
rect 17052 31736 17080 31844
rect 17126 31764 17132 31816
rect 17184 31804 17190 31816
rect 17221 31807 17279 31813
rect 17221 31804 17233 31807
rect 17184 31776 17233 31804
rect 17184 31764 17190 31776
rect 17221 31773 17233 31776
rect 17267 31773 17279 31807
rect 17221 31767 17279 31773
rect 17310 31764 17316 31816
rect 17368 31764 17374 31816
rect 17402 31764 17408 31816
rect 17460 31804 17466 31816
rect 17497 31807 17555 31813
rect 17497 31804 17509 31807
rect 17460 31776 17509 31804
rect 17460 31764 17466 31776
rect 17497 31773 17509 31776
rect 17543 31773 17555 31807
rect 18046 31804 18052 31816
rect 17497 31767 17555 31773
rect 17604 31776 18052 31804
rect 17604 31736 17632 31776
rect 18046 31764 18052 31776
rect 18104 31804 18110 31816
rect 18187 31807 18245 31813
rect 18187 31804 18199 31807
rect 18104 31776 18199 31804
rect 18104 31764 18110 31776
rect 18187 31773 18199 31776
rect 18233 31773 18245 31807
rect 18187 31767 18245 31773
rect 18322 31764 18328 31816
rect 18380 31764 18386 31816
rect 18432 31813 18460 31844
rect 18708 31844 18889 31872
rect 18417 31807 18475 31813
rect 18417 31773 18429 31807
rect 18463 31804 18475 31807
rect 18463 31776 18517 31804
rect 18463 31773 18475 31776
rect 18417 31767 18475 31773
rect 16408 31708 16712 31736
rect 17052 31708 17632 31736
rect 16684 31680 16712 31708
rect 10962 31668 10968 31680
rect 8260 31640 10968 31668
rect 8260 31628 8266 31640
rect 10962 31628 10968 31640
rect 11020 31628 11026 31680
rect 12529 31671 12587 31677
rect 12529 31637 12541 31671
rect 12575 31668 12587 31671
rect 13446 31668 13452 31680
rect 12575 31640 13452 31668
rect 12575 31637 12587 31640
rect 12529 31631 12587 31637
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 16666 31628 16672 31680
rect 16724 31668 16730 31680
rect 17310 31668 17316 31680
rect 16724 31640 17316 31668
rect 16724 31628 16730 31640
rect 17310 31628 17316 31640
rect 17368 31628 17374 31680
rect 17405 31671 17463 31677
rect 17405 31637 17417 31671
rect 17451 31668 17463 31671
rect 17678 31668 17684 31680
rect 17451 31640 17684 31668
rect 17451 31637 17463 31640
rect 17405 31631 17463 31637
rect 17678 31628 17684 31640
rect 17736 31628 17742 31680
rect 18432 31668 18460 31767
rect 18598 31764 18604 31816
rect 18656 31764 18662 31816
rect 18708 31813 18736 31844
rect 18877 31841 18889 31844
rect 18923 31841 18935 31875
rect 18877 31835 18935 31841
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31773 18751 31807
rect 18693 31767 18751 31773
rect 18782 31764 18788 31816
rect 18840 31764 18846 31816
rect 18969 31807 19027 31813
rect 18969 31773 18981 31807
rect 19015 31804 19027 31807
rect 19426 31804 19432 31816
rect 19015 31776 19432 31804
rect 19015 31773 19027 31776
rect 18969 31767 19027 31773
rect 19426 31764 19432 31776
rect 19484 31764 19490 31816
rect 20717 31807 20775 31813
rect 20717 31773 20729 31807
rect 20763 31804 20775 31807
rect 20806 31804 20812 31816
rect 20763 31776 20812 31804
rect 20763 31773 20775 31776
rect 20717 31767 20775 31773
rect 20806 31764 20812 31776
rect 20864 31764 20870 31816
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31773 20959 31807
rect 20901 31767 20959 31773
rect 19610 31696 19616 31748
rect 19668 31736 19674 31748
rect 20916 31736 20944 31767
rect 20990 31764 20996 31816
rect 21048 31764 21054 31816
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31773 21143 31807
rect 21192 31804 21220 31912
rect 21269 31909 21281 31943
rect 21315 31940 21327 31943
rect 21450 31940 21456 31952
rect 21315 31912 21456 31940
rect 21315 31909 21327 31912
rect 21269 31903 21327 31909
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 22066 31872 22094 31980
rect 25038 31968 25044 32020
rect 25096 32008 25102 32020
rect 25225 32011 25283 32017
rect 25225 32008 25237 32011
rect 25096 31980 25237 32008
rect 25096 31968 25102 31980
rect 25225 31977 25237 31980
rect 25271 31977 25283 32011
rect 25225 31971 25283 31977
rect 26694 31968 26700 32020
rect 26752 32008 26758 32020
rect 27522 32008 27528 32020
rect 26752 31980 27528 32008
rect 26752 31968 26758 31980
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 28534 31968 28540 32020
rect 28592 31968 28598 32020
rect 30650 32008 30656 32020
rect 29012 31980 30656 32008
rect 27801 31943 27859 31949
rect 27801 31909 27813 31943
rect 27847 31940 27859 31943
rect 28626 31940 28632 31952
rect 27847 31912 28632 31940
rect 27847 31909 27859 31912
rect 27801 31903 27859 31909
rect 28626 31900 28632 31912
rect 28684 31900 28690 31952
rect 24029 31875 24087 31881
rect 24029 31872 24041 31875
rect 22066 31844 24041 31872
rect 24029 31841 24041 31844
rect 24075 31872 24087 31875
rect 25498 31872 25504 31884
rect 24075 31844 25504 31872
rect 24075 31841 24087 31844
rect 24029 31835 24087 31841
rect 25498 31832 25504 31844
rect 25556 31832 25562 31884
rect 25682 31832 25688 31884
rect 25740 31832 25746 31884
rect 25774 31832 25780 31884
rect 25832 31832 25838 31884
rect 29012 31881 29040 31980
rect 30650 31968 30656 31980
rect 30708 31968 30714 32020
rect 31021 32011 31079 32017
rect 31021 31977 31033 32011
rect 31067 32008 31079 32011
rect 32122 32008 32128 32020
rect 31067 31980 32128 32008
rect 31067 31977 31079 31980
rect 31021 31971 31079 31977
rect 32122 31968 32128 31980
rect 32180 31968 32186 32020
rect 35342 31968 35348 32020
rect 35400 32008 35406 32020
rect 35437 32011 35495 32017
rect 35437 32008 35449 32011
rect 35400 31980 35449 32008
rect 35400 31968 35406 31980
rect 35437 31977 35449 31980
rect 35483 31977 35495 32011
rect 35437 31971 35495 31977
rect 37642 31968 37648 32020
rect 37700 32008 37706 32020
rect 37829 32011 37887 32017
rect 37829 32008 37841 32011
rect 37700 31980 37841 32008
rect 37700 31968 37706 31980
rect 37829 31977 37841 31980
rect 37875 31977 37887 32011
rect 41325 32011 41383 32017
rect 41325 32008 41337 32011
rect 37829 31971 37887 31977
rect 39224 31980 41337 32008
rect 33778 31900 33784 31952
rect 33836 31940 33842 31952
rect 33965 31943 34023 31949
rect 33965 31940 33977 31943
rect 33836 31912 33977 31940
rect 33836 31900 33842 31912
rect 33965 31909 33977 31912
rect 34011 31909 34023 31943
rect 33965 31903 34023 31909
rect 26421 31875 26479 31881
rect 26421 31841 26433 31875
rect 26467 31841 26479 31875
rect 26421 31835 26479 31841
rect 28997 31875 29055 31881
rect 28997 31841 29009 31875
rect 29043 31841 29055 31875
rect 28997 31835 29055 31841
rect 29089 31875 29147 31881
rect 29089 31841 29101 31875
rect 29135 31841 29147 31875
rect 29089 31835 29147 31841
rect 21361 31807 21419 31813
rect 21361 31804 21373 31807
rect 21192 31776 21373 31804
rect 21085 31767 21143 31773
rect 21361 31773 21373 31776
rect 21407 31773 21419 31807
rect 21361 31767 21419 31773
rect 21100 31736 21128 31767
rect 21542 31764 21548 31816
rect 21600 31764 21606 31816
rect 21634 31764 21640 31816
rect 21692 31764 21698 31816
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 23750 31764 23756 31816
rect 23808 31764 23814 31816
rect 23842 31764 23848 31816
rect 23900 31764 23906 31816
rect 24118 31764 24124 31816
rect 24176 31764 24182 31816
rect 26436 31804 26464 31835
rect 26970 31804 26976 31816
rect 26436 31776 26976 31804
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 27522 31764 27528 31816
rect 27580 31804 27586 31816
rect 29104 31804 29132 31835
rect 29454 31832 29460 31884
rect 29512 31872 29518 31884
rect 29549 31875 29607 31881
rect 29549 31872 29561 31875
rect 29512 31844 29561 31872
rect 29512 31832 29518 31844
rect 29549 31841 29561 31844
rect 29595 31841 29607 31875
rect 33980 31872 34008 31903
rect 34238 31900 34244 31952
rect 34296 31940 34302 31952
rect 34296 31912 38424 31940
rect 34296 31900 34302 31912
rect 35253 31875 35311 31881
rect 35253 31872 35265 31875
rect 33980 31844 35265 31872
rect 29549 31835 29607 31841
rect 35253 31841 35265 31844
rect 35299 31841 35311 31875
rect 35253 31835 35311 31841
rect 35802 31832 35808 31884
rect 35860 31872 35866 31884
rect 35989 31875 36047 31881
rect 35989 31872 36001 31875
rect 35860 31844 36001 31872
rect 35860 31832 35866 31844
rect 35989 31841 36001 31844
rect 36035 31841 36047 31875
rect 35989 31835 36047 31841
rect 36814 31832 36820 31884
rect 36872 31832 36878 31884
rect 38286 31832 38292 31884
rect 38344 31832 38350 31884
rect 38396 31881 38424 31912
rect 38381 31875 38439 31881
rect 38381 31841 38393 31875
rect 38427 31872 38439 31875
rect 39022 31872 39028 31884
rect 38427 31844 39028 31872
rect 38427 31841 38439 31844
rect 38381 31835 38439 31841
rect 39022 31832 39028 31844
rect 39080 31832 39086 31884
rect 39224 31881 39252 31980
rect 41325 31977 41337 31980
rect 41371 31977 41383 32011
rect 41325 31971 41383 31977
rect 41230 31900 41236 31952
rect 41288 31940 41294 31952
rect 41288 31912 41920 31940
rect 41288 31900 41294 31912
rect 41892 31881 41920 31912
rect 39209 31875 39267 31881
rect 39209 31841 39221 31875
rect 39255 31841 39267 31875
rect 39209 31835 39267 31841
rect 41877 31875 41935 31881
rect 41877 31841 41889 31875
rect 41923 31841 41935 31875
rect 41877 31835 41935 31841
rect 29816 31807 29874 31813
rect 27580 31776 29316 31804
rect 27580 31764 27586 31776
rect 21450 31736 21456 31748
rect 19668 31708 21066 31736
rect 21100 31708 21456 31736
rect 19668 31696 19674 31708
rect 20714 31668 20720 31680
rect 18432 31640 20720 31668
rect 20714 31628 20720 31640
rect 20772 31628 20778 31680
rect 21038 31668 21066 31708
rect 21450 31696 21456 31708
rect 21508 31696 21514 31748
rect 26234 31696 26240 31748
rect 26292 31736 26298 31748
rect 26666 31739 26724 31745
rect 26666 31736 26678 31739
rect 26292 31708 26678 31736
rect 26292 31696 26298 31708
rect 26666 31705 26678 31708
rect 26712 31705 26724 31739
rect 29288 31736 29316 31776
rect 29816 31773 29828 31807
rect 29862 31804 29874 31807
rect 30374 31804 30380 31816
rect 29862 31776 30380 31804
rect 29862 31773 29874 31776
rect 29816 31767 29874 31773
rect 30374 31764 30380 31776
rect 30432 31764 30438 31816
rect 31202 31764 31208 31816
rect 31260 31804 31266 31816
rect 32401 31807 32459 31813
rect 32401 31804 32413 31807
rect 31260 31776 32413 31804
rect 31260 31764 31266 31776
rect 32401 31773 32413 31776
rect 32447 31804 32459 31807
rect 32585 31807 32643 31813
rect 32585 31804 32597 31807
rect 32447 31776 32597 31804
rect 32447 31773 32459 31776
rect 32401 31767 32459 31773
rect 32585 31773 32597 31776
rect 32631 31773 32643 31807
rect 32585 31767 32643 31773
rect 32852 31807 32910 31813
rect 32852 31773 32864 31807
rect 32898 31804 32910 31807
rect 33318 31804 33324 31816
rect 32898 31776 33324 31804
rect 32898 31773 32910 31776
rect 32852 31767 32910 31773
rect 33318 31764 33324 31776
rect 33376 31764 33382 31816
rect 33410 31764 33416 31816
rect 33468 31804 33474 31816
rect 34057 31807 34115 31813
rect 34057 31804 34069 31807
rect 33468 31776 34069 31804
rect 33468 31764 33474 31776
rect 34057 31773 34069 31776
rect 34103 31773 34115 31807
rect 34057 31767 34115 31773
rect 35897 31807 35955 31813
rect 35897 31773 35909 31807
rect 35943 31804 35955 31807
rect 36265 31807 36323 31813
rect 36265 31804 36277 31807
rect 35943 31776 36277 31804
rect 35943 31773 35955 31776
rect 35897 31767 35955 31773
rect 36265 31773 36277 31776
rect 36311 31773 36323 31807
rect 36265 31767 36323 31773
rect 37366 31764 37372 31816
rect 37424 31804 37430 31816
rect 39853 31807 39911 31813
rect 39853 31804 39865 31807
rect 37424 31776 39865 31804
rect 37424 31764 37430 31776
rect 39853 31773 39865 31776
rect 39899 31804 39911 31807
rect 40402 31804 40408 31816
rect 39899 31776 40408 31804
rect 39899 31773 39911 31776
rect 39853 31767 39911 31773
rect 40402 31764 40408 31776
rect 40460 31764 40466 31816
rect 30190 31736 30196 31748
rect 29288 31708 30196 31736
rect 26666 31699 26724 31705
rect 30190 31696 30196 31708
rect 30248 31696 30254 31748
rect 32122 31696 32128 31748
rect 32180 31745 32186 31748
rect 32180 31699 32192 31745
rect 40098 31739 40156 31745
rect 40098 31736 40110 31739
rect 39684 31708 40110 31736
rect 32180 31696 32186 31699
rect 22370 31668 22376 31680
rect 21038 31640 22376 31668
rect 22370 31628 22376 31640
rect 22428 31628 22434 31680
rect 23474 31628 23480 31680
rect 23532 31668 23538 31680
rect 23569 31671 23627 31677
rect 23569 31668 23581 31671
rect 23532 31640 23581 31668
rect 23532 31628 23538 31640
rect 23569 31637 23581 31640
rect 23615 31637 23627 31671
rect 23569 31631 23627 31637
rect 25590 31628 25596 31680
rect 25648 31628 25654 31680
rect 28905 31671 28963 31677
rect 28905 31637 28917 31671
rect 28951 31668 28963 31671
rect 30006 31668 30012 31680
rect 28951 31640 30012 31668
rect 28951 31637 28963 31640
rect 28905 31631 28963 31637
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 30929 31671 30987 31677
rect 30929 31637 30941 31671
rect 30975 31668 30987 31671
rect 31570 31668 31576 31680
rect 30975 31640 31576 31668
rect 30975 31637 30987 31640
rect 30929 31631 30987 31637
rect 31570 31628 31576 31640
rect 31628 31628 31634 31680
rect 32582 31628 32588 31680
rect 32640 31668 32646 31680
rect 32858 31668 32864 31680
rect 32640 31640 32864 31668
rect 32640 31628 32646 31640
rect 32858 31628 32864 31640
rect 32916 31628 32922 31680
rect 34514 31628 34520 31680
rect 34572 31668 34578 31680
rect 34701 31671 34759 31677
rect 34701 31668 34713 31671
rect 34572 31640 34713 31668
rect 34572 31628 34578 31640
rect 34701 31637 34713 31640
rect 34747 31637 34759 31671
rect 34701 31631 34759 31637
rect 35805 31671 35863 31677
rect 35805 31637 35817 31671
rect 35851 31668 35863 31671
rect 35986 31668 35992 31680
rect 35851 31640 35992 31668
rect 35851 31637 35863 31640
rect 35805 31631 35863 31637
rect 35986 31628 35992 31640
rect 36044 31628 36050 31680
rect 36078 31628 36084 31680
rect 36136 31668 36142 31680
rect 38197 31671 38255 31677
rect 38197 31668 38209 31671
rect 36136 31640 38209 31668
rect 36136 31628 36142 31640
rect 38197 31637 38209 31640
rect 38243 31637 38255 31671
rect 38197 31631 38255 31637
rect 38286 31628 38292 31680
rect 38344 31668 38350 31680
rect 39684 31677 39712 31708
rect 40098 31705 40110 31708
rect 40144 31705 40156 31739
rect 40098 31699 40156 31705
rect 39301 31671 39359 31677
rect 39301 31668 39313 31671
rect 38344 31640 39313 31668
rect 38344 31628 38350 31640
rect 39301 31637 39313 31640
rect 39347 31637 39359 31671
rect 39301 31631 39359 31637
rect 39669 31671 39727 31677
rect 39669 31637 39681 31671
rect 39715 31637 39727 31671
rect 39669 31631 39727 31637
rect 1104 31578 42504 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 42504 31578
rect 1104 31504 42504 31526
rect 2590 31424 2596 31476
rect 2648 31424 2654 31476
rect 3602 31424 3608 31476
rect 3660 31464 3666 31476
rect 3907 31467 3965 31473
rect 3907 31464 3919 31467
rect 3660 31436 3919 31464
rect 3660 31424 3666 31436
rect 3907 31433 3919 31436
rect 3953 31464 3965 31467
rect 4062 31464 4068 31476
rect 3953 31436 4068 31464
rect 3953 31433 3965 31436
rect 3907 31427 3965 31433
rect 4062 31424 4068 31436
rect 4120 31464 4126 31476
rect 5166 31464 5172 31476
rect 4120 31436 5172 31464
rect 4120 31424 4126 31436
rect 5166 31424 5172 31436
rect 5224 31424 5230 31476
rect 5350 31473 5356 31476
rect 5337 31467 5356 31473
rect 5337 31433 5349 31467
rect 5337 31427 5356 31433
rect 5350 31424 5356 31427
rect 5408 31424 5414 31476
rect 5813 31467 5871 31473
rect 5813 31464 5825 31467
rect 5552 31436 5825 31464
rect 2866 31356 2872 31408
rect 2924 31396 2930 31408
rect 3510 31396 3516 31408
rect 2924 31368 3516 31396
rect 2924 31356 2930 31368
rect 3510 31356 3516 31368
rect 3568 31396 3574 31408
rect 5552 31405 5580 31436
rect 5813 31433 5825 31436
rect 5859 31464 5871 31467
rect 5902 31464 5908 31476
rect 5859 31436 5908 31464
rect 5859 31433 5871 31436
rect 5813 31427 5871 31433
rect 5902 31424 5908 31436
rect 5960 31424 5966 31476
rect 7190 31424 7196 31476
rect 7248 31464 7254 31476
rect 7561 31467 7619 31473
rect 7561 31464 7573 31467
rect 7248 31436 7573 31464
rect 7248 31424 7254 31436
rect 7561 31433 7573 31436
rect 7607 31433 7619 31467
rect 8662 31464 8668 31476
rect 7561 31427 7619 31433
rect 7852 31436 8668 31464
rect 3697 31399 3755 31405
rect 3697 31396 3709 31399
rect 3568 31368 3709 31396
rect 3568 31356 3574 31368
rect 3697 31365 3709 31368
rect 3743 31365 3755 31399
rect 3697 31359 3755 31365
rect 5537 31399 5595 31405
rect 5537 31365 5549 31399
rect 5583 31365 5595 31399
rect 5537 31359 5595 31365
rect 5629 31399 5687 31405
rect 5629 31365 5641 31399
rect 5675 31396 5687 31399
rect 6086 31396 6092 31408
rect 5675 31368 6092 31396
rect 5675 31365 5687 31368
rect 5629 31359 5687 31365
rect 6086 31356 6092 31368
rect 6144 31356 6150 31408
rect 2501 31331 2559 31337
rect 2501 31297 2513 31331
rect 2547 31328 2559 31331
rect 3234 31328 3240 31340
rect 2547 31300 3240 31328
rect 2547 31297 2559 31300
rect 2501 31291 2559 31297
rect 3234 31288 3240 31300
rect 3292 31288 3298 31340
rect 5810 31328 5816 31340
rect 3620 31300 5816 31328
rect 2777 31263 2835 31269
rect 2777 31229 2789 31263
rect 2823 31260 2835 31263
rect 2961 31263 3019 31269
rect 2961 31260 2973 31263
rect 2823 31232 2973 31260
rect 2823 31229 2835 31232
rect 2777 31223 2835 31229
rect 2961 31229 2973 31232
rect 3007 31229 3019 31263
rect 2961 31223 3019 31229
rect 3142 31220 3148 31272
rect 3200 31260 3206 31272
rect 3513 31263 3571 31269
rect 3513 31260 3525 31263
rect 3200 31232 3525 31260
rect 3200 31220 3206 31232
rect 3513 31229 3525 31232
rect 3559 31229 3571 31263
rect 3513 31223 3571 31229
rect 3050 31152 3056 31204
rect 3108 31192 3114 31204
rect 3620 31192 3648 31300
rect 5810 31288 5816 31300
rect 5868 31288 5874 31340
rect 5905 31331 5963 31337
rect 5905 31297 5917 31331
rect 5951 31328 5963 31331
rect 6362 31328 6368 31340
rect 5951 31300 6368 31328
rect 5951 31297 5963 31300
rect 5905 31291 5963 31297
rect 6362 31288 6368 31300
rect 6420 31288 6426 31340
rect 6457 31331 6515 31337
rect 6457 31297 6469 31331
rect 6503 31297 6515 31331
rect 6457 31291 6515 31297
rect 4614 31220 4620 31272
rect 4672 31260 4678 31272
rect 6472 31260 6500 31291
rect 7742 31288 7748 31340
rect 7800 31288 7806 31340
rect 7852 31337 7880 31436
rect 8662 31424 8668 31436
rect 8720 31424 8726 31476
rect 12345 31467 12403 31473
rect 12345 31433 12357 31467
rect 12391 31464 12403 31467
rect 13814 31464 13820 31476
rect 12391 31436 13820 31464
rect 12391 31433 12403 31436
rect 12345 31427 12403 31433
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 15286 31464 15292 31476
rect 14384 31436 15292 31464
rect 8018 31356 8024 31408
rect 8076 31396 8082 31408
rect 8113 31399 8171 31405
rect 8113 31396 8125 31399
rect 8076 31368 8125 31396
rect 8076 31356 8082 31368
rect 8113 31365 8125 31368
rect 8159 31365 8171 31399
rect 10962 31396 10968 31408
rect 10810 31368 10968 31396
rect 8113 31359 8171 31365
rect 10962 31356 10968 31368
rect 11020 31356 11026 31408
rect 14384 31396 14412 31436
rect 15286 31424 15292 31436
rect 15344 31424 15350 31476
rect 15378 31424 15384 31476
rect 15436 31464 15442 31476
rect 15473 31467 15531 31473
rect 15473 31464 15485 31467
rect 15436 31436 15485 31464
rect 15436 31424 15442 31436
rect 15473 31433 15485 31436
rect 15519 31433 15531 31467
rect 15473 31427 15531 31433
rect 15930 31424 15936 31476
rect 15988 31424 15994 31476
rect 17034 31424 17040 31476
rect 17092 31424 17098 31476
rect 17129 31467 17187 31473
rect 17129 31433 17141 31467
rect 17175 31464 17187 31467
rect 17310 31464 17316 31476
rect 17175 31436 17316 31464
rect 17175 31433 17187 31436
rect 17129 31427 17187 31433
rect 17310 31424 17316 31436
rect 17368 31424 17374 31476
rect 18049 31467 18107 31473
rect 18049 31433 18061 31467
rect 18095 31464 18107 31467
rect 19058 31464 19064 31476
rect 18095 31436 19064 31464
rect 18095 31433 18107 31436
rect 18049 31427 18107 31433
rect 19058 31424 19064 31436
rect 19116 31424 19122 31476
rect 19610 31424 19616 31476
rect 19668 31424 19674 31476
rect 21361 31467 21419 31473
rect 21361 31433 21373 31467
rect 21407 31464 21419 31467
rect 21634 31464 21640 31476
rect 21407 31436 21640 31464
rect 21407 31433 21419 31436
rect 21361 31427 21419 31433
rect 21634 31424 21640 31436
rect 21692 31424 21698 31476
rect 23842 31424 23848 31476
rect 23900 31464 23906 31476
rect 24765 31467 24823 31473
rect 24765 31464 24777 31467
rect 23900 31436 24777 31464
rect 23900 31424 23906 31436
rect 24765 31433 24777 31436
rect 24811 31433 24823 31467
rect 25130 31464 25136 31476
rect 24765 31427 24823 31433
rect 24964 31436 25136 31464
rect 14306 31368 14412 31396
rect 15028 31368 18368 31396
rect 7837 31331 7895 31337
rect 7837 31297 7849 31331
rect 7883 31297 7895 31331
rect 7837 31291 7895 31297
rect 7926 31288 7932 31340
rect 7984 31328 7990 31340
rect 8205 31331 8263 31337
rect 8205 31328 8217 31331
rect 7984 31300 8217 31328
rect 7984 31288 7990 31300
rect 8205 31297 8217 31300
rect 8251 31297 8263 31331
rect 11514 31328 11520 31340
rect 8205 31291 8263 31297
rect 11072 31300 11520 31328
rect 6914 31260 6920 31272
rect 4672 31232 6920 31260
rect 4672 31220 4678 31232
rect 6914 31220 6920 31232
rect 6972 31260 6978 31272
rect 9309 31263 9367 31269
rect 9309 31260 9321 31263
rect 6972 31232 9321 31260
rect 6972 31220 6978 31232
rect 9309 31229 9321 31232
rect 9355 31229 9367 31263
rect 9309 31223 9367 31229
rect 9585 31263 9643 31269
rect 9585 31229 9597 31263
rect 9631 31260 9643 31263
rect 10134 31260 10140 31272
rect 9631 31232 10140 31260
rect 9631 31229 9643 31232
rect 9585 31223 9643 31229
rect 10134 31220 10140 31232
rect 10192 31220 10198 31272
rect 11072 31269 11100 31300
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 15028 31337 15056 31368
rect 15013 31331 15071 31337
rect 15013 31297 15025 31331
rect 15059 31297 15071 31331
rect 15013 31291 15071 31297
rect 16117 31331 16175 31337
rect 16117 31297 16129 31331
rect 16163 31297 16175 31331
rect 16117 31291 16175 31297
rect 11057 31263 11115 31269
rect 11057 31229 11069 31263
rect 11103 31229 11115 31263
rect 11057 31223 11115 31229
rect 12066 31220 12072 31272
rect 12124 31220 12130 31272
rect 14737 31263 14795 31269
rect 14737 31229 14749 31263
rect 14783 31260 14795 31263
rect 14783 31232 15148 31260
rect 14783 31229 14795 31232
rect 14737 31223 14795 31229
rect 3108 31164 3648 31192
rect 3108 31152 3114 31164
rect 4890 31152 4896 31204
rect 4948 31192 4954 31204
rect 6086 31192 6092 31204
rect 4948 31164 6092 31192
rect 4948 31152 4954 31164
rect 1670 31084 1676 31136
rect 1728 31124 1734 31136
rect 2133 31127 2191 31133
rect 2133 31124 2145 31127
rect 1728 31096 2145 31124
rect 1728 31084 1734 31096
rect 2133 31093 2145 31096
rect 2179 31093 2191 31127
rect 2133 31087 2191 31093
rect 2958 31084 2964 31136
rect 3016 31124 3022 31136
rect 3326 31124 3332 31136
rect 3016 31096 3332 31124
rect 3016 31084 3022 31096
rect 3326 31084 3332 31096
rect 3384 31124 3390 31136
rect 3881 31127 3939 31133
rect 3881 31124 3893 31127
rect 3384 31096 3893 31124
rect 3384 31084 3390 31096
rect 3881 31093 3893 31096
rect 3927 31093 3939 31127
rect 3881 31087 3939 31093
rect 4062 31084 4068 31136
rect 4120 31084 4126 31136
rect 5368 31133 5396 31164
rect 6086 31152 6092 31164
rect 6144 31152 6150 31204
rect 11885 31195 11943 31201
rect 11885 31161 11897 31195
rect 11931 31192 11943 31195
rect 13722 31192 13728 31204
rect 11931 31164 13728 31192
rect 11931 31161 11943 31164
rect 11885 31155 11943 31161
rect 13722 31152 13728 31164
rect 13780 31152 13786 31204
rect 15120 31192 15148 31232
rect 15194 31220 15200 31272
rect 15252 31220 15258 31272
rect 15381 31263 15439 31269
rect 15381 31229 15393 31263
rect 15427 31260 15439 31263
rect 16132 31260 16160 31291
rect 16206 31288 16212 31340
rect 16264 31288 16270 31340
rect 16301 31331 16359 31337
rect 16301 31297 16313 31331
rect 16347 31328 16359 31331
rect 16390 31328 16396 31340
rect 16347 31300 16396 31328
rect 16347 31297 16359 31300
rect 16301 31291 16359 31297
rect 16390 31288 16396 31300
rect 16448 31288 16454 31340
rect 16485 31331 16543 31337
rect 16485 31297 16497 31331
rect 16531 31328 16543 31331
rect 16850 31328 16856 31340
rect 16531 31300 16856 31328
rect 16531 31297 16543 31300
rect 16485 31291 16543 31297
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 17310 31288 17316 31340
rect 17368 31288 17374 31340
rect 17494 31288 17500 31340
rect 17552 31288 17558 31340
rect 17681 31331 17739 31337
rect 17681 31297 17693 31331
rect 17727 31297 17739 31331
rect 17681 31291 17739 31297
rect 17221 31263 17279 31269
rect 15427 31232 15608 31260
rect 16132 31232 16252 31260
rect 15427 31229 15439 31232
rect 15381 31223 15439 31229
rect 15470 31192 15476 31204
rect 15120 31164 15476 31192
rect 15470 31152 15476 31164
rect 15528 31152 15534 31204
rect 5353 31127 5411 31133
rect 5353 31093 5365 31127
rect 5399 31093 5411 31127
rect 5353 31087 5411 31093
rect 5626 31084 5632 31136
rect 5684 31084 5690 31136
rect 5810 31084 5816 31136
rect 5868 31124 5874 31136
rect 8202 31124 8208 31136
rect 5868 31096 8208 31124
rect 5868 31084 5874 31096
rect 8202 31084 8208 31096
rect 8260 31084 8266 31136
rect 11974 31084 11980 31136
rect 12032 31124 12038 31136
rect 12158 31124 12164 31136
rect 12032 31096 12164 31124
rect 12032 31084 12038 31096
rect 12158 31084 12164 31096
rect 12216 31084 12222 31136
rect 13265 31127 13323 31133
rect 13265 31093 13277 31127
rect 13311 31124 13323 31127
rect 14366 31124 14372 31136
rect 13311 31096 14372 31124
rect 13311 31093 13323 31096
rect 13265 31087 13323 31093
rect 14366 31084 14372 31096
rect 14424 31124 14430 31136
rect 15580 31124 15608 31232
rect 15654 31124 15660 31136
rect 14424 31096 15660 31124
rect 14424 31084 14430 31096
rect 15654 31084 15660 31096
rect 15712 31084 15718 31136
rect 15746 31084 15752 31136
rect 15804 31124 15810 31136
rect 15841 31127 15899 31133
rect 15841 31124 15853 31127
rect 15804 31096 15853 31124
rect 15804 31084 15810 31096
rect 15841 31093 15853 31096
rect 15887 31093 15899 31127
rect 16224 31124 16252 31232
rect 17221 31229 17233 31263
rect 17267 31260 17279 31263
rect 17328 31260 17356 31288
rect 17267 31232 17356 31260
rect 17696 31260 17724 31291
rect 17770 31288 17776 31340
rect 17828 31288 17834 31340
rect 17862 31288 17868 31340
rect 17920 31288 17926 31340
rect 18340 31337 18368 31368
rect 18325 31331 18383 31337
rect 18325 31297 18337 31331
rect 18371 31328 18383 31331
rect 18874 31328 18880 31340
rect 18371 31300 18880 31328
rect 18371 31297 18383 31300
rect 18325 31291 18383 31297
rect 18874 31288 18880 31300
rect 18932 31288 18938 31340
rect 19628 31328 19656 31424
rect 19794 31356 19800 31408
rect 19852 31396 19858 31408
rect 19852 31368 20760 31396
rect 19852 31356 19858 31368
rect 19306 31300 19656 31328
rect 19306 31260 19334 31300
rect 19702 31288 19708 31340
rect 19760 31288 19766 31340
rect 19981 31331 20039 31337
rect 19981 31297 19993 31331
rect 20027 31297 20039 31331
rect 19981 31291 20039 31297
rect 20073 31331 20131 31337
rect 20073 31297 20085 31331
rect 20119 31328 20131 31331
rect 20162 31328 20168 31340
rect 20119 31300 20168 31328
rect 20119 31297 20131 31300
rect 20073 31291 20131 31297
rect 17696 31232 19334 31260
rect 17267 31229 17279 31232
rect 17221 31223 17279 31229
rect 16390 31152 16396 31204
rect 16448 31192 16454 31204
rect 17696 31192 17724 31232
rect 19426 31220 19432 31272
rect 19484 31260 19490 31272
rect 19996 31260 20024 31291
rect 20162 31288 20168 31300
rect 20220 31288 20226 31340
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31297 20315 31331
rect 20257 31291 20315 31297
rect 19484 31232 20024 31260
rect 19484 31220 19490 31232
rect 16448 31164 17724 31192
rect 19996 31192 20024 31232
rect 20070 31192 20076 31204
rect 19996 31164 20076 31192
rect 16448 31152 16454 31164
rect 20070 31152 20076 31164
rect 20128 31152 20134 31204
rect 20272 31192 20300 31291
rect 20346 31288 20352 31340
rect 20404 31288 20410 31340
rect 20732 31337 20760 31368
rect 20990 31356 20996 31408
rect 21048 31356 21054 31408
rect 21085 31399 21143 31405
rect 21085 31365 21097 31399
rect 21131 31396 21143 31399
rect 21726 31396 21732 31408
rect 21131 31368 21732 31396
rect 21131 31365 21143 31368
rect 21085 31359 21143 31365
rect 21726 31356 21732 31368
rect 21784 31356 21790 31408
rect 23201 31399 23259 31405
rect 23201 31365 23213 31399
rect 23247 31396 23259 31399
rect 23474 31396 23480 31408
rect 23247 31368 23480 31396
rect 23247 31365 23259 31368
rect 23201 31359 23259 31365
rect 23474 31356 23480 31368
rect 23532 31356 23538 31408
rect 24964 31396 24992 31436
rect 25130 31424 25136 31436
rect 25188 31424 25194 31476
rect 25314 31424 25320 31476
rect 25372 31424 25378 31476
rect 26145 31467 26203 31473
rect 26145 31433 26157 31467
rect 26191 31464 26203 31467
rect 26234 31464 26240 31476
rect 26191 31436 26240 31464
rect 26191 31433 26203 31436
rect 26145 31427 26203 31433
rect 26234 31424 26240 31436
rect 26292 31424 26298 31476
rect 28261 31467 28319 31473
rect 28261 31433 28273 31467
rect 28307 31464 28319 31467
rect 29638 31464 29644 31476
rect 28307 31436 29644 31464
rect 28307 31433 28319 31436
rect 28261 31427 28319 31433
rect 29638 31424 29644 31436
rect 29696 31424 29702 31476
rect 29733 31467 29791 31473
rect 29733 31433 29745 31467
rect 29779 31433 29791 31467
rect 29733 31427 29791 31433
rect 24426 31368 24992 31396
rect 25041 31399 25099 31405
rect 25041 31365 25053 31399
rect 25087 31396 25099 31399
rect 25332 31396 25360 31424
rect 25087 31368 25360 31396
rect 27341 31399 27399 31405
rect 25087 31365 25099 31368
rect 25041 31359 25099 31365
rect 27341 31365 27353 31399
rect 27387 31396 27399 31399
rect 27706 31396 27712 31408
rect 27387 31368 27712 31396
rect 27387 31365 27399 31368
rect 27341 31359 27399 31365
rect 27706 31356 27712 31368
rect 27764 31356 27770 31408
rect 29396 31399 29454 31405
rect 29396 31365 29408 31399
rect 29442 31396 29454 31399
rect 29748 31396 29776 31427
rect 30374 31424 30380 31476
rect 30432 31464 30438 31476
rect 30561 31467 30619 31473
rect 30561 31464 30573 31467
rect 30432 31436 30573 31464
rect 30432 31424 30438 31436
rect 30561 31433 30573 31436
rect 30607 31433 30619 31467
rect 30561 31427 30619 31433
rect 32585 31467 32643 31473
rect 32585 31433 32597 31467
rect 32631 31464 32643 31467
rect 32766 31464 32772 31476
rect 32631 31436 32772 31464
rect 32631 31433 32643 31436
rect 32585 31427 32643 31433
rect 32766 31424 32772 31436
rect 32824 31424 32830 31476
rect 33318 31424 33324 31476
rect 33376 31424 33382 31476
rect 33781 31467 33839 31473
rect 33781 31433 33793 31467
rect 33827 31464 33839 31467
rect 34514 31464 34520 31476
rect 33827 31436 34520 31464
rect 33827 31433 33839 31436
rect 33781 31427 33839 31433
rect 34514 31424 34520 31436
rect 34572 31424 34578 31476
rect 41966 31464 41972 31476
rect 40328 31436 41972 31464
rect 29442 31368 29776 31396
rect 29442 31365 29454 31368
rect 29396 31359 29454 31365
rect 35342 31356 35348 31408
rect 35400 31396 35406 31408
rect 35400 31368 36384 31396
rect 35400 31356 35406 31368
rect 20898 31337 20904 31340
rect 20717 31331 20775 31337
rect 20717 31297 20729 31331
rect 20763 31297 20775 31331
rect 20717 31291 20775 31297
rect 20865 31331 20904 31337
rect 20865 31297 20877 31331
rect 20865 31291 20904 31297
rect 20732 31260 20760 31291
rect 20898 31288 20904 31291
rect 20956 31288 20962 31340
rect 21223 31331 21281 31337
rect 21223 31297 21235 31331
rect 21269 31328 21281 31331
rect 21634 31328 21640 31340
rect 21269 31300 21640 31328
rect 21269 31297 21281 31300
rect 21223 31291 21281 31297
rect 21634 31288 21640 31300
rect 21692 31288 21698 31340
rect 24946 31288 24952 31340
rect 25004 31288 25010 31340
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31328 25191 31331
rect 25222 31328 25228 31340
rect 25179 31300 25228 31328
rect 25179 31297 25191 31300
rect 25133 31291 25191 31297
rect 25222 31288 25228 31300
rect 25280 31288 25286 31340
rect 25317 31331 25375 31337
rect 25317 31297 25329 31331
rect 25363 31297 25375 31331
rect 25317 31291 25375 31297
rect 27433 31331 27491 31337
rect 27433 31297 27445 31331
rect 27479 31328 27491 31331
rect 28810 31328 28816 31340
rect 27479 31300 28816 31328
rect 27479 31297 27491 31300
rect 27433 31291 27491 31297
rect 22462 31260 22468 31272
rect 20732 31232 22468 31260
rect 22462 31220 22468 31232
rect 22520 31220 22526 31272
rect 22922 31220 22928 31272
rect 22980 31220 22986 31272
rect 23842 31260 23848 31272
rect 23032 31232 23848 31260
rect 20714 31192 20720 31204
rect 20272 31164 20720 31192
rect 16669 31127 16727 31133
rect 16669 31124 16681 31127
rect 16224 31096 16681 31124
rect 15841 31087 15899 31093
rect 16669 31093 16681 31096
rect 16715 31124 16727 31127
rect 16850 31124 16856 31136
rect 16715 31096 16856 31124
rect 16715 31093 16727 31096
rect 16669 31087 16727 31093
rect 16850 31084 16856 31096
rect 16908 31084 16914 31136
rect 17034 31084 17040 31136
rect 17092 31124 17098 31136
rect 18322 31124 18328 31136
rect 17092 31096 18328 31124
rect 17092 31084 17098 31096
rect 18322 31084 18328 31096
rect 18380 31084 18386 31136
rect 19886 31084 19892 31136
rect 19944 31124 19950 31136
rect 20272 31124 20300 31164
rect 20714 31152 20720 31164
rect 20772 31152 20778 31204
rect 21082 31152 21088 31204
rect 21140 31192 21146 31204
rect 23032 31192 23060 31232
rect 23842 31220 23848 31232
rect 23900 31220 23906 31272
rect 24394 31220 24400 31272
rect 24452 31260 24458 31272
rect 25332 31260 25360 31291
rect 28810 31288 28816 31300
rect 28868 31288 28874 31340
rect 29546 31288 29552 31340
rect 29604 31328 29610 31340
rect 29641 31331 29699 31337
rect 29641 31328 29653 31331
rect 29604 31300 29653 31328
rect 29604 31288 29610 31300
rect 29641 31297 29653 31300
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 30098 31288 30104 31340
rect 30156 31288 30162 31340
rect 30193 31331 30251 31337
rect 30193 31297 30205 31331
rect 30239 31328 30251 31331
rect 30558 31328 30564 31340
rect 30239 31300 30564 31328
rect 30239 31297 30251 31300
rect 30193 31291 30251 31297
rect 30558 31288 30564 31300
rect 30616 31288 30622 31340
rect 30742 31288 30748 31340
rect 30800 31328 30806 31340
rect 30929 31331 30987 31337
rect 30929 31328 30941 31331
rect 30800 31300 30941 31328
rect 30800 31288 30806 31300
rect 30929 31297 30941 31300
rect 30975 31297 30987 31331
rect 30929 31291 30987 31297
rect 32490 31288 32496 31340
rect 32548 31288 32554 31340
rect 33689 31331 33747 31337
rect 33689 31297 33701 31331
rect 33735 31328 33747 31331
rect 34146 31328 34152 31340
rect 33735 31300 34152 31328
rect 33735 31297 33747 31300
rect 33689 31291 33747 31297
rect 34146 31288 34152 31300
rect 34204 31288 34210 31340
rect 34606 31288 34612 31340
rect 34664 31328 34670 31340
rect 35069 31331 35127 31337
rect 35069 31328 35081 31331
rect 34664 31300 35081 31328
rect 34664 31288 34670 31300
rect 35069 31297 35081 31300
rect 35115 31297 35127 31331
rect 35069 31291 35127 31297
rect 35161 31331 35219 31337
rect 35161 31297 35173 31331
rect 35207 31297 35219 31331
rect 35161 31291 35219 31297
rect 35437 31331 35495 31337
rect 35437 31297 35449 31331
rect 35483 31328 35495 31331
rect 35986 31328 35992 31340
rect 35483 31300 35992 31328
rect 35483 31297 35495 31300
rect 35437 31291 35495 31297
rect 24452 31232 25360 31260
rect 26789 31263 26847 31269
rect 24452 31220 24458 31232
rect 26789 31229 26801 31263
rect 26835 31229 26847 31263
rect 26789 31223 26847 31229
rect 21140 31164 23060 31192
rect 21140 31152 21146 31164
rect 24210 31152 24216 31204
rect 24268 31192 24274 31204
rect 24578 31192 24584 31204
rect 24268 31164 24584 31192
rect 24268 31152 24274 31164
rect 24578 31152 24584 31164
rect 24636 31192 24642 31204
rect 24673 31195 24731 31201
rect 24673 31192 24685 31195
rect 24636 31164 24685 31192
rect 24636 31152 24642 31164
rect 24673 31161 24685 31164
rect 24719 31161 24731 31195
rect 26804 31192 26832 31223
rect 27522 31220 27528 31272
rect 27580 31220 27586 31272
rect 30282 31220 30288 31272
rect 30340 31220 30346 31272
rect 31018 31220 31024 31272
rect 31076 31220 31082 31272
rect 31113 31263 31171 31269
rect 31113 31229 31125 31263
rect 31159 31260 31171 31263
rect 32674 31260 32680 31272
rect 31159 31232 32680 31260
rect 31159 31229 31171 31232
rect 31113 31223 31171 31229
rect 26973 31195 27031 31201
rect 26973 31192 26985 31195
rect 26804 31164 26985 31192
rect 24673 31155 24731 31161
rect 26973 31161 26985 31164
rect 27019 31161 27031 31195
rect 30300 31192 30328 31220
rect 31128 31192 31156 31223
rect 32674 31220 32680 31232
rect 32732 31220 32738 31272
rect 33965 31263 34023 31269
rect 33965 31229 33977 31263
rect 34011 31260 34023 31263
rect 34238 31260 34244 31272
rect 34011 31232 34244 31260
rect 34011 31229 34023 31232
rect 33965 31223 34023 31229
rect 34238 31220 34244 31232
rect 34296 31220 34302 31272
rect 34514 31220 34520 31272
rect 34572 31260 34578 31272
rect 34790 31260 34796 31272
rect 34572 31232 34796 31260
rect 34572 31220 34578 31232
rect 34790 31220 34796 31232
rect 34848 31220 34854 31272
rect 35176 31260 35204 31291
rect 35986 31288 35992 31300
rect 36044 31288 36050 31340
rect 36262 31260 36268 31272
rect 35176 31232 36268 31260
rect 36262 31220 36268 31232
rect 36320 31220 36326 31272
rect 36356 31260 36384 31368
rect 36630 31356 36636 31408
rect 36688 31396 36694 31408
rect 36998 31396 37004 31408
rect 36688 31368 37004 31396
rect 36688 31356 36694 31368
rect 36998 31356 37004 31368
rect 37056 31396 37062 31408
rect 40037 31399 40095 31405
rect 40037 31396 40049 31399
rect 37056 31368 40049 31396
rect 37056 31356 37062 31368
rect 40037 31365 40049 31368
rect 40083 31365 40095 31399
rect 40037 31359 40095 31365
rect 37274 31288 37280 31340
rect 37332 31288 37338 31340
rect 37458 31288 37464 31340
rect 37516 31328 37522 31340
rect 37553 31331 37611 31337
rect 37553 31328 37565 31331
rect 37516 31300 37565 31328
rect 37516 31288 37522 31300
rect 37553 31297 37565 31300
rect 37599 31297 37611 31331
rect 37553 31291 37611 31297
rect 37645 31331 37703 31337
rect 37645 31297 37657 31331
rect 37691 31328 37703 31331
rect 37826 31328 37832 31340
rect 37691 31300 37832 31328
rect 37691 31297 37703 31300
rect 37645 31291 37703 31297
rect 37826 31288 37832 31300
rect 37884 31288 37890 31340
rect 39945 31331 40003 31337
rect 39945 31297 39957 31331
rect 39991 31297 40003 31331
rect 39945 31291 40003 31297
rect 39960 31260 39988 31291
rect 40126 31288 40132 31340
rect 40184 31288 40190 31340
rect 40328 31337 40356 31436
rect 41966 31424 41972 31436
rect 42024 31464 42030 31476
rect 42153 31467 42211 31473
rect 42153 31464 42165 31467
rect 42024 31436 42165 31464
rect 42024 31424 42030 31436
rect 42153 31433 42165 31436
rect 42199 31433 42211 31467
rect 42153 31427 42211 31433
rect 40313 31331 40371 31337
rect 40313 31297 40325 31331
rect 40359 31297 40371 31331
rect 40313 31291 40371 31297
rect 40402 31288 40408 31340
rect 40460 31288 40466 31340
rect 41782 31288 41788 31340
rect 41840 31288 41846 31340
rect 36356 31232 39988 31260
rect 40681 31263 40739 31269
rect 40681 31229 40693 31263
rect 40727 31260 40739 31263
rect 41046 31260 41052 31272
rect 40727 31232 41052 31260
rect 40727 31229 40739 31232
rect 40681 31223 40739 31229
rect 41046 31220 41052 31232
rect 41104 31220 41110 31272
rect 30300 31164 31156 31192
rect 26973 31155 27031 31161
rect 34330 31152 34336 31204
rect 34388 31192 34394 31204
rect 35345 31195 35403 31201
rect 35345 31192 35357 31195
rect 34388 31164 35357 31192
rect 34388 31152 34394 31164
rect 35345 31161 35357 31164
rect 35391 31192 35403 31195
rect 37369 31195 37427 31201
rect 37369 31192 37381 31195
rect 35391 31164 37381 31192
rect 35391 31161 35403 31164
rect 35345 31155 35403 31161
rect 37369 31161 37381 31164
rect 37415 31192 37427 31195
rect 37734 31192 37740 31204
rect 37415 31164 37740 31192
rect 37415 31161 37427 31164
rect 37369 31155 37427 31161
rect 37734 31152 37740 31164
rect 37792 31152 37798 31204
rect 19944 31096 20300 31124
rect 19944 31084 19950 31096
rect 20530 31084 20536 31136
rect 20588 31084 20594 31136
rect 20806 31084 20812 31136
rect 20864 31124 20870 31136
rect 24302 31124 24308 31136
rect 20864 31096 24308 31124
rect 20864 31084 20870 31096
rect 24302 31084 24308 31096
rect 24360 31084 24366 31136
rect 32125 31127 32183 31133
rect 32125 31093 32137 31127
rect 32171 31124 32183 31127
rect 32766 31124 32772 31136
rect 32171 31096 32772 31124
rect 32171 31093 32183 31096
rect 32125 31087 32183 31093
rect 32766 31084 32772 31096
rect 32824 31084 32830 31136
rect 34790 31084 34796 31136
rect 34848 31124 34854 31136
rect 34885 31127 34943 31133
rect 34885 31124 34897 31127
rect 34848 31096 34897 31124
rect 34848 31084 34854 31096
rect 34885 31093 34897 31096
rect 34931 31093 34943 31127
rect 34885 31087 34943 31093
rect 37642 31084 37648 31136
rect 37700 31124 37706 31136
rect 37829 31127 37887 31133
rect 37829 31124 37841 31127
rect 37700 31096 37841 31124
rect 37700 31084 37706 31096
rect 37829 31093 37841 31096
rect 37875 31093 37887 31127
rect 37829 31087 37887 31093
rect 39761 31127 39819 31133
rect 39761 31093 39773 31127
rect 39807 31124 39819 31127
rect 40862 31124 40868 31136
rect 39807 31096 40868 31124
rect 39807 31093 39819 31096
rect 39761 31087 39819 31093
rect 40862 31084 40868 31096
rect 40920 31084 40926 31136
rect 1104 31034 42504 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 42504 31034
rect 1104 30960 42504 30982
rect 3142 30880 3148 30932
rect 3200 30880 3206 30932
rect 3234 30880 3240 30932
rect 3292 30880 3298 30932
rect 3510 30880 3516 30932
rect 3568 30920 3574 30932
rect 4798 30920 4804 30932
rect 3568 30892 4804 30920
rect 3568 30880 3574 30892
rect 4798 30880 4804 30892
rect 4856 30880 4862 30932
rect 5261 30923 5319 30929
rect 5261 30889 5273 30923
rect 5307 30920 5319 30923
rect 5626 30920 5632 30932
rect 5307 30892 5632 30920
rect 5307 30889 5319 30892
rect 5261 30883 5319 30889
rect 5626 30880 5632 30892
rect 5684 30880 5690 30932
rect 10778 30880 10784 30932
rect 10836 30880 10842 30932
rect 12621 30923 12679 30929
rect 12621 30889 12633 30923
rect 12667 30920 12679 30923
rect 12894 30920 12900 30932
rect 12667 30892 12900 30920
rect 12667 30889 12679 30892
rect 12621 30883 12679 30889
rect 12894 30880 12900 30892
rect 12952 30880 12958 30932
rect 14458 30880 14464 30932
rect 14516 30920 14522 30932
rect 15010 30920 15016 30932
rect 14516 30892 15016 30920
rect 14516 30880 14522 30892
rect 15010 30880 15016 30892
rect 15068 30880 15074 30932
rect 15838 30880 15844 30932
rect 15896 30920 15902 30932
rect 16117 30923 16175 30929
rect 16117 30920 16129 30923
rect 15896 30892 16129 30920
rect 15896 30880 15902 30892
rect 16117 30889 16129 30892
rect 16163 30889 16175 30923
rect 16117 30883 16175 30889
rect 16206 30880 16212 30932
rect 16264 30920 16270 30932
rect 16390 30920 16396 30932
rect 16264 30892 16396 30920
rect 16264 30880 16270 30892
rect 16390 30880 16396 30892
rect 16448 30920 16454 30932
rect 17402 30920 17408 30932
rect 16448 30892 17408 30920
rect 16448 30880 16454 30892
rect 17402 30880 17408 30892
rect 17460 30880 17466 30932
rect 18049 30923 18107 30929
rect 18049 30889 18061 30923
rect 18095 30920 18107 30923
rect 18782 30920 18788 30932
rect 18095 30892 18788 30920
rect 18095 30889 18107 30892
rect 18049 30883 18107 30889
rect 18782 30880 18788 30892
rect 18840 30880 18846 30932
rect 19426 30880 19432 30932
rect 19484 30880 19490 30932
rect 19794 30920 19800 30932
rect 19536 30892 19800 30920
rect 2746 30824 3740 30852
rect 1397 30787 1455 30793
rect 1397 30753 1409 30787
rect 1443 30784 1455 30787
rect 2746 30784 2774 30824
rect 1443 30756 2774 30784
rect 3712 30784 3740 30824
rect 3786 30812 3792 30864
rect 3844 30812 3850 30864
rect 4709 30855 4767 30861
rect 4709 30821 4721 30855
rect 4755 30852 4767 30855
rect 5534 30852 5540 30864
rect 4755 30824 5540 30852
rect 4755 30821 4767 30824
rect 4709 30815 4767 30821
rect 5534 30812 5540 30824
rect 5592 30812 5598 30864
rect 4614 30784 4620 30796
rect 3712 30756 4620 30784
rect 1443 30753 1455 30756
rect 1397 30747 1455 30753
rect 4614 30744 4620 30756
rect 4672 30744 4678 30796
rect 4801 30787 4859 30793
rect 4801 30753 4813 30787
rect 4847 30784 4859 30787
rect 4890 30784 4896 30796
rect 4847 30756 4896 30784
rect 4847 30753 4859 30756
rect 4801 30747 4859 30753
rect 4890 30744 4896 30756
rect 4948 30744 4954 30796
rect 5166 30744 5172 30796
rect 5224 30744 5230 30796
rect 6914 30744 6920 30796
rect 6972 30744 6978 30796
rect 10502 30744 10508 30796
rect 10560 30744 10566 30796
rect 10870 30744 10876 30796
rect 10928 30744 10934 30796
rect 12912 30784 12940 30880
rect 19536 30852 19564 30892
rect 19794 30880 19800 30892
rect 19852 30880 19858 30932
rect 19889 30923 19947 30929
rect 19889 30889 19901 30923
rect 19935 30920 19947 30923
rect 20346 30920 20352 30932
rect 19935 30892 20352 30920
rect 19935 30889 19947 30892
rect 19889 30883 19947 30889
rect 19904 30852 19932 30883
rect 20346 30880 20352 30892
rect 20404 30880 20410 30932
rect 20622 30880 20628 30932
rect 20680 30880 20686 30932
rect 23569 30923 23627 30929
rect 23569 30889 23581 30923
rect 23615 30920 23627 30923
rect 23658 30920 23664 30932
rect 23615 30892 23664 30920
rect 23615 30889 23627 30892
rect 23569 30883 23627 30889
rect 23658 30880 23664 30892
rect 23716 30880 23722 30932
rect 23750 30880 23756 30932
rect 23808 30920 23814 30932
rect 24397 30923 24455 30929
rect 24397 30920 24409 30923
rect 23808 30892 24409 30920
rect 23808 30880 23814 30892
rect 24397 30889 24409 30892
rect 24443 30889 24455 30923
rect 24946 30920 24952 30932
rect 24397 30883 24455 30889
rect 24504 30892 24952 30920
rect 16408 30824 19564 30852
rect 19812 30824 19932 30852
rect 13265 30787 13323 30793
rect 13265 30784 13277 30787
rect 12912 30756 13277 30784
rect 13265 30753 13277 30756
rect 13311 30753 13323 30787
rect 13265 30747 13323 30753
rect 14366 30744 14372 30796
rect 14424 30744 14430 30796
rect 15654 30744 15660 30796
rect 15712 30784 15718 30796
rect 15841 30787 15899 30793
rect 15841 30784 15853 30787
rect 15712 30756 15853 30784
rect 15712 30744 15718 30756
rect 15841 30753 15853 30756
rect 15887 30753 15899 30787
rect 16408 30784 16436 30824
rect 15841 30747 15899 30753
rect 16316 30756 16436 30784
rect 16316 30728 16344 30756
rect 16574 30744 16580 30796
rect 16632 30784 16638 30796
rect 18414 30784 18420 30796
rect 16632 30756 17080 30784
rect 16632 30744 16638 30756
rect 3421 30719 3479 30725
rect 3421 30685 3433 30719
rect 3467 30685 3479 30719
rect 3421 30679 3479 30685
rect 1670 30608 1676 30660
rect 1728 30608 1734 30660
rect 3050 30648 3056 30660
rect 2898 30620 3056 30648
rect 3050 30608 3056 30620
rect 3108 30608 3114 30660
rect 3436 30648 3464 30679
rect 3510 30676 3516 30728
rect 3568 30676 3574 30728
rect 4062 30716 4068 30728
rect 3712 30688 4068 30716
rect 3712 30648 3740 30688
rect 4062 30676 4068 30688
rect 4120 30676 4126 30728
rect 4246 30676 4252 30728
rect 4304 30716 4310 30728
rect 4525 30719 4583 30725
rect 4525 30716 4537 30719
rect 4304 30688 4537 30716
rect 4304 30676 4310 30688
rect 4525 30685 4537 30688
rect 4571 30685 4583 30719
rect 4525 30679 4583 30685
rect 5626 30676 5632 30728
rect 5684 30676 5690 30728
rect 5905 30719 5963 30725
rect 5905 30685 5917 30719
rect 5951 30716 5963 30719
rect 5994 30716 6000 30728
rect 5951 30688 6000 30716
rect 5951 30685 5963 30688
rect 5905 30679 5963 30685
rect 5994 30676 6000 30688
rect 6052 30676 6058 30728
rect 6086 30676 6092 30728
rect 6144 30676 6150 30728
rect 10594 30676 10600 30728
rect 10652 30676 10658 30728
rect 13446 30676 13452 30728
rect 13504 30676 13510 30728
rect 13633 30719 13691 30725
rect 13633 30685 13645 30719
rect 13679 30716 13691 30719
rect 13814 30716 13820 30728
rect 13679 30688 13820 30716
rect 13679 30685 13691 30688
rect 13633 30679 13691 30685
rect 13814 30676 13820 30688
rect 13872 30716 13878 30728
rect 14182 30716 14188 30728
rect 13872 30688 14188 30716
rect 13872 30676 13878 30688
rect 14182 30676 14188 30688
rect 14240 30676 14246 30728
rect 15562 30676 15568 30728
rect 15620 30676 15626 30728
rect 15749 30719 15807 30725
rect 15749 30685 15761 30719
rect 15795 30716 15807 30719
rect 16114 30716 16120 30728
rect 15795 30688 16120 30716
rect 15795 30685 15807 30688
rect 15749 30679 15807 30685
rect 16114 30676 16120 30688
rect 16172 30676 16178 30728
rect 16298 30676 16304 30728
rect 16356 30676 16362 30728
rect 16393 30719 16451 30725
rect 16393 30685 16405 30719
rect 16439 30685 16451 30719
rect 16393 30679 16451 30685
rect 3436 30620 3740 30648
rect 3789 30651 3847 30657
rect 3789 30617 3801 30651
rect 3835 30648 3847 30651
rect 5077 30651 5135 30657
rect 3835 30620 4108 30648
rect 3835 30617 3847 30620
rect 3789 30611 3847 30617
rect 4080 30592 4108 30620
rect 5077 30617 5089 30651
rect 5123 30648 5135 30651
rect 5258 30648 5264 30660
rect 5123 30620 5264 30648
rect 5123 30617 5135 30620
rect 5077 30611 5135 30617
rect 5258 30608 5264 30620
rect 5316 30608 5322 30660
rect 5537 30651 5595 30657
rect 5537 30617 5549 30651
rect 5583 30617 5595 30651
rect 5537 30611 5595 30617
rect 3142 30540 3148 30592
rect 3200 30580 3206 30592
rect 3973 30583 4031 30589
rect 3973 30580 3985 30583
rect 3200 30552 3985 30580
rect 3200 30540 3206 30552
rect 3973 30549 3985 30552
rect 4019 30549 4031 30583
rect 3973 30543 4031 30549
rect 4062 30540 4068 30592
rect 4120 30540 4126 30592
rect 4341 30583 4399 30589
rect 4341 30549 4353 30583
rect 4387 30580 4399 30583
rect 4614 30580 4620 30592
rect 4387 30552 4620 30580
rect 4387 30549 4399 30552
rect 4341 30543 4399 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 5442 30540 5448 30592
rect 5500 30540 5506 30592
rect 5552 30580 5580 30611
rect 6178 30608 6184 30660
rect 6236 30608 6242 30660
rect 11146 30608 11152 30660
rect 11204 30608 11210 30660
rect 11256 30620 11638 30648
rect 5813 30583 5871 30589
rect 5813 30580 5825 30583
rect 5552 30552 5825 30580
rect 5813 30549 5825 30552
rect 5859 30549 5871 30583
rect 5813 30543 5871 30549
rect 10137 30583 10195 30589
rect 10137 30549 10149 30583
rect 10183 30580 10195 30583
rect 10686 30580 10692 30592
rect 10183 30552 10692 30580
rect 10183 30549 10195 30552
rect 10137 30543 10195 30549
rect 10686 30540 10692 30552
rect 10744 30540 10750 30592
rect 10962 30540 10968 30592
rect 11020 30580 11026 30592
rect 11256 30580 11284 30620
rect 15102 30608 15108 30660
rect 15160 30648 15166 30660
rect 16408 30648 16436 30679
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 17052 30716 17080 30756
rect 17512 30756 18420 30784
rect 17512 30716 17540 30756
rect 18414 30744 18420 30756
rect 18472 30744 18478 30796
rect 18874 30744 18880 30796
rect 18932 30744 18938 30796
rect 18975 30756 19656 30784
rect 17052 30688 17540 30716
rect 17589 30697 17647 30703
rect 17589 30663 17601 30697
rect 17635 30663 17647 30697
rect 17678 30676 17684 30728
rect 17736 30676 17742 30728
rect 17770 30676 17776 30728
rect 17828 30716 17834 30728
rect 17865 30719 17923 30725
rect 17865 30716 17877 30719
rect 17828 30688 17877 30716
rect 17828 30676 17834 30688
rect 17865 30685 17877 30688
rect 17911 30685 17923 30719
rect 17865 30679 17923 30685
rect 18138 30676 18144 30728
rect 18196 30676 18202 30728
rect 18506 30676 18512 30728
rect 18564 30716 18570 30728
rect 18975 30716 19003 30756
rect 18564 30688 19003 30716
rect 19245 30719 19303 30725
rect 18564 30676 18570 30688
rect 19245 30685 19257 30719
rect 19291 30685 19303 30719
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 19245 30679 19303 30685
rect 19352 30688 19441 30716
rect 17034 30648 17040 30660
rect 15160 30620 16344 30648
rect 16408 30620 17040 30648
rect 15160 30608 15166 30620
rect 11020 30552 11284 30580
rect 11020 30540 11026 30552
rect 12710 30540 12716 30592
rect 12768 30540 12774 30592
rect 13541 30583 13599 30589
rect 13541 30549 13553 30583
rect 13587 30580 13599 30583
rect 13722 30580 13728 30592
rect 13587 30552 13728 30580
rect 13587 30549 13599 30552
rect 13541 30543 13599 30549
rect 13722 30540 13728 30552
rect 13780 30540 13786 30592
rect 15194 30540 15200 30592
rect 15252 30580 15258 30592
rect 15381 30583 15439 30589
rect 15381 30580 15393 30583
rect 15252 30552 15393 30580
rect 15252 30540 15258 30552
rect 15381 30549 15393 30552
rect 15427 30549 15439 30583
rect 16316 30580 16344 30620
rect 17034 30608 17040 30620
rect 17092 30608 17098 30660
rect 17126 30608 17132 30660
rect 17184 30608 17190 30660
rect 17589 30657 17647 30663
rect 16482 30580 16488 30592
rect 16316 30552 16488 30580
rect 15381 30543 15439 30549
rect 16482 30540 16488 30552
rect 16540 30580 16546 30592
rect 16853 30583 16911 30589
rect 16853 30580 16865 30583
rect 16540 30552 16865 30580
rect 16540 30540 16546 30552
rect 16853 30549 16865 30552
rect 16899 30580 16911 30583
rect 17402 30580 17408 30592
rect 16899 30552 17408 30580
rect 16899 30549 16911 30552
rect 16853 30543 16911 30549
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 17604 30580 17632 30657
rect 17696 30648 17724 30676
rect 19260 30648 19288 30679
rect 17696 30620 19288 30648
rect 18690 30580 18696 30592
rect 17604 30552 18696 30580
rect 18690 30540 18696 30552
rect 18748 30580 18754 30592
rect 19352 30580 19380 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19518 30608 19524 30660
rect 19576 30608 19582 30660
rect 18748 30552 19380 30580
rect 19628 30580 19656 30756
rect 19812 30716 19840 30824
rect 21634 30812 21640 30864
rect 21692 30852 21698 30864
rect 24504 30852 24532 30892
rect 24946 30880 24952 30892
rect 25004 30920 25010 30932
rect 25004 30892 25452 30920
rect 25004 30880 25010 30892
rect 21692 30824 24532 30852
rect 21692 30812 21698 30824
rect 24578 30812 24584 30864
rect 24636 30852 24642 30864
rect 24636 30824 25360 30852
rect 24636 30812 24642 30824
rect 20070 30744 20076 30796
rect 20128 30784 20134 30796
rect 20806 30784 20812 30796
rect 20128 30756 20300 30784
rect 20128 30744 20134 30756
rect 20272 30725 20300 30756
rect 20456 30756 20812 30784
rect 19981 30719 20039 30725
rect 19981 30716 19993 30719
rect 19812 30688 19993 30716
rect 19981 30685 19993 30688
rect 20027 30685 20039 30719
rect 20165 30719 20223 30725
rect 20165 30713 20177 30719
rect 19981 30679 20039 30685
rect 20088 30685 20177 30713
rect 20211 30685 20223 30719
rect 19705 30651 19763 30657
rect 19705 30617 19717 30651
rect 19751 30648 19763 30651
rect 19794 30648 19800 30660
rect 19751 30620 19800 30648
rect 19751 30617 19763 30620
rect 19705 30611 19763 30617
rect 19794 30608 19800 30620
rect 19852 30608 19858 30660
rect 19886 30608 19892 30660
rect 19944 30648 19950 30660
rect 20088 30648 20116 30685
rect 20165 30679 20223 30685
rect 20257 30719 20315 30725
rect 20257 30685 20269 30719
rect 20303 30685 20315 30719
rect 20257 30679 20315 30685
rect 20346 30676 20352 30728
rect 20404 30725 20410 30728
rect 20404 30719 20427 30725
rect 20415 30685 20427 30719
rect 20404 30679 20427 30685
rect 20404 30676 20410 30679
rect 20456 30648 20484 30756
rect 20806 30744 20812 30756
rect 20864 30744 20870 30796
rect 20993 30787 21051 30793
rect 20993 30753 21005 30787
rect 21039 30784 21051 30787
rect 21082 30784 21088 30796
rect 21039 30756 21088 30784
rect 21039 30753 21051 30756
rect 20993 30747 21051 30753
rect 21082 30744 21088 30756
rect 21140 30784 21146 30796
rect 21910 30784 21916 30796
rect 21140 30756 21916 30784
rect 21140 30744 21146 30756
rect 21910 30744 21916 30756
rect 21968 30744 21974 30796
rect 24765 30787 24823 30793
rect 24765 30753 24777 30787
rect 24811 30784 24823 30787
rect 24946 30784 24952 30796
rect 24811 30756 24952 30784
rect 24811 30753 24823 30756
rect 24765 30747 24823 30753
rect 24946 30744 24952 30756
rect 25004 30784 25010 30796
rect 25332 30793 25360 30824
rect 25133 30787 25191 30793
rect 25133 30784 25145 30787
rect 25004 30756 25145 30784
rect 25004 30744 25010 30756
rect 25133 30753 25145 30756
rect 25179 30753 25191 30787
rect 25133 30747 25191 30753
rect 25317 30787 25375 30793
rect 25317 30753 25329 30787
rect 25363 30753 25375 30787
rect 25317 30747 25375 30753
rect 20714 30676 20720 30728
rect 20772 30716 20778 30728
rect 21545 30719 21603 30725
rect 21545 30716 21557 30719
rect 20772 30688 21557 30716
rect 20772 30676 20778 30688
rect 21545 30685 21557 30688
rect 21591 30685 21603 30719
rect 21545 30679 21603 30685
rect 22005 30719 22063 30725
rect 22005 30685 22017 30719
rect 22051 30716 22063 30719
rect 22094 30716 22100 30728
rect 22051 30688 22100 30716
rect 22051 30685 22063 30688
rect 22005 30679 22063 30685
rect 22094 30676 22100 30688
rect 22152 30676 22158 30728
rect 23750 30676 23756 30728
rect 23808 30676 23814 30728
rect 24026 30676 24032 30728
rect 24084 30716 24090 30728
rect 24121 30719 24179 30725
rect 24121 30716 24133 30719
rect 24084 30688 24133 30716
rect 24084 30676 24090 30688
rect 24121 30685 24133 30688
rect 24167 30716 24179 30719
rect 24394 30716 24400 30728
rect 24167 30688 24400 30716
rect 24167 30685 24179 30688
rect 24121 30679 24179 30685
rect 24394 30676 24400 30688
rect 24452 30676 24458 30728
rect 24578 30676 24584 30728
rect 24636 30676 24642 30728
rect 24670 30676 24676 30728
rect 24728 30676 24734 30728
rect 24854 30676 24860 30728
rect 24912 30676 24918 30728
rect 25041 30719 25099 30725
rect 25041 30685 25053 30719
rect 25087 30685 25099 30719
rect 25424 30716 25452 30892
rect 31018 30880 31024 30932
rect 31076 30880 31082 30932
rect 32122 30880 32128 30932
rect 32180 30920 32186 30932
rect 32217 30923 32275 30929
rect 32217 30920 32229 30923
rect 32180 30892 32229 30920
rect 32180 30880 32186 30892
rect 32217 30889 32229 30892
rect 32263 30889 32275 30923
rect 32217 30883 32275 30889
rect 34790 30880 34796 30932
rect 34848 30880 34854 30932
rect 35986 30880 35992 30932
rect 36044 30920 36050 30932
rect 36449 30923 36507 30929
rect 36449 30920 36461 30923
rect 36044 30892 36461 30920
rect 36044 30880 36050 30892
rect 36449 30889 36461 30892
rect 36495 30889 36507 30923
rect 36449 30883 36507 30889
rect 37277 30923 37335 30929
rect 37277 30889 37289 30923
rect 37323 30920 37335 30923
rect 37458 30920 37464 30932
rect 37323 30892 37464 30920
rect 37323 30889 37335 30892
rect 37277 30883 37335 30889
rect 37458 30880 37464 30892
rect 37516 30880 37522 30932
rect 41046 30880 41052 30932
rect 41104 30880 41110 30932
rect 30834 30852 30840 30864
rect 30484 30824 30840 30852
rect 28258 30784 28264 30796
rect 27448 30756 28264 30784
rect 26050 30716 26056 30728
rect 25424 30688 26056 30716
rect 25041 30679 25099 30685
rect 19944 30620 20116 30648
rect 20364 30620 20484 30648
rect 22189 30651 22247 30657
rect 19944 30608 19950 30620
rect 20364 30580 20392 30620
rect 22189 30617 22201 30651
rect 22235 30648 22247 30651
rect 22646 30648 22652 30660
rect 22235 30620 22652 30648
rect 22235 30617 22247 30620
rect 22189 30611 22247 30617
rect 22646 30608 22652 30620
rect 22704 30608 22710 30660
rect 23842 30608 23848 30660
rect 23900 30608 23906 30660
rect 23937 30651 23995 30657
rect 23937 30617 23949 30651
rect 23983 30648 23995 30651
rect 24688 30648 24716 30676
rect 25056 30648 25084 30679
rect 26050 30676 26056 30688
rect 26108 30716 26114 30728
rect 27448 30725 27476 30756
rect 28258 30744 28264 30756
rect 28316 30744 28322 30796
rect 30484 30793 30512 30824
rect 30834 30812 30840 30824
rect 30892 30852 30898 30864
rect 32490 30852 32496 30864
rect 30892 30824 32496 30852
rect 30892 30812 30898 30824
rect 32490 30812 32496 30824
rect 32548 30812 32554 30864
rect 30469 30787 30527 30793
rect 30469 30753 30481 30787
rect 30515 30753 30527 30787
rect 30469 30747 30527 30753
rect 31570 30744 31576 30796
rect 31628 30744 31634 30796
rect 32766 30744 32772 30796
rect 32824 30744 32830 30796
rect 34698 30744 34704 30796
rect 34756 30744 34762 30796
rect 34808 30784 34836 30880
rect 34977 30787 35035 30793
rect 34977 30784 34989 30787
rect 34808 30756 34989 30784
rect 34977 30753 34989 30756
rect 35023 30753 35035 30787
rect 34977 30747 35035 30753
rect 36170 30744 36176 30796
rect 36228 30744 36234 30796
rect 36354 30744 36360 30796
rect 36412 30784 36418 30796
rect 36412 30756 37136 30784
rect 36412 30744 36418 30756
rect 27295 30719 27353 30725
rect 27295 30716 27307 30719
rect 26108 30688 27307 30716
rect 26108 30676 26114 30688
rect 27295 30685 27307 30688
rect 27341 30685 27353 30719
rect 27295 30679 27353 30685
rect 27433 30719 27491 30725
rect 27433 30685 27445 30719
rect 27479 30685 27491 30719
rect 27433 30679 27491 30685
rect 27614 30676 27620 30728
rect 27672 30725 27678 30728
rect 27672 30719 27711 30725
rect 27699 30685 27711 30719
rect 27672 30679 27711 30685
rect 27801 30719 27859 30725
rect 27801 30685 27813 30719
rect 27847 30716 27859 30719
rect 28074 30716 28080 30728
rect 27847 30688 28080 30716
rect 27847 30685 27859 30688
rect 27801 30679 27859 30685
rect 27672 30676 27678 30679
rect 28074 30676 28080 30688
rect 28132 30676 28138 30728
rect 28902 30676 28908 30728
rect 28960 30716 28966 30728
rect 28960 30688 29684 30716
rect 28960 30676 28966 30688
rect 23983 30620 24164 30648
rect 24688 30620 25084 30648
rect 23983 30617 23995 30620
rect 23937 30611 23995 30617
rect 24136 30592 24164 30620
rect 25222 30608 25228 30660
rect 25280 30648 25286 30660
rect 27525 30651 27583 30657
rect 27525 30648 27537 30651
rect 25280 30620 27537 30648
rect 25280 30608 25286 30620
rect 27525 30617 27537 30620
rect 27571 30617 27583 30651
rect 27525 30611 27583 30617
rect 28721 30651 28779 30657
rect 28721 30617 28733 30651
rect 28767 30617 28779 30651
rect 28721 30611 28779 30617
rect 19628 30552 20392 30580
rect 18748 30540 18754 30552
rect 20438 30540 20444 30592
rect 20496 30580 20502 30592
rect 21085 30583 21143 30589
rect 21085 30580 21097 30583
rect 20496 30552 21097 30580
rect 20496 30540 20502 30552
rect 21085 30549 21097 30552
rect 21131 30549 21143 30583
rect 21085 30543 21143 30549
rect 21450 30540 21456 30592
rect 21508 30540 21514 30592
rect 21637 30583 21695 30589
rect 21637 30549 21649 30583
rect 21683 30580 21695 30583
rect 21726 30580 21732 30592
rect 21683 30552 21732 30580
rect 21683 30549 21695 30552
rect 21637 30543 21695 30549
rect 21726 30540 21732 30552
rect 21784 30540 21790 30592
rect 21818 30540 21824 30592
rect 21876 30540 21882 30592
rect 22370 30540 22376 30592
rect 22428 30580 22434 30592
rect 24118 30580 24124 30592
rect 22428 30552 24124 30580
rect 22428 30540 22434 30552
rect 24118 30540 24124 30552
rect 24176 30540 24182 30592
rect 25317 30583 25375 30589
rect 25317 30549 25329 30583
rect 25363 30580 25375 30583
rect 25958 30580 25964 30592
rect 25363 30552 25964 30580
rect 25363 30549 25375 30552
rect 25317 30543 25375 30549
rect 25958 30540 25964 30552
rect 26016 30540 26022 30592
rect 27154 30540 27160 30592
rect 27212 30540 27218 30592
rect 28350 30540 28356 30592
rect 28408 30580 28414 30592
rect 28445 30583 28503 30589
rect 28445 30580 28457 30583
rect 28408 30552 28457 30580
rect 28408 30540 28414 30552
rect 28445 30549 28457 30552
rect 28491 30580 28503 30583
rect 28736 30580 28764 30611
rect 29178 30608 29184 30660
rect 29236 30648 29242 30660
rect 29549 30651 29607 30657
rect 29549 30648 29561 30651
rect 29236 30620 29561 30648
rect 29236 30608 29242 30620
rect 29549 30617 29561 30620
rect 29595 30617 29607 30651
rect 29549 30611 29607 30617
rect 28491 30552 28764 30580
rect 28491 30549 28503 30552
rect 28445 30543 28503 30549
rect 29086 30540 29092 30592
rect 29144 30540 29150 30592
rect 29656 30580 29684 30688
rect 29730 30676 29736 30728
rect 29788 30716 29794 30728
rect 29825 30719 29883 30725
rect 29825 30716 29837 30719
rect 29788 30688 29837 30716
rect 29788 30676 29794 30688
rect 29825 30685 29837 30688
rect 29871 30685 29883 30719
rect 29825 30679 29883 30685
rect 30009 30719 30067 30725
rect 30009 30685 30021 30719
rect 30055 30716 30067 30719
rect 30374 30716 30380 30728
rect 30055 30688 30380 30716
rect 30055 30685 30067 30688
rect 30009 30679 30067 30685
rect 30374 30676 30380 30688
rect 30432 30676 30438 30728
rect 30558 30676 30564 30728
rect 30616 30676 30622 30728
rect 30745 30719 30803 30725
rect 30745 30685 30757 30719
rect 30791 30685 30803 30719
rect 36188 30716 36216 30744
rect 36633 30719 36691 30725
rect 36633 30716 36645 30719
rect 36188 30688 36645 30716
rect 30745 30679 30803 30685
rect 36633 30685 36645 30688
rect 36679 30685 36691 30719
rect 36633 30679 36691 30685
rect 36781 30719 36839 30725
rect 36781 30685 36793 30719
rect 36827 30716 36839 30719
rect 36827 30685 36860 30716
rect 36781 30679 36860 30685
rect 29917 30651 29975 30657
rect 29917 30617 29929 30651
rect 29963 30648 29975 30651
rect 30760 30648 30788 30679
rect 33778 30648 33784 30660
rect 29963 30620 30788 30648
rect 30852 30620 33784 30648
rect 29963 30617 29975 30620
rect 29917 30611 29975 30617
rect 30852 30580 30880 30620
rect 33778 30608 33784 30620
rect 33836 30648 33842 30660
rect 34330 30648 34336 30660
rect 33836 30620 34336 30648
rect 33836 30608 33842 30620
rect 34330 30608 34336 30620
rect 34388 30608 34394 30660
rect 36202 30620 36676 30648
rect 36648 30592 36676 30620
rect 29656 30552 30880 30580
rect 30929 30583 30987 30589
rect 30929 30549 30941 30583
rect 30975 30580 30987 30583
rect 31570 30580 31576 30592
rect 30975 30552 31576 30580
rect 30975 30549 30987 30552
rect 30929 30543 30987 30549
rect 31570 30540 31576 30552
rect 31628 30540 31634 30592
rect 36630 30540 36636 30592
rect 36688 30540 36694 30592
rect 36832 30580 36860 30679
rect 36998 30676 37004 30728
rect 37056 30676 37062 30728
rect 37108 30725 37136 30756
rect 37642 30744 37648 30796
rect 37700 30744 37706 30796
rect 40402 30744 40408 30796
rect 40460 30744 40466 30796
rect 37098 30719 37156 30725
rect 37098 30685 37110 30719
rect 37144 30685 37156 30719
rect 37098 30679 37156 30685
rect 37366 30676 37372 30728
rect 37424 30676 37430 30728
rect 40313 30719 40371 30725
rect 40313 30716 40325 30719
rect 39132 30688 40325 30716
rect 36906 30608 36912 30660
rect 36964 30608 36970 30660
rect 38930 30648 38936 30660
rect 38870 30620 38936 30648
rect 38930 30608 38936 30620
rect 38988 30608 38994 30660
rect 37918 30580 37924 30592
rect 36832 30552 37924 30580
rect 37918 30540 37924 30552
rect 37976 30540 37982 30592
rect 38286 30540 38292 30592
rect 38344 30580 38350 30592
rect 39132 30589 39160 30688
rect 40313 30685 40325 30688
rect 40359 30685 40371 30719
rect 40313 30679 40371 30685
rect 40862 30676 40868 30728
rect 40920 30676 40926 30728
rect 40034 30608 40040 30660
rect 40092 30648 40098 30660
rect 40681 30651 40739 30657
rect 40681 30648 40693 30651
rect 40092 30620 40693 30648
rect 40092 30608 40098 30620
rect 40681 30617 40693 30620
rect 40727 30617 40739 30651
rect 40681 30611 40739 30617
rect 39117 30583 39175 30589
rect 39117 30580 39129 30583
rect 38344 30552 39129 30580
rect 38344 30540 38350 30552
rect 39117 30549 39129 30552
rect 39163 30549 39175 30583
rect 39117 30543 39175 30549
rect 39666 30540 39672 30592
rect 39724 30580 39730 30592
rect 39853 30583 39911 30589
rect 39853 30580 39865 30583
rect 39724 30552 39865 30580
rect 39724 30540 39730 30552
rect 39853 30549 39865 30552
rect 39899 30549 39911 30583
rect 39853 30543 39911 30549
rect 40221 30583 40279 30589
rect 40221 30549 40233 30583
rect 40267 30580 40279 30583
rect 40310 30580 40316 30592
rect 40267 30552 40316 30580
rect 40267 30549 40279 30552
rect 40221 30543 40279 30549
rect 40310 30540 40316 30552
rect 40368 30580 40374 30592
rect 40586 30580 40592 30592
rect 40368 30552 40592 30580
rect 40368 30540 40374 30552
rect 40586 30540 40592 30552
rect 40644 30540 40650 30592
rect 1104 30490 42504 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 42504 30490
rect 1104 30416 42504 30438
rect 3053 30379 3111 30385
rect 3053 30345 3065 30379
rect 3099 30376 3111 30379
rect 3142 30376 3148 30388
rect 3099 30348 3148 30376
rect 3099 30345 3111 30348
rect 3053 30339 3111 30345
rect 3142 30336 3148 30348
rect 3200 30336 3206 30388
rect 3234 30336 3240 30388
rect 3292 30376 3298 30388
rect 4062 30376 4068 30388
rect 3292 30348 4068 30376
rect 3292 30336 3298 30348
rect 4062 30336 4068 30348
rect 4120 30336 4126 30388
rect 4157 30379 4215 30385
rect 4157 30345 4169 30379
rect 4203 30376 4215 30379
rect 5626 30376 5632 30388
rect 4203 30348 4936 30376
rect 4203 30345 4215 30348
rect 4157 30339 4215 30345
rect 2866 30268 2872 30320
rect 2924 30268 2930 30320
rect 3605 30311 3663 30317
rect 3605 30308 3617 30311
rect 3472 30280 3617 30308
rect 2958 30200 2964 30252
rect 3016 30240 3022 30252
rect 3145 30243 3203 30249
rect 3145 30240 3157 30243
rect 3016 30212 3157 30240
rect 3016 30200 3022 30212
rect 3145 30209 3157 30212
rect 3191 30209 3203 30243
rect 3145 30203 3203 30209
rect 3326 30200 3332 30252
rect 3384 30240 3390 30252
rect 3472 30249 3500 30280
rect 3605 30277 3617 30280
rect 3651 30277 3663 30311
rect 3605 30271 3663 30277
rect 3786 30268 3792 30320
rect 3844 30268 3850 30320
rect 4341 30311 4399 30317
rect 4341 30277 4353 30311
rect 4387 30308 4399 30311
rect 4908 30308 4936 30348
rect 5552 30348 5632 30376
rect 5552 30308 5580 30348
rect 5626 30336 5632 30348
rect 5684 30336 5690 30388
rect 6086 30336 6092 30388
rect 6144 30376 6150 30388
rect 6365 30379 6423 30385
rect 6365 30376 6377 30379
rect 6144 30348 6377 30376
rect 6144 30336 6150 30348
rect 6365 30345 6377 30348
rect 6411 30345 6423 30379
rect 6365 30339 6423 30345
rect 6914 30336 6920 30388
rect 6972 30376 6978 30388
rect 11057 30379 11115 30385
rect 6972 30348 8156 30376
rect 6972 30336 6978 30348
rect 4387 30280 4844 30308
rect 4908 30280 5580 30308
rect 5746 30311 5804 30317
rect 4387 30277 4399 30280
rect 4341 30271 4399 30277
rect 3421 30243 3500 30249
rect 3421 30240 3433 30243
rect 3384 30212 3433 30240
rect 3384 30200 3390 30212
rect 3421 30209 3433 30212
rect 3467 30212 3500 30243
rect 3529 30243 3587 30249
rect 3467 30209 3479 30212
rect 3421 30203 3479 30209
rect 3529 30209 3541 30243
rect 3575 30240 3587 30243
rect 3973 30243 4031 30249
rect 3973 30240 3985 30243
rect 3575 30238 3648 30240
rect 3575 30212 3740 30238
rect 3575 30209 3587 30212
rect 3620 30210 3740 30212
rect 3529 30203 3587 30209
rect 3712 30116 3740 30210
rect 3912 30212 3985 30240
rect 3694 30064 3700 30116
rect 3752 30064 3758 30116
rect 3786 29996 3792 30048
rect 3844 29996 3850 30048
rect 3912 30036 3940 30212
rect 3973 30209 3985 30212
rect 4019 30209 4031 30243
rect 3973 30203 4031 30209
rect 4062 30200 4068 30252
rect 4120 30240 4126 30252
rect 4157 30243 4215 30249
rect 4157 30240 4169 30243
rect 4120 30212 4169 30240
rect 4120 30200 4126 30212
rect 4157 30209 4169 30212
rect 4203 30209 4215 30243
rect 4157 30203 4215 30209
rect 4246 30200 4252 30252
rect 4304 30200 4310 30252
rect 4430 30200 4436 30252
rect 4488 30200 4494 30252
rect 4522 30200 4528 30252
rect 4580 30200 4586 30252
rect 4706 30200 4712 30252
rect 4764 30200 4770 30252
rect 4816 30249 4844 30280
rect 5746 30277 5758 30311
rect 5792 30308 5804 30311
rect 6104 30308 6132 30336
rect 5792 30280 6132 30308
rect 5792 30277 5804 30280
rect 5746 30271 5804 30277
rect 6270 30268 6276 30320
rect 6328 30308 6334 30320
rect 6546 30308 6552 30320
rect 6328 30280 6552 30308
rect 6328 30268 6334 30280
rect 6546 30268 6552 30280
rect 6604 30308 6610 30320
rect 6604 30280 6670 30308
rect 6604 30268 6610 30280
rect 4801 30243 4859 30249
rect 4801 30209 4813 30243
rect 4847 30209 4859 30243
rect 4801 30203 4859 30209
rect 4890 30200 4896 30252
rect 4948 30200 4954 30252
rect 8128 30249 8156 30348
rect 11057 30345 11069 30379
rect 11103 30345 11115 30379
rect 11057 30339 11115 30345
rect 10134 30268 10140 30320
rect 10192 30268 10198 30320
rect 11072 30308 11100 30339
rect 11146 30336 11152 30388
rect 11204 30376 11210 30388
rect 11517 30379 11575 30385
rect 11517 30376 11529 30379
rect 11204 30348 11529 30376
rect 11204 30336 11210 30348
rect 11517 30345 11529 30348
rect 11563 30345 11575 30379
rect 11517 30339 11575 30345
rect 15286 30336 15292 30388
rect 15344 30336 15350 30388
rect 15654 30336 15660 30388
rect 15712 30376 15718 30388
rect 16209 30379 16267 30385
rect 16209 30376 16221 30379
rect 15712 30348 16221 30376
rect 15712 30336 15718 30348
rect 16209 30345 16221 30348
rect 16255 30345 16267 30379
rect 17770 30376 17776 30388
rect 16209 30339 16267 30345
rect 16960 30348 17776 30376
rect 11885 30311 11943 30317
rect 11072 30280 11836 30308
rect 5629 30243 5687 30249
rect 5629 30240 5641 30243
rect 5000 30212 5641 30240
rect 4448 30172 4476 30200
rect 5000 30172 5028 30212
rect 5629 30209 5641 30212
rect 5675 30209 5687 30243
rect 5629 30203 5687 30209
rect 8113 30243 8171 30249
rect 8113 30209 8125 30243
rect 8159 30209 8171 30243
rect 8113 30203 8171 30209
rect 10410 30200 10416 30252
rect 10468 30200 10474 30252
rect 10686 30240 10692 30252
rect 10520 30212 10692 30240
rect 4448 30144 5028 30172
rect 5261 30175 5319 30181
rect 5261 30141 5273 30175
rect 5307 30141 5319 30175
rect 5261 30135 5319 30141
rect 5537 30175 5595 30181
rect 5537 30141 5549 30175
rect 5583 30141 5595 30175
rect 5537 30135 5595 30141
rect 4246 30064 4252 30116
rect 4304 30104 4310 30116
rect 5276 30104 5304 30135
rect 4304 30076 5304 30104
rect 5552 30104 5580 30135
rect 7834 30132 7840 30184
rect 7892 30132 7898 30184
rect 8941 30175 8999 30181
rect 8941 30141 8953 30175
rect 8987 30172 8999 30175
rect 9030 30172 9036 30184
rect 8987 30144 9036 30172
rect 8987 30141 8999 30144
rect 8941 30135 8999 30141
rect 9030 30132 9036 30144
rect 9088 30132 9094 30184
rect 10321 30175 10379 30181
rect 10321 30141 10333 30175
rect 10367 30172 10379 30175
rect 10520 30172 10548 30212
rect 10686 30200 10692 30212
rect 10744 30240 10750 30252
rect 10873 30243 10931 30249
rect 10873 30240 10885 30243
rect 10744 30212 10885 30240
rect 10744 30200 10750 30212
rect 10873 30209 10885 30212
rect 10919 30209 10931 30243
rect 10873 30203 10931 30209
rect 10962 30200 10968 30252
rect 11020 30240 11026 30252
rect 11057 30243 11115 30249
rect 11057 30240 11069 30243
rect 11020 30212 11069 30240
rect 11020 30200 11026 30212
rect 11057 30209 11069 30212
rect 11103 30209 11115 30243
rect 11808 30240 11836 30280
rect 11885 30277 11897 30311
rect 11931 30308 11943 30311
rect 12710 30308 12716 30320
rect 11931 30280 12716 30308
rect 11931 30277 11943 30280
rect 11885 30271 11943 30277
rect 12710 30268 12716 30280
rect 12768 30268 12774 30320
rect 15304 30308 15332 30336
rect 15746 30308 15752 30320
rect 14214 30280 15752 30308
rect 15746 30268 15752 30280
rect 15804 30268 15810 30320
rect 16393 30311 16451 30317
rect 16393 30277 16405 30311
rect 16439 30308 16451 30311
rect 16482 30308 16488 30320
rect 16439 30280 16488 30308
rect 16439 30277 16451 30280
rect 16393 30271 16451 30277
rect 16482 30268 16488 30280
rect 16540 30308 16546 30320
rect 16960 30308 16988 30348
rect 17770 30336 17776 30348
rect 17828 30336 17834 30388
rect 18690 30336 18696 30388
rect 18748 30336 18754 30388
rect 19705 30379 19763 30385
rect 19705 30345 19717 30379
rect 19751 30376 19763 30379
rect 20162 30376 20168 30388
rect 19751 30348 20168 30376
rect 19751 30345 19763 30348
rect 19705 30339 19763 30345
rect 20162 30336 20168 30348
rect 20220 30336 20226 30388
rect 20530 30336 20536 30388
rect 20588 30376 20594 30388
rect 20625 30379 20683 30385
rect 20625 30376 20637 30379
rect 20588 30348 20637 30376
rect 20588 30336 20594 30348
rect 20625 30345 20637 30348
rect 20671 30345 20683 30379
rect 20625 30339 20683 30345
rect 20714 30336 20720 30388
rect 20772 30376 20778 30388
rect 20993 30379 21051 30385
rect 20993 30376 21005 30379
rect 20772 30348 21005 30376
rect 20772 30336 20778 30348
rect 20993 30345 21005 30348
rect 21039 30345 21051 30379
rect 22094 30376 22100 30388
rect 20993 30339 21051 30345
rect 21652 30348 22100 30376
rect 16540 30280 16988 30308
rect 16540 30268 16546 30280
rect 17034 30268 17040 30320
rect 17092 30308 17098 30320
rect 17313 30311 17371 30317
rect 17313 30308 17325 30311
rect 17092 30280 17325 30308
rect 17092 30268 17098 30280
rect 17313 30277 17325 30280
rect 17359 30277 17371 30311
rect 17313 30271 17371 30277
rect 17402 30268 17408 30320
rect 17460 30308 17466 30320
rect 17460 30280 17812 30308
rect 17460 30268 17466 30280
rect 11808 30212 12112 30240
rect 11057 30203 11115 30209
rect 10367 30144 10548 30172
rect 10367 30141 10379 30144
rect 10321 30135 10379 30141
rect 10594 30132 10600 30184
rect 10652 30172 10658 30184
rect 10781 30175 10839 30181
rect 10781 30172 10793 30175
rect 10652 30144 10793 30172
rect 10652 30132 10658 30144
rect 10781 30141 10793 30144
rect 10827 30172 10839 30175
rect 10980 30172 11008 30200
rect 10827 30144 11008 30172
rect 10827 30141 10839 30144
rect 10781 30135 10839 30141
rect 11146 30132 11152 30184
rect 11204 30172 11210 30184
rect 12084 30181 12112 30212
rect 14826 30200 14832 30252
rect 14884 30200 14890 30252
rect 15010 30200 15016 30252
rect 15068 30200 15074 30252
rect 15194 30200 15200 30252
rect 15252 30200 15258 30252
rect 15286 30200 15292 30252
rect 15344 30200 15350 30252
rect 15396 30212 15884 30240
rect 11977 30175 12035 30181
rect 11977 30172 11989 30175
rect 11204 30144 11989 30172
rect 11204 30132 11210 30144
rect 11977 30141 11989 30144
rect 12023 30141 12035 30175
rect 11977 30135 12035 30141
rect 12069 30175 12127 30181
rect 12069 30141 12081 30175
rect 12115 30172 12127 30175
rect 12250 30172 12256 30184
rect 12115 30144 12256 30172
rect 12115 30141 12127 30144
rect 12069 30135 12127 30141
rect 12250 30132 12256 30144
rect 12308 30132 12314 30184
rect 12713 30175 12771 30181
rect 12713 30172 12725 30175
rect 12406 30144 12725 30172
rect 5626 30104 5632 30116
rect 5552 30076 5632 30104
rect 4304 30064 4310 30076
rect 5626 30064 5632 30076
rect 5684 30064 5690 30116
rect 10870 30064 10876 30116
rect 10928 30104 10934 30116
rect 12406 30104 12434 30144
rect 12713 30141 12725 30144
rect 12759 30141 12771 30175
rect 12713 30135 12771 30141
rect 12986 30132 12992 30184
rect 13044 30132 13050 30184
rect 14737 30175 14795 30181
rect 14737 30141 14749 30175
rect 14783 30172 14795 30175
rect 14918 30172 14924 30184
rect 14783 30144 14924 30172
rect 14783 30141 14795 30144
rect 14737 30135 14795 30141
rect 14918 30132 14924 30144
rect 14976 30132 14982 30184
rect 15105 30175 15163 30181
rect 15105 30141 15117 30175
rect 15151 30172 15163 30175
rect 15396 30172 15424 30212
rect 15151 30144 15424 30172
rect 15151 30141 15163 30144
rect 15105 30135 15163 30141
rect 15470 30132 15476 30184
rect 15528 30132 15534 30184
rect 15856 30172 15884 30212
rect 15930 30200 15936 30252
rect 15988 30200 15994 30252
rect 16114 30200 16120 30252
rect 16172 30200 16178 30252
rect 17497 30243 17555 30249
rect 17497 30240 17509 30243
rect 17420 30212 17509 30240
rect 17420 30184 17448 30212
rect 17497 30209 17509 30212
rect 17543 30209 17555 30243
rect 17497 30203 17555 30209
rect 17681 30243 17739 30249
rect 17681 30209 17693 30243
rect 17727 30209 17739 30243
rect 17681 30203 17739 30209
rect 17034 30172 17040 30184
rect 15856 30144 17040 30172
rect 17034 30132 17040 30144
rect 17092 30132 17098 30184
rect 17402 30132 17408 30184
rect 17460 30132 17466 30184
rect 10928 30076 12434 30104
rect 10928 30064 10934 30076
rect 15562 30064 15568 30116
rect 15620 30104 15626 30116
rect 16393 30107 16451 30113
rect 16393 30104 16405 30107
rect 15620 30076 16405 30104
rect 15620 30064 15626 30076
rect 16393 30073 16405 30076
rect 16439 30073 16451 30107
rect 17696 30104 17724 30203
rect 17784 30172 17812 30280
rect 17954 30268 17960 30320
rect 18012 30308 18018 30320
rect 18141 30311 18199 30317
rect 18141 30308 18153 30311
rect 18012 30280 18153 30308
rect 18012 30268 18018 30280
rect 18141 30277 18153 30280
rect 18187 30308 18199 30311
rect 18187 30280 19104 30308
rect 18187 30277 18199 30280
rect 18141 30271 18199 30277
rect 18230 30200 18236 30252
rect 18288 30200 18294 30252
rect 19076 30249 19104 30280
rect 19610 30268 19616 30320
rect 19668 30308 19674 30320
rect 19668 30280 20944 30308
rect 19668 30268 19674 30280
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19337 30243 19395 30249
rect 19337 30240 19349 30243
rect 19107 30212 19349 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 19337 30209 19349 30212
rect 19383 30209 19395 30243
rect 19337 30203 19395 30209
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30209 19579 30243
rect 19521 30203 19579 30209
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30240 20315 30243
rect 20622 30240 20628 30252
rect 20303 30212 20628 30240
rect 20303 30209 20315 30212
rect 20257 30203 20315 30209
rect 17957 30175 18015 30181
rect 17957 30172 17969 30175
rect 17784 30144 17969 30172
rect 17957 30141 17969 30144
rect 18003 30172 18015 30175
rect 18506 30172 18512 30184
rect 18003 30144 18512 30172
rect 18003 30141 18015 30144
rect 17957 30135 18015 30141
rect 18506 30132 18512 30144
rect 18564 30132 18570 30184
rect 18966 30132 18972 30184
rect 19024 30172 19030 30184
rect 19536 30172 19564 30203
rect 20622 30200 20628 30212
rect 20680 30200 20686 30252
rect 20916 30249 20944 30280
rect 20901 30243 20959 30249
rect 20901 30209 20913 30243
rect 20947 30209 20959 30243
rect 20901 30203 20959 30209
rect 21082 30200 21088 30252
rect 21140 30200 21146 30252
rect 21652 30249 21680 30348
rect 22094 30336 22100 30348
rect 22152 30376 22158 30388
rect 22370 30376 22376 30388
rect 22152 30348 22376 30376
rect 22152 30336 22158 30348
rect 22370 30336 22376 30348
rect 22428 30336 22434 30388
rect 22646 30336 22652 30388
rect 22704 30376 22710 30388
rect 24305 30379 24363 30385
rect 22704 30348 23428 30376
rect 22704 30336 22710 30348
rect 21726 30268 21732 30320
rect 21784 30308 21790 30320
rect 22741 30311 22799 30317
rect 21784 30280 22232 30308
rect 21784 30268 21790 30280
rect 21453 30243 21511 30249
rect 21453 30209 21465 30243
rect 21499 30209 21511 30243
rect 21453 30203 21511 30209
rect 21637 30243 21695 30249
rect 21637 30209 21649 30243
rect 21683 30209 21695 30243
rect 21637 30203 21695 30209
rect 19024 30144 19564 30172
rect 19024 30132 19030 30144
rect 19794 30132 19800 30184
rect 19852 30172 19858 30184
rect 21100 30172 21128 30200
rect 19852 30144 21128 30172
rect 19852 30132 19858 30144
rect 20254 30104 20260 30116
rect 16393 30067 16451 30073
rect 17420 30076 20260 30104
rect 3970 30036 3976 30048
rect 3912 30008 3976 30036
rect 3970 29996 3976 30008
rect 4028 29996 4034 30048
rect 4062 29996 4068 30048
rect 4120 30036 4126 30048
rect 4522 30036 4528 30048
rect 4120 30008 4528 30036
rect 4120 29996 4126 30008
rect 4522 29996 4528 30008
rect 4580 29996 4586 30048
rect 5169 30039 5227 30045
rect 5169 30005 5181 30039
rect 5215 30036 5227 30039
rect 5350 30036 5356 30048
rect 5215 30008 5356 30036
rect 5215 30005 5227 30008
rect 5169 29999 5227 30005
rect 5350 29996 5356 30008
rect 5408 29996 5414 30048
rect 5534 29996 5540 30048
rect 5592 30036 5598 30048
rect 5905 30039 5963 30045
rect 5905 30036 5917 30039
rect 5592 30008 5917 30036
rect 5592 29996 5598 30008
rect 5905 30005 5917 30008
rect 5951 30005 5963 30039
rect 5905 29999 5963 30005
rect 9306 29996 9312 30048
rect 9364 30036 9370 30048
rect 9493 30039 9551 30045
rect 9493 30036 9505 30039
rect 9364 30008 9505 30036
rect 9364 29996 9370 30008
rect 9493 30005 9505 30008
rect 9539 30005 9551 30039
rect 9493 29999 9551 30005
rect 15286 29996 15292 30048
rect 15344 30036 15350 30048
rect 15841 30039 15899 30045
rect 15841 30036 15853 30039
rect 15344 30008 15853 30036
rect 15344 29996 15350 30008
rect 15841 30005 15853 30008
rect 15887 30036 15899 30039
rect 16298 30036 16304 30048
rect 15887 30008 16304 30036
rect 15887 30005 15899 30008
rect 15841 29999 15899 30005
rect 16298 29996 16304 30008
rect 16356 29996 16362 30048
rect 16942 29996 16948 30048
rect 17000 30036 17006 30048
rect 17420 30036 17448 30076
rect 20254 30064 20260 30076
rect 20312 30104 20318 30116
rect 20809 30107 20867 30113
rect 20312 30076 20668 30104
rect 20312 30064 20318 30076
rect 17000 30008 17448 30036
rect 17000 29996 17006 30008
rect 17954 29996 17960 30048
rect 18012 30036 18018 30048
rect 18598 30036 18604 30048
rect 18012 30008 18604 30036
rect 18012 29996 18018 30008
rect 18598 29996 18604 30008
rect 18656 29996 18662 30048
rect 20640 30045 20668 30076
rect 20809 30073 20821 30107
rect 20855 30104 20867 30107
rect 21174 30104 21180 30116
rect 20855 30076 21180 30104
rect 20855 30073 20867 30076
rect 20809 30067 20867 30073
rect 21174 30064 21180 30076
rect 21232 30064 21238 30116
rect 20625 30039 20683 30045
rect 20625 30005 20637 30039
rect 20671 30005 20683 30039
rect 21468 30036 21496 30203
rect 21818 30200 21824 30252
rect 21876 30200 21882 30252
rect 22204 30249 22232 30280
rect 22741 30277 22753 30311
rect 22787 30308 22799 30311
rect 22830 30308 22836 30320
rect 22787 30280 22836 30308
rect 22787 30277 22799 30280
rect 22741 30271 22799 30277
rect 22830 30268 22836 30280
rect 22888 30268 22894 30320
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22097 30243 22155 30249
rect 22097 30209 22109 30243
rect 22143 30209 22155 30243
rect 22097 30203 22155 30209
rect 22189 30243 22247 30249
rect 22189 30209 22201 30243
rect 22235 30209 22247 30243
rect 22189 30203 22247 30209
rect 21545 30175 21603 30181
rect 21545 30141 21557 30175
rect 21591 30172 21603 30175
rect 21910 30172 21916 30184
rect 21591 30144 21916 30172
rect 21591 30141 21603 30144
rect 21545 30135 21603 30141
rect 21910 30132 21916 30144
rect 21968 30172 21974 30184
rect 22020 30172 22048 30203
rect 21968 30144 22048 30172
rect 21968 30132 21974 30144
rect 22002 30064 22008 30116
rect 22060 30104 22066 30116
rect 22112 30104 22140 30203
rect 22370 30200 22376 30252
rect 22428 30240 22434 30252
rect 23400 30249 23428 30348
rect 24305 30345 24317 30379
rect 24351 30376 24363 30379
rect 24578 30376 24584 30388
rect 24351 30348 24584 30376
rect 24351 30345 24363 30348
rect 24305 30339 24363 30345
rect 24578 30336 24584 30348
rect 24636 30376 24642 30388
rect 25225 30379 25283 30385
rect 25225 30376 25237 30379
rect 24636 30348 25237 30376
rect 24636 30336 24642 30348
rect 25225 30345 25237 30348
rect 25271 30345 25283 30379
rect 25225 30339 25283 30345
rect 25317 30379 25375 30385
rect 25317 30345 25329 30379
rect 25363 30376 25375 30379
rect 25590 30376 25596 30388
rect 25363 30348 25596 30376
rect 25363 30345 25375 30348
rect 25317 30339 25375 30345
rect 25590 30336 25596 30348
rect 25648 30336 25654 30388
rect 30469 30379 30527 30385
rect 30469 30345 30481 30379
rect 30515 30376 30527 30379
rect 30558 30376 30564 30388
rect 30515 30348 30564 30376
rect 30515 30345 30527 30348
rect 30469 30339 30527 30345
rect 30558 30336 30564 30348
rect 30616 30336 30622 30388
rect 30834 30336 30840 30388
rect 30892 30336 30898 30388
rect 34790 30336 34796 30388
rect 34848 30376 34854 30388
rect 34848 30348 35572 30376
rect 34848 30336 34854 30348
rect 23569 30311 23627 30317
rect 23569 30277 23581 30311
rect 23615 30308 23627 30311
rect 24670 30308 24676 30320
rect 23615 30280 24676 30308
rect 23615 30277 23627 30280
rect 23569 30271 23627 30277
rect 24670 30268 24676 30280
rect 24728 30308 24734 30320
rect 24728 30280 24992 30308
rect 24728 30268 24734 30280
rect 23201 30243 23259 30249
rect 23201 30240 23213 30243
rect 22428 30212 23213 30240
rect 22428 30200 22434 30212
rect 23201 30209 23213 30212
rect 23247 30209 23259 30243
rect 23201 30203 23259 30209
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 23934 30200 23940 30252
rect 23992 30240 23998 30252
rect 24964 30249 24992 30280
rect 25424 30280 26280 30308
rect 25424 30249 25452 30280
rect 26252 30252 26280 30280
rect 26878 30268 26884 30320
rect 26936 30308 26942 30320
rect 27249 30311 27307 30317
rect 27249 30308 27261 30311
rect 26936 30280 27261 30308
rect 26936 30268 26942 30280
rect 27249 30277 27261 30280
rect 27295 30277 27307 30311
rect 27249 30271 27307 30277
rect 28810 30268 28816 30320
rect 28868 30268 28874 30320
rect 30098 30268 30104 30320
rect 30156 30268 30162 30320
rect 30301 30311 30359 30317
rect 30301 30308 30313 30311
rect 30208 30280 30313 30308
rect 24213 30243 24271 30249
rect 24213 30240 24225 30243
rect 23992 30212 24225 30240
rect 23992 30200 23998 30212
rect 24213 30209 24225 30212
rect 24259 30209 24271 30243
rect 24213 30203 24271 30209
rect 24949 30243 25007 30249
rect 24949 30209 24961 30243
rect 24995 30209 25007 30243
rect 24949 30203 25007 30209
rect 25409 30243 25467 30249
rect 25409 30209 25421 30243
rect 25455 30209 25467 30243
rect 25409 30203 25467 30209
rect 25774 30200 25780 30252
rect 25832 30200 25838 30252
rect 25958 30200 25964 30252
rect 26016 30200 26022 30252
rect 26234 30200 26240 30252
rect 26292 30200 26298 30252
rect 26421 30243 26479 30249
rect 26421 30209 26433 30243
rect 26467 30240 26479 30243
rect 26513 30243 26571 30249
rect 26513 30240 26525 30243
rect 26467 30212 26525 30240
rect 26467 30209 26479 30212
rect 26421 30203 26479 30209
rect 26513 30209 26525 30212
rect 26559 30209 26571 30243
rect 26513 30203 26571 30209
rect 28350 30200 28356 30252
rect 28408 30200 28414 30252
rect 28626 30200 28632 30252
rect 28684 30240 28690 30252
rect 29365 30243 29423 30249
rect 29365 30240 29377 30243
rect 28684 30212 29377 30240
rect 28684 30200 28690 30212
rect 29365 30209 29377 30212
rect 29411 30209 29423 30243
rect 29365 30203 29423 30209
rect 29546 30200 29552 30252
rect 29604 30200 29610 30252
rect 29730 30200 29736 30252
rect 29788 30200 29794 30252
rect 29822 30200 29828 30252
rect 29880 30240 29886 30252
rect 30208 30240 30236 30280
rect 30301 30277 30313 30280
rect 30347 30308 30359 30311
rect 30929 30311 30987 30317
rect 30929 30308 30941 30311
rect 30347 30280 30941 30308
rect 30347 30277 30359 30280
rect 30301 30271 30359 30277
rect 30929 30277 30941 30280
rect 30975 30277 30987 30311
rect 30929 30271 30987 30277
rect 32490 30268 32496 30320
rect 32548 30308 32554 30320
rect 32548 30280 33732 30308
rect 32548 30268 32554 30280
rect 30561 30243 30619 30249
rect 30561 30240 30573 30243
rect 29880 30212 30236 30240
rect 30300 30212 30573 30240
rect 29880 30200 29886 30212
rect 22465 30175 22523 30181
rect 22465 30141 22477 30175
rect 22511 30172 22523 30175
rect 23109 30175 23167 30181
rect 23109 30172 23121 30175
rect 22511 30144 23121 30172
rect 22511 30141 22523 30144
rect 22465 30135 22523 30141
rect 23109 30141 23121 30144
rect 23155 30141 23167 30175
rect 23109 30135 23167 30141
rect 22060 30076 22140 30104
rect 22060 30064 22066 30076
rect 22186 30064 22192 30116
rect 22244 30104 22250 30116
rect 22557 30107 22615 30113
rect 22557 30104 22569 30107
rect 22244 30076 22569 30104
rect 22244 30064 22250 30076
rect 22557 30073 22569 30076
rect 22603 30073 22615 30107
rect 23124 30104 23152 30135
rect 24302 30132 24308 30184
rect 24360 30172 24366 30184
rect 24397 30175 24455 30181
rect 24397 30172 24409 30175
rect 24360 30144 24409 30172
rect 24360 30132 24366 30144
rect 24397 30141 24409 30144
rect 24443 30141 24455 30175
rect 24397 30135 24455 30141
rect 26786 30132 26792 30184
rect 26844 30132 26850 30184
rect 26970 30132 26976 30184
rect 27028 30132 27034 30184
rect 29748 30172 29776 30200
rect 27080 30144 29776 30172
rect 24946 30104 24952 30116
rect 23124 30076 24952 30104
rect 22557 30067 22615 30073
rect 24946 30064 24952 30076
rect 25004 30104 25010 30116
rect 25041 30107 25099 30113
rect 25041 30104 25053 30107
rect 25004 30076 25053 30104
rect 25004 30064 25010 30076
rect 25041 30073 25053 30076
rect 25087 30073 25099 30107
rect 25041 30067 25099 30073
rect 25685 30107 25743 30113
rect 25685 30073 25697 30107
rect 25731 30104 25743 30107
rect 26602 30104 26608 30116
rect 25731 30076 26608 30104
rect 25731 30073 25743 30076
rect 25685 30067 25743 30073
rect 26602 30064 26608 30076
rect 26660 30064 26666 30116
rect 26804 30104 26832 30132
rect 27080 30104 27108 30144
rect 30190 30132 30196 30184
rect 30248 30172 30254 30184
rect 30300 30172 30328 30212
rect 30561 30209 30573 30212
rect 30607 30209 30619 30243
rect 30561 30203 30619 30209
rect 30742 30200 30748 30252
rect 30800 30240 30806 30252
rect 31478 30240 31484 30252
rect 30800 30212 31484 30240
rect 30800 30200 30806 30212
rect 31478 30200 31484 30212
rect 31536 30200 31542 30252
rect 31570 30200 31576 30252
rect 31628 30200 31634 30252
rect 31662 30200 31668 30252
rect 31720 30200 31726 30252
rect 33704 30249 33732 30280
rect 34054 30268 34060 30320
rect 34112 30268 34118 30320
rect 35544 30317 35572 30348
rect 36262 30336 36268 30388
rect 36320 30336 36326 30388
rect 36906 30376 36912 30388
rect 36648 30348 36912 30376
rect 35324 30311 35382 30317
rect 35324 30277 35336 30311
rect 35370 30277 35382 30311
rect 35324 30271 35382 30277
rect 35529 30311 35587 30317
rect 35529 30277 35541 30311
rect 35575 30308 35587 30311
rect 35986 30308 35992 30320
rect 35575 30280 35992 30308
rect 35575 30277 35587 30280
rect 35529 30271 35587 30277
rect 31941 30243 31999 30249
rect 31941 30209 31953 30243
rect 31987 30240 31999 30243
rect 33137 30243 33195 30249
rect 33137 30240 33149 30243
rect 31987 30212 33149 30240
rect 31987 30209 31999 30212
rect 31941 30203 31999 30209
rect 33137 30209 33149 30212
rect 33183 30209 33195 30243
rect 33137 30203 33195 30209
rect 33689 30243 33747 30249
rect 33689 30209 33701 30243
rect 33735 30209 33747 30243
rect 33689 30203 33747 30209
rect 34701 30243 34759 30249
rect 34701 30209 34713 30243
rect 34747 30240 34759 30243
rect 35344 30240 35372 30271
rect 35986 30268 35992 30280
rect 36044 30268 36050 30320
rect 36648 30317 36676 30348
rect 36906 30336 36912 30348
rect 36964 30336 36970 30388
rect 37826 30336 37832 30388
rect 37884 30336 37890 30388
rect 37918 30336 37924 30388
rect 37976 30376 37982 30388
rect 38562 30376 38568 30388
rect 37976 30348 38568 30376
rect 37976 30336 37982 30348
rect 38562 30336 38568 30348
rect 38620 30336 38626 30388
rect 36633 30311 36691 30317
rect 36633 30277 36645 30311
rect 36679 30277 36691 30311
rect 36633 30271 36691 30277
rect 37642 30268 37648 30320
rect 37700 30268 37706 30320
rect 38289 30311 38347 30317
rect 38289 30277 38301 30311
rect 38335 30308 38347 30311
rect 38838 30308 38844 30320
rect 38335 30280 38844 30308
rect 38335 30277 38347 30280
rect 38289 30271 38347 30277
rect 38838 30268 38844 30280
rect 38896 30268 38902 30320
rect 39574 30268 39580 30320
rect 39632 30308 39638 30320
rect 40126 30308 40132 30320
rect 39632 30280 40132 30308
rect 39632 30268 39638 30280
rect 40126 30268 40132 30280
rect 40184 30308 40190 30320
rect 40589 30311 40647 30317
rect 40589 30308 40601 30311
rect 40184 30280 40601 30308
rect 40184 30268 40190 30280
rect 40589 30277 40601 30280
rect 40635 30277 40647 30311
rect 40589 30271 40647 30277
rect 40788 30280 41414 30308
rect 35618 30240 35624 30252
rect 34747 30212 35296 30240
rect 35344 30212 35624 30240
rect 34747 30209 34759 30212
rect 34701 30203 34759 30209
rect 30248 30144 30328 30172
rect 30248 30132 30254 30144
rect 30374 30132 30380 30184
rect 30432 30172 30438 30184
rect 31113 30175 31171 30181
rect 31113 30172 31125 30175
rect 30432 30144 31125 30172
rect 30432 30132 30438 30144
rect 31113 30141 31125 30144
rect 31159 30172 31171 30175
rect 31159 30144 31754 30172
rect 31159 30141 31171 30144
rect 31113 30135 31171 30141
rect 26804 30076 27108 30104
rect 29454 30064 29460 30116
rect 29512 30104 29518 30116
rect 29733 30107 29791 30113
rect 29733 30104 29745 30107
rect 29512 30076 29745 30104
rect 29512 30064 29518 30076
rect 29733 30073 29745 30076
rect 29779 30104 29791 30107
rect 29779 30076 30788 30104
rect 29779 30073 29791 30076
rect 29733 30067 29791 30073
rect 22646 30036 22652 30048
rect 21468 30008 22652 30036
rect 20625 29999 20683 30005
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 22738 29996 22744 30048
rect 22796 29996 22802 30048
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 23845 30039 23903 30045
rect 23845 30036 23857 30039
rect 23808 30008 23857 30036
rect 23808 29996 23814 30008
rect 23845 30005 23857 30008
rect 23891 30005 23903 30039
rect 23845 29999 23903 30005
rect 26697 30039 26755 30045
rect 26697 30005 26709 30039
rect 26743 30036 26755 30039
rect 27062 30036 27068 30048
rect 26743 30008 27068 30036
rect 26743 30005 26755 30008
rect 26697 29999 26755 30005
rect 27062 29996 27068 30008
rect 27120 29996 27126 30048
rect 27706 29996 27712 30048
rect 27764 30036 27770 30048
rect 28721 30039 28779 30045
rect 28721 30036 28733 30039
rect 27764 30008 28733 30036
rect 27764 29996 27770 30008
rect 28721 30005 28733 30008
rect 28767 30005 28779 30039
rect 28721 29999 28779 30005
rect 30282 29996 30288 30048
rect 30340 29996 30346 30048
rect 30760 30036 30788 30076
rect 30834 30064 30840 30116
rect 30892 30104 30898 30116
rect 31726 30104 31754 30144
rect 32214 30132 32220 30184
rect 32272 30132 32278 30184
rect 32493 30175 32551 30181
rect 32493 30141 32505 30175
rect 32539 30172 32551 30175
rect 33410 30172 33416 30184
rect 32539 30144 33416 30172
rect 32539 30141 32551 30144
rect 32493 30135 32551 30141
rect 33410 30132 33416 30144
rect 33468 30132 33474 30184
rect 34146 30132 34152 30184
rect 34204 30172 34210 30184
rect 34330 30172 34336 30184
rect 34204 30144 34336 30172
rect 34204 30132 34210 30144
rect 34330 30132 34336 30144
rect 34388 30172 34394 30184
rect 34388 30144 34744 30172
rect 34388 30132 34394 30144
rect 34238 30104 34244 30116
rect 30892 30076 31616 30104
rect 31726 30076 34244 30104
rect 30892 30064 30898 30076
rect 31018 30036 31024 30048
rect 30760 30008 31024 30036
rect 31018 29996 31024 30008
rect 31076 29996 31082 30048
rect 31389 30039 31447 30045
rect 31389 30005 31401 30039
rect 31435 30036 31447 30039
rect 31478 30036 31484 30048
rect 31435 30008 31484 30036
rect 31435 30005 31447 30008
rect 31389 29999 31447 30005
rect 31478 29996 31484 30008
rect 31536 29996 31542 30048
rect 31588 30036 31616 30076
rect 34238 30064 34244 30076
rect 34296 30064 34302 30116
rect 34422 30064 34428 30116
rect 34480 30064 34486 30116
rect 34716 30104 34744 30144
rect 34790 30132 34796 30184
rect 34848 30132 34854 30184
rect 34882 30132 34888 30184
rect 34940 30132 34946 30184
rect 34977 30175 35035 30181
rect 34977 30141 34989 30175
rect 35023 30141 35035 30175
rect 35268 30172 35296 30212
rect 35618 30200 35624 30212
rect 35676 30200 35682 30252
rect 35805 30243 35863 30249
rect 35805 30209 35817 30243
rect 35851 30209 35863 30243
rect 35805 30203 35863 30209
rect 35526 30172 35532 30184
rect 35268 30144 35532 30172
rect 34977 30135 35035 30141
rect 34992 30104 35020 30135
rect 35526 30132 35532 30144
rect 35584 30172 35590 30184
rect 35820 30172 35848 30203
rect 36354 30200 36360 30252
rect 36412 30249 36418 30252
rect 36412 30243 36461 30249
rect 36412 30209 36415 30243
rect 36449 30209 36461 30243
rect 36412 30203 36461 30209
rect 36412 30200 36418 30203
rect 36538 30200 36544 30252
rect 36596 30200 36602 30252
rect 36722 30200 36728 30252
rect 36780 30249 36786 30252
rect 36780 30243 36819 30249
rect 36807 30209 36819 30243
rect 36780 30203 36819 30209
rect 36920 30243 36978 30249
rect 36920 30209 36932 30243
rect 36966 30240 36978 30243
rect 36966 30212 37044 30240
rect 36966 30209 36978 30212
rect 36920 30203 36978 30209
rect 36780 30200 36786 30203
rect 35584 30144 35848 30172
rect 35584 30132 35590 30144
rect 34716 30076 35020 30104
rect 31849 30039 31907 30045
rect 31849 30036 31861 30039
rect 31588 30008 31861 30036
rect 31849 30005 31861 30008
rect 31895 30005 31907 30039
rect 31849 29999 31907 30005
rect 33870 29996 33876 30048
rect 33928 29996 33934 30048
rect 34057 30039 34115 30045
rect 34057 30005 34069 30039
rect 34103 30036 34115 30039
rect 34517 30039 34575 30045
rect 34517 30036 34529 30039
rect 34103 30008 34529 30036
rect 34103 30005 34115 30008
rect 34057 29999 34115 30005
rect 34517 30005 34529 30008
rect 34563 30005 34575 30039
rect 34992 30036 35020 30076
rect 35158 30064 35164 30116
rect 35216 30064 35222 30116
rect 35820 30104 35848 30144
rect 35894 30132 35900 30184
rect 35952 30172 35958 30184
rect 35989 30175 36047 30181
rect 35989 30172 36001 30175
rect 35952 30144 36001 30172
rect 35952 30132 35958 30144
rect 35989 30141 36001 30144
rect 36035 30172 36047 30175
rect 36078 30172 36084 30184
rect 36035 30144 36084 30172
rect 36035 30141 36047 30144
rect 35989 30135 36047 30141
rect 36078 30132 36084 30144
rect 36136 30132 36142 30184
rect 36170 30132 36176 30184
rect 36228 30172 36234 30184
rect 37016 30172 37044 30212
rect 38102 30200 38108 30252
rect 38160 30200 38166 30252
rect 38381 30243 38439 30249
rect 38381 30209 38393 30243
rect 38427 30209 38439 30243
rect 38381 30203 38439 30209
rect 36228 30144 37044 30172
rect 36228 30132 36234 30144
rect 37826 30132 37832 30184
rect 37884 30172 37890 30184
rect 38396 30172 38424 30203
rect 38562 30200 38568 30252
rect 38620 30240 38626 30252
rect 39025 30243 39083 30249
rect 39025 30240 39037 30243
rect 38620 30212 39037 30240
rect 38620 30200 38626 30212
rect 39025 30209 39037 30212
rect 39071 30209 39083 30243
rect 39025 30203 39083 30209
rect 39206 30200 39212 30252
rect 39264 30200 39270 30252
rect 39301 30243 39359 30249
rect 39301 30209 39313 30243
rect 39347 30209 39359 30243
rect 39301 30203 39359 30209
rect 39393 30243 39451 30249
rect 39393 30209 39405 30243
rect 39439 30240 39451 30243
rect 39666 30240 39672 30252
rect 39439 30212 39672 30240
rect 39439 30209 39451 30212
rect 39393 30203 39451 30209
rect 37884 30144 38424 30172
rect 37884 30132 37890 30144
rect 37277 30107 37335 30113
rect 37277 30104 37289 30107
rect 35820 30076 37289 30104
rect 37277 30073 37289 30076
rect 37323 30073 37335 30107
rect 37277 30067 37335 30073
rect 38378 30064 38384 30116
rect 38436 30104 38442 30116
rect 39316 30104 39344 30203
rect 39666 30200 39672 30212
rect 39724 30200 39730 30252
rect 40218 30200 40224 30252
rect 40276 30240 40282 30252
rect 40405 30243 40463 30249
rect 40405 30240 40417 30243
rect 40276 30212 40417 30240
rect 40276 30200 40282 30212
rect 40405 30209 40417 30212
rect 40451 30209 40463 30243
rect 40405 30203 40463 30209
rect 40494 30200 40500 30252
rect 40552 30200 40558 30252
rect 40788 30249 40816 30280
rect 40773 30243 40831 30249
rect 40773 30209 40785 30243
rect 40819 30209 40831 30243
rect 40773 30203 40831 30209
rect 40862 30200 40868 30252
rect 40920 30200 40926 30252
rect 41049 30243 41107 30249
rect 41049 30209 41061 30243
rect 41095 30209 41107 30243
rect 41386 30240 41414 30280
rect 41874 30240 41880 30252
rect 41386 30212 41880 30240
rect 41049 30203 41107 30209
rect 41064 30172 41092 30203
rect 41874 30200 41880 30212
rect 41932 30200 41938 30252
rect 40236 30144 41092 30172
rect 38436 30076 39344 30104
rect 39577 30107 39635 30113
rect 38436 30064 38442 30076
rect 39577 30073 39589 30107
rect 39623 30104 39635 30107
rect 40034 30104 40040 30116
rect 39623 30076 40040 30104
rect 39623 30073 39635 30076
rect 39577 30067 39635 30073
rect 40034 30064 40040 30076
rect 40092 30064 40098 30116
rect 40236 30113 40264 30144
rect 40221 30107 40279 30113
rect 40221 30073 40233 30107
rect 40267 30073 40279 30107
rect 40221 30067 40279 30073
rect 35345 30039 35403 30045
rect 35345 30036 35357 30039
rect 34992 30008 35357 30036
rect 34517 29999 34575 30005
rect 35345 30005 35357 30008
rect 35391 30005 35403 30039
rect 35345 29999 35403 30005
rect 37645 30039 37703 30045
rect 37645 30005 37657 30039
rect 37691 30036 37703 30039
rect 37921 30039 37979 30045
rect 37921 30036 37933 30039
rect 37691 30008 37933 30036
rect 37691 30005 37703 30008
rect 37645 29999 37703 30005
rect 37921 30005 37933 30008
rect 37967 30005 37979 30039
rect 37921 29999 37979 30005
rect 40678 29996 40684 30048
rect 40736 30036 40742 30048
rect 41233 30039 41291 30045
rect 41233 30036 41245 30039
rect 40736 30008 41245 30036
rect 40736 29996 40742 30008
rect 41233 30005 41245 30008
rect 41279 30005 41291 30039
rect 41233 29999 41291 30005
rect 42058 29996 42064 30048
rect 42116 29996 42122 30048
rect 1104 29946 42504 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 42504 29946
rect 1104 29872 42504 29894
rect 3418 29792 3424 29844
rect 3476 29832 3482 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 3476 29804 3801 29832
rect 3476 29792 3482 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 3789 29795 3847 29801
rect 5534 29792 5540 29844
rect 5592 29792 5598 29844
rect 5721 29835 5779 29841
rect 5721 29801 5733 29835
rect 5767 29832 5779 29835
rect 7834 29832 7840 29844
rect 5767 29804 7840 29832
rect 5767 29801 5779 29804
rect 5721 29795 5779 29801
rect 7834 29792 7840 29804
rect 7892 29792 7898 29844
rect 17402 29792 17408 29844
rect 17460 29832 17466 29844
rect 17678 29832 17684 29844
rect 17460 29804 17684 29832
rect 17460 29792 17466 29804
rect 17678 29792 17684 29804
rect 17736 29792 17742 29844
rect 20254 29792 20260 29844
rect 20312 29832 20318 29844
rect 22189 29835 22247 29841
rect 20312 29804 22140 29832
rect 20312 29792 20318 29804
rect 3510 29764 3516 29776
rect 3160 29736 3516 29764
rect 1762 29588 1768 29640
rect 1820 29628 1826 29640
rect 2682 29628 2688 29640
rect 1820 29600 2688 29628
rect 1820 29588 1826 29600
rect 2682 29588 2688 29600
rect 2740 29588 2746 29640
rect 2866 29588 2872 29640
rect 2924 29588 2930 29640
rect 3160 29637 3188 29736
rect 3510 29724 3516 29736
rect 3568 29764 3574 29776
rect 3970 29764 3976 29776
rect 3568 29736 3976 29764
rect 3568 29724 3574 29736
rect 3970 29724 3976 29736
rect 4028 29724 4034 29776
rect 22002 29764 22008 29776
rect 21652 29736 22008 29764
rect 3786 29696 3792 29708
rect 3344 29668 3792 29696
rect 3140 29631 3198 29637
rect 3140 29597 3152 29631
rect 3186 29597 3198 29631
rect 3140 29591 3198 29597
rect 3234 29588 3240 29640
rect 3292 29588 3298 29640
rect 3344 29637 3372 29668
rect 3786 29656 3792 29668
rect 3844 29656 3850 29708
rect 4249 29699 4307 29705
rect 4249 29665 4261 29699
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 3329 29631 3387 29637
rect 3329 29597 3341 29631
rect 3375 29597 3387 29631
rect 3457 29631 3515 29637
rect 3457 29628 3469 29631
rect 3329 29591 3387 29597
rect 3436 29597 3469 29628
rect 3503 29597 3515 29631
rect 3436 29591 3515 29597
rect 2777 29563 2835 29569
rect 2777 29529 2789 29563
rect 2823 29560 2835 29563
rect 3436 29560 3464 29591
rect 3602 29588 3608 29640
rect 3660 29588 3666 29640
rect 3970 29588 3976 29640
rect 4028 29588 4034 29640
rect 4062 29588 4068 29640
rect 4120 29588 4126 29640
rect 4264 29572 4292 29659
rect 5074 29656 5080 29708
rect 5132 29696 5138 29708
rect 5445 29699 5503 29705
rect 5445 29696 5457 29699
rect 5132 29668 5457 29696
rect 5132 29656 5138 29668
rect 5445 29665 5457 29668
rect 5491 29665 5503 29699
rect 5445 29659 5503 29665
rect 8665 29699 8723 29705
rect 8665 29665 8677 29699
rect 8711 29696 8723 29699
rect 9582 29696 9588 29708
rect 8711 29668 9588 29696
rect 8711 29665 8723 29668
rect 8665 29659 8723 29665
rect 9582 29656 9588 29668
rect 9640 29656 9646 29708
rect 12894 29656 12900 29708
rect 12952 29696 12958 29708
rect 13081 29699 13139 29705
rect 13081 29696 13093 29699
rect 12952 29668 13093 29696
rect 12952 29656 12958 29668
rect 13081 29665 13093 29668
rect 13127 29696 13139 29699
rect 13170 29696 13176 29708
rect 13127 29668 13176 29696
rect 13127 29665 13139 29668
rect 13081 29659 13139 29665
rect 13170 29656 13176 29668
rect 13228 29656 13234 29708
rect 17770 29656 17776 29708
rect 17828 29696 17834 29708
rect 21174 29696 21180 29708
rect 17828 29668 21180 29696
rect 17828 29656 17834 29668
rect 21174 29656 21180 29668
rect 21232 29656 21238 29708
rect 4338 29588 4344 29640
rect 4396 29588 4402 29640
rect 5350 29588 5356 29640
rect 5408 29588 5414 29640
rect 9306 29588 9312 29640
rect 9364 29588 9370 29640
rect 10226 29588 10232 29640
rect 10284 29628 10290 29640
rect 10321 29631 10379 29637
rect 10321 29628 10333 29631
rect 10284 29600 10333 29628
rect 10284 29588 10290 29600
rect 10321 29597 10333 29600
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 10689 29631 10747 29637
rect 10689 29597 10701 29631
rect 10735 29628 10747 29631
rect 11054 29628 11060 29640
rect 10735 29600 11060 29628
rect 10735 29597 10747 29600
rect 10689 29591 10747 29597
rect 11054 29588 11060 29600
rect 11112 29588 11118 29640
rect 20349 29631 20407 29637
rect 20349 29597 20361 29631
rect 20395 29597 20407 29631
rect 20349 29591 20407 29597
rect 4246 29560 4252 29572
rect 2823 29532 3188 29560
rect 2823 29529 2835 29532
rect 2777 29523 2835 29529
rect 2958 29452 2964 29504
rect 3016 29452 3022 29504
rect 3160 29492 3188 29532
rect 3436 29532 4252 29560
rect 3436 29492 3464 29532
rect 4246 29520 4252 29532
rect 4304 29520 4310 29572
rect 8389 29563 8447 29569
rect 8389 29529 8401 29563
rect 8435 29560 8447 29563
rect 8662 29560 8668 29572
rect 8435 29532 8668 29560
rect 8435 29529 8447 29532
rect 8389 29523 8447 29529
rect 8662 29520 8668 29532
rect 8720 29520 8726 29572
rect 12710 29520 12716 29572
rect 12768 29520 12774 29572
rect 12897 29563 12955 29569
rect 12897 29529 12909 29563
rect 12943 29529 12955 29563
rect 20364 29560 20392 29591
rect 20622 29588 20628 29640
rect 20680 29628 20686 29640
rect 21652 29637 21680 29736
rect 22002 29724 22008 29736
rect 22060 29724 22066 29776
rect 22112 29764 22140 29804
rect 22189 29801 22201 29835
rect 22235 29832 22247 29835
rect 22738 29832 22744 29844
rect 22235 29804 22744 29832
rect 22235 29801 22247 29804
rect 22189 29795 22247 29801
rect 22738 29792 22744 29804
rect 22796 29792 22802 29844
rect 24673 29835 24731 29841
rect 24673 29801 24685 29835
rect 24719 29832 24731 29835
rect 24854 29832 24860 29844
rect 24719 29804 24860 29832
rect 24719 29801 24731 29804
rect 24673 29795 24731 29801
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 26878 29792 26884 29844
rect 26936 29792 26942 29844
rect 27341 29835 27399 29841
rect 27341 29801 27353 29835
rect 27387 29832 27399 29835
rect 28902 29832 28908 29844
rect 27387 29804 28908 29832
rect 27387 29801 27399 29804
rect 27341 29795 27399 29801
rect 28902 29792 28908 29804
rect 28960 29792 28966 29844
rect 30742 29792 30748 29844
rect 30800 29792 30806 29844
rect 31662 29792 31668 29844
rect 31720 29832 31726 29844
rect 33045 29835 33103 29841
rect 33045 29832 33057 29835
rect 31720 29804 33057 29832
rect 31720 29792 31726 29804
rect 33045 29801 33057 29804
rect 33091 29801 33103 29835
rect 33045 29795 33103 29801
rect 34606 29792 34612 29844
rect 34664 29832 34670 29844
rect 34793 29835 34851 29841
rect 34793 29832 34805 29835
rect 34664 29804 34805 29832
rect 34664 29792 34670 29804
rect 34793 29801 34805 29804
rect 34839 29801 34851 29835
rect 34793 29795 34851 29801
rect 34974 29792 34980 29844
rect 35032 29832 35038 29844
rect 35032 29804 35480 29832
rect 35032 29792 35038 29804
rect 22830 29764 22836 29776
rect 22112 29736 22836 29764
rect 22830 29724 22836 29736
rect 22888 29764 22894 29776
rect 25958 29764 25964 29776
rect 22888 29736 25084 29764
rect 22888 29724 22894 29736
rect 21818 29656 21824 29708
rect 21876 29696 21882 29708
rect 21876 29668 22048 29696
rect 21876 29656 21882 29668
rect 21637 29631 21695 29637
rect 21637 29628 21649 29631
rect 20680 29600 21649 29628
rect 20680 29588 20686 29600
rect 21637 29597 21649 29600
rect 21683 29597 21695 29631
rect 21637 29591 21695 29597
rect 21726 29588 21732 29640
rect 21784 29588 21790 29640
rect 21910 29588 21916 29640
rect 21968 29588 21974 29640
rect 22020 29637 22048 29668
rect 23014 29656 23020 29708
rect 23072 29696 23078 29708
rect 23072 29668 23152 29696
rect 23072 29656 23078 29668
rect 22005 29631 22063 29637
rect 22005 29597 22017 29631
rect 22051 29597 22063 29631
rect 22005 29591 22063 29597
rect 22738 29588 22744 29640
rect 22796 29588 22802 29640
rect 23124 29637 23152 29668
rect 22834 29631 22892 29637
rect 22834 29597 22846 29631
rect 22880 29597 22892 29631
rect 22834 29591 22892 29597
rect 23109 29631 23167 29637
rect 23109 29597 23121 29631
rect 23155 29597 23167 29631
rect 23109 29591 23167 29597
rect 20364 29532 20668 29560
rect 12897 29523 12955 29529
rect 3160 29464 3464 29492
rect 3602 29452 3608 29504
rect 3660 29492 3666 29504
rect 4062 29492 4068 29504
rect 3660 29464 4068 29492
rect 3660 29452 3666 29464
rect 4062 29452 4068 29464
rect 4120 29452 4126 29504
rect 8018 29452 8024 29504
rect 8076 29452 8082 29504
rect 8478 29452 8484 29504
rect 8536 29452 8542 29504
rect 8938 29452 8944 29504
rect 8996 29452 9002 29504
rect 9398 29452 9404 29504
rect 9456 29452 9462 29504
rect 9766 29452 9772 29504
rect 9824 29452 9830 29504
rect 10042 29452 10048 29504
rect 10100 29492 10106 29504
rect 10597 29495 10655 29501
rect 10597 29492 10609 29495
rect 10100 29464 10609 29492
rect 10100 29452 10106 29464
rect 10597 29461 10609 29464
rect 10643 29461 10655 29495
rect 10597 29455 10655 29461
rect 12434 29452 12440 29504
rect 12492 29492 12498 29504
rect 12912 29492 12940 29523
rect 12492 29464 12940 29492
rect 12492 29452 12498 29464
rect 18046 29452 18052 29504
rect 18104 29492 18110 29504
rect 20530 29492 20536 29504
rect 18104 29464 20536 29492
rect 18104 29452 18110 29464
rect 20530 29452 20536 29464
rect 20588 29452 20594 29504
rect 20640 29492 20668 29532
rect 20806 29520 20812 29572
rect 20864 29520 20870 29572
rect 20990 29520 20996 29572
rect 21048 29560 21054 29572
rect 21542 29560 21548 29572
rect 21048 29532 21548 29560
rect 21048 29520 21054 29532
rect 21542 29520 21548 29532
rect 21600 29520 21606 29572
rect 22278 29520 22284 29572
rect 22336 29560 22342 29572
rect 22848 29560 22876 29591
rect 23198 29588 23204 29640
rect 23256 29637 23262 29640
rect 23256 29631 23305 29637
rect 23256 29597 23259 29631
rect 23293 29628 23305 29631
rect 23382 29628 23388 29640
rect 23293 29600 23388 29628
rect 23293 29597 23305 29600
rect 23256 29591 23305 29597
rect 23256 29588 23262 29591
rect 23382 29588 23388 29600
rect 23440 29588 23446 29640
rect 24854 29588 24860 29640
rect 24912 29588 24918 29640
rect 22336 29532 22876 29560
rect 23017 29563 23075 29569
rect 22336 29520 22342 29532
rect 23017 29529 23029 29563
rect 23063 29560 23075 29563
rect 24118 29560 24124 29572
rect 23063 29532 24124 29560
rect 23063 29529 23075 29532
rect 23017 29523 23075 29529
rect 24118 29520 24124 29532
rect 24176 29560 24182 29572
rect 24670 29560 24676 29572
rect 24176 29532 24676 29560
rect 24176 29520 24182 29532
rect 24670 29520 24676 29532
rect 24728 29520 24734 29572
rect 25056 29569 25084 29736
rect 25424 29736 25964 29764
rect 25424 29705 25452 29736
rect 25958 29724 25964 29736
rect 26016 29724 26022 29776
rect 27798 29724 27804 29776
rect 27856 29764 27862 29776
rect 27982 29764 27988 29776
rect 27856 29736 27988 29764
rect 27856 29724 27862 29736
rect 27982 29724 27988 29736
rect 28040 29724 28046 29776
rect 29454 29764 29460 29776
rect 28184 29736 29460 29764
rect 25409 29699 25467 29705
rect 25409 29665 25421 29699
rect 25455 29665 25467 29699
rect 25774 29696 25780 29708
rect 25409 29659 25467 29665
rect 25516 29668 25780 29696
rect 25133 29631 25191 29637
rect 25133 29597 25145 29631
rect 25179 29628 25191 29631
rect 25424 29628 25452 29659
rect 25516 29637 25544 29668
rect 25774 29656 25780 29668
rect 25832 29696 25838 29708
rect 26053 29699 26111 29705
rect 26053 29696 26065 29699
rect 25832 29668 26065 29696
rect 25832 29656 25838 29668
rect 26053 29665 26065 29668
rect 26099 29665 26111 29699
rect 26053 29659 26111 29665
rect 26602 29656 26608 29708
rect 26660 29696 26666 29708
rect 28184 29705 28212 29736
rect 29454 29724 29460 29736
rect 29512 29724 29518 29776
rect 30760 29764 30788 29792
rect 30484 29736 30788 29764
rect 28169 29699 28227 29705
rect 26660 29668 28120 29696
rect 26660 29656 26666 29668
rect 25179 29600 25452 29628
rect 25501 29631 25559 29637
rect 25179 29597 25191 29600
rect 25133 29591 25191 29597
rect 25501 29597 25513 29631
rect 25547 29597 25559 29631
rect 25501 29591 25559 29597
rect 25590 29588 25596 29640
rect 25648 29628 25654 29640
rect 25961 29631 26019 29637
rect 25961 29628 25973 29631
rect 25648 29600 25973 29628
rect 25648 29588 25654 29600
rect 25961 29597 25973 29600
rect 26007 29597 26019 29631
rect 25961 29591 26019 29597
rect 27062 29588 27068 29640
rect 27120 29588 27126 29640
rect 27154 29588 27160 29640
rect 27212 29588 27218 29640
rect 27433 29631 27491 29637
rect 27433 29628 27445 29631
rect 27255 29600 27445 29628
rect 25041 29563 25099 29569
rect 25041 29529 25053 29563
rect 25087 29560 25099 29563
rect 25087 29532 26188 29560
rect 25087 29529 25099 29532
rect 25041 29523 25099 29529
rect 21008 29492 21036 29520
rect 20640 29464 21036 29492
rect 21174 29452 21180 29504
rect 21232 29492 21238 29504
rect 23198 29492 23204 29504
rect 21232 29464 23204 29492
rect 21232 29452 21238 29464
rect 23198 29452 23204 29464
rect 23256 29452 23262 29504
rect 23385 29495 23443 29501
rect 23385 29461 23397 29495
rect 23431 29492 23443 29495
rect 24394 29492 24400 29504
rect 23431 29464 24400 29492
rect 23431 29461 23443 29464
rect 23385 29455 23443 29461
rect 24394 29452 24400 29464
rect 24452 29452 24458 29504
rect 25774 29452 25780 29504
rect 25832 29492 25838 29504
rect 25869 29495 25927 29501
rect 25869 29492 25881 29495
rect 25832 29464 25881 29492
rect 25832 29452 25838 29464
rect 25869 29461 25881 29464
rect 25915 29461 25927 29495
rect 26160 29492 26188 29532
rect 26234 29520 26240 29572
rect 26292 29560 26298 29572
rect 27255 29560 27283 29600
rect 27433 29597 27445 29600
rect 27479 29628 27491 29631
rect 27706 29628 27712 29640
rect 27479 29600 27712 29628
rect 27479 29597 27491 29600
rect 27433 29591 27491 29597
rect 27706 29588 27712 29600
rect 27764 29628 27770 29640
rect 27985 29631 28043 29637
rect 27985 29628 27997 29631
rect 27764 29600 27997 29628
rect 27764 29588 27770 29600
rect 27985 29597 27997 29600
rect 28031 29597 28043 29631
rect 28092 29628 28120 29668
rect 28169 29665 28181 29699
rect 28215 29665 28227 29699
rect 28169 29659 28227 29665
rect 28994 29656 29000 29708
rect 29052 29696 29058 29708
rect 29089 29699 29147 29705
rect 29089 29696 29101 29699
rect 29052 29668 29101 29696
rect 29052 29656 29058 29668
rect 29089 29665 29101 29668
rect 29135 29665 29147 29699
rect 29089 29659 29147 29665
rect 29638 29656 29644 29708
rect 29696 29696 29702 29708
rect 30377 29699 30435 29705
rect 30377 29696 30389 29699
rect 29696 29668 30389 29696
rect 29696 29656 29702 29668
rect 30377 29665 30389 29668
rect 30423 29665 30435 29699
rect 30377 29659 30435 29665
rect 29273 29631 29331 29637
rect 29273 29628 29285 29631
rect 28092 29600 29285 29628
rect 27985 29591 28043 29597
rect 29273 29597 29285 29600
rect 29319 29597 29331 29631
rect 29273 29591 29331 29597
rect 28994 29560 29000 29572
rect 26292 29532 27283 29560
rect 27356 29532 29000 29560
rect 26292 29520 26298 29532
rect 27356 29492 27384 29532
rect 28994 29520 29000 29532
rect 29052 29520 29058 29572
rect 29288 29560 29316 29591
rect 29362 29588 29368 29640
rect 29420 29588 29426 29640
rect 29822 29588 29828 29640
rect 29880 29588 29886 29640
rect 30009 29631 30067 29637
rect 30009 29597 30021 29631
rect 30055 29628 30067 29631
rect 30190 29628 30196 29640
rect 30055 29600 30196 29628
rect 30055 29597 30067 29600
rect 30009 29591 30067 29597
rect 30190 29588 30196 29600
rect 30248 29588 30254 29640
rect 30282 29588 30288 29640
rect 30340 29628 30346 29640
rect 30484 29628 30512 29736
rect 32490 29724 32496 29776
rect 32548 29764 32554 29776
rect 32953 29767 33011 29773
rect 32953 29764 32965 29767
rect 32548 29736 32965 29764
rect 32548 29724 32554 29736
rect 32953 29733 32965 29736
rect 32999 29733 33011 29767
rect 35342 29764 35348 29776
rect 32953 29727 33011 29733
rect 33152 29736 35348 29764
rect 30929 29699 30987 29705
rect 30929 29696 30941 29699
rect 30576 29668 30941 29696
rect 30576 29637 30604 29668
rect 30929 29665 30941 29668
rect 30975 29665 30987 29699
rect 30929 29659 30987 29665
rect 31478 29656 31484 29708
rect 31536 29656 31542 29708
rect 30340 29600 30512 29628
rect 30561 29631 30619 29637
rect 30340 29588 30346 29600
rect 30561 29597 30573 29631
rect 30607 29597 30619 29631
rect 30561 29591 30619 29597
rect 30650 29588 30656 29640
rect 30708 29628 30714 29640
rect 30837 29631 30895 29637
rect 30837 29628 30849 29631
rect 30708 29600 30849 29628
rect 30708 29588 30714 29600
rect 30837 29597 30849 29600
rect 30883 29597 30895 29631
rect 30837 29591 30895 29597
rect 31021 29631 31079 29637
rect 31021 29597 31033 29631
rect 31067 29597 31079 29631
rect 31021 29591 31079 29597
rect 29840 29560 29868 29588
rect 31036 29560 31064 29591
rect 31110 29588 31116 29640
rect 31168 29628 31174 29640
rect 31205 29631 31263 29637
rect 31205 29628 31217 29631
rect 31168 29600 31217 29628
rect 31168 29588 31174 29600
rect 31205 29597 31217 29600
rect 31251 29597 31263 29631
rect 31205 29591 31263 29597
rect 33152 29622 33180 29736
rect 35342 29724 35348 29736
rect 35400 29724 35406 29776
rect 35452 29764 35480 29804
rect 35526 29792 35532 29844
rect 35584 29832 35590 29844
rect 37185 29835 37243 29841
rect 37185 29832 37197 29835
rect 35584 29804 37197 29832
rect 35584 29792 35590 29804
rect 37185 29801 37197 29804
rect 37231 29801 37243 29835
rect 37185 29795 37243 29801
rect 37274 29792 37280 29844
rect 37332 29832 37338 29844
rect 37369 29835 37427 29841
rect 37369 29832 37381 29835
rect 37332 29804 37381 29832
rect 37332 29792 37338 29804
rect 37369 29801 37381 29804
rect 37415 29832 37427 29835
rect 38102 29832 38108 29844
rect 37415 29804 38108 29832
rect 37415 29801 37427 29804
rect 37369 29795 37427 29801
rect 38102 29792 38108 29804
rect 38160 29792 38166 29844
rect 38286 29792 38292 29844
rect 38344 29832 38350 29844
rect 40402 29832 40408 29844
rect 38344 29804 40408 29832
rect 38344 29792 38350 29804
rect 40402 29792 40408 29804
rect 40460 29792 40466 29844
rect 41874 29792 41880 29844
rect 41932 29832 41938 29844
rect 42153 29835 42211 29841
rect 42153 29832 42165 29835
rect 41932 29804 42165 29832
rect 41932 29792 41938 29804
rect 42153 29801 42165 29804
rect 42199 29801 42211 29835
rect 42153 29795 42211 29801
rect 35452 29736 36216 29764
rect 33410 29656 33416 29708
rect 33468 29696 33474 29708
rect 33468 29668 33732 29696
rect 33468 29656 33474 29668
rect 33224 29631 33282 29637
rect 33224 29622 33236 29631
rect 33152 29597 33236 29622
rect 33270 29597 33282 29631
rect 33594 29628 33600 29640
rect 33555 29600 33600 29628
rect 33152 29594 33282 29597
rect 33224 29591 33282 29594
rect 33594 29588 33600 29600
rect 33652 29588 33658 29640
rect 33704 29637 33732 29668
rect 34882 29656 34888 29708
rect 34940 29696 34946 29708
rect 35437 29699 35495 29705
rect 34940 29668 35204 29696
rect 34940 29656 34946 29668
rect 33689 29631 33747 29637
rect 33689 29597 33701 29631
rect 33735 29628 33747 29631
rect 34698 29628 34704 29640
rect 33735 29600 34704 29628
rect 33735 29597 33747 29600
rect 33689 29591 33747 29597
rect 34698 29588 34704 29600
rect 34756 29588 34762 29640
rect 35066 29588 35072 29640
rect 35124 29588 35130 29640
rect 35176 29628 35204 29668
rect 35437 29665 35449 29699
rect 35483 29696 35495 29699
rect 35526 29696 35532 29708
rect 35483 29668 35532 29696
rect 35483 29665 35495 29668
rect 35437 29659 35495 29665
rect 35526 29656 35532 29668
rect 35584 29656 35590 29708
rect 35636 29705 35664 29736
rect 35621 29699 35679 29705
rect 35621 29665 35633 29699
rect 35667 29665 35679 29699
rect 35621 29659 35679 29665
rect 35897 29699 35955 29705
rect 35897 29665 35909 29699
rect 35943 29665 35955 29699
rect 35897 29659 35955 29665
rect 35345 29631 35403 29637
rect 35345 29628 35357 29631
rect 35176 29600 35357 29628
rect 35345 29597 35357 29600
rect 35391 29628 35403 29631
rect 35802 29628 35808 29640
rect 35391 29600 35808 29628
rect 35391 29597 35403 29600
rect 35345 29591 35403 29597
rect 35802 29588 35808 29600
rect 35860 29588 35866 29640
rect 35912 29628 35940 29659
rect 35986 29656 35992 29708
rect 36044 29696 36050 29708
rect 36081 29699 36139 29705
rect 36081 29696 36093 29699
rect 36044 29668 36093 29696
rect 36044 29656 36050 29668
rect 36081 29665 36093 29668
rect 36127 29665 36139 29699
rect 36188 29696 36216 29736
rect 36538 29724 36544 29776
rect 36596 29764 36602 29776
rect 37090 29764 37096 29776
rect 36596 29736 37096 29764
rect 36596 29724 36602 29736
rect 37090 29724 37096 29736
rect 37148 29764 37154 29776
rect 37148 29736 38516 29764
rect 37148 29724 37154 29736
rect 37642 29696 37648 29708
rect 36188 29668 37648 29696
rect 36081 29659 36139 29665
rect 37642 29656 37648 29668
rect 37700 29656 37706 29708
rect 37752 29668 38240 29696
rect 36173 29631 36231 29637
rect 35912 29600 36124 29628
rect 33042 29560 33048 29572
rect 29288 29532 29868 29560
rect 30484 29532 31064 29560
rect 32706 29532 33048 29560
rect 26160 29464 27384 29492
rect 27525 29495 27583 29501
rect 25869 29455 25927 29461
rect 27525 29461 27537 29495
rect 27571 29492 27583 29495
rect 27706 29492 27712 29504
rect 27571 29464 27712 29492
rect 27571 29461 27583 29464
rect 27525 29455 27583 29461
rect 27706 29452 27712 29464
rect 27764 29452 27770 29504
rect 27890 29452 27896 29504
rect 27948 29452 27954 29504
rect 29089 29495 29147 29501
rect 29089 29461 29101 29495
rect 29135 29492 29147 29495
rect 29454 29492 29460 29504
rect 29135 29464 29460 29492
rect 29135 29461 29147 29464
rect 29089 29455 29147 29461
rect 29454 29452 29460 29464
rect 29512 29452 29518 29504
rect 29730 29452 29736 29504
rect 29788 29492 29794 29504
rect 30484 29492 30512 29532
rect 33042 29520 33048 29532
rect 33100 29520 33106 29572
rect 33321 29563 33379 29569
rect 33321 29560 33333 29563
rect 33152 29532 33333 29560
rect 29788 29464 30512 29492
rect 29788 29452 29794 29464
rect 30558 29452 30564 29504
rect 30616 29492 30622 29504
rect 30745 29495 30803 29501
rect 30745 29492 30757 29495
rect 30616 29464 30757 29492
rect 30616 29452 30622 29464
rect 30745 29461 30757 29464
rect 30791 29461 30803 29495
rect 30745 29455 30803 29461
rect 31018 29452 31024 29504
rect 31076 29492 31082 29504
rect 31754 29492 31760 29504
rect 31076 29464 31760 29492
rect 31076 29452 31082 29464
rect 31754 29452 31760 29464
rect 31812 29452 31818 29504
rect 32950 29452 32956 29504
rect 33008 29492 33014 29504
rect 33152 29492 33180 29532
rect 33321 29529 33333 29532
rect 33367 29529 33379 29563
rect 33321 29523 33379 29529
rect 33413 29563 33471 29569
rect 33413 29529 33425 29563
rect 33459 29560 33471 29563
rect 34146 29560 34152 29572
rect 33459 29532 34152 29560
rect 33459 29529 33471 29532
rect 33413 29523 33471 29529
rect 34146 29520 34152 29532
rect 34204 29520 34210 29572
rect 34793 29563 34851 29569
rect 34793 29529 34805 29563
rect 34839 29560 34851 29563
rect 34882 29560 34888 29572
rect 34839 29532 34888 29560
rect 34839 29529 34851 29532
rect 34793 29523 34851 29529
rect 34882 29520 34888 29532
rect 34940 29520 34946 29572
rect 34977 29563 35035 29569
rect 34977 29529 34989 29563
rect 35023 29560 35035 29563
rect 35986 29560 35992 29572
rect 35023 29532 35992 29560
rect 35023 29529 35035 29532
rect 34977 29523 35035 29529
rect 35986 29520 35992 29532
rect 36044 29520 36050 29572
rect 36096 29560 36124 29600
rect 36173 29597 36185 29631
rect 36219 29628 36231 29631
rect 36446 29628 36452 29640
rect 36219 29600 36452 29628
rect 36219 29597 36231 29600
rect 36173 29591 36231 29597
rect 36446 29588 36452 29600
rect 36504 29588 36510 29640
rect 37274 29628 37280 29640
rect 36556 29600 37280 29628
rect 36556 29560 36584 29600
rect 37274 29588 37280 29600
rect 37332 29588 37338 29640
rect 37752 29628 37780 29668
rect 38212 29640 38240 29668
rect 37476 29600 37780 29628
rect 37476 29560 37504 29600
rect 37826 29588 37832 29640
rect 37884 29588 37890 29640
rect 37921 29631 37979 29637
rect 37921 29597 37933 29631
rect 37967 29597 37979 29631
rect 37921 29591 37979 29597
rect 36096 29532 36584 29560
rect 37108 29532 37504 29560
rect 37553 29563 37611 29569
rect 33008 29464 33180 29492
rect 33008 29452 33014 29464
rect 33226 29452 33232 29504
rect 33284 29492 33290 29504
rect 33594 29492 33600 29504
rect 33284 29464 33600 29492
rect 33284 29452 33290 29464
rect 33594 29452 33600 29464
rect 33652 29452 33658 29504
rect 35434 29452 35440 29504
rect 35492 29492 35498 29504
rect 35621 29495 35679 29501
rect 35621 29492 35633 29495
rect 35492 29464 35633 29492
rect 35492 29452 35498 29464
rect 35621 29461 35633 29464
rect 35667 29461 35679 29495
rect 35621 29455 35679 29461
rect 36541 29495 36599 29501
rect 36541 29461 36553 29495
rect 36587 29492 36599 29495
rect 37108 29492 37136 29532
rect 37553 29529 37565 29563
rect 37599 29560 37611 29563
rect 37936 29560 37964 29591
rect 38194 29588 38200 29640
rect 38252 29588 38258 29640
rect 38378 29588 38384 29640
rect 38436 29588 38442 29640
rect 38488 29637 38516 29736
rect 38654 29656 38660 29708
rect 38712 29696 38718 29708
rect 39298 29696 39304 29708
rect 38712 29668 39304 29696
rect 38712 29656 38718 29668
rect 39298 29656 39304 29668
rect 39356 29656 39362 29708
rect 40678 29656 40684 29708
rect 40736 29656 40742 29708
rect 38473 29631 38531 29637
rect 38473 29597 38485 29631
rect 38519 29597 38531 29631
rect 38473 29591 38531 29597
rect 38565 29631 38623 29637
rect 38565 29597 38577 29631
rect 38611 29628 38623 29631
rect 40218 29628 40224 29640
rect 38611 29600 40224 29628
rect 38611 29597 38623 29600
rect 38565 29591 38623 29597
rect 40218 29588 40224 29600
rect 40276 29588 40282 29640
rect 40402 29588 40408 29640
rect 40460 29588 40466 29640
rect 38838 29560 38844 29572
rect 37599 29532 38844 29560
rect 37599 29529 37611 29532
rect 37553 29523 37611 29529
rect 38838 29520 38844 29532
rect 38896 29520 38902 29572
rect 39853 29563 39911 29569
rect 39853 29529 39865 29563
rect 39899 29529 39911 29563
rect 39853 29523 39911 29529
rect 36587 29464 37136 29492
rect 36587 29461 36599 29464
rect 36541 29455 36599 29461
rect 37182 29452 37188 29504
rect 37240 29492 37246 29504
rect 37343 29495 37401 29501
rect 37343 29492 37355 29495
rect 37240 29464 37355 29492
rect 37240 29452 37246 29464
rect 37343 29461 37355 29464
rect 37389 29461 37401 29495
rect 37343 29455 37401 29461
rect 37645 29495 37703 29501
rect 37645 29461 37657 29495
rect 37691 29492 37703 29495
rect 37918 29492 37924 29504
rect 37691 29464 37924 29492
rect 37691 29461 37703 29464
rect 37645 29455 37703 29461
rect 37918 29452 37924 29464
rect 37976 29452 37982 29504
rect 38749 29495 38807 29501
rect 38749 29461 38761 29495
rect 38795 29492 38807 29495
rect 39868 29492 39896 29523
rect 40034 29520 40040 29572
rect 40092 29520 40098 29572
rect 41414 29520 41420 29572
rect 41472 29520 41478 29572
rect 38795 29464 39896 29492
rect 38795 29461 38807 29464
rect 38749 29455 38807 29461
rect 40218 29452 40224 29504
rect 40276 29452 40282 29504
rect 1104 29402 42504 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 42504 29402
rect 1104 29328 42504 29350
rect 5166 29288 5172 29300
rect 1412 29260 5172 29288
rect 1412 29161 1440 29260
rect 5166 29248 5172 29260
rect 5224 29248 5230 29300
rect 5442 29248 5448 29300
rect 5500 29248 5506 29300
rect 8938 29288 8944 29300
rect 8036 29260 8944 29288
rect 3050 29220 3056 29232
rect 2898 29192 3056 29220
rect 3050 29180 3056 29192
rect 3108 29180 3114 29232
rect 3234 29180 3240 29232
rect 3292 29220 3298 29232
rect 7184 29223 7242 29229
rect 3292 29192 4108 29220
rect 3292 29180 3298 29192
rect 1397 29155 1455 29161
rect 1397 29121 1409 29155
rect 1443 29121 1455 29155
rect 1397 29115 1455 29121
rect 3421 29155 3479 29161
rect 3421 29121 3433 29155
rect 3467 29152 3479 29155
rect 3786 29152 3792 29164
rect 3467 29124 3792 29152
rect 3467 29121 3479 29124
rect 3421 29115 3479 29121
rect 3786 29112 3792 29124
rect 3844 29112 3850 29164
rect 4080 29161 4108 29192
rect 7184 29189 7196 29223
rect 7230 29220 7242 29223
rect 8036 29220 8064 29260
rect 8938 29248 8944 29260
rect 8996 29248 9002 29300
rect 9769 29291 9827 29297
rect 9769 29257 9781 29291
rect 9815 29288 9827 29291
rect 10226 29288 10232 29300
rect 9815 29260 10232 29288
rect 9815 29257 9827 29260
rect 9769 29251 9827 29257
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 10686 29248 10692 29300
rect 10744 29248 10750 29300
rect 10962 29248 10968 29300
rect 11020 29248 11026 29300
rect 12621 29291 12679 29297
rect 12621 29257 12633 29291
rect 12667 29288 12679 29291
rect 12986 29288 12992 29300
rect 12667 29260 12992 29288
rect 12667 29257 12679 29260
rect 12621 29251 12679 29257
rect 12986 29248 12992 29260
rect 13044 29248 13050 29300
rect 14274 29248 14280 29300
rect 14332 29248 14338 29300
rect 14826 29248 14832 29300
rect 14884 29288 14890 29300
rect 15013 29291 15071 29297
rect 15013 29288 15025 29291
rect 14884 29260 15025 29288
rect 14884 29248 14890 29260
rect 15013 29257 15025 29260
rect 15059 29257 15071 29291
rect 15013 29251 15071 29257
rect 15470 29248 15476 29300
rect 15528 29248 15534 29300
rect 16022 29248 16028 29300
rect 16080 29248 16086 29300
rect 16942 29248 16948 29300
rect 17000 29248 17006 29300
rect 17034 29248 17040 29300
rect 17092 29288 17098 29300
rect 18233 29291 18291 29297
rect 18233 29288 18245 29291
rect 17092 29260 18245 29288
rect 17092 29248 17098 29260
rect 18233 29257 18245 29260
rect 18279 29288 18291 29291
rect 18785 29291 18843 29297
rect 18279 29260 18644 29288
rect 18279 29257 18291 29260
rect 18233 29251 18291 29257
rect 10778 29220 10784 29232
rect 7230 29192 8064 29220
rect 8404 29192 10784 29220
rect 7230 29189 7242 29192
rect 7184 29183 7242 29189
rect 8404 29164 8432 29192
rect 10778 29180 10784 29192
rect 10836 29180 10842 29232
rect 12710 29220 12716 29232
rect 10888 29192 12716 29220
rect 4065 29155 4123 29161
rect 4065 29121 4077 29155
rect 4111 29121 4123 29155
rect 4065 29115 4123 29121
rect 4246 29112 4252 29164
rect 4304 29112 4310 29164
rect 5350 29112 5356 29164
rect 5408 29152 5414 29164
rect 5445 29155 5503 29161
rect 5445 29152 5457 29155
rect 5408 29124 5457 29152
rect 5408 29112 5414 29124
rect 5445 29121 5457 29124
rect 5491 29121 5503 29155
rect 5445 29115 5503 29121
rect 5629 29155 5687 29161
rect 5629 29121 5641 29155
rect 5675 29152 5687 29155
rect 5718 29152 5724 29164
rect 5675 29124 5724 29152
rect 5675 29121 5687 29124
rect 5629 29115 5687 29121
rect 5718 29112 5724 29124
rect 5776 29112 5782 29164
rect 6914 29112 6920 29164
rect 6972 29112 6978 29164
rect 8386 29112 8392 29164
rect 8444 29112 8450 29164
rect 8656 29155 8714 29161
rect 8656 29121 8668 29155
rect 8702 29152 8714 29155
rect 9122 29152 9128 29164
rect 8702 29124 9128 29152
rect 8702 29121 8714 29124
rect 8656 29115 8714 29121
rect 9122 29112 9128 29124
rect 9180 29112 9186 29164
rect 9861 29155 9919 29161
rect 9861 29121 9873 29155
rect 9907 29121 9919 29155
rect 9861 29115 9919 29121
rect 1670 29044 1676 29096
rect 1728 29044 1734 29096
rect 3145 29087 3203 29093
rect 3145 29053 3157 29087
rect 3191 29084 3203 29087
rect 3234 29084 3240 29096
rect 3191 29056 3240 29084
rect 3191 29053 3203 29056
rect 3145 29047 3203 29053
rect 3234 29044 3240 29056
rect 3292 29044 3298 29096
rect 3510 29044 3516 29096
rect 3568 29044 3574 29096
rect 3602 29044 3608 29096
rect 3660 29044 3666 29096
rect 3697 29087 3755 29093
rect 3697 29053 3709 29087
rect 3743 29084 3755 29087
rect 3881 29087 3939 29093
rect 3881 29084 3893 29087
rect 3743 29056 3893 29084
rect 3743 29053 3755 29056
rect 3697 29047 3755 29053
rect 3881 29053 3893 29056
rect 3927 29053 3939 29087
rect 3881 29047 3939 29053
rect 4338 29044 4344 29096
rect 4396 29084 4402 29096
rect 4798 29084 4804 29096
rect 4396 29056 4804 29084
rect 4396 29044 4402 29056
rect 4798 29044 4804 29056
rect 4856 29044 4862 29096
rect 9876 29084 9904 29115
rect 10042 29112 10048 29164
rect 10100 29112 10106 29164
rect 10226 29112 10232 29164
rect 10284 29112 10290 29164
rect 10686 29112 10692 29164
rect 10744 29112 10750 29164
rect 10888 29161 10916 29192
rect 11164 29161 11192 29192
rect 12710 29180 12716 29192
rect 12768 29220 12774 29232
rect 13170 29220 13176 29232
rect 12768 29192 13176 29220
rect 12768 29180 12774 29192
rect 13170 29180 13176 29192
rect 13228 29220 13234 29232
rect 15378 29220 15384 29232
rect 13228 29192 13768 29220
rect 13228 29180 13234 29192
rect 10873 29155 10931 29161
rect 10873 29121 10885 29155
rect 10919 29121 10931 29155
rect 10873 29115 10931 29121
rect 10965 29155 11023 29161
rect 10965 29121 10977 29155
rect 11011 29121 11023 29155
rect 10965 29115 11023 29121
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29121 11207 29155
rect 11149 29115 11207 29121
rect 12805 29155 12863 29161
rect 12805 29121 12817 29155
rect 12851 29121 12863 29155
rect 12805 29115 12863 29121
rect 9876 29056 10272 29084
rect 10244 29028 10272 29056
rect 10502 29044 10508 29096
rect 10560 29084 10566 29096
rect 10980 29084 11008 29115
rect 10560 29056 11008 29084
rect 12820 29084 12848 29115
rect 13078 29112 13084 29164
rect 13136 29112 13142 29164
rect 13265 29155 13323 29161
rect 13265 29121 13277 29155
rect 13311 29152 13323 29155
rect 13357 29155 13415 29161
rect 13357 29152 13369 29155
rect 13311 29124 13369 29152
rect 13311 29121 13323 29124
rect 13265 29115 13323 29121
rect 13357 29121 13369 29124
rect 13403 29152 13415 29155
rect 13446 29152 13452 29164
rect 13403 29124 13452 29152
rect 13403 29121 13415 29124
rect 13357 29115 13415 29121
rect 13446 29112 13452 29124
rect 13504 29112 13510 29164
rect 12820 29056 13676 29084
rect 10560 29044 10566 29056
rect 8297 29019 8355 29025
rect 8297 28985 8309 29019
rect 8343 29016 8355 29019
rect 10137 29019 10195 29025
rect 10137 29016 10149 29019
rect 8343 28988 8432 29016
rect 8343 28985 8355 28988
rect 8297 28979 8355 28985
rect 3234 28908 3240 28960
rect 3292 28908 3298 28960
rect 4614 28908 4620 28960
rect 4672 28948 4678 28960
rect 4890 28948 4896 28960
rect 4672 28920 4896 28948
rect 4672 28908 4678 28920
rect 4890 28908 4896 28920
rect 4948 28908 4954 28960
rect 8404 28948 8432 28988
rect 9324 28988 10149 29016
rect 9030 28948 9036 28960
rect 8404 28920 9036 28948
rect 9030 28908 9036 28920
rect 9088 28948 9094 28960
rect 9324 28948 9352 28988
rect 10137 28985 10149 28988
rect 10183 28985 10195 29019
rect 10137 28979 10195 28985
rect 10226 28976 10232 29028
rect 10284 29016 10290 29028
rect 12526 29016 12532 29028
rect 10284 28988 12532 29016
rect 10284 28976 10290 28988
rect 12526 28976 12532 28988
rect 12584 28976 12590 29028
rect 12710 28976 12716 29028
rect 12768 29016 12774 29028
rect 13262 29016 13268 29028
rect 12768 28988 13268 29016
rect 12768 28976 12774 28988
rect 13262 28976 13268 28988
rect 13320 29016 13326 29028
rect 13495 29019 13553 29025
rect 13495 29016 13507 29019
rect 13320 28988 13507 29016
rect 13320 28976 13326 28988
rect 13495 28985 13507 28988
rect 13541 28985 13553 29019
rect 13495 28979 13553 28985
rect 13648 28960 13676 29056
rect 13740 29016 13768 29192
rect 14936 29192 15384 29220
rect 13817 29155 13875 29161
rect 13817 29121 13829 29155
rect 13863 29152 13875 29155
rect 14182 29152 14188 29164
rect 13863 29124 14188 29152
rect 13863 29121 13875 29124
rect 13817 29115 13875 29121
rect 14182 29112 14188 29124
rect 14240 29112 14246 29164
rect 14936 29161 14964 29192
rect 15378 29180 15384 29192
rect 15436 29220 15442 29232
rect 15562 29220 15568 29232
rect 15436 29192 15568 29220
rect 15436 29180 15442 29192
rect 15562 29180 15568 29192
rect 15620 29180 15626 29232
rect 14921 29155 14979 29161
rect 14921 29121 14933 29155
rect 14967 29121 14979 29155
rect 14921 29115 14979 29121
rect 15197 29155 15255 29161
rect 15197 29121 15209 29155
rect 15243 29152 15255 29155
rect 16040 29152 16068 29248
rect 16117 29223 16175 29229
rect 16117 29189 16129 29223
rect 16163 29220 16175 29223
rect 16206 29220 16212 29232
rect 16163 29192 16212 29220
rect 16163 29189 16175 29192
rect 16117 29183 16175 29189
rect 16206 29180 16212 29192
rect 16264 29180 16270 29232
rect 17865 29223 17923 29229
rect 17865 29220 17877 29223
rect 17052 29192 17877 29220
rect 17052 29164 17080 29192
rect 17865 29189 17877 29192
rect 17911 29189 17923 29223
rect 17865 29183 17923 29189
rect 15243 29124 16068 29152
rect 15243 29121 15255 29124
rect 15197 29115 15255 29121
rect 16666 29112 16672 29164
rect 16724 29112 16730 29164
rect 16945 29155 17003 29161
rect 16945 29121 16957 29155
rect 16991 29152 17003 29155
rect 17034 29152 17040 29164
rect 16991 29124 17040 29152
rect 16991 29121 17003 29124
rect 16945 29115 17003 29121
rect 17034 29112 17040 29124
rect 17092 29112 17098 29164
rect 17126 29112 17132 29164
rect 17184 29112 17190 29164
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29152 17371 29155
rect 17359 29124 17448 29152
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 17420 29096 17448 29124
rect 17586 29112 17592 29164
rect 17644 29112 17650 29164
rect 17747 29155 17805 29161
rect 17747 29121 17759 29155
rect 17793 29152 17805 29155
rect 17793 29124 17908 29152
rect 17793 29121 17805 29124
rect 17747 29115 17805 29121
rect 15286 29044 15292 29096
rect 15344 29044 15350 29096
rect 15565 29087 15623 29093
rect 15565 29053 15577 29087
rect 15611 29053 15623 29087
rect 15565 29047 15623 29053
rect 15580 29016 15608 29047
rect 15654 29044 15660 29096
rect 15712 29044 15718 29096
rect 17402 29044 17408 29096
rect 17460 29044 17466 29096
rect 17880 29084 17908 29124
rect 17954 29112 17960 29164
rect 18012 29112 18018 29164
rect 18049 29155 18107 29161
rect 18049 29121 18061 29155
rect 18095 29152 18107 29155
rect 18230 29152 18236 29164
rect 18095 29124 18236 29152
rect 18095 29121 18107 29124
rect 18049 29115 18107 29121
rect 18230 29112 18236 29124
rect 18288 29112 18294 29164
rect 18616 29161 18644 29260
rect 18785 29257 18797 29291
rect 18831 29288 18843 29291
rect 19242 29288 19248 29300
rect 18831 29260 19248 29288
rect 18831 29257 18843 29260
rect 18785 29251 18843 29257
rect 19242 29248 19248 29260
rect 19300 29248 19306 29300
rect 23198 29248 23204 29300
rect 23256 29288 23262 29300
rect 26786 29288 26792 29300
rect 23256 29260 26792 29288
rect 23256 29248 23262 29260
rect 21634 29220 21640 29232
rect 20548 29192 21640 29220
rect 20548 29164 20576 29192
rect 21634 29180 21640 29192
rect 21692 29220 21698 29232
rect 22097 29223 22155 29229
rect 22097 29220 22109 29223
rect 21692 29192 22109 29220
rect 21692 29180 21698 29192
rect 22097 29189 22109 29192
rect 22143 29189 22155 29223
rect 22097 29183 22155 29189
rect 22189 29223 22247 29229
rect 22189 29189 22201 29223
rect 22235 29220 22247 29223
rect 22370 29220 22376 29232
rect 22235 29192 22376 29220
rect 22235 29189 22247 29192
rect 22189 29183 22247 29189
rect 22370 29180 22376 29192
rect 22428 29180 22434 29232
rect 22833 29223 22891 29229
rect 22833 29189 22845 29223
rect 22879 29220 22891 29223
rect 22922 29220 22928 29232
rect 22879 29192 22928 29220
rect 22879 29189 22891 29192
rect 22833 29183 22891 29189
rect 22922 29180 22928 29192
rect 22980 29180 22986 29232
rect 23569 29223 23627 29229
rect 23569 29189 23581 29223
rect 23615 29220 23627 29223
rect 24486 29220 24492 29232
rect 23615 29192 24492 29220
rect 23615 29189 23627 29192
rect 23569 29183 23627 29189
rect 24486 29180 24492 29192
rect 24544 29180 24550 29232
rect 18601 29155 18659 29161
rect 18601 29121 18613 29155
rect 18647 29121 18659 29155
rect 18601 29115 18659 29121
rect 20254 29112 20260 29164
rect 20312 29112 20318 29164
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29152 20499 29155
rect 20530 29152 20536 29164
rect 20487 29124 20536 29152
rect 20487 29121 20499 29124
rect 20441 29115 20499 29121
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 21910 29112 21916 29164
rect 21968 29112 21974 29164
rect 22281 29155 22339 29161
rect 22281 29121 22293 29155
rect 22327 29121 22339 29155
rect 22388 29152 22416 29180
rect 23382 29152 23388 29164
rect 22388 29124 23388 29152
rect 22281 29115 22339 29121
rect 18138 29084 18144 29096
rect 17880 29056 18144 29084
rect 18138 29044 18144 29056
rect 18196 29044 18202 29096
rect 18325 29087 18383 29093
rect 18325 29053 18337 29087
rect 18371 29084 18383 29087
rect 18690 29084 18696 29096
rect 18371 29056 18696 29084
rect 18371 29053 18383 29056
rect 18325 29047 18383 29053
rect 18690 29044 18696 29056
rect 18748 29044 18754 29096
rect 18782 29044 18788 29096
rect 18840 29084 18846 29096
rect 22296 29084 22324 29115
rect 23382 29112 23388 29124
rect 23440 29112 23446 29164
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29152 24087 29155
rect 24302 29152 24308 29164
rect 24075 29124 24308 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 24302 29112 24308 29124
rect 24360 29112 24366 29164
rect 25774 29112 25780 29164
rect 25832 29112 25838 29164
rect 25976 29161 26004 29260
rect 26786 29248 26792 29260
rect 26844 29248 26850 29300
rect 27985 29291 28043 29297
rect 27985 29257 27997 29291
rect 28031 29288 28043 29291
rect 28442 29288 28448 29300
rect 28031 29260 28448 29288
rect 28031 29257 28043 29260
rect 27985 29251 28043 29257
rect 28442 29248 28448 29260
rect 28500 29248 28506 29300
rect 32490 29248 32496 29300
rect 32548 29288 32554 29300
rect 32677 29291 32735 29297
rect 32677 29288 32689 29291
rect 32548 29260 32689 29288
rect 32548 29248 32554 29260
rect 32677 29257 32689 29260
rect 32723 29257 32735 29291
rect 32677 29251 32735 29257
rect 32769 29291 32827 29297
rect 32769 29257 32781 29291
rect 32815 29288 32827 29291
rect 32858 29288 32864 29300
rect 32815 29260 32864 29288
rect 32815 29257 32827 29260
rect 32769 29251 32827 29257
rect 32858 29248 32864 29260
rect 32916 29248 32922 29300
rect 34146 29288 34152 29300
rect 33060 29260 34152 29288
rect 27709 29223 27767 29229
rect 27709 29189 27721 29223
rect 27755 29220 27767 29223
rect 29178 29220 29184 29232
rect 27755 29192 29184 29220
rect 27755 29189 27767 29192
rect 27709 29183 27767 29189
rect 29178 29180 29184 29192
rect 29236 29180 29242 29232
rect 30926 29180 30932 29232
rect 30984 29220 30990 29232
rect 31205 29223 31263 29229
rect 31205 29220 31217 29223
rect 30984 29192 31217 29220
rect 30984 29180 30990 29192
rect 31205 29189 31217 29192
rect 31251 29189 31263 29223
rect 31205 29183 31263 29189
rect 31297 29223 31355 29229
rect 31297 29189 31309 29223
rect 31343 29220 31355 29223
rect 31343 29192 32260 29220
rect 31343 29189 31355 29192
rect 31297 29183 31355 29189
rect 25961 29155 26019 29161
rect 25961 29121 25973 29155
rect 26007 29121 26019 29155
rect 25961 29115 26019 29121
rect 26418 29112 26424 29164
rect 26476 29152 26482 29164
rect 27433 29155 27491 29161
rect 27433 29152 27445 29155
rect 26476 29124 27445 29152
rect 26476 29112 26482 29124
rect 27433 29121 27445 29124
rect 27479 29152 27491 29155
rect 27522 29152 27528 29164
rect 27479 29124 27528 29152
rect 27479 29121 27491 29124
rect 27433 29115 27491 29121
rect 27522 29112 27528 29124
rect 27580 29112 27586 29164
rect 27617 29155 27675 29161
rect 27617 29121 27629 29155
rect 27663 29152 27675 29155
rect 27663 29124 27752 29152
rect 27663 29121 27675 29124
rect 27617 29115 27675 29121
rect 18840 29056 22324 29084
rect 18840 29044 18846 29056
rect 23474 29044 23480 29096
rect 23532 29084 23538 29096
rect 23753 29087 23811 29093
rect 23753 29084 23765 29087
rect 23532 29056 23765 29084
rect 23532 29044 23538 29056
rect 23753 29053 23765 29056
rect 23799 29084 23811 29087
rect 23799 29056 27660 29084
rect 23799 29053 23811 29056
rect 23753 29047 23811 29053
rect 18800 29016 18828 29044
rect 27632 29028 27660 29056
rect 13740 28988 18828 29016
rect 20441 29019 20499 29025
rect 20441 28985 20453 29019
rect 20487 29016 20499 29019
rect 21174 29016 21180 29028
rect 20487 28988 21180 29016
rect 20487 28985 20499 28988
rect 20441 28979 20499 28985
rect 21174 28976 21180 28988
rect 21232 28976 21238 29028
rect 22465 29019 22523 29025
rect 22465 28985 22477 29019
rect 22511 29016 22523 29019
rect 24578 29016 24584 29028
rect 22511 28988 24584 29016
rect 22511 28985 22523 28988
rect 22465 28979 22523 28985
rect 24578 28976 24584 28988
rect 24636 28976 24642 29028
rect 24670 28976 24676 29028
rect 24728 29016 24734 29028
rect 24728 28988 27568 29016
rect 24728 28976 24734 28988
rect 9088 28920 9352 28948
rect 9088 28908 9094 28920
rect 10318 28908 10324 28960
rect 10376 28908 10382 28960
rect 10594 28908 10600 28960
rect 10652 28908 10658 28960
rect 13630 28908 13636 28960
rect 13688 28908 13694 28960
rect 13722 28908 13728 28960
rect 13780 28908 13786 28960
rect 13906 28908 13912 28960
rect 13964 28948 13970 28960
rect 16298 28948 16304 28960
rect 13964 28920 16304 28948
rect 13964 28908 13970 28920
rect 16298 28908 16304 28920
rect 16356 28908 16362 28960
rect 16390 28908 16396 28960
rect 16448 28948 16454 28960
rect 16758 28948 16764 28960
rect 16448 28920 16764 28948
rect 16448 28908 16454 28920
rect 16758 28908 16764 28920
rect 16816 28908 16822 28960
rect 18417 28951 18475 28957
rect 18417 28917 18429 28951
rect 18463 28948 18475 28951
rect 18506 28948 18512 28960
rect 18463 28920 18512 28948
rect 18463 28917 18475 28920
rect 18417 28911 18475 28917
rect 18506 28908 18512 28920
rect 18564 28908 18570 28960
rect 21082 28908 21088 28960
rect 21140 28948 21146 28960
rect 22002 28948 22008 28960
rect 21140 28920 22008 28948
rect 21140 28908 21146 28920
rect 22002 28908 22008 28920
rect 22060 28948 22066 28960
rect 25222 28948 25228 28960
rect 22060 28920 25228 28948
rect 22060 28908 22066 28920
rect 25222 28908 25228 28920
rect 25280 28908 25286 28960
rect 25314 28908 25320 28960
rect 25372 28948 25378 28960
rect 25777 28951 25835 28957
rect 25777 28948 25789 28951
rect 25372 28920 25789 28948
rect 25372 28908 25378 28920
rect 25777 28917 25789 28920
rect 25823 28917 25835 28951
rect 27540 28948 27568 28988
rect 27614 28976 27620 29028
rect 27672 28976 27678 29028
rect 27724 29016 27752 29124
rect 27798 29112 27804 29164
rect 27856 29112 27862 29164
rect 29454 29112 29460 29164
rect 29512 29112 29518 29164
rect 29638 29112 29644 29164
rect 29696 29112 29702 29164
rect 30466 29112 30472 29164
rect 30524 29112 30530 29164
rect 30561 29155 30619 29161
rect 30561 29121 30573 29155
rect 30607 29152 30619 29155
rect 30837 29155 30895 29161
rect 30607 29124 30696 29152
rect 30607 29121 30619 29124
rect 30561 29115 30619 29121
rect 30668 29095 30696 29124
rect 30837 29121 30849 29155
rect 30883 29152 30895 29155
rect 30883 29124 30972 29152
rect 30883 29121 30895 29124
rect 30837 29115 30895 29121
rect 30668 29084 30788 29095
rect 30944 29084 30972 29124
rect 31018 29112 31024 29164
rect 31076 29161 31082 29164
rect 31076 29155 31125 29161
rect 31076 29121 31079 29155
rect 31113 29121 31125 29155
rect 31478 29152 31484 29164
rect 31439 29124 31484 29152
rect 31076 29115 31125 29121
rect 31076 29112 31082 29115
rect 31478 29112 31484 29124
rect 31536 29112 31542 29164
rect 31573 29155 31631 29161
rect 31573 29121 31585 29155
rect 31619 29152 31631 29155
rect 31662 29152 31668 29164
rect 31619 29124 31668 29152
rect 31619 29121 31631 29124
rect 31573 29115 31631 29121
rect 31662 29112 31668 29124
rect 31720 29112 31726 29164
rect 32232 29152 32260 29192
rect 32306 29180 32312 29232
rect 32364 29220 32370 29232
rect 32950 29220 32956 29232
rect 32364 29192 32956 29220
rect 32364 29180 32370 29192
rect 32950 29180 32956 29192
rect 33008 29180 33014 29232
rect 32766 29152 32772 29164
rect 32232 29124 32772 29152
rect 32766 29112 32772 29124
rect 32824 29152 32830 29164
rect 33060 29152 33088 29260
rect 34146 29248 34152 29260
rect 34204 29288 34210 29300
rect 34422 29288 34428 29300
rect 34204 29260 34428 29288
rect 34204 29248 34210 29260
rect 34422 29248 34428 29260
rect 34480 29248 34486 29300
rect 34882 29248 34888 29300
rect 34940 29248 34946 29300
rect 36354 29248 36360 29300
rect 36412 29288 36418 29300
rect 36538 29288 36544 29300
rect 36412 29260 36544 29288
rect 36412 29248 36418 29260
rect 36538 29248 36544 29260
rect 36596 29248 36602 29300
rect 38105 29291 38163 29297
rect 38105 29288 38117 29291
rect 37476 29260 38117 29288
rect 33134 29180 33140 29232
rect 33192 29220 33198 29232
rect 33413 29223 33471 29229
rect 33413 29220 33425 29223
rect 33192 29192 33425 29220
rect 33192 29180 33198 29192
rect 33413 29189 33425 29192
rect 33459 29189 33471 29223
rect 33413 29183 33471 29189
rect 33505 29223 33563 29229
rect 33505 29189 33517 29223
rect 33551 29220 33563 29223
rect 34606 29220 34612 29232
rect 33551 29192 34612 29220
rect 33551 29189 33563 29192
rect 33505 29183 33563 29189
rect 32824 29124 33088 29152
rect 32824 29112 32830 29124
rect 33226 29112 33232 29164
rect 33284 29112 33290 29164
rect 33597 29155 33655 29161
rect 33597 29152 33609 29155
rect 33336 29124 33609 29152
rect 30668 29067 30880 29084
rect 30760 29056 30880 29067
rect 30944 29056 31616 29084
rect 27798 29016 27804 29028
rect 27724 28988 27804 29016
rect 27798 28976 27804 28988
rect 27856 28976 27862 29028
rect 27982 28976 27988 29028
rect 28040 29016 28046 29028
rect 29638 29016 29644 29028
rect 28040 28988 29644 29016
rect 28040 28976 28046 28988
rect 29638 28976 29644 28988
rect 29696 28976 29702 29028
rect 30285 29019 30343 29025
rect 30285 28985 30297 29019
rect 30331 29016 30343 29019
rect 30466 29016 30472 29028
rect 30331 28988 30472 29016
rect 30331 28985 30343 28988
rect 30285 28979 30343 28985
rect 30466 28976 30472 28988
rect 30524 28976 30530 29028
rect 30650 28976 30656 29028
rect 30708 29016 30714 29028
rect 30745 29019 30803 29025
rect 30745 29016 30757 29019
rect 30708 28988 30757 29016
rect 30708 28976 30714 28988
rect 30745 28985 30757 28988
rect 30791 28985 30803 29019
rect 30852 29016 30880 29056
rect 31588 29028 31616 29056
rect 31754 29044 31760 29096
rect 31812 29084 31818 29096
rect 32585 29087 32643 29093
rect 32585 29084 32597 29087
rect 31812 29056 32597 29084
rect 31812 29044 31818 29056
rect 32585 29053 32597 29056
rect 32631 29084 32643 29087
rect 33042 29084 33048 29096
rect 32631 29056 33048 29084
rect 32631 29053 32643 29056
rect 32585 29047 32643 29053
rect 33042 29044 33048 29056
rect 33100 29044 33106 29096
rect 33336 29084 33364 29124
rect 33597 29121 33609 29124
rect 33643 29121 33655 29155
rect 33597 29115 33655 29121
rect 33704 29084 33732 29192
rect 34606 29180 34612 29192
rect 34664 29180 34670 29232
rect 35986 29220 35992 29232
rect 35176 29192 35992 29220
rect 33870 29112 33876 29164
rect 33928 29152 33934 29164
rect 34057 29155 34115 29161
rect 34057 29152 34069 29155
rect 33928 29124 34069 29152
rect 33928 29112 33934 29124
rect 34057 29121 34069 29124
rect 34103 29121 34115 29155
rect 34057 29115 34115 29121
rect 34146 29112 34152 29164
rect 34204 29112 34210 29164
rect 34330 29112 34336 29164
rect 34388 29152 34394 29164
rect 34425 29155 34483 29161
rect 34425 29152 34437 29155
rect 34388 29124 34437 29152
rect 34388 29112 34394 29124
rect 34425 29121 34437 29124
rect 34471 29152 34483 29155
rect 34514 29152 34520 29164
rect 34471 29124 34520 29152
rect 34471 29121 34483 29124
rect 34425 29115 34483 29121
rect 34514 29112 34520 29124
rect 34572 29112 34578 29164
rect 35066 29112 35072 29164
rect 35124 29112 35130 29164
rect 35176 29161 35204 29192
rect 35986 29180 35992 29192
rect 36044 29180 36050 29232
rect 35161 29155 35219 29161
rect 35161 29121 35173 29155
rect 35207 29121 35219 29155
rect 35161 29115 35219 29121
rect 35345 29155 35403 29161
rect 35345 29121 35357 29155
rect 35391 29121 35403 29155
rect 35345 29115 35403 29121
rect 33152 29056 33364 29084
rect 33520 29056 33732 29084
rect 33152 29028 33180 29056
rect 30929 29019 30987 29025
rect 30929 29016 30941 29019
rect 30852 28988 30941 29016
rect 30745 28979 30803 28985
rect 30929 28985 30941 28988
rect 30975 28985 30987 29019
rect 30929 28979 30987 28985
rect 27816 28948 27844 28976
rect 27540 28920 27844 28948
rect 29457 28951 29515 28957
rect 25777 28911 25835 28917
rect 29457 28917 29469 28951
rect 29503 28948 29515 28951
rect 29730 28948 29736 28960
rect 29503 28920 29736 28948
rect 29503 28917 29515 28920
rect 29457 28911 29515 28917
rect 29730 28908 29736 28920
rect 29788 28908 29794 28960
rect 30760 28948 30788 28979
rect 31570 28976 31576 29028
rect 31628 28976 31634 29028
rect 33134 28976 33140 29028
rect 33192 28976 33198 29028
rect 33520 29016 33548 29056
rect 33778 29044 33784 29096
rect 33836 29084 33842 29096
rect 34885 29087 34943 29093
rect 33836 29056 34192 29084
rect 33836 29044 33842 29056
rect 33873 29019 33931 29025
rect 33873 29016 33885 29019
rect 33244 28988 33548 29016
rect 33612 28988 33885 29016
rect 30834 28948 30840 28960
rect 30760 28920 30840 28948
rect 30834 28908 30840 28920
rect 30892 28908 30898 28960
rect 32950 28908 32956 28960
rect 33008 28948 33014 28960
rect 33244 28948 33272 28988
rect 33008 28920 33272 28948
rect 33008 28908 33014 28920
rect 33318 28908 33324 28960
rect 33376 28948 33382 28960
rect 33612 28948 33640 28988
rect 33873 28985 33885 28988
rect 33919 28985 33931 29019
rect 33873 28979 33931 28985
rect 33962 28976 33968 29028
rect 34020 28976 34026 29028
rect 33376 28920 33640 28948
rect 33781 28951 33839 28957
rect 33376 28908 33382 28920
rect 33781 28917 33793 28951
rect 33827 28948 33839 28951
rect 33980 28948 34008 28976
rect 33827 28920 34008 28948
rect 34164 28948 34192 29056
rect 34885 29053 34897 29087
rect 34931 29084 34943 29087
rect 34974 29084 34980 29096
rect 34931 29056 34980 29084
rect 34931 29053 34943 29056
rect 34885 29047 34943 29053
rect 34974 29044 34980 29056
rect 35032 29044 35038 29096
rect 35084 29084 35112 29112
rect 35360 29084 35388 29115
rect 35434 29112 35440 29164
rect 35492 29152 35498 29164
rect 35529 29155 35587 29161
rect 35529 29152 35541 29155
rect 35492 29124 35541 29152
rect 35492 29112 35498 29124
rect 35529 29121 35541 29124
rect 35575 29121 35587 29155
rect 35529 29115 35587 29121
rect 37277 29155 37335 29161
rect 37277 29121 37289 29155
rect 37323 29152 37335 29155
rect 37476 29152 37504 29260
rect 38105 29257 38117 29260
rect 38151 29288 38163 29291
rect 38838 29288 38844 29300
rect 38151 29260 38844 29288
rect 38151 29257 38163 29260
rect 38105 29251 38163 29257
rect 38838 29248 38844 29260
rect 38896 29248 38902 29300
rect 39577 29291 39635 29297
rect 39577 29257 39589 29291
rect 39623 29288 39635 29291
rect 40034 29288 40040 29300
rect 39623 29260 40040 29288
rect 39623 29257 39635 29260
rect 39577 29251 39635 29257
rect 40034 29248 40040 29260
rect 40092 29248 40098 29300
rect 37918 29180 37924 29232
rect 37976 29180 37982 29232
rect 39206 29220 39212 29232
rect 37323 29124 37504 29152
rect 37323 29121 37335 29124
rect 37277 29115 37335 29121
rect 37550 29112 37556 29164
rect 37608 29112 37614 29164
rect 37645 29155 37703 29161
rect 37645 29121 37657 29155
rect 37691 29152 37703 29155
rect 37691 29124 37964 29152
rect 38102 29146 38108 29198
rect 38160 29152 38166 29198
rect 38304 29192 39212 29220
rect 38197 29155 38255 29161
rect 38197 29152 38209 29155
rect 38160 29146 38209 29152
rect 38120 29124 38209 29146
rect 37691 29121 37703 29124
rect 37645 29115 37703 29121
rect 37182 29084 37188 29096
rect 35084 29056 35388 29084
rect 35452 29056 37188 29084
rect 34238 28976 34244 29028
rect 34296 29016 34302 29028
rect 35452 29016 35480 29056
rect 37182 29044 37188 29056
rect 37240 29084 37246 29096
rect 37826 29084 37832 29096
rect 37240 29056 37832 29084
rect 37240 29044 37246 29056
rect 37826 29044 37832 29056
rect 37884 29044 37890 29096
rect 34296 28988 35480 29016
rect 35529 29019 35587 29025
rect 34296 28976 34302 28988
rect 35529 28985 35541 29019
rect 35575 29016 35587 29019
rect 36354 29016 36360 29028
rect 35575 28988 36360 29016
rect 35575 28985 35587 28988
rect 35529 28979 35587 28985
rect 36354 28976 36360 28988
rect 36412 28976 36418 29028
rect 37369 29019 37427 29025
rect 37369 28985 37381 29019
rect 37415 29016 37427 29019
rect 37734 29016 37740 29028
rect 37415 28988 37740 29016
rect 37415 28985 37427 28988
rect 37369 28979 37427 28985
rect 37734 28976 37740 28988
rect 37792 28976 37798 29028
rect 37936 29025 37964 29124
rect 38197 29121 38209 29124
rect 38243 29121 38255 29155
rect 38197 29115 38255 29121
rect 38102 29044 38108 29096
rect 38160 29084 38166 29096
rect 38304 29084 38332 29192
rect 39206 29180 39212 29192
rect 39264 29180 39270 29232
rect 39301 29223 39359 29229
rect 39301 29189 39313 29223
rect 39347 29220 39359 29223
rect 39850 29220 39856 29232
rect 39347 29192 39856 29220
rect 39347 29189 39359 29192
rect 39301 29183 39359 29189
rect 39850 29180 39856 29192
rect 39908 29180 39914 29232
rect 39945 29223 40003 29229
rect 39945 29189 39957 29223
rect 39991 29220 40003 29223
rect 40218 29220 40224 29232
rect 39991 29192 40224 29220
rect 39991 29189 40003 29192
rect 39945 29183 40003 29189
rect 40218 29180 40224 29192
rect 40276 29180 40282 29232
rect 41966 29220 41972 29232
rect 41170 29192 41972 29220
rect 41966 29180 41972 29192
rect 42024 29180 42030 29232
rect 39025 29155 39083 29161
rect 39025 29121 39037 29155
rect 39071 29152 39083 29155
rect 39114 29152 39120 29164
rect 39071 29124 39120 29152
rect 39071 29121 39083 29124
rect 39025 29115 39083 29121
rect 39114 29112 39120 29124
rect 39172 29112 39178 29164
rect 39393 29155 39451 29161
rect 39393 29121 39405 29155
rect 39439 29152 39451 29155
rect 39574 29152 39580 29164
rect 39439 29124 39580 29152
rect 39439 29121 39451 29124
rect 39393 29115 39451 29121
rect 39408 29084 39436 29115
rect 39574 29112 39580 29124
rect 39632 29112 39638 29164
rect 41877 29155 41935 29161
rect 41877 29152 41889 29155
rect 41432 29124 41889 29152
rect 38160 29056 38332 29084
rect 39040 29056 39436 29084
rect 39669 29087 39727 29093
rect 38160 29044 38166 29056
rect 39040 29028 39068 29056
rect 39669 29053 39681 29087
rect 39715 29084 39727 29087
rect 39715 29056 39804 29084
rect 39715 29053 39727 29056
rect 39669 29047 39727 29053
rect 37921 29019 37979 29025
rect 37921 28985 37933 29019
rect 37967 28985 37979 29019
rect 37921 28979 37979 28985
rect 39022 28976 39028 29028
rect 39080 28976 39086 29028
rect 34333 28951 34391 28957
rect 34333 28948 34345 28951
rect 34164 28920 34345 28948
rect 33827 28917 33839 28920
rect 33781 28911 33839 28917
rect 34333 28917 34345 28920
rect 34379 28917 34391 28951
rect 34333 28911 34391 28917
rect 34422 28908 34428 28960
rect 34480 28948 34486 28960
rect 35710 28948 35716 28960
rect 34480 28920 35716 28948
rect 34480 28908 34486 28920
rect 35710 28908 35716 28920
rect 35768 28948 35774 28960
rect 36906 28948 36912 28960
rect 35768 28920 36912 28948
rect 35768 28908 35774 28920
rect 36906 28908 36912 28920
rect 36964 28908 36970 28960
rect 37642 28908 37648 28960
rect 37700 28948 37706 28960
rect 37829 28951 37887 28957
rect 37829 28948 37841 28951
rect 37700 28920 37841 28948
rect 37700 28908 37706 28920
rect 37829 28917 37841 28920
rect 37875 28917 37887 28951
rect 39776 28948 39804 29056
rect 39942 29044 39948 29096
rect 40000 29084 40006 29096
rect 41432 29093 41460 29124
rect 41877 29121 41889 29124
rect 41923 29121 41935 29155
rect 41877 29115 41935 29121
rect 41417 29087 41475 29093
rect 41417 29084 41429 29087
rect 40000 29056 41429 29084
rect 40000 29044 40006 29056
rect 41417 29053 41429 29056
rect 41463 29053 41475 29087
rect 41417 29047 41475 29053
rect 42058 28976 42064 29028
rect 42116 28976 42122 29028
rect 40402 28948 40408 28960
rect 39776 28920 40408 28948
rect 37829 28911 37887 28917
rect 40402 28908 40408 28920
rect 40460 28908 40466 28960
rect 1104 28858 42504 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 42504 28858
rect 1104 28784 42504 28806
rect 1670 28704 1676 28756
rect 1728 28744 1734 28756
rect 2593 28747 2651 28753
rect 2593 28744 2605 28747
rect 1728 28716 2605 28744
rect 1728 28704 1734 28716
rect 2593 28713 2605 28716
rect 2639 28713 2651 28747
rect 2593 28707 2651 28713
rect 2961 28747 3019 28753
rect 2961 28713 2973 28747
rect 3007 28744 3019 28747
rect 3234 28744 3240 28756
rect 3007 28716 3240 28744
rect 3007 28713 3019 28716
rect 2961 28707 3019 28713
rect 3234 28704 3240 28716
rect 3292 28704 3298 28756
rect 4617 28747 4675 28753
rect 4617 28713 4629 28747
rect 4663 28744 4675 28747
rect 5258 28744 5264 28756
rect 4663 28716 5264 28744
rect 4663 28713 4675 28716
rect 4617 28707 4675 28713
rect 5258 28704 5264 28716
rect 5316 28704 5322 28756
rect 6917 28747 6975 28753
rect 6917 28713 6929 28747
rect 6963 28744 6975 28747
rect 7098 28744 7104 28756
rect 6963 28716 7104 28744
rect 6963 28713 6975 28716
rect 6917 28707 6975 28713
rect 7098 28704 7104 28716
rect 7156 28704 7162 28756
rect 9122 28704 9128 28756
rect 9180 28704 9186 28756
rect 9674 28704 9680 28756
rect 9732 28704 9738 28756
rect 12437 28747 12495 28753
rect 12437 28713 12449 28747
rect 12483 28744 12495 28747
rect 12802 28744 12808 28756
rect 12483 28716 12808 28744
rect 12483 28713 12495 28716
rect 12437 28707 12495 28713
rect 12802 28704 12808 28716
rect 12860 28704 12866 28756
rect 13630 28704 13636 28756
rect 13688 28744 13694 28756
rect 16574 28744 16580 28756
rect 13688 28716 16580 28744
rect 13688 28704 13694 28716
rect 16574 28704 16580 28716
rect 16632 28704 16638 28756
rect 17034 28744 17040 28756
rect 16776 28716 17040 28744
rect 3510 28636 3516 28688
rect 3568 28676 3574 28688
rect 4709 28679 4767 28685
rect 4709 28676 4721 28679
rect 3568 28648 4721 28676
rect 3568 28636 3574 28648
rect 2777 28543 2835 28549
rect 2777 28509 2789 28543
rect 2823 28540 2835 28543
rect 2958 28540 2964 28552
rect 2823 28512 2964 28540
rect 2823 28509 2835 28512
rect 2777 28503 2835 28509
rect 2958 28500 2964 28512
rect 3016 28500 3022 28552
rect 3050 28500 3056 28552
rect 3108 28500 3114 28552
rect 4080 28549 4108 28648
rect 4709 28645 4721 28648
rect 4755 28645 4767 28679
rect 4709 28639 4767 28645
rect 8757 28679 8815 28685
rect 8757 28645 8769 28679
rect 8803 28676 8815 28679
rect 9692 28676 9720 28704
rect 16776 28688 16804 28716
rect 17034 28704 17040 28716
rect 17092 28704 17098 28756
rect 17313 28747 17371 28753
rect 17313 28713 17325 28747
rect 17359 28713 17371 28747
rect 17313 28707 17371 28713
rect 10318 28676 10324 28688
rect 8803 28648 10324 28676
rect 8803 28645 8815 28648
rect 8757 28639 8815 28645
rect 10318 28636 10324 28648
rect 10376 28636 10382 28688
rect 12069 28679 12127 28685
rect 12069 28645 12081 28679
rect 12115 28676 12127 28679
rect 12115 28648 12434 28676
rect 12115 28645 12127 28648
rect 12069 28639 12127 28645
rect 4614 28568 4620 28620
rect 4672 28608 4678 28620
rect 5166 28608 5172 28620
rect 4672 28580 5172 28608
rect 4672 28568 4678 28580
rect 5166 28568 5172 28580
rect 5224 28568 5230 28620
rect 9582 28568 9588 28620
rect 9640 28608 9646 28620
rect 9677 28611 9735 28617
rect 9677 28608 9689 28611
rect 9640 28580 9689 28608
rect 9640 28568 9646 28580
rect 9677 28577 9689 28580
rect 9723 28608 9735 28611
rect 9723 28580 10272 28608
rect 9723 28577 9735 28580
rect 9677 28571 9735 28577
rect 4065 28543 4123 28549
rect 4065 28509 4077 28543
rect 4111 28509 4123 28543
rect 4065 28503 4123 28509
rect 4433 28543 4491 28549
rect 4433 28509 4445 28543
rect 4479 28540 4491 28543
rect 4709 28543 4767 28549
rect 4709 28540 4721 28543
rect 4479 28512 4721 28540
rect 4479 28509 4491 28512
rect 4433 28503 4491 28509
rect 4709 28509 4721 28512
rect 4755 28540 4767 28543
rect 4755 28512 4844 28540
rect 4755 28509 4767 28512
rect 4709 28503 4767 28509
rect 3878 28432 3884 28484
rect 3936 28472 3942 28484
rect 4249 28475 4307 28481
rect 4249 28472 4261 28475
rect 3936 28444 4261 28472
rect 3936 28432 3942 28444
rect 4249 28441 4261 28444
rect 4295 28441 4307 28475
rect 4249 28435 4307 28441
rect 4338 28432 4344 28484
rect 4396 28432 4402 28484
rect 4816 28404 4844 28512
rect 4890 28500 4896 28552
rect 4948 28500 4954 28552
rect 6546 28500 6552 28552
rect 6604 28500 6610 28552
rect 7377 28543 7435 28549
rect 7377 28509 7389 28543
rect 7423 28540 7435 28543
rect 8386 28540 8392 28552
rect 7423 28512 8392 28540
rect 7423 28509 7435 28512
rect 7377 28503 7435 28509
rect 8386 28500 8392 28512
rect 8444 28500 8450 28552
rect 9493 28543 9551 28549
rect 9493 28509 9505 28543
rect 9539 28540 9551 28543
rect 9766 28540 9772 28552
rect 9539 28512 9772 28540
rect 9539 28509 9551 28512
rect 9493 28503 9551 28509
rect 9766 28500 9772 28512
rect 9824 28500 9830 28552
rect 9953 28543 10011 28549
rect 9953 28509 9965 28543
rect 9999 28540 10011 28543
rect 10042 28540 10048 28552
rect 9999 28512 10048 28540
rect 9999 28509 10011 28512
rect 9953 28503 10011 28509
rect 10042 28500 10048 28512
rect 10100 28500 10106 28552
rect 10134 28500 10140 28552
rect 10192 28500 10198 28552
rect 5445 28475 5503 28481
rect 5445 28441 5457 28475
rect 5491 28472 5503 28475
rect 5534 28472 5540 28484
rect 5491 28444 5540 28472
rect 5491 28441 5503 28444
rect 5445 28435 5503 28441
rect 5534 28432 5540 28444
rect 5592 28432 5598 28484
rect 7644 28475 7702 28481
rect 7644 28441 7656 28475
rect 7690 28472 7702 28475
rect 8018 28472 8024 28484
rect 7690 28444 8024 28472
rect 7690 28441 7702 28444
rect 7644 28435 7702 28441
rect 8018 28432 8024 28444
rect 8076 28432 8082 28484
rect 5718 28404 5724 28416
rect 4816 28376 5724 28404
rect 5718 28364 5724 28376
rect 5776 28364 5782 28416
rect 9585 28407 9643 28413
rect 9585 28373 9597 28407
rect 9631 28404 9643 28407
rect 10045 28407 10103 28413
rect 10045 28404 10057 28407
rect 9631 28376 10057 28404
rect 9631 28373 9643 28376
rect 9585 28367 9643 28373
rect 10045 28373 10057 28376
rect 10091 28373 10103 28407
rect 10244 28404 10272 28580
rect 10594 28568 10600 28620
rect 10652 28608 10658 28620
rect 12406 28608 12434 28648
rect 12526 28636 12532 28688
rect 12584 28676 12590 28688
rect 13722 28676 13728 28688
rect 12584 28648 13728 28676
rect 12584 28636 12590 28648
rect 13722 28636 13728 28648
rect 13780 28636 13786 28688
rect 15841 28679 15899 28685
rect 15841 28645 15853 28679
rect 15887 28676 15899 28679
rect 16206 28676 16212 28688
rect 15887 28648 16212 28676
rect 15887 28645 15899 28648
rect 15841 28639 15899 28645
rect 16206 28636 16212 28648
rect 16264 28636 16270 28688
rect 16393 28679 16451 28685
rect 16393 28645 16405 28679
rect 16439 28676 16451 28679
rect 16482 28676 16488 28688
rect 16439 28648 16488 28676
rect 16439 28645 16451 28648
rect 16393 28639 16451 28645
rect 16482 28636 16488 28648
rect 16540 28636 16546 28688
rect 16758 28636 16764 28688
rect 16816 28636 16822 28688
rect 16942 28685 16948 28688
rect 16899 28679 16948 28685
rect 16899 28645 16911 28679
rect 16945 28645 16948 28679
rect 16899 28639 16948 28645
rect 16942 28636 16948 28639
rect 17000 28676 17006 28688
rect 17126 28676 17132 28688
rect 17000 28648 17132 28676
rect 17000 28636 17006 28648
rect 17126 28636 17132 28648
rect 17184 28676 17190 28688
rect 17328 28676 17356 28707
rect 17862 28704 17868 28756
rect 17920 28744 17926 28756
rect 18690 28744 18696 28756
rect 17920 28716 18696 28744
rect 17920 28704 17926 28716
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 20990 28704 20996 28756
rect 21048 28704 21054 28756
rect 22462 28704 22468 28756
rect 22520 28744 22526 28756
rect 22520 28716 24900 28744
rect 22520 28704 22526 28716
rect 24872 28688 24900 28716
rect 25498 28704 25504 28756
rect 25556 28744 25562 28756
rect 25593 28747 25651 28753
rect 25593 28744 25605 28747
rect 25556 28716 25605 28744
rect 25556 28704 25562 28716
rect 25593 28713 25605 28716
rect 25639 28744 25651 28747
rect 30009 28747 30067 28753
rect 30009 28744 30021 28747
rect 25639 28716 30021 28744
rect 25639 28713 25651 28716
rect 25593 28707 25651 28713
rect 30009 28713 30021 28716
rect 30055 28744 30067 28747
rect 30650 28744 30656 28756
rect 30055 28716 30656 28744
rect 30055 28713 30067 28716
rect 30009 28707 30067 28713
rect 30650 28704 30656 28716
rect 30708 28704 30714 28756
rect 32493 28747 32551 28753
rect 32493 28713 32505 28747
rect 32539 28744 32551 28747
rect 32766 28744 32772 28756
rect 32539 28716 32772 28744
rect 32539 28713 32551 28716
rect 32493 28707 32551 28713
rect 32766 28704 32772 28716
rect 32824 28704 32830 28756
rect 33042 28704 33048 28756
rect 33100 28744 33106 28756
rect 33502 28744 33508 28756
rect 33100 28716 33508 28744
rect 33100 28704 33106 28716
rect 33502 28704 33508 28716
rect 33560 28704 33566 28756
rect 34514 28704 34520 28756
rect 34572 28704 34578 28756
rect 34698 28704 34704 28756
rect 34756 28744 34762 28756
rect 35434 28744 35440 28756
rect 34756 28716 35440 28744
rect 34756 28704 34762 28716
rect 35434 28704 35440 28716
rect 35492 28744 35498 28756
rect 36170 28744 36176 28756
rect 35492 28716 36176 28744
rect 35492 28704 35498 28716
rect 36170 28704 36176 28716
rect 36228 28704 36234 28756
rect 36633 28747 36691 28753
rect 36633 28713 36645 28747
rect 36679 28744 36691 28747
rect 37734 28744 37740 28756
rect 36679 28716 37740 28744
rect 36679 28713 36691 28716
rect 36633 28707 36691 28713
rect 37734 28704 37740 28716
rect 37792 28704 37798 28756
rect 17184 28648 18092 28676
rect 17184 28636 17190 28648
rect 14369 28611 14427 28617
rect 14369 28608 14381 28611
rect 10652 28580 11744 28608
rect 12406 28580 14381 28608
rect 10652 28568 10658 28580
rect 10965 28543 11023 28549
rect 10965 28509 10977 28543
rect 11011 28509 11023 28543
rect 10965 28503 11023 28509
rect 11149 28543 11207 28549
rect 11149 28509 11161 28543
rect 11195 28540 11207 28543
rect 11606 28540 11612 28552
rect 11195 28512 11612 28540
rect 11195 28509 11207 28512
rect 11149 28503 11207 28509
rect 10980 28472 11008 28503
rect 11606 28500 11612 28512
rect 11664 28500 11670 28552
rect 11716 28549 11744 28580
rect 14369 28577 14381 28580
rect 14415 28577 14427 28611
rect 16666 28608 16672 28620
rect 14369 28571 14427 28577
rect 16132 28580 16672 28608
rect 11701 28543 11759 28549
rect 11701 28509 11713 28543
rect 11747 28509 11759 28543
rect 11701 28503 11759 28509
rect 11793 28543 11851 28549
rect 11793 28509 11805 28543
rect 11839 28509 11851 28543
rect 11793 28503 11851 28509
rect 11977 28543 12035 28549
rect 11977 28509 11989 28543
rect 12023 28540 12035 28543
rect 12066 28540 12072 28552
rect 12023 28512 12072 28540
rect 12023 28509 12035 28512
rect 11977 28503 12035 28509
rect 11808 28472 11836 28503
rect 12066 28500 12072 28512
rect 12124 28500 12130 28552
rect 12250 28500 12256 28552
rect 12308 28500 12314 28552
rect 12437 28543 12495 28549
rect 12437 28509 12449 28543
rect 12483 28540 12495 28543
rect 12526 28540 12532 28552
rect 12483 28512 12532 28540
rect 12483 28509 12495 28512
rect 12437 28503 12495 28509
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 12710 28500 12716 28552
rect 12768 28500 12774 28552
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28540 12863 28543
rect 13262 28540 13268 28552
rect 12851 28512 13268 28540
rect 12851 28509 12863 28512
rect 12805 28503 12863 28509
rect 13262 28500 13268 28512
rect 13320 28540 13326 28552
rect 13538 28540 13544 28552
rect 13320 28512 13544 28540
rect 13320 28500 13326 28512
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 14090 28500 14096 28552
rect 14148 28500 14154 28552
rect 12986 28472 12992 28484
rect 10980 28444 11744 28472
rect 11808 28444 12992 28472
rect 10962 28404 10968 28416
rect 10244 28376 10968 28404
rect 10045 28367 10103 28373
rect 10962 28364 10968 28376
rect 11020 28404 11026 28416
rect 11057 28407 11115 28413
rect 11057 28404 11069 28407
rect 11020 28376 11069 28404
rect 11020 28364 11026 28376
rect 11057 28373 11069 28376
rect 11103 28373 11115 28407
rect 11057 28367 11115 28373
rect 11333 28407 11391 28413
rect 11333 28373 11345 28407
rect 11379 28404 11391 28407
rect 11514 28404 11520 28416
rect 11379 28376 11520 28404
rect 11379 28373 11391 28376
rect 11333 28367 11391 28373
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 11716 28404 11744 28444
rect 12986 28432 12992 28444
rect 13044 28432 13050 28484
rect 13078 28432 13084 28484
rect 13136 28432 13142 28484
rect 13170 28432 13176 28484
rect 13228 28432 13234 28484
rect 13633 28475 13691 28481
rect 13633 28472 13645 28475
rect 13280 28444 13645 28472
rect 11974 28404 11980 28416
rect 11716 28376 11980 28404
rect 11974 28364 11980 28376
rect 12032 28404 12038 28416
rect 12250 28404 12256 28416
rect 12032 28376 12256 28404
rect 12032 28364 12038 28376
rect 12250 28364 12256 28376
rect 12308 28364 12314 28416
rect 12526 28364 12532 28416
rect 12584 28364 12590 28416
rect 12894 28364 12900 28416
rect 12952 28404 12958 28416
rect 13280 28404 13308 28444
rect 13633 28441 13645 28444
rect 13679 28441 13691 28475
rect 13633 28435 13691 28441
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 14458 28472 14464 28484
rect 13872 28444 14464 28472
rect 13872 28432 13878 28444
rect 14458 28432 14464 28444
rect 14516 28432 14522 28484
rect 15746 28472 15752 28484
rect 15594 28444 15752 28472
rect 12952 28376 13308 28404
rect 12952 28364 12958 28376
rect 13354 28364 13360 28416
rect 13412 28404 13418 28416
rect 13541 28407 13599 28413
rect 13541 28404 13553 28407
rect 13412 28376 13553 28404
rect 13412 28364 13418 28376
rect 13541 28373 13553 28376
rect 13587 28404 13599 28407
rect 13906 28404 13912 28416
rect 13587 28376 13912 28404
rect 13587 28373 13599 28376
rect 13541 28367 13599 28373
rect 13906 28364 13912 28376
rect 13964 28364 13970 28416
rect 15194 28364 15200 28416
rect 15252 28404 15258 28416
rect 15672 28404 15700 28444
rect 15746 28432 15752 28444
rect 15804 28432 15810 28484
rect 15252 28376 15700 28404
rect 15252 28364 15258 28376
rect 15930 28364 15936 28416
rect 15988 28404 15994 28416
rect 16132 28413 16160 28580
rect 16666 28568 16672 28580
rect 16724 28608 16730 28620
rect 18064 28617 18092 28648
rect 18782 28636 18788 28688
rect 18840 28636 18846 28688
rect 24854 28636 24860 28688
rect 24912 28676 24918 28688
rect 24912 28648 26464 28676
rect 24912 28636 24918 28648
rect 18049 28611 18107 28617
rect 16724 28580 17448 28608
rect 16724 28568 16730 28580
rect 16206 28500 16212 28552
rect 16264 28500 16270 28552
rect 17420 28549 17448 28580
rect 18049 28577 18061 28611
rect 18095 28608 18107 28611
rect 18095 28580 18552 28608
rect 18095 28577 18107 28580
rect 18049 28571 18107 28577
rect 17129 28543 17187 28549
rect 17129 28509 17141 28543
rect 17175 28540 17187 28543
rect 17405 28543 17463 28549
rect 17175 28512 17209 28540
rect 17175 28509 17187 28512
rect 17129 28503 17187 28509
rect 17405 28509 17417 28543
rect 17451 28509 17463 28543
rect 17405 28503 17463 28509
rect 16298 28432 16304 28484
rect 16356 28472 16362 28484
rect 17037 28475 17095 28481
rect 17037 28472 17049 28475
rect 16356 28444 17049 28472
rect 16356 28432 16362 28444
rect 17037 28441 17049 28444
rect 17083 28472 17095 28475
rect 17144 28472 17172 28503
rect 17678 28500 17684 28552
rect 17736 28540 17742 28552
rect 17773 28543 17831 28549
rect 17773 28540 17785 28543
rect 17736 28512 17785 28540
rect 17736 28500 17742 28512
rect 17773 28509 17785 28512
rect 17819 28509 17831 28543
rect 17773 28503 17831 28509
rect 18230 28500 18236 28552
rect 18288 28500 18294 28552
rect 18524 28549 18552 28580
rect 18874 28568 18880 28620
rect 18932 28608 18938 28620
rect 19245 28611 19303 28617
rect 19245 28608 19257 28611
rect 18932 28580 19257 28608
rect 18932 28568 18938 28580
rect 19245 28577 19257 28580
rect 19291 28577 19303 28611
rect 19245 28571 19303 28577
rect 22830 28568 22836 28620
rect 22888 28608 22894 28620
rect 24121 28611 24179 28617
rect 24121 28608 24133 28611
rect 22888 28580 24133 28608
rect 22888 28568 22894 28580
rect 24121 28577 24133 28580
rect 24167 28577 24179 28611
rect 24121 28571 24179 28577
rect 18509 28543 18567 28549
rect 18509 28509 18521 28543
rect 18555 28540 18567 28543
rect 18598 28540 18604 28552
rect 18555 28512 18604 28540
rect 18555 28509 18567 28512
rect 18509 28503 18567 28509
rect 18598 28500 18604 28512
rect 18656 28500 18662 28552
rect 18782 28500 18788 28552
rect 18840 28500 18846 28552
rect 21174 28500 21180 28552
rect 21232 28500 21238 28552
rect 21634 28500 21640 28552
rect 21692 28540 21698 28552
rect 21775 28543 21833 28549
rect 21775 28540 21787 28543
rect 21692 28512 21787 28540
rect 21692 28500 21698 28512
rect 21775 28509 21787 28512
rect 21821 28509 21833 28543
rect 21775 28503 21833 28509
rect 21910 28500 21916 28552
rect 21968 28500 21974 28552
rect 22002 28500 22008 28552
rect 22060 28500 22066 28552
rect 22188 28543 22246 28549
rect 22188 28509 22200 28543
rect 22234 28509 22246 28543
rect 22188 28503 22246 28509
rect 22281 28543 22339 28549
rect 22281 28509 22293 28543
rect 22327 28540 22339 28543
rect 22462 28540 22468 28552
rect 22327 28512 22468 28540
rect 22327 28509 22339 28512
rect 22281 28503 22339 28509
rect 17494 28472 17500 28484
rect 17083 28444 17500 28472
rect 17083 28441 17095 28444
rect 17037 28435 17095 28441
rect 17494 28432 17500 28444
rect 17552 28472 17558 28484
rect 18046 28472 18052 28484
rect 17552 28444 18052 28472
rect 17552 28432 17558 28444
rect 18046 28432 18052 28444
rect 18104 28432 18110 28484
rect 19426 28432 19432 28484
rect 19484 28472 19490 28484
rect 19521 28475 19579 28481
rect 19521 28472 19533 28475
rect 19484 28444 19533 28472
rect 19484 28432 19490 28444
rect 19521 28441 19533 28444
rect 19567 28441 19579 28475
rect 19521 28435 19579 28441
rect 19978 28432 19984 28484
rect 20036 28432 20042 28484
rect 21545 28475 21603 28481
rect 21545 28441 21557 28475
rect 21591 28472 21603 28475
rect 22020 28472 22048 28500
rect 21591 28444 22048 28472
rect 22204 28472 22232 28503
rect 22462 28500 22468 28512
rect 22520 28500 22526 28552
rect 24136 28540 24164 28571
rect 25222 28568 25228 28620
rect 25280 28608 25286 28620
rect 25280 28580 26188 28608
rect 25280 28568 25286 28580
rect 24397 28543 24455 28549
rect 24397 28540 24409 28543
rect 24136 28512 24409 28540
rect 24397 28509 24409 28512
rect 24443 28540 24455 28543
rect 24946 28540 24952 28552
rect 24443 28512 24952 28540
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 24946 28500 24952 28512
rect 25004 28500 25010 28552
rect 25314 28500 25320 28552
rect 25372 28500 25378 28552
rect 25409 28543 25467 28549
rect 25409 28509 25421 28543
rect 25455 28509 25467 28543
rect 25409 28503 25467 28509
rect 22204 28444 22324 28472
rect 21591 28441 21603 28444
rect 21545 28435 21603 28441
rect 22296 28416 22324 28444
rect 22554 28432 22560 28484
rect 22612 28472 22618 28484
rect 23845 28475 23903 28481
rect 22612 28444 22678 28472
rect 22612 28432 22618 28444
rect 23845 28441 23857 28475
rect 23891 28472 23903 28475
rect 24762 28472 24768 28484
rect 23891 28444 24768 28472
rect 23891 28441 23903 28444
rect 23845 28435 23903 28441
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 25424 28472 25452 28503
rect 25682 28500 25688 28552
rect 25740 28500 25746 28552
rect 25958 28549 25964 28552
rect 25956 28540 25964 28549
rect 25919 28512 25964 28540
rect 25956 28503 25964 28512
rect 25958 28500 25964 28503
rect 26016 28500 26022 28552
rect 26050 28500 26056 28552
rect 26108 28500 26114 28552
rect 25424 28444 25820 28472
rect 16117 28407 16175 28413
rect 16117 28404 16129 28407
rect 15988 28376 16129 28404
rect 15988 28364 15994 28376
rect 16117 28373 16129 28376
rect 16163 28373 16175 28407
rect 16117 28367 16175 28373
rect 17586 28364 17592 28416
rect 17644 28364 17650 28416
rect 18417 28407 18475 28413
rect 18417 28373 18429 28407
rect 18463 28404 18475 28407
rect 18506 28404 18512 28416
rect 18463 28376 18512 28404
rect 18463 28373 18475 28376
rect 18417 28367 18475 28373
rect 18506 28364 18512 28376
rect 18564 28364 18570 28416
rect 21637 28407 21695 28413
rect 21637 28373 21649 28407
rect 21683 28404 21695 28407
rect 21910 28404 21916 28416
rect 21683 28376 21916 28404
rect 21683 28373 21695 28376
rect 21637 28367 21695 28373
rect 21910 28364 21916 28376
rect 21968 28364 21974 28416
rect 22278 28364 22284 28416
rect 22336 28364 22342 28416
rect 22373 28407 22431 28413
rect 22373 28373 22385 28407
rect 22419 28404 22431 28407
rect 23014 28404 23020 28416
rect 22419 28376 23020 28404
rect 22419 28373 22431 28376
rect 22373 28367 22431 28373
rect 23014 28364 23020 28376
rect 23072 28364 23078 28416
rect 25133 28407 25191 28413
rect 25133 28373 25145 28407
rect 25179 28404 25191 28407
rect 25222 28404 25228 28416
rect 25179 28376 25228 28404
rect 25179 28373 25191 28376
rect 25133 28367 25191 28373
rect 25222 28364 25228 28376
rect 25280 28364 25286 28416
rect 25792 28413 25820 28444
rect 25777 28407 25835 28413
rect 25777 28373 25789 28407
rect 25823 28373 25835 28407
rect 26068 28404 26096 28500
rect 26160 28481 26188 28580
rect 26326 28540 26332 28552
rect 26287 28512 26332 28540
rect 26326 28500 26332 28512
rect 26384 28500 26390 28552
rect 26436 28549 26464 28648
rect 29362 28636 29368 28688
rect 29420 28676 29426 28688
rect 29420 28648 30144 28676
rect 29420 28636 29426 28648
rect 26970 28568 26976 28620
rect 27028 28608 27034 28620
rect 27617 28611 27675 28617
rect 27617 28608 27629 28611
rect 27028 28580 27629 28608
rect 27028 28568 27034 28580
rect 27617 28577 27629 28580
rect 27663 28577 27675 28611
rect 27617 28571 27675 28577
rect 27893 28611 27951 28617
rect 27893 28577 27905 28611
rect 27939 28608 27951 28611
rect 29549 28611 29607 28617
rect 29549 28608 29561 28611
rect 27939 28580 29561 28608
rect 27939 28577 27951 28580
rect 27893 28571 27951 28577
rect 29549 28577 29561 28580
rect 29595 28577 29607 28611
rect 29549 28571 29607 28577
rect 26421 28543 26479 28549
rect 26421 28509 26433 28543
rect 26467 28540 26479 28543
rect 27338 28540 27344 28552
rect 26467 28512 27344 28540
rect 26467 28509 26479 28512
rect 26421 28503 26479 28509
rect 27338 28500 27344 28512
rect 27396 28500 27402 28552
rect 29730 28500 29736 28552
rect 29788 28500 29794 28552
rect 29822 28500 29828 28552
rect 29880 28500 29886 28552
rect 30116 28549 30144 28648
rect 31202 28636 31208 28688
rect 31260 28676 31266 28688
rect 31662 28676 31668 28688
rect 31260 28648 31668 28676
rect 31260 28636 31266 28648
rect 31662 28636 31668 28648
rect 31720 28676 31726 28688
rect 32674 28676 32680 28688
rect 31720 28648 32680 28676
rect 31720 28636 31726 28648
rect 32674 28636 32680 28648
rect 32732 28636 32738 28688
rect 34790 28636 34796 28688
rect 34848 28676 34854 28688
rect 35526 28676 35532 28688
rect 34848 28648 35532 28676
rect 34848 28636 34854 28648
rect 32769 28611 32827 28617
rect 32769 28577 32781 28611
rect 32815 28608 32827 28611
rect 35250 28608 35256 28620
rect 32815 28580 35256 28608
rect 32815 28577 32827 28580
rect 32769 28571 32827 28577
rect 35250 28568 35256 28580
rect 35308 28568 35314 28620
rect 30101 28543 30159 28549
rect 30101 28509 30113 28543
rect 30147 28540 30159 28543
rect 30190 28540 30196 28552
rect 30147 28512 30196 28540
rect 30147 28509 30159 28512
rect 30101 28503 30159 28509
rect 30190 28500 30196 28512
rect 30248 28500 30254 28552
rect 31110 28500 31116 28552
rect 31168 28500 31174 28552
rect 31294 28500 31300 28552
rect 31352 28500 31358 28552
rect 35360 28549 35388 28648
rect 35526 28636 35532 28648
rect 35584 28636 35590 28688
rect 36081 28679 36139 28685
rect 36081 28645 36093 28679
rect 36127 28676 36139 28679
rect 36127 28648 36384 28676
rect 36127 28645 36139 28648
rect 36081 28639 36139 28645
rect 36356 28608 36384 28648
rect 36538 28636 36544 28688
rect 36596 28676 36602 28688
rect 36722 28676 36728 28688
rect 36596 28648 36728 28676
rect 36596 28636 36602 28648
rect 36722 28636 36728 28648
rect 36780 28636 36786 28688
rect 36356 28580 36492 28608
rect 32033 28543 32091 28549
rect 32033 28540 32045 28543
rect 31726 28512 32045 28540
rect 26145 28475 26203 28481
rect 26145 28441 26157 28475
rect 26191 28472 26203 28475
rect 26191 28444 28212 28472
rect 26191 28441 26203 28444
rect 26145 28435 26203 28441
rect 27246 28404 27252 28416
rect 26068 28376 27252 28404
rect 25777 28367 25835 28373
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 27338 28364 27344 28416
rect 27396 28404 27402 28416
rect 28074 28404 28080 28416
rect 27396 28376 28080 28404
rect 27396 28364 27402 28376
rect 28074 28364 28080 28376
rect 28132 28364 28138 28416
rect 28184 28404 28212 28444
rect 28350 28432 28356 28484
rect 28408 28432 28414 28484
rect 29362 28472 29368 28484
rect 29196 28444 29368 28472
rect 29196 28404 29224 28444
rect 29362 28432 29368 28444
rect 29420 28432 29426 28484
rect 29914 28432 29920 28484
rect 29972 28472 29978 28484
rect 31128 28472 31156 28500
rect 31726 28472 31754 28512
rect 32033 28509 32045 28512
rect 32079 28509 32091 28543
rect 34977 28543 35035 28549
rect 34977 28540 34989 28543
rect 32033 28503 32091 28509
rect 34348 28512 34989 28540
rect 29972 28444 31064 28472
rect 31128 28444 31754 28472
rect 29972 28432 29978 28444
rect 31036 28416 31064 28444
rect 32398 28432 32404 28484
rect 32456 28432 32462 28484
rect 33045 28475 33103 28481
rect 33045 28441 33057 28475
rect 33091 28472 33103 28475
rect 33318 28472 33324 28484
rect 33091 28444 33324 28472
rect 33091 28441 33103 28444
rect 33045 28435 33103 28441
rect 33318 28432 33324 28444
rect 33376 28432 33382 28484
rect 34054 28432 34060 28484
rect 34112 28432 34118 28484
rect 28184 28376 29224 28404
rect 29270 28364 29276 28416
rect 29328 28404 29334 28416
rect 30742 28404 30748 28416
rect 29328 28376 30748 28404
rect 29328 28364 29334 28376
rect 30742 28364 30748 28376
rect 30800 28364 30806 28416
rect 31018 28364 31024 28416
rect 31076 28404 31082 28416
rect 31662 28404 31668 28416
rect 31076 28376 31668 28404
rect 31076 28364 31082 28376
rect 31662 28364 31668 28376
rect 31720 28364 31726 28416
rect 33410 28364 33416 28416
rect 33468 28404 33474 28416
rect 34348 28404 34376 28512
rect 34977 28509 34989 28512
rect 35023 28509 35035 28543
rect 34977 28503 35035 28509
rect 35345 28543 35403 28549
rect 35345 28509 35357 28543
rect 35391 28509 35403 28543
rect 35345 28503 35403 28509
rect 35434 28500 35440 28552
rect 35492 28500 35498 28552
rect 35585 28543 35643 28549
rect 35585 28509 35597 28543
rect 35631 28540 35643 28543
rect 35631 28509 35664 28540
rect 35585 28503 35664 28509
rect 35066 28432 35072 28484
rect 35124 28432 35130 28484
rect 35158 28432 35164 28484
rect 35216 28432 35222 28484
rect 33468 28376 34376 28404
rect 34793 28407 34851 28413
rect 33468 28364 33474 28376
rect 34793 28373 34805 28407
rect 34839 28404 34851 28407
rect 35434 28404 35440 28416
rect 34839 28376 35440 28404
rect 34839 28373 34851 28376
rect 34793 28367 34851 28373
rect 35434 28364 35440 28376
rect 35492 28364 35498 28416
rect 35636 28404 35664 28503
rect 35710 28500 35716 28552
rect 35768 28500 35774 28552
rect 35802 28500 35808 28552
rect 35860 28500 35866 28552
rect 35943 28543 36001 28549
rect 35943 28509 35955 28543
rect 35989 28540 36001 28543
rect 35989 28512 36313 28540
rect 35989 28509 36001 28512
rect 35943 28503 36001 28509
rect 35986 28404 35992 28416
rect 35636 28376 35992 28404
rect 35986 28364 35992 28376
rect 36044 28364 36050 28416
rect 36170 28364 36176 28416
rect 36228 28364 36234 28416
rect 36285 28404 36313 28512
rect 36354 28500 36360 28552
rect 36412 28500 36418 28552
rect 36464 28549 36492 28580
rect 37366 28568 37372 28620
rect 37424 28568 37430 28620
rect 37642 28568 37648 28620
rect 37700 28568 37706 28620
rect 38838 28568 38844 28620
rect 38896 28608 38902 28620
rect 39114 28608 39120 28620
rect 38896 28580 39120 28608
rect 38896 28568 38902 28580
rect 39114 28568 39120 28580
rect 39172 28568 39178 28620
rect 36449 28543 36507 28549
rect 36449 28509 36461 28543
rect 36495 28509 36507 28543
rect 36449 28503 36507 28509
rect 36725 28543 36783 28549
rect 36725 28509 36737 28543
rect 36771 28540 36783 28543
rect 36998 28540 37004 28552
rect 36771 28512 37004 28540
rect 36771 28509 36783 28512
rect 36725 28503 36783 28509
rect 36998 28500 37004 28512
rect 37056 28500 37062 28552
rect 41414 28540 41420 28552
rect 39592 28512 41420 28540
rect 39592 28484 39620 28512
rect 41414 28500 41420 28512
rect 41472 28500 41478 28552
rect 41509 28543 41567 28549
rect 41509 28509 41521 28543
rect 41555 28509 41567 28543
rect 41509 28503 41567 28509
rect 38930 28472 38936 28484
rect 38870 28444 38936 28472
rect 38930 28432 38936 28444
rect 38988 28472 38994 28484
rect 39574 28472 39580 28484
rect 38988 28444 39580 28472
rect 38988 28432 38994 28444
rect 39574 28432 39580 28444
rect 39632 28432 39638 28484
rect 39850 28432 39856 28484
rect 39908 28472 39914 28484
rect 40313 28475 40371 28481
rect 40313 28472 40325 28475
rect 39908 28444 40325 28472
rect 39908 28432 39914 28444
rect 40313 28441 40325 28444
rect 40359 28441 40371 28475
rect 40313 28435 40371 28441
rect 40494 28432 40500 28484
rect 40552 28432 40558 28484
rect 41524 28472 41552 28503
rect 41874 28500 41880 28552
rect 41932 28500 41938 28552
rect 40604 28444 42564 28472
rect 36354 28404 36360 28416
rect 36285 28376 36360 28404
rect 36354 28364 36360 28376
rect 36412 28404 36418 28416
rect 36722 28404 36728 28416
rect 36412 28376 36728 28404
rect 36412 28364 36418 28376
rect 36722 28364 36728 28376
rect 36780 28404 36786 28416
rect 37734 28404 37740 28416
rect 36780 28376 37740 28404
rect 36780 28364 36786 28376
rect 37734 28364 37740 28376
rect 37792 28364 37798 28416
rect 39114 28364 39120 28416
rect 39172 28364 39178 28416
rect 39758 28364 39764 28416
rect 39816 28404 39822 28416
rect 40604 28404 40632 28444
rect 39816 28376 40632 28404
rect 39816 28364 39822 28376
rect 40678 28364 40684 28416
rect 40736 28364 40742 28416
rect 41690 28364 41696 28416
rect 41748 28364 41754 28416
rect 42058 28364 42064 28416
rect 42116 28364 42122 28416
rect 1104 28314 42504 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 42504 28314
rect 1104 28240 42504 28262
rect 3970 28160 3976 28212
rect 4028 28200 4034 28212
rect 4338 28200 4344 28212
rect 4028 28172 4344 28200
rect 4028 28160 4034 28172
rect 4338 28160 4344 28172
rect 4396 28200 4402 28212
rect 5350 28200 5356 28212
rect 4396 28172 5356 28200
rect 4396 28160 4402 28172
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 5534 28160 5540 28212
rect 5592 28160 5598 28212
rect 8478 28160 8484 28212
rect 8536 28160 8542 28212
rect 8662 28160 8668 28212
rect 8720 28160 8726 28212
rect 9398 28160 9404 28212
rect 9456 28160 9462 28212
rect 11606 28160 11612 28212
rect 11664 28200 11670 28212
rect 11885 28203 11943 28209
rect 11885 28200 11897 28203
rect 11664 28172 11897 28200
rect 11664 28160 11670 28172
rect 11885 28169 11897 28172
rect 11931 28169 11943 28203
rect 12526 28200 12532 28212
rect 11885 28163 11943 28169
rect 12268 28172 12532 28200
rect 3050 28092 3056 28144
rect 3108 28132 3114 28144
rect 5442 28132 5448 28144
rect 3108 28104 5448 28132
rect 3108 28092 3114 28104
rect 3878 28024 3884 28076
rect 3936 28064 3942 28076
rect 4433 28067 4491 28073
rect 4433 28064 4445 28067
rect 3936 28036 4445 28064
rect 3936 28024 3942 28036
rect 4433 28033 4445 28036
rect 4479 28033 4491 28067
rect 4433 28027 4491 28033
rect 4540 27869 4568 28104
rect 5442 28092 5448 28104
rect 5500 28132 5506 28144
rect 5626 28132 5632 28144
rect 5500 28104 5632 28132
rect 5500 28092 5506 28104
rect 5626 28092 5632 28104
rect 5684 28092 5690 28144
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28064 4675 28067
rect 5997 28067 6055 28073
rect 5997 28064 6009 28067
rect 4663 28036 6009 28064
rect 4663 28033 4675 28036
rect 4617 28027 4675 28033
rect 5997 28033 6009 28036
rect 6043 28064 6055 28067
rect 6457 28067 6515 28073
rect 6457 28064 6469 28067
rect 6043 28036 6469 28064
rect 6043 28033 6055 28036
rect 5997 28027 6055 28033
rect 6457 28033 6469 28036
rect 6503 28033 6515 28067
rect 6457 28027 6515 28033
rect 6549 28067 6607 28073
rect 6549 28033 6561 28067
rect 6595 28064 6607 28067
rect 7098 28064 7104 28076
rect 6595 28036 7104 28064
rect 6595 28033 6607 28036
rect 6549 28027 6607 28033
rect 7098 28024 7104 28036
rect 7156 28024 7162 28076
rect 9309 28067 9367 28073
rect 9309 28033 9321 28067
rect 9355 28064 9367 28067
rect 9674 28064 9680 28076
rect 9355 28036 9680 28064
rect 9355 28033 9367 28036
rect 9309 28027 9367 28033
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 11974 28024 11980 28076
rect 12032 28024 12038 28076
rect 12066 28024 12072 28076
rect 12124 28024 12130 28076
rect 4890 27956 4896 28008
rect 4948 27956 4954 28008
rect 5258 27956 5264 28008
rect 5316 27956 5322 28008
rect 5353 27999 5411 28005
rect 5353 27965 5365 27999
rect 5399 27965 5411 27999
rect 5353 27959 5411 27965
rect 5166 27888 5172 27940
rect 5224 27928 5230 27940
rect 5368 27928 5396 27959
rect 5718 27956 5724 28008
rect 5776 27996 5782 28008
rect 5905 27999 5963 28005
rect 5905 27996 5917 27999
rect 5776 27968 5917 27996
rect 5776 27956 5782 27968
rect 5905 27965 5917 27968
rect 5951 27965 5963 27999
rect 5905 27959 5963 27965
rect 8021 27999 8079 28005
rect 8021 27965 8033 27999
rect 8067 27996 8079 27999
rect 8110 27996 8116 28008
rect 8067 27968 8116 27996
rect 8067 27965 8079 27968
rect 8021 27959 8079 27965
rect 8110 27956 8116 27968
rect 8168 27996 8174 28008
rect 9861 27999 9919 28005
rect 9861 27996 9873 27999
rect 8168 27968 9873 27996
rect 8168 27956 8174 27968
rect 9861 27965 9873 27968
rect 9907 27996 9919 27999
rect 10134 27996 10140 28008
rect 9907 27968 10140 27996
rect 9907 27965 9919 27968
rect 9861 27959 9919 27965
rect 10134 27956 10140 27968
rect 10192 27956 10198 28008
rect 12268 27996 12296 28172
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 12802 28160 12808 28212
rect 12860 28160 12866 28212
rect 12986 28160 12992 28212
rect 13044 28200 13050 28212
rect 13541 28203 13599 28209
rect 13541 28200 13553 28203
rect 13044 28172 13553 28200
rect 13044 28160 13050 28172
rect 13541 28169 13553 28172
rect 13587 28169 13599 28203
rect 15289 28203 15347 28209
rect 15289 28200 15301 28203
rect 13541 28163 13599 28169
rect 15120 28172 15301 28200
rect 12342 28092 12348 28144
rect 12400 28132 12406 28144
rect 12400 28104 12664 28132
rect 12400 28092 12406 28104
rect 12547 28067 12605 28073
rect 12547 28033 12559 28067
rect 12593 28064 12605 28067
rect 12636 28064 12664 28104
rect 12894 28092 12900 28144
rect 12952 28132 12958 28144
rect 13081 28135 13139 28141
rect 13081 28132 13093 28135
rect 12952 28104 13093 28132
rect 12952 28092 12958 28104
rect 13081 28101 13093 28104
rect 13127 28101 13139 28135
rect 13081 28095 13139 28101
rect 13371 28104 13584 28132
rect 12986 28073 12992 28076
rect 12984 28064 12992 28073
rect 12593 28036 12664 28064
rect 12947 28036 12992 28064
rect 12593 28033 12605 28036
rect 12547 28027 12605 28033
rect 12984 28027 12992 28036
rect 12986 28024 12992 28027
rect 13044 28024 13050 28076
rect 13170 28024 13176 28076
rect 13228 28024 13234 28076
rect 13371 28073 13399 28104
rect 13556 28076 13584 28104
rect 14292 28104 14688 28132
rect 13356 28067 13414 28073
rect 13356 28033 13368 28067
rect 13402 28033 13414 28067
rect 13356 28027 13414 28033
rect 13449 28067 13507 28073
rect 13449 28033 13461 28067
rect 13495 28033 13507 28067
rect 13449 28027 13507 28033
rect 12345 27999 12403 28005
rect 12345 27996 12357 27999
rect 12268 27968 12357 27996
rect 12345 27965 12357 27968
rect 12391 27965 12403 27999
rect 13464 27996 13492 28027
rect 13538 28024 13544 28076
rect 13596 28024 13602 28076
rect 13630 28024 13636 28076
rect 13688 28064 13694 28076
rect 13725 28067 13783 28073
rect 13725 28064 13737 28067
rect 13688 28036 13737 28064
rect 13688 28024 13694 28036
rect 13725 28033 13737 28036
rect 13771 28033 13783 28067
rect 13725 28027 13783 28033
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28064 13875 28067
rect 13906 28064 13912 28076
rect 13863 28036 13912 28064
rect 13863 28033 13875 28036
rect 13817 28027 13875 28033
rect 13906 28024 13912 28036
rect 13964 28024 13970 28076
rect 13998 28024 14004 28076
rect 14056 28024 14062 28076
rect 14292 28073 14320 28104
rect 14277 28067 14335 28073
rect 14277 28033 14289 28067
rect 14323 28033 14335 28067
rect 14277 28027 14335 28033
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28064 14519 28067
rect 14550 28064 14556 28076
rect 14507 28036 14556 28064
rect 14507 28033 14519 28036
rect 14461 28027 14519 28033
rect 14550 28024 14556 28036
rect 14608 28024 14614 28076
rect 14660 28073 14688 28104
rect 14918 28092 14924 28144
rect 14976 28092 14982 28144
rect 15120 28141 15148 28172
rect 15289 28169 15301 28172
rect 15335 28200 15347 28203
rect 16482 28200 16488 28212
rect 15335 28172 16488 28200
rect 15335 28169 15347 28172
rect 15289 28163 15347 28169
rect 16482 28160 16488 28172
rect 16540 28160 16546 28212
rect 16574 28160 16580 28212
rect 16632 28200 16638 28212
rect 16669 28203 16727 28209
rect 16669 28200 16681 28203
rect 16632 28172 16681 28200
rect 16632 28160 16638 28172
rect 16669 28169 16681 28172
rect 16715 28169 16727 28203
rect 18417 28203 18475 28209
rect 16669 28163 16727 28169
rect 17236 28172 18368 28200
rect 15105 28135 15163 28141
rect 15105 28101 15117 28135
rect 15151 28101 15163 28135
rect 15105 28095 15163 28101
rect 15657 28135 15715 28141
rect 15657 28101 15669 28135
rect 15703 28132 15715 28135
rect 15838 28132 15844 28144
rect 15703 28104 15844 28132
rect 15703 28101 15715 28104
rect 15657 28095 15715 28101
rect 15838 28092 15844 28104
rect 15896 28092 15902 28144
rect 15930 28092 15936 28144
rect 15988 28132 15994 28144
rect 16853 28135 16911 28141
rect 16853 28132 16865 28135
rect 15988 28104 16865 28132
rect 15988 28092 15994 28104
rect 16853 28101 16865 28104
rect 16899 28101 16911 28135
rect 17236 28132 17264 28172
rect 16853 28095 16911 28101
rect 16960 28104 17264 28132
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28064 14703 28067
rect 14737 28067 14795 28073
rect 14737 28064 14749 28067
rect 14691 28036 14749 28064
rect 14691 28033 14703 28036
rect 14645 28027 14703 28033
rect 14737 28033 14749 28036
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 15194 28024 15200 28076
rect 15252 28024 15258 28076
rect 15473 28067 15531 28073
rect 15473 28033 15485 28067
rect 15519 28064 15531 28067
rect 16114 28064 16120 28076
rect 15519 28036 16120 28064
rect 15519 28033 15531 28036
rect 15473 28027 15531 28033
rect 14366 27996 14372 28008
rect 12345 27959 12403 27965
rect 12544 27968 14372 27996
rect 5629 27931 5687 27937
rect 5629 27928 5641 27931
rect 5224 27900 5641 27928
rect 5224 27888 5230 27900
rect 5629 27897 5641 27900
rect 5675 27897 5687 27931
rect 5629 27891 5687 27897
rect 8389 27931 8447 27937
rect 8389 27897 8401 27931
rect 8435 27897 8447 27931
rect 8389 27891 8447 27897
rect 9585 27931 9643 27937
rect 9585 27897 9597 27931
rect 9631 27928 9643 27931
rect 10042 27928 10048 27940
rect 9631 27900 10048 27928
rect 9631 27897 9643 27900
rect 9585 27891 9643 27897
rect 4525 27863 4583 27869
rect 4525 27829 4537 27863
rect 4571 27829 4583 27863
rect 4525 27823 4583 27829
rect 4801 27863 4859 27869
rect 4801 27829 4813 27863
rect 4847 27860 4859 27863
rect 5258 27860 5264 27872
rect 4847 27832 5264 27860
rect 4847 27829 4859 27832
rect 4801 27823 4859 27829
rect 5258 27820 5264 27832
rect 5316 27820 5322 27872
rect 8404 27860 8432 27891
rect 10042 27888 10048 27900
rect 10100 27928 10106 27940
rect 10686 27928 10692 27940
rect 10100 27900 10692 27928
rect 10100 27888 10106 27900
rect 10686 27888 10692 27900
rect 10744 27888 10750 27940
rect 10502 27860 10508 27872
rect 8404 27832 10508 27860
rect 10502 27820 10508 27832
rect 10560 27820 10566 27872
rect 12544 27869 12572 27968
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 15488 27996 15516 28027
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 16298 28024 16304 28076
rect 16356 28024 16362 28076
rect 16960 28064 16988 28104
rect 16408 28036 16988 28064
rect 17037 28067 17095 28073
rect 14660 27968 15516 27996
rect 16025 27999 16083 28005
rect 12710 27888 12716 27940
rect 12768 27888 12774 27940
rect 14660 27872 14688 27968
rect 16025 27965 16037 27999
rect 16071 27965 16083 27999
rect 16025 27959 16083 27965
rect 16040 27928 16068 27959
rect 16206 27956 16212 28008
rect 16264 27996 16270 28008
rect 16408 27996 16436 28036
rect 17037 28033 17049 28067
rect 17083 28064 17095 28067
rect 17126 28064 17132 28076
rect 17083 28036 17132 28064
rect 17083 28033 17095 28036
rect 17037 28027 17095 28033
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 17236 28073 17264 28104
rect 17313 28135 17371 28141
rect 17313 28101 17325 28135
rect 17359 28132 17371 28135
rect 18230 28132 18236 28144
rect 17359 28104 18236 28132
rect 17359 28101 17371 28104
rect 17313 28095 17371 28101
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28033 17279 28067
rect 17221 28027 17279 28033
rect 17402 28024 17408 28076
rect 17460 28024 17466 28076
rect 17512 28073 17540 28104
rect 18230 28092 18236 28104
rect 18288 28092 18294 28144
rect 17497 28067 17555 28073
rect 17497 28033 17509 28067
rect 17543 28033 17555 28067
rect 17497 28027 17555 28033
rect 17678 28024 17684 28076
rect 17736 28024 17742 28076
rect 17773 28067 17831 28073
rect 17773 28033 17785 28067
rect 17819 28033 17831 28067
rect 17773 28027 17831 28033
rect 17957 28067 18015 28073
rect 17957 28033 17969 28067
rect 18003 28033 18015 28067
rect 17957 28027 18015 28033
rect 16264 27968 16436 27996
rect 16264 27956 16270 27968
rect 16482 27956 16488 28008
rect 16540 27996 16546 28008
rect 17589 27999 17647 28005
rect 17589 27996 17601 27999
rect 16540 27968 17601 27996
rect 16540 27956 16546 27968
rect 17589 27965 17601 27968
rect 17635 27996 17647 27999
rect 17788 27996 17816 28027
rect 17635 27968 17816 27996
rect 17635 27965 17647 27968
rect 17589 27959 17647 27965
rect 16298 27928 16304 27940
rect 16040 27900 16304 27928
rect 16298 27888 16304 27900
rect 16356 27928 16362 27940
rect 16758 27928 16764 27940
rect 16356 27900 16764 27928
rect 16356 27888 16362 27900
rect 16758 27888 16764 27900
rect 16816 27888 16822 27940
rect 17972 27928 18000 28027
rect 18046 28024 18052 28076
rect 18104 28024 18110 28076
rect 18141 28067 18199 28073
rect 18141 28033 18153 28067
rect 18187 28064 18199 28067
rect 18340 28064 18368 28172
rect 18417 28169 18429 28203
rect 18463 28169 18475 28203
rect 18417 28163 18475 28169
rect 18432 28132 18460 28163
rect 19426 28160 19432 28212
rect 19484 28160 19490 28212
rect 22830 28200 22836 28212
rect 22066 28172 22836 28200
rect 18782 28132 18788 28144
rect 18432 28104 18788 28132
rect 18782 28092 18788 28104
rect 18840 28132 18846 28144
rect 19337 28135 19395 28141
rect 18840 28104 19196 28132
rect 18840 28092 18846 28104
rect 18187 28036 18368 28064
rect 18187 28033 18199 28036
rect 18141 28027 18199 28033
rect 18598 28024 18604 28076
rect 18656 28024 18662 28076
rect 19168 28073 19196 28104
rect 19337 28101 19349 28135
rect 19383 28132 19395 28135
rect 20806 28132 20812 28144
rect 19383 28104 20812 28132
rect 19383 28101 19395 28104
rect 19337 28095 19395 28101
rect 20806 28092 20812 28104
rect 20864 28092 20870 28144
rect 22066 28132 22094 28172
rect 22830 28160 22836 28172
rect 22888 28160 22894 28212
rect 23382 28160 23388 28212
rect 23440 28200 23446 28212
rect 23569 28203 23627 28209
rect 23569 28200 23581 28203
rect 23440 28172 23581 28200
rect 23440 28160 23446 28172
rect 23569 28169 23581 28172
rect 23615 28169 23627 28203
rect 23569 28163 23627 28169
rect 24762 28160 24768 28212
rect 24820 28160 24826 28212
rect 25130 28160 25136 28212
rect 25188 28200 25194 28212
rect 25188 28172 25360 28200
rect 25188 28160 25194 28172
rect 21836 28104 22094 28132
rect 19061 28067 19119 28073
rect 19061 28033 19073 28067
rect 19107 28033 19119 28067
rect 19061 28027 19119 28033
rect 19153 28067 19211 28073
rect 19153 28033 19165 28067
rect 19199 28064 19211 28067
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 19199 28036 19625 28064
rect 19199 28033 19211 28036
rect 19153 28027 19211 28033
rect 19613 28033 19625 28036
rect 19659 28033 19671 28067
rect 19613 28027 19671 28033
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28064 19763 28067
rect 20349 28067 20407 28073
rect 20349 28064 20361 28067
rect 19751 28036 20361 28064
rect 19751 28033 19763 28036
rect 19705 28027 19763 28033
rect 20349 28033 20361 28036
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 18693 27999 18751 28005
rect 18693 27996 18705 27999
rect 18248 27968 18705 27996
rect 18248 27940 18276 27968
rect 18693 27965 18705 27968
rect 18739 27996 18751 27999
rect 19076 27996 19104 28027
rect 20990 28024 20996 28076
rect 21048 28024 21054 28076
rect 19797 27999 19855 28005
rect 19797 27996 19809 27999
rect 18739 27968 19809 27996
rect 18739 27965 18751 27968
rect 18693 27959 18751 27965
rect 19797 27965 19809 27968
rect 19843 27965 19855 27999
rect 19797 27959 19855 27965
rect 19889 27999 19947 28005
rect 19889 27965 19901 27999
rect 19935 27965 19947 27999
rect 19889 27959 19947 27965
rect 18230 27928 18236 27940
rect 17604 27900 17908 27928
rect 17972 27900 18236 27928
rect 12529 27863 12587 27869
rect 12529 27829 12541 27863
rect 12575 27829 12587 27863
rect 12529 27823 12587 27829
rect 13906 27820 13912 27872
rect 13964 27860 13970 27872
rect 14001 27863 14059 27869
rect 14001 27860 14013 27863
rect 13964 27832 14013 27860
rect 13964 27820 13970 27832
rect 14001 27829 14013 27832
rect 14047 27860 14059 27863
rect 14185 27863 14243 27869
rect 14185 27860 14197 27863
rect 14047 27832 14197 27860
rect 14047 27829 14059 27832
rect 14001 27823 14059 27829
rect 14185 27829 14197 27832
rect 14231 27829 14243 27863
rect 14185 27823 14243 27829
rect 14642 27820 14648 27872
rect 14700 27820 14706 27872
rect 15746 27820 15752 27872
rect 15804 27820 15810 27872
rect 15838 27820 15844 27872
rect 15896 27860 15902 27872
rect 15933 27863 15991 27869
rect 15933 27860 15945 27863
rect 15896 27832 15945 27860
rect 15896 27820 15902 27832
rect 15933 27829 15945 27832
rect 15979 27829 15991 27863
rect 16776 27860 16804 27888
rect 17604 27872 17632 27900
rect 17586 27860 17592 27872
rect 16776 27832 17592 27860
rect 15933 27823 15991 27829
rect 17586 27820 17592 27832
rect 17644 27820 17650 27872
rect 17770 27820 17776 27872
rect 17828 27820 17834 27872
rect 17880 27860 17908 27900
rect 18230 27888 18236 27900
rect 18288 27888 18294 27940
rect 18049 27863 18107 27869
rect 18049 27860 18061 27863
rect 17880 27832 18061 27860
rect 18049 27829 18061 27832
rect 18095 27829 18107 27863
rect 18049 27823 18107 27829
rect 18506 27820 18512 27872
rect 18564 27860 18570 27872
rect 19242 27860 19248 27872
rect 18564 27832 19248 27860
rect 18564 27820 18570 27832
rect 19242 27820 19248 27832
rect 19300 27860 19306 27872
rect 19904 27860 19932 27959
rect 21358 27956 21364 28008
rect 21416 27996 21422 28008
rect 21836 28005 21864 28104
rect 23842 28092 23848 28144
rect 23900 28132 23906 28144
rect 23900 28104 24348 28132
rect 23900 28092 23906 28104
rect 24118 28064 24124 28076
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21416 27968 21833 27996
rect 21416 27956 21422 27968
rect 21821 27965 21833 27968
rect 21867 27965 21879 27999
rect 21821 27959 21879 27965
rect 22094 27956 22100 28008
rect 22152 27956 22158 28008
rect 22554 27956 22560 28008
rect 22612 27996 22618 28008
rect 22830 27996 22836 28008
rect 22612 27968 22836 27996
rect 22612 27956 22618 27968
rect 22830 27956 22836 27968
rect 22888 27996 22894 28008
rect 23216 27996 23244 28050
rect 22888 27968 23244 27996
rect 23492 28036 24124 28064
rect 22888 27956 22894 27968
rect 23492 27860 23520 28036
rect 24118 28024 24124 28036
rect 24176 28024 24182 28076
rect 24320 28073 24348 28104
rect 24394 28092 24400 28144
rect 24452 28092 24458 28144
rect 24578 28092 24584 28144
rect 24636 28092 24642 28144
rect 25222 28092 25228 28144
rect 25280 28092 25286 28144
rect 25332 28132 25360 28172
rect 25590 28160 25596 28212
rect 25648 28200 25654 28212
rect 26050 28200 26056 28212
rect 25648 28172 26056 28200
rect 25648 28160 25654 28172
rect 26050 28160 26056 28172
rect 26108 28200 26114 28212
rect 26697 28203 26755 28209
rect 26697 28200 26709 28203
rect 26108 28172 26709 28200
rect 26108 28160 26114 28172
rect 26697 28169 26709 28172
rect 26743 28169 26755 28203
rect 28350 28200 28356 28212
rect 26697 28163 26755 28169
rect 27540 28172 28356 28200
rect 25682 28132 25688 28144
rect 25332 28104 25688 28132
rect 25682 28092 25688 28104
rect 25740 28092 25746 28144
rect 24305 28067 24363 28073
rect 24305 28033 24317 28067
rect 24351 28064 24363 28067
rect 24762 28064 24768 28076
rect 24351 28036 24768 28064
rect 24351 28033 24363 28036
rect 24305 28027 24363 28033
rect 24762 28024 24768 28036
rect 24820 28024 24826 28076
rect 24946 28024 24952 28076
rect 25004 28024 25010 28076
rect 27540 28064 27568 28172
rect 28350 28160 28356 28172
rect 28408 28160 28414 28212
rect 28902 28160 28908 28212
rect 28960 28160 28966 28212
rect 29362 28200 29368 28212
rect 29196 28172 29368 28200
rect 27709 28135 27767 28141
rect 27709 28101 27721 28135
rect 27755 28132 27767 28135
rect 28920 28132 28948 28160
rect 29196 28141 29224 28172
rect 29362 28160 29368 28172
rect 29420 28160 29426 28212
rect 29549 28203 29607 28209
rect 29549 28169 29561 28203
rect 29595 28200 29607 28203
rect 29822 28200 29828 28212
rect 29595 28172 29828 28200
rect 29595 28169 29607 28172
rect 29549 28163 29607 28169
rect 29822 28160 29828 28172
rect 29880 28160 29886 28212
rect 31110 28200 31116 28212
rect 30024 28172 31116 28200
rect 27755 28104 28948 28132
rect 29181 28135 29239 28141
rect 27755 28101 27767 28104
rect 27709 28095 27767 28101
rect 29181 28101 29193 28135
rect 29227 28101 29239 28135
rect 29181 28095 29239 28101
rect 29270 28092 29276 28144
rect 29328 28092 29334 28144
rect 29638 28092 29644 28144
rect 29696 28132 29702 28144
rect 29733 28135 29791 28141
rect 29733 28132 29745 28135
rect 29696 28104 29745 28132
rect 29696 28092 29702 28104
rect 29733 28101 29745 28104
rect 29779 28101 29791 28135
rect 29733 28095 29791 28101
rect 29914 28092 29920 28144
rect 29972 28092 29978 28144
rect 26252 28036 27568 28064
rect 25682 27956 25688 28008
rect 25740 27996 25746 28008
rect 26252 27996 26280 28036
rect 27614 28024 27620 28076
rect 27672 28024 27678 28076
rect 27798 28024 27804 28076
rect 27856 28024 27862 28076
rect 27985 28067 28043 28073
rect 27985 28033 27997 28067
rect 28031 28033 28043 28067
rect 27985 28027 28043 28033
rect 28000 27996 28028 28027
rect 28074 28024 28080 28076
rect 28132 28064 28138 28076
rect 28810 28064 28816 28076
rect 28132 28036 28816 28064
rect 28132 28024 28138 28036
rect 28810 28024 28816 28036
rect 28868 28064 28874 28076
rect 28905 28067 28963 28073
rect 28905 28064 28917 28067
rect 28868 28036 28917 28064
rect 28868 28024 28874 28036
rect 28905 28033 28917 28036
rect 28951 28033 28963 28067
rect 28905 28027 28963 28033
rect 29053 28067 29111 28073
rect 29053 28033 29065 28067
rect 29099 28064 29111 28067
rect 29411 28067 29469 28073
rect 29099 28036 29316 28064
rect 29099 28033 29111 28036
rect 29053 28027 29111 28033
rect 29288 28008 29316 28036
rect 29411 28033 29423 28067
rect 29457 28064 29469 28067
rect 29932 28064 29960 28092
rect 29457 28036 29960 28064
rect 29457 28033 29469 28036
rect 29411 28027 29469 28033
rect 25740 27968 26280 27996
rect 26344 27968 28028 27996
rect 25740 27956 25746 27968
rect 26344 27940 26372 27968
rect 29270 27956 29276 28008
rect 29328 27956 29334 28008
rect 30024 27996 30052 28172
rect 31110 28160 31116 28172
rect 31168 28160 31174 28212
rect 31294 28160 31300 28212
rect 31352 28200 31358 28212
rect 34514 28200 34520 28212
rect 31352 28172 34520 28200
rect 31352 28160 31358 28172
rect 34514 28160 34520 28172
rect 34572 28160 34578 28212
rect 34790 28160 34796 28212
rect 34848 28200 34854 28212
rect 35342 28200 35348 28212
rect 34848 28172 35348 28200
rect 34848 28160 34854 28172
rect 35342 28160 35348 28172
rect 35400 28160 35406 28212
rect 36170 28200 36176 28212
rect 35544 28172 36176 28200
rect 30098 28092 30104 28144
rect 30156 28132 30162 28144
rect 30926 28132 30932 28144
rect 30156 28104 30932 28132
rect 30156 28092 30162 28104
rect 30926 28092 30932 28104
rect 30984 28092 30990 28144
rect 32493 28135 32551 28141
rect 32493 28101 32505 28135
rect 32539 28132 32551 28135
rect 32582 28132 32588 28144
rect 32539 28104 32588 28132
rect 32539 28101 32551 28104
rect 32493 28095 32551 28101
rect 31938 28024 31944 28076
rect 31996 28064 32002 28076
rect 32508 28064 32536 28095
rect 32582 28092 32588 28104
rect 32640 28092 32646 28144
rect 32674 28092 32680 28144
rect 32732 28132 32738 28144
rect 33689 28135 33747 28141
rect 32732 28104 33456 28132
rect 32732 28092 32738 28104
rect 31996 28036 32536 28064
rect 31996 28024 32002 28036
rect 32766 28024 32772 28076
rect 32824 28024 32830 28076
rect 32953 28067 33011 28073
rect 32953 28033 32965 28067
rect 32999 28033 33011 28067
rect 32953 28027 33011 28033
rect 30193 27999 30251 28005
rect 30193 27996 30205 27999
rect 30024 27968 30205 27996
rect 30193 27965 30205 27968
rect 30239 27965 30251 27999
rect 30193 27959 30251 27965
rect 30466 27956 30472 28008
rect 30524 27956 30530 28008
rect 30926 27956 30932 28008
rect 30984 27996 30990 28008
rect 30984 27968 31523 27996
rect 30984 27956 30990 27968
rect 24302 27888 24308 27940
rect 24360 27888 24366 27940
rect 26326 27888 26332 27940
rect 26384 27888 26390 27940
rect 27798 27888 27804 27940
rect 27856 27928 27862 27940
rect 27982 27928 27988 27940
rect 27856 27900 27988 27928
rect 27856 27888 27862 27900
rect 27982 27888 27988 27900
rect 28040 27888 28046 27940
rect 28350 27888 28356 27940
rect 28408 27928 28414 27940
rect 30098 27928 30104 27940
rect 28408 27900 30104 27928
rect 28408 27888 28414 27900
rect 30098 27888 30104 27900
rect 30156 27888 30162 27940
rect 31495 27928 31523 27968
rect 31662 27956 31668 28008
rect 31720 27996 31726 28008
rect 32968 27996 32996 28027
rect 33042 28024 33048 28076
rect 33100 28024 33106 28076
rect 33137 28067 33195 28073
rect 33137 28033 33149 28067
rect 33183 28064 33195 28067
rect 33318 28064 33324 28076
rect 33183 28036 33324 28064
rect 33183 28033 33195 28036
rect 33137 28027 33195 28033
rect 33318 28024 33324 28036
rect 33376 28024 33382 28076
rect 33428 28073 33456 28104
rect 33689 28101 33701 28135
rect 33735 28132 33747 28135
rect 34422 28132 34428 28144
rect 33735 28104 34428 28132
rect 33735 28101 33747 28104
rect 33689 28095 33747 28101
rect 34422 28092 34428 28104
rect 34480 28092 34486 28144
rect 35544 28141 35572 28172
rect 36170 28160 36176 28172
rect 36228 28160 36234 28212
rect 36262 28160 36268 28212
rect 36320 28200 36326 28212
rect 36320 28172 37320 28200
rect 36320 28160 36326 28172
rect 35529 28135 35587 28141
rect 35529 28101 35541 28135
rect 35575 28101 35587 28135
rect 35529 28095 35587 28101
rect 33413 28067 33471 28073
rect 33413 28033 33425 28067
rect 33459 28033 33471 28067
rect 33413 28027 33471 28033
rect 33502 28024 33508 28076
rect 33560 28064 33566 28076
rect 33560 28036 33605 28064
rect 33560 28024 33566 28036
rect 33778 28024 33784 28076
rect 33836 28024 33842 28076
rect 33962 28073 33968 28076
rect 33919 28067 33968 28073
rect 33919 28033 33931 28067
rect 33965 28033 33968 28067
rect 33919 28027 33968 28033
rect 33962 28024 33968 28027
rect 34020 28024 34026 28076
rect 34330 28024 34336 28076
rect 34388 28024 34394 28076
rect 35250 28024 35256 28076
rect 35308 28024 35314 28076
rect 36630 28024 36636 28076
rect 36688 28024 36694 28076
rect 37292 28073 37320 28172
rect 37458 28160 37464 28212
rect 37516 28160 37522 28212
rect 37550 28160 37556 28212
rect 37608 28200 37614 28212
rect 37921 28203 37979 28209
rect 37921 28200 37933 28203
rect 37608 28172 37933 28200
rect 37608 28160 37614 28172
rect 37921 28169 37933 28172
rect 37967 28169 37979 28203
rect 37921 28163 37979 28169
rect 40313 28203 40371 28209
rect 40313 28169 40325 28203
rect 40359 28200 40371 28203
rect 40494 28200 40500 28212
rect 40359 28172 40500 28200
rect 40359 28169 40371 28172
rect 40313 28163 40371 28169
rect 40494 28160 40500 28172
rect 40552 28160 40558 28212
rect 42153 28203 42211 28209
rect 42153 28169 42165 28203
rect 42199 28200 42211 28203
rect 42536 28200 42564 28444
rect 42199 28172 42564 28200
rect 42199 28169 42211 28172
rect 42153 28163 42211 28169
rect 37476 28132 37504 28160
rect 37645 28135 37703 28141
rect 37645 28132 37657 28135
rect 37476 28104 37657 28132
rect 37645 28101 37657 28104
rect 37691 28132 37703 28135
rect 39482 28132 39488 28144
rect 37691 28104 39488 28132
rect 37691 28101 37703 28104
rect 37645 28095 37703 28101
rect 39482 28092 39488 28104
rect 39540 28092 39546 28144
rect 40034 28092 40040 28144
rect 40092 28092 40098 28144
rect 40678 28092 40684 28144
rect 40736 28092 40742 28144
rect 41414 28092 41420 28144
rect 41472 28092 41478 28144
rect 37458 28073 37464 28076
rect 37277 28067 37335 28073
rect 37277 28033 37289 28067
rect 37323 28033 37335 28067
rect 37277 28027 37335 28033
rect 37425 28067 37464 28073
rect 37425 28033 37437 28067
rect 37425 28027 37464 28033
rect 37458 28024 37464 28027
rect 37516 28024 37522 28076
rect 37553 28067 37611 28073
rect 37553 28033 37565 28067
rect 37599 28033 37611 28067
rect 37553 28027 37611 28033
rect 34609 27999 34667 28005
rect 31720 27968 33088 27996
rect 31720 27956 31726 27968
rect 33060 27940 33088 27968
rect 34609 27965 34621 27999
rect 34655 27965 34667 27999
rect 34609 27959 34667 27965
rect 32217 27931 32275 27937
rect 32217 27928 32229 27931
rect 31495 27900 32229 27928
rect 32217 27897 32229 27900
rect 32263 27897 32275 27931
rect 32217 27891 32275 27897
rect 33042 27888 33048 27940
rect 33100 27888 33106 27940
rect 34057 27931 34115 27937
rect 34057 27897 34069 27931
rect 34103 27928 34115 27931
rect 34146 27928 34152 27940
rect 34103 27900 34152 27928
rect 34103 27897 34115 27900
rect 34057 27891 34115 27897
rect 34146 27888 34152 27900
rect 34204 27888 34210 27940
rect 34624 27928 34652 27959
rect 35158 27956 35164 28008
rect 35216 27996 35222 28008
rect 36262 27996 36268 28008
rect 35216 27968 36268 27996
rect 35216 27956 35222 27968
rect 36262 27956 36268 27968
rect 36320 27956 36326 28008
rect 36648 27928 36676 28024
rect 36906 27956 36912 28008
rect 36964 27996 36970 28008
rect 37568 27996 37596 28027
rect 37734 28024 37740 28076
rect 37792 28073 37798 28076
rect 37792 28067 37819 28073
rect 37807 28033 37819 28067
rect 37792 28027 37819 28033
rect 37792 28024 37806 28027
rect 38930 28024 38936 28076
rect 38988 28024 38994 28076
rect 39758 28024 39764 28076
rect 39816 28024 39822 28076
rect 39945 28067 40003 28073
rect 39945 28033 39957 28067
rect 39991 28033 40003 28067
rect 39945 28027 40003 28033
rect 40129 28067 40187 28073
rect 40129 28033 40141 28067
rect 40175 28064 40187 28067
rect 40218 28064 40224 28076
rect 40175 28036 40224 28064
rect 40175 28033 40187 28036
rect 40129 28027 40187 28033
rect 36964 27968 37596 27996
rect 36964 27956 36970 27968
rect 37778 27928 37806 28024
rect 37918 27956 37924 28008
rect 37976 27996 37982 28008
rect 39960 27996 39988 28027
rect 40218 28024 40224 28036
rect 40276 28024 40282 28076
rect 40310 27996 40316 28008
rect 37976 27968 40316 27996
rect 37976 27956 37982 27968
rect 40310 27956 40316 27968
rect 40368 27956 40374 28008
rect 40402 27956 40408 28008
rect 40460 27956 40466 28008
rect 40218 27928 40224 27940
rect 34624 27900 35388 27928
rect 36648 27900 36952 27928
rect 37778 27900 40224 27928
rect 19300 27832 23520 27860
rect 19300 27820 19306 27832
rect 26878 27820 26884 27872
rect 26936 27860 26942 27872
rect 27433 27863 27491 27869
rect 27433 27860 27445 27863
rect 26936 27832 27445 27860
rect 26936 27820 26942 27832
rect 27433 27829 27445 27832
rect 27479 27829 27491 27863
rect 27433 27823 27491 27829
rect 27614 27820 27620 27872
rect 27672 27860 27678 27872
rect 30834 27860 30840 27872
rect 27672 27832 30840 27860
rect 27672 27820 27678 27832
rect 30834 27820 30840 27832
rect 30892 27820 30898 27872
rect 31754 27820 31760 27872
rect 31812 27860 31818 27872
rect 31941 27863 31999 27869
rect 31941 27860 31953 27863
rect 31812 27832 31953 27860
rect 31812 27820 31818 27832
rect 31941 27829 31953 27832
rect 31987 27829 31999 27863
rect 31941 27823 31999 27829
rect 33321 27863 33379 27869
rect 33321 27829 33333 27863
rect 33367 27860 33379 27863
rect 34698 27860 34704 27872
rect 33367 27832 34704 27860
rect 33367 27829 33379 27832
rect 33321 27823 33379 27829
rect 34698 27820 34704 27832
rect 34756 27820 34762 27872
rect 35360 27860 35388 27900
rect 36924 27872 36952 27900
rect 40218 27888 40224 27900
rect 40276 27888 40282 27940
rect 35618 27860 35624 27872
rect 35360 27832 35624 27860
rect 35618 27820 35624 27832
rect 35676 27820 35682 27872
rect 36906 27820 36912 27872
rect 36964 27820 36970 27872
rect 36998 27820 37004 27872
rect 37056 27820 37062 27872
rect 39022 27820 39028 27872
rect 39080 27820 39086 27872
rect 1104 27770 42504 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 42504 27770
rect 1104 27696 42504 27718
rect 3970 27616 3976 27668
rect 4028 27656 4034 27668
rect 4065 27659 4123 27665
rect 4065 27656 4077 27659
rect 4028 27628 4077 27656
rect 4028 27616 4034 27628
rect 4065 27625 4077 27628
rect 4111 27656 4123 27659
rect 4338 27656 4344 27668
rect 4111 27628 4344 27656
rect 4111 27625 4123 27628
rect 4065 27619 4123 27625
rect 4338 27616 4344 27628
rect 4396 27616 4402 27668
rect 4801 27659 4859 27665
rect 4801 27625 4813 27659
rect 4847 27656 4859 27659
rect 4890 27656 4896 27668
rect 4847 27628 4896 27656
rect 4847 27625 4859 27628
rect 4801 27619 4859 27625
rect 4890 27616 4896 27628
rect 4948 27616 4954 27668
rect 12066 27616 12072 27668
rect 12124 27656 12130 27668
rect 12124 27628 14228 27656
rect 12124 27616 12130 27628
rect 14200 27600 14228 27628
rect 14918 27616 14924 27668
rect 14976 27656 14982 27668
rect 15838 27656 15844 27668
rect 14976 27628 15844 27656
rect 14976 27616 14982 27628
rect 15838 27616 15844 27628
rect 15896 27656 15902 27668
rect 16942 27656 16948 27668
rect 15896 27628 16948 27656
rect 15896 27616 15902 27628
rect 16942 27616 16948 27628
rect 17000 27616 17006 27668
rect 17770 27616 17776 27668
rect 17828 27656 17834 27668
rect 19334 27656 19340 27668
rect 17828 27628 19340 27656
rect 17828 27616 17834 27628
rect 19334 27616 19340 27628
rect 19392 27616 19398 27668
rect 21174 27616 21180 27668
rect 21232 27656 21238 27668
rect 21232 27628 22048 27656
rect 21232 27616 21238 27628
rect 5166 27548 5172 27600
rect 5224 27548 5230 27600
rect 13265 27591 13323 27597
rect 13265 27557 13277 27591
rect 13311 27588 13323 27591
rect 13998 27588 14004 27600
rect 13311 27560 14004 27588
rect 13311 27557 13323 27560
rect 13265 27551 13323 27557
rect 13998 27548 14004 27560
rect 14056 27548 14062 27600
rect 14182 27548 14188 27600
rect 14240 27588 14246 27600
rect 15657 27591 15715 27597
rect 15657 27588 15669 27591
rect 14240 27560 15669 27588
rect 14240 27548 14246 27560
rect 15657 27557 15669 27560
rect 15703 27557 15715 27591
rect 15657 27551 15715 27557
rect 16022 27548 16028 27600
rect 16080 27588 16086 27600
rect 16117 27591 16175 27597
rect 16117 27588 16129 27591
rect 16080 27560 16129 27588
rect 16080 27548 16086 27560
rect 16117 27557 16129 27560
rect 16163 27557 16175 27591
rect 16117 27551 16175 27557
rect 17221 27591 17279 27597
rect 17221 27557 17233 27591
rect 17267 27588 17279 27591
rect 18690 27588 18696 27600
rect 17267 27560 18696 27588
rect 17267 27557 17279 27560
rect 17221 27551 17279 27557
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 21266 27548 21272 27600
rect 21324 27588 21330 27600
rect 21821 27591 21879 27597
rect 21821 27588 21833 27591
rect 21324 27560 21833 27588
rect 21324 27548 21330 27560
rect 21821 27557 21833 27560
rect 21867 27557 21879 27591
rect 22020 27588 22048 27628
rect 22094 27616 22100 27668
rect 22152 27656 22158 27668
rect 22281 27659 22339 27665
rect 22281 27656 22293 27659
rect 22152 27628 22293 27656
rect 22152 27616 22158 27628
rect 22281 27625 22293 27628
rect 22327 27625 22339 27659
rect 32398 27656 32404 27668
rect 22281 27619 22339 27625
rect 22388 27628 32404 27656
rect 22388 27588 22416 27628
rect 32398 27616 32404 27628
rect 32456 27616 32462 27668
rect 33042 27616 33048 27668
rect 33100 27656 33106 27668
rect 33962 27656 33968 27668
rect 33100 27628 33968 27656
rect 33100 27616 33106 27628
rect 33962 27616 33968 27628
rect 34020 27656 34026 27668
rect 34790 27656 34796 27668
rect 34020 27628 34796 27656
rect 34020 27616 34026 27628
rect 34790 27616 34796 27628
rect 34848 27656 34854 27668
rect 34848 27628 35204 27656
rect 34848 27616 34854 27628
rect 22020 27560 22416 27588
rect 21821 27551 21879 27557
rect 22738 27548 22744 27600
rect 22796 27588 22802 27600
rect 22925 27591 22983 27597
rect 22925 27588 22937 27591
rect 22796 27560 22937 27588
rect 22796 27548 22802 27560
rect 22925 27557 22937 27560
rect 22971 27557 22983 27591
rect 24210 27588 24216 27600
rect 22925 27551 22983 27557
rect 23032 27560 24216 27588
rect 3896 27492 4752 27520
rect 3896 27461 3924 27492
rect 4724 27464 4752 27492
rect 4798 27480 4804 27532
rect 4856 27520 4862 27532
rect 5077 27523 5135 27529
rect 5077 27520 5089 27523
rect 4856 27492 5089 27520
rect 4856 27480 4862 27492
rect 5077 27489 5089 27492
rect 5123 27489 5135 27523
rect 5077 27483 5135 27489
rect 12250 27480 12256 27532
rect 12308 27520 12314 27532
rect 14090 27520 14096 27532
rect 12308 27492 14096 27520
rect 12308 27480 12314 27492
rect 14090 27480 14096 27492
rect 14148 27480 14154 27532
rect 16206 27520 16212 27532
rect 15396 27492 16212 27520
rect 3881 27455 3939 27461
rect 3881 27421 3893 27455
rect 3927 27421 3939 27455
rect 3881 27415 3939 27421
rect 4062 27412 4068 27464
rect 4120 27412 4126 27464
rect 4706 27412 4712 27464
rect 4764 27452 4770 27464
rect 4985 27455 5043 27461
rect 4985 27452 4997 27455
rect 4764 27424 4997 27452
rect 4764 27412 4770 27424
rect 4985 27421 4997 27424
rect 5031 27421 5043 27455
rect 4985 27415 5043 27421
rect 5258 27412 5264 27464
rect 5316 27412 5322 27464
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27452 10011 27455
rect 10778 27452 10784 27464
rect 9999 27424 10784 27452
rect 9999 27421 10011 27424
rect 9953 27415 10011 27421
rect 10778 27412 10784 27424
rect 10836 27412 10842 27464
rect 12618 27452 12624 27464
rect 11440 27424 12624 27452
rect 11440 27396 11468 27424
rect 12618 27412 12624 27424
rect 12676 27412 12682 27464
rect 12989 27455 13047 27461
rect 12989 27421 13001 27455
rect 13035 27421 13047 27455
rect 12989 27415 13047 27421
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27452 13231 27455
rect 13262 27452 13268 27464
rect 13219 27424 13268 27452
rect 13219 27421 13231 27424
rect 13173 27415 13231 27421
rect 10220 27387 10278 27393
rect 10220 27353 10232 27387
rect 10266 27384 10278 27387
rect 10410 27384 10416 27396
rect 10266 27356 10416 27384
rect 10266 27353 10278 27356
rect 10220 27347 10278 27353
rect 10410 27344 10416 27356
rect 10468 27344 10474 27396
rect 11422 27344 11428 27396
rect 11480 27344 11486 27396
rect 13004 27384 13032 27415
rect 13262 27412 13268 27424
rect 13320 27412 13326 27464
rect 15396 27461 15424 27492
rect 16206 27480 16212 27492
rect 16264 27520 16270 27532
rect 18138 27520 18144 27532
rect 16264 27492 18144 27520
rect 16264 27480 16270 27492
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27421 13415 27455
rect 13357 27415 13415 27421
rect 15381 27455 15439 27461
rect 15381 27421 15393 27455
rect 15427 27421 15439 27455
rect 15381 27415 15439 27421
rect 12268 27356 13032 27384
rect 13372 27384 13400 27415
rect 15470 27412 15476 27464
rect 15528 27412 15534 27464
rect 15565 27455 15623 27461
rect 15565 27421 15577 27455
rect 15611 27452 15623 27455
rect 15746 27452 15752 27464
rect 15611 27424 15752 27452
rect 15611 27421 15623 27424
rect 15565 27415 15623 27421
rect 15746 27412 15752 27424
rect 15804 27452 15810 27464
rect 16025 27455 16083 27461
rect 16025 27452 16037 27455
rect 15804 27424 16037 27452
rect 15804 27412 15810 27424
rect 16025 27421 16037 27424
rect 16071 27421 16083 27455
rect 16025 27415 16083 27421
rect 16114 27412 16120 27464
rect 16172 27412 16178 27464
rect 16390 27412 16396 27464
rect 16448 27412 16454 27464
rect 17052 27461 17080 27492
rect 18138 27480 18144 27492
rect 18196 27520 18202 27532
rect 18196 27492 18368 27520
rect 18196 27480 18202 27492
rect 17037 27455 17095 27461
rect 17037 27421 17049 27455
rect 17083 27421 17095 27455
rect 17037 27415 17095 27421
rect 17126 27412 17132 27464
rect 17184 27452 17190 27464
rect 17221 27455 17279 27461
rect 17221 27452 17233 27455
rect 17184 27424 17233 27452
rect 17184 27412 17190 27424
rect 17221 27421 17233 27424
rect 17267 27452 17279 27455
rect 17267 27424 17448 27452
rect 17267 27421 17279 27424
rect 17221 27415 17279 27421
rect 15488 27384 15516 27412
rect 13372 27356 15516 27384
rect 15841 27387 15899 27393
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 5442 27316 5448 27328
rect 4580 27288 5448 27316
rect 4580 27276 4586 27288
rect 5442 27276 5448 27288
rect 5500 27276 5506 27328
rect 5718 27276 5724 27328
rect 5776 27316 5782 27328
rect 10594 27316 10600 27328
rect 5776 27288 10600 27316
rect 5776 27276 5782 27288
rect 10594 27276 10600 27288
rect 10652 27276 10658 27328
rect 11333 27319 11391 27325
rect 11333 27285 11345 27319
rect 11379 27316 11391 27319
rect 12268 27316 12296 27356
rect 11379 27288 12296 27316
rect 11379 27285 11391 27288
rect 11333 27279 11391 27285
rect 12342 27276 12348 27328
rect 12400 27316 12406 27328
rect 12437 27319 12495 27325
rect 12437 27316 12449 27319
rect 12400 27288 12449 27316
rect 12400 27276 12406 27288
rect 12437 27285 12449 27288
rect 12483 27285 12495 27319
rect 12437 27279 12495 27285
rect 12802 27276 12808 27328
rect 12860 27316 12866 27328
rect 13372 27316 13400 27356
rect 15841 27353 15853 27387
rect 15887 27384 15899 27387
rect 15930 27384 15936 27396
rect 15887 27356 15936 27384
rect 15887 27353 15899 27356
rect 15841 27347 15899 27353
rect 15930 27344 15936 27356
rect 15988 27344 15994 27396
rect 16301 27387 16359 27393
rect 16301 27353 16313 27387
rect 16347 27384 16359 27387
rect 16482 27384 16488 27396
rect 16347 27356 16488 27384
rect 16347 27353 16359 27356
rect 16301 27347 16359 27353
rect 16482 27344 16488 27356
rect 16540 27344 16546 27396
rect 16666 27344 16672 27396
rect 16724 27384 16730 27396
rect 17313 27387 17371 27393
rect 17313 27384 17325 27387
rect 16724 27356 17325 27384
rect 16724 27344 16730 27356
rect 17313 27353 17325 27356
rect 17359 27353 17371 27387
rect 17313 27347 17371 27353
rect 17420 27328 17448 27424
rect 17586 27412 17592 27464
rect 17644 27412 17650 27464
rect 18230 27452 18236 27464
rect 17696 27424 18236 27452
rect 17497 27387 17555 27393
rect 17497 27353 17509 27387
rect 17543 27384 17555 27387
rect 17696 27384 17724 27424
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 18340 27461 18368 27492
rect 18782 27480 18788 27532
rect 18840 27520 18846 27532
rect 18840 27492 22508 27520
rect 18840 27480 18846 27492
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 19518 27412 19524 27464
rect 19576 27452 19582 27464
rect 20530 27452 20536 27464
rect 19576 27424 20536 27452
rect 19576 27412 19582 27424
rect 20530 27412 20536 27424
rect 20588 27452 20594 27464
rect 21361 27455 21419 27461
rect 21361 27452 21373 27455
rect 20588 27424 21373 27452
rect 20588 27412 20594 27424
rect 21361 27421 21373 27424
rect 21407 27452 21419 27455
rect 21450 27452 21456 27464
rect 21407 27424 21456 27452
rect 21407 27421 21419 27424
rect 21361 27415 21419 27421
rect 21450 27412 21456 27424
rect 21508 27412 21514 27464
rect 21729 27455 21787 27461
rect 21729 27421 21741 27455
rect 21775 27421 21787 27455
rect 21729 27415 21787 27421
rect 17543 27356 17724 27384
rect 17543 27353 17555 27356
rect 17497 27347 17555 27353
rect 17770 27344 17776 27396
rect 17828 27344 17834 27396
rect 17862 27344 17868 27396
rect 17920 27344 17926 27396
rect 18417 27387 18475 27393
rect 18417 27353 18429 27387
rect 18463 27353 18475 27387
rect 18417 27347 18475 27353
rect 12860 27288 13400 27316
rect 12860 27276 12866 27288
rect 14734 27276 14740 27328
rect 14792 27316 14798 27328
rect 15473 27319 15531 27325
rect 15473 27316 15485 27319
rect 14792 27288 15485 27316
rect 14792 27276 14798 27288
rect 15473 27285 15485 27288
rect 15519 27285 15531 27319
rect 15473 27279 15531 27285
rect 17402 27276 17408 27328
rect 17460 27276 17466 27328
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 18432 27316 18460 27347
rect 19610 27344 19616 27396
rect 19668 27384 19674 27396
rect 20901 27387 20959 27393
rect 20901 27384 20913 27387
rect 19668 27356 20913 27384
rect 19668 27344 19674 27356
rect 20901 27353 20913 27356
rect 20947 27353 20959 27387
rect 20901 27347 20959 27353
rect 21174 27344 21180 27396
rect 21232 27344 21238 27396
rect 21744 27384 21772 27415
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 22005 27455 22063 27461
rect 22005 27452 22017 27455
rect 21968 27424 22017 27452
rect 21968 27412 21974 27424
rect 22005 27421 22017 27424
rect 22051 27421 22063 27455
rect 22005 27415 22063 27421
rect 22097 27455 22155 27461
rect 22097 27421 22109 27455
rect 22143 27452 22155 27455
rect 22186 27452 22192 27464
rect 22143 27424 22192 27452
rect 22143 27421 22155 27424
rect 22097 27415 22155 27421
rect 22186 27412 22192 27424
rect 22244 27412 22250 27464
rect 22370 27412 22376 27464
rect 22428 27412 22434 27464
rect 22480 27384 22508 27492
rect 22557 27455 22615 27461
rect 22557 27421 22569 27455
rect 22603 27452 22615 27455
rect 22756 27452 22784 27548
rect 22603 27424 22784 27452
rect 22833 27455 22891 27461
rect 22603 27421 22615 27424
rect 22557 27415 22615 27421
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 23032 27452 23060 27560
rect 24210 27548 24216 27560
rect 24268 27588 24274 27600
rect 24268 27560 27292 27588
rect 24268 27548 24274 27560
rect 25884 27529 25912 27560
rect 25869 27523 25927 27529
rect 23124 27492 24624 27520
rect 23124 27461 23152 27492
rect 22879 27424 23060 27452
rect 23109 27455 23167 27461
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 23109 27421 23121 27455
rect 23155 27421 23167 27455
rect 23109 27415 23167 27421
rect 23124 27384 23152 27415
rect 23290 27412 23296 27464
rect 23348 27412 23354 27464
rect 24118 27412 24124 27464
rect 24176 27452 24182 27464
rect 24596 27461 24624 27492
rect 25869 27489 25881 27523
rect 25915 27489 25927 27523
rect 25869 27483 25927 27489
rect 26050 27480 26056 27532
rect 26108 27480 26114 27532
rect 27264 27520 27292 27560
rect 28902 27548 28908 27600
rect 28960 27548 28966 27600
rect 29178 27548 29184 27600
rect 29236 27588 29242 27600
rect 29822 27588 29828 27600
rect 29236 27560 29828 27588
rect 29236 27548 29242 27560
rect 29822 27548 29828 27560
rect 29880 27588 29886 27600
rect 32677 27591 32735 27597
rect 29880 27560 32628 27588
rect 29880 27548 29886 27560
rect 27264 27492 29132 27520
rect 24397 27455 24455 27461
rect 24397 27452 24409 27455
rect 24176 27424 24409 27452
rect 24176 27412 24182 27424
rect 24397 27421 24409 27424
rect 24443 27421 24455 27455
rect 24397 27415 24455 27421
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27452 24639 27455
rect 24670 27452 24676 27464
rect 24627 27424 24676 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 24670 27412 24676 27424
rect 24728 27412 24734 27464
rect 24762 27412 24768 27464
rect 24820 27452 24826 27464
rect 26602 27452 26608 27464
rect 24820 27424 26608 27452
rect 24820 27412 24826 27424
rect 26602 27412 26608 27424
rect 26660 27412 26666 27464
rect 26878 27412 26884 27464
rect 26936 27412 26942 27464
rect 27157 27455 27215 27461
rect 27157 27421 27169 27455
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 21744 27356 22416 27384
rect 22480 27356 23152 27384
rect 24489 27387 24547 27393
rect 17644 27288 18460 27316
rect 17644 27276 17650 27288
rect 20346 27276 20352 27328
rect 20404 27316 20410 27328
rect 20625 27319 20683 27325
rect 20625 27316 20637 27319
rect 20404 27288 20637 27316
rect 20404 27276 20410 27288
rect 20625 27285 20637 27288
rect 20671 27285 20683 27319
rect 21192 27316 21220 27344
rect 21818 27316 21824 27328
rect 21192 27288 21824 27316
rect 20625 27279 20683 27285
rect 21818 27276 21824 27288
rect 21876 27276 21882 27328
rect 22388 27316 22416 27356
rect 24489 27353 24501 27387
rect 24535 27384 24547 27387
rect 24535 27356 26648 27384
rect 24535 27353 24547 27356
rect 24489 27347 24547 27353
rect 22741 27319 22799 27325
rect 22741 27316 22753 27319
rect 22388 27288 22753 27316
rect 22741 27285 22753 27288
rect 22787 27316 22799 27319
rect 23382 27316 23388 27328
rect 22787 27288 23388 27316
rect 22787 27285 22799 27288
rect 22741 27279 22799 27285
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 24578 27276 24584 27328
rect 24636 27316 24642 27328
rect 25682 27316 25688 27328
rect 24636 27288 25688 27316
rect 24636 27276 24642 27288
rect 25682 27276 25688 27288
rect 25740 27276 25746 27328
rect 25866 27276 25872 27328
rect 25924 27316 25930 27328
rect 26145 27319 26203 27325
rect 26145 27316 26157 27319
rect 25924 27288 26157 27316
rect 25924 27276 25930 27288
rect 26145 27285 26157 27288
rect 26191 27285 26203 27319
rect 26145 27279 26203 27285
rect 26510 27276 26516 27328
rect 26568 27276 26574 27328
rect 26620 27316 26648 27356
rect 26694 27344 26700 27396
rect 26752 27344 26758 27396
rect 27062 27344 27068 27396
rect 27120 27344 27126 27396
rect 27172 27384 27200 27415
rect 27338 27384 27344 27396
rect 27172 27356 27344 27384
rect 27338 27344 27344 27356
rect 27396 27344 27402 27396
rect 27430 27344 27436 27396
rect 27488 27344 27494 27396
rect 27890 27344 27896 27396
rect 27948 27344 27954 27396
rect 29104 27384 29132 27492
rect 30190 27480 30196 27532
rect 30248 27480 30254 27532
rect 30285 27523 30343 27529
rect 30285 27489 30297 27523
rect 30331 27520 30343 27523
rect 31849 27523 31907 27529
rect 31849 27520 31861 27523
rect 30331 27492 31861 27520
rect 30331 27489 30343 27492
rect 30285 27483 30343 27489
rect 31849 27489 31861 27492
rect 31895 27489 31907 27523
rect 31849 27483 31907 27489
rect 29178 27412 29184 27464
rect 29236 27452 29242 27464
rect 30006 27452 30012 27464
rect 29236 27424 30012 27452
rect 29236 27412 29242 27424
rect 30006 27412 30012 27424
rect 30064 27452 30070 27464
rect 30101 27455 30159 27461
rect 30101 27452 30113 27455
rect 30064 27424 30113 27452
rect 30064 27412 30070 27424
rect 30101 27421 30113 27424
rect 30147 27421 30159 27455
rect 30101 27415 30159 27421
rect 30300 27384 30328 27483
rect 30834 27412 30840 27464
rect 30892 27452 30898 27464
rect 31478 27452 31484 27464
rect 30892 27424 31484 27452
rect 30892 27412 30898 27424
rect 31478 27412 31484 27424
rect 31536 27452 31542 27464
rect 32125 27455 32183 27461
rect 32125 27452 32137 27455
rect 31536 27424 32137 27452
rect 31536 27412 31542 27424
rect 32125 27421 32137 27424
rect 32171 27421 32183 27455
rect 32493 27455 32551 27461
rect 32493 27452 32505 27455
rect 32125 27415 32183 27421
rect 32232 27424 32505 27452
rect 32232 27384 32260 27424
rect 32493 27421 32505 27424
rect 32539 27421 32551 27455
rect 32493 27415 32551 27421
rect 29104 27356 30328 27384
rect 31312 27356 32260 27384
rect 31312 27328 31340 27356
rect 32306 27344 32312 27396
rect 32364 27344 32370 27396
rect 32401 27387 32459 27393
rect 32401 27353 32413 27387
rect 32447 27384 32459 27387
rect 32600 27384 32628 27560
rect 32677 27557 32689 27591
rect 32723 27588 32735 27591
rect 35066 27588 35072 27600
rect 32723 27560 35072 27588
rect 32723 27557 32735 27560
rect 32677 27551 32735 27557
rect 35066 27548 35072 27560
rect 35124 27548 35130 27600
rect 33870 27480 33876 27532
rect 33928 27520 33934 27532
rect 34422 27520 34428 27532
rect 33928 27492 34428 27520
rect 33928 27480 33934 27492
rect 34422 27480 34428 27492
rect 34480 27480 34486 27532
rect 35176 27520 35204 27628
rect 35250 27548 35256 27600
rect 35308 27588 35314 27600
rect 39850 27588 39856 27600
rect 35308 27560 39856 27588
rect 35308 27548 35314 27560
rect 39850 27548 39856 27560
rect 39908 27548 39914 27600
rect 34624 27492 35112 27520
rect 35176 27492 35356 27520
rect 34624 27464 34652 27492
rect 33594 27412 33600 27464
rect 33652 27452 33658 27464
rect 34149 27455 34207 27461
rect 34149 27452 34161 27455
rect 33652 27424 34161 27452
rect 33652 27412 33658 27424
rect 34149 27421 34161 27424
rect 34195 27421 34207 27455
rect 34149 27415 34207 27421
rect 34241 27455 34299 27461
rect 34241 27421 34253 27455
rect 34287 27452 34299 27455
rect 34606 27452 34612 27464
rect 34287 27424 34612 27452
rect 34287 27421 34299 27424
rect 34241 27415 34299 27421
rect 34606 27412 34612 27424
rect 34664 27412 34670 27464
rect 34698 27412 34704 27464
rect 34756 27412 34762 27464
rect 35084 27461 35112 27492
rect 34794 27455 34852 27461
rect 34794 27421 34806 27455
rect 34840 27421 34852 27455
rect 34794 27415 34852 27421
rect 35069 27455 35127 27461
rect 35069 27421 35081 27455
rect 35115 27421 35127 27455
rect 35069 27415 35127 27421
rect 32950 27384 32956 27396
rect 32447 27356 32956 27384
rect 32447 27353 32459 27356
rect 32401 27347 32459 27353
rect 32950 27344 32956 27356
rect 33008 27344 33014 27396
rect 33502 27344 33508 27396
rect 33560 27384 33566 27396
rect 33962 27384 33968 27396
rect 33560 27356 33968 27384
rect 33560 27344 33566 27356
rect 33962 27344 33968 27356
rect 34020 27384 34026 27396
rect 34809 27384 34837 27415
rect 35158 27412 35164 27464
rect 35216 27461 35222 27464
rect 35216 27452 35224 27461
rect 35328 27452 35356 27492
rect 35434 27480 35440 27532
rect 35492 27520 35498 27532
rect 35492 27492 35848 27520
rect 35492 27480 35498 27492
rect 35820 27461 35848 27492
rect 36078 27480 36084 27532
rect 36136 27520 36142 27532
rect 36998 27520 37004 27532
rect 36136 27492 37004 27520
rect 36136 27480 36142 27492
rect 35986 27461 35992 27464
rect 35713 27455 35771 27461
rect 35713 27452 35725 27455
rect 35216 27424 35261 27452
rect 35328 27424 35725 27452
rect 35216 27415 35224 27424
rect 35713 27421 35725 27424
rect 35759 27421 35771 27455
rect 35713 27415 35771 27421
rect 35805 27455 35863 27461
rect 35805 27421 35817 27455
rect 35851 27421 35863 27455
rect 35805 27415 35863 27421
rect 35953 27455 35992 27461
rect 35953 27421 35965 27455
rect 35953 27415 35992 27421
rect 35216 27412 35222 27415
rect 35986 27412 35992 27415
rect 36044 27412 36050 27464
rect 36188 27461 36216 27492
rect 36998 27480 37004 27492
rect 37056 27480 37062 27532
rect 37274 27480 37280 27532
rect 37332 27520 37338 27532
rect 38286 27520 38292 27532
rect 37332 27492 38292 27520
rect 37332 27480 37338 27492
rect 38286 27480 38292 27492
rect 38344 27520 38350 27532
rect 38841 27523 38899 27529
rect 38841 27520 38853 27523
rect 38344 27492 38853 27520
rect 38344 27480 38350 27492
rect 38841 27489 38853 27492
rect 38887 27489 38899 27523
rect 38841 27483 38899 27489
rect 38930 27480 38936 27532
rect 38988 27520 38994 27532
rect 39114 27520 39120 27532
rect 38988 27492 39120 27520
rect 38988 27480 38994 27492
rect 39114 27480 39120 27492
rect 39172 27480 39178 27532
rect 40144 27492 40724 27520
rect 36173 27455 36231 27461
rect 36173 27421 36185 27455
rect 36219 27421 36231 27455
rect 36173 27415 36231 27421
rect 36262 27412 36268 27464
rect 36320 27461 36326 27464
rect 36320 27452 36328 27461
rect 36320 27424 36365 27452
rect 36320 27415 36328 27424
rect 36320 27412 36326 27415
rect 36446 27412 36452 27464
rect 36504 27452 36510 27464
rect 40144 27461 40172 27492
rect 40129 27455 40187 27461
rect 36504 27424 39528 27452
rect 36504 27412 36510 27424
rect 34020 27356 34837 27384
rect 34977 27387 35035 27393
rect 34020 27344 34026 27356
rect 34977 27353 34989 27387
rect 35023 27384 35035 27387
rect 35618 27384 35624 27396
rect 35023 27356 35624 27384
rect 35023 27353 35035 27356
rect 34977 27347 35035 27353
rect 35618 27344 35624 27356
rect 35676 27384 35682 27396
rect 36081 27387 36139 27393
rect 36081 27384 36093 27387
rect 35676 27356 36093 27384
rect 35676 27344 35682 27356
rect 36081 27353 36093 27356
rect 36127 27384 36139 27387
rect 38102 27384 38108 27396
rect 36127 27356 38108 27384
rect 36127 27353 36139 27356
rect 36081 27347 36139 27353
rect 38102 27344 38108 27356
rect 38160 27344 38166 27396
rect 39043 27387 39101 27393
rect 39043 27353 39055 27387
rect 39089 27384 39101 27387
rect 39089 27356 39160 27384
rect 39089 27353 39101 27356
rect 39043 27347 39101 27353
rect 28074 27316 28080 27328
rect 26620 27288 28080 27316
rect 28074 27276 28080 27288
rect 28132 27276 28138 27328
rect 29733 27319 29791 27325
rect 29733 27285 29745 27319
rect 29779 27316 29791 27319
rect 29914 27316 29920 27328
rect 29779 27288 29920 27316
rect 29779 27285 29791 27288
rect 29733 27279 29791 27285
rect 29914 27276 29920 27288
rect 29972 27276 29978 27328
rect 31294 27276 31300 27328
rect 31352 27276 31358 27328
rect 31386 27276 31392 27328
rect 31444 27316 31450 27328
rect 31665 27319 31723 27325
rect 31665 27316 31677 27319
rect 31444 27288 31677 27316
rect 31444 27276 31450 27288
rect 31665 27285 31677 27288
rect 31711 27285 31723 27319
rect 31665 27279 31723 27285
rect 31754 27276 31760 27328
rect 31812 27276 31818 27328
rect 33781 27319 33839 27325
rect 33781 27285 33793 27319
rect 33827 27316 33839 27319
rect 34054 27316 34060 27328
rect 33827 27288 34060 27316
rect 33827 27285 33839 27288
rect 33781 27279 33839 27285
rect 34054 27276 34060 27288
rect 34112 27276 34118 27328
rect 35345 27319 35403 27325
rect 35345 27285 35357 27319
rect 35391 27316 35403 27319
rect 35434 27316 35440 27328
rect 35391 27288 35440 27316
rect 35391 27285 35403 27288
rect 35345 27279 35403 27285
rect 35434 27276 35440 27288
rect 35492 27276 35498 27328
rect 35529 27319 35587 27325
rect 35529 27285 35541 27319
rect 35575 27316 35587 27319
rect 36354 27316 36360 27328
rect 35575 27288 36360 27316
rect 35575 27285 35587 27288
rect 35529 27279 35587 27285
rect 36354 27276 36360 27288
rect 36412 27276 36418 27328
rect 36449 27319 36507 27325
rect 36449 27285 36461 27319
rect 36495 27316 36507 27319
rect 37826 27316 37832 27328
rect 36495 27288 37832 27316
rect 36495 27285 36507 27288
rect 36449 27279 36507 27285
rect 37826 27276 37832 27288
rect 37884 27276 37890 27328
rect 38010 27276 38016 27328
rect 38068 27316 38074 27328
rect 38197 27319 38255 27325
rect 38197 27316 38209 27319
rect 38068 27288 38209 27316
rect 38068 27276 38074 27288
rect 38197 27285 38209 27288
rect 38243 27285 38255 27319
rect 38197 27279 38255 27285
rect 38470 27276 38476 27328
rect 38528 27316 38534 27328
rect 38565 27319 38623 27325
rect 38565 27316 38577 27319
rect 38528 27288 38577 27316
rect 38528 27276 38534 27288
rect 38565 27285 38577 27288
rect 38611 27285 38623 27319
rect 38565 27279 38623 27285
rect 38657 27319 38715 27325
rect 38657 27285 38669 27319
rect 38703 27316 38715 27319
rect 38746 27316 38752 27328
rect 38703 27288 38752 27316
rect 38703 27285 38715 27288
rect 38657 27279 38715 27285
rect 38746 27276 38752 27288
rect 38804 27276 38810 27328
rect 38930 27276 38936 27328
rect 38988 27316 38994 27328
rect 39132 27316 39160 27356
rect 39206 27344 39212 27396
rect 39264 27344 39270 27396
rect 39500 27384 39528 27424
rect 40129 27421 40141 27455
rect 40175 27421 40187 27455
rect 40405 27455 40463 27461
rect 40405 27452 40417 27455
rect 40129 27415 40187 27421
rect 40236 27424 40417 27452
rect 40236 27384 40264 27424
rect 40405 27421 40417 27424
rect 40451 27421 40463 27455
rect 40405 27415 40463 27421
rect 40497 27455 40555 27461
rect 40497 27421 40509 27455
rect 40543 27421 40555 27455
rect 40497 27415 40555 27421
rect 39500 27356 40264 27384
rect 40310 27344 40316 27396
rect 40368 27344 40374 27396
rect 40512 27384 40540 27415
rect 40420 27356 40540 27384
rect 40696 27384 40724 27492
rect 40770 27412 40776 27464
rect 40828 27412 40834 27464
rect 41325 27455 41383 27461
rect 41325 27452 41337 27455
rect 40880 27424 41337 27452
rect 40880 27384 40908 27424
rect 41325 27421 41337 27424
rect 41371 27452 41383 27455
rect 41598 27452 41604 27464
rect 41371 27424 41604 27452
rect 41371 27421 41383 27424
rect 41325 27415 41383 27421
rect 41598 27412 41604 27424
rect 41656 27412 41662 27464
rect 41693 27455 41751 27461
rect 41693 27421 41705 27455
rect 41739 27421 41751 27455
rect 41693 27415 41751 27421
rect 40696 27356 40908 27384
rect 40957 27387 41015 27393
rect 38988 27288 39160 27316
rect 38988 27276 38994 27288
rect 39390 27276 39396 27328
rect 39448 27276 39454 27328
rect 40218 27276 40224 27328
rect 40276 27316 40282 27328
rect 40420 27316 40448 27356
rect 40957 27353 40969 27387
rect 41003 27353 41015 27387
rect 40957 27347 41015 27353
rect 40276 27288 40448 27316
rect 40681 27319 40739 27325
rect 40276 27276 40282 27288
rect 40681 27285 40693 27319
rect 40727 27316 40739 27319
rect 40972 27316 41000 27347
rect 41046 27344 41052 27396
rect 41104 27384 41110 27396
rect 41708 27384 41736 27415
rect 41104 27356 41736 27384
rect 41104 27344 41110 27356
rect 40727 27288 41000 27316
rect 40727 27285 40739 27288
rect 40681 27279 40739 27285
rect 41138 27276 41144 27328
rect 41196 27276 41202 27328
rect 41506 27276 41512 27328
rect 41564 27276 41570 27328
rect 41874 27276 41880 27328
rect 41932 27276 41938 27328
rect 1104 27226 42504 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 42504 27226
rect 1104 27152 42504 27174
rect 3050 27072 3056 27124
rect 3108 27072 3114 27124
rect 3605 27115 3663 27121
rect 3605 27081 3617 27115
rect 3651 27112 3663 27115
rect 4798 27112 4804 27124
rect 3651 27084 4804 27112
rect 3651 27081 3663 27084
rect 3605 27075 3663 27081
rect 4798 27072 4804 27084
rect 4856 27072 4862 27124
rect 8110 27112 8116 27124
rect 7208 27084 8116 27112
rect 2869 27047 2927 27053
rect 2869 27013 2881 27047
rect 2915 27013 2927 27047
rect 2869 27007 2927 27013
rect 3237 27047 3295 27053
rect 3237 27013 3249 27047
rect 3283 27044 3295 27047
rect 3510 27044 3516 27056
rect 3283 27016 3516 27044
rect 3283 27013 3295 27016
rect 3237 27007 3295 27013
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 1762 26976 1768 26988
rect 1719 26948 1768 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 2884 26976 2912 27007
rect 3510 27004 3516 27016
rect 3568 27004 3574 27056
rect 7208 27053 7236 27084
rect 8110 27072 8116 27084
rect 8168 27072 8174 27124
rect 10137 27115 10195 27121
rect 10137 27081 10149 27115
rect 10183 27112 10195 27115
rect 10226 27112 10232 27124
rect 10183 27084 10232 27112
rect 10183 27081 10195 27084
rect 10137 27075 10195 27081
rect 10226 27072 10232 27084
rect 10284 27072 10290 27124
rect 10410 27072 10416 27124
rect 10468 27072 10474 27124
rect 10594 27072 10600 27124
rect 10652 27112 10658 27124
rect 12802 27112 12808 27124
rect 10652 27084 12808 27112
rect 10652 27072 10658 27084
rect 12802 27072 12808 27084
rect 12860 27072 12866 27124
rect 12897 27115 12955 27121
rect 12897 27081 12909 27115
rect 12943 27112 12955 27115
rect 13170 27112 13176 27124
rect 12943 27084 13176 27112
rect 12943 27081 12955 27084
rect 12897 27075 12955 27081
rect 13170 27072 13176 27084
rect 13228 27072 13234 27124
rect 14369 27115 14427 27121
rect 14369 27081 14381 27115
rect 14415 27112 14427 27115
rect 14415 27084 14780 27112
rect 14415 27081 14427 27084
rect 14369 27075 14427 27081
rect 7193 27047 7251 27053
rect 7193 27013 7205 27047
rect 7239 27013 7251 27047
rect 7193 27007 7251 27013
rect 8202 27004 8208 27056
rect 8260 27004 8266 27056
rect 10873 27047 10931 27053
rect 10873 27044 10885 27047
rect 10152 27016 10885 27044
rect 10152 26988 10180 27016
rect 10873 27013 10885 27016
rect 10919 27044 10931 27047
rect 13541 27047 13599 27053
rect 13541 27044 13553 27047
rect 10919 27016 12726 27044
rect 10919 27013 10931 27016
rect 10873 27007 10931 27013
rect 3326 26976 3332 26988
rect 2884 26948 3332 26976
rect 3326 26936 3332 26948
rect 3384 26976 3390 26988
rect 3421 26979 3479 26985
rect 3421 26976 3433 26979
rect 3384 26948 3433 26976
rect 3384 26936 3390 26948
rect 3421 26945 3433 26948
rect 3467 26945 3479 26979
rect 3421 26939 3479 26945
rect 3878 26936 3884 26988
rect 3936 26976 3942 26988
rect 3973 26979 4031 26985
rect 3973 26976 3985 26979
rect 3936 26948 3985 26976
rect 3936 26936 3942 26948
rect 3973 26945 3985 26948
rect 4019 26945 4031 26979
rect 3973 26939 4031 26945
rect 4065 26979 4123 26985
rect 4065 26945 4077 26979
rect 4111 26945 4123 26979
rect 4065 26939 4123 26945
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26945 4307 26979
rect 4249 26939 4307 26945
rect 2501 26843 2559 26849
rect 2501 26809 2513 26843
rect 2547 26840 2559 26843
rect 2590 26840 2596 26852
rect 2547 26812 2596 26840
rect 2547 26809 2559 26812
rect 2501 26803 2559 26809
rect 2590 26800 2596 26812
rect 2648 26800 2654 26852
rect 4080 26840 4108 26939
rect 4264 26908 4292 26939
rect 4338 26936 4344 26988
rect 4396 26936 4402 26988
rect 4522 26936 4528 26988
rect 4580 26976 4586 26988
rect 4709 26979 4767 26985
rect 4709 26976 4721 26979
rect 4580 26948 4721 26976
rect 4580 26936 4586 26948
rect 4709 26945 4721 26948
rect 4755 26945 4767 26979
rect 4985 26979 5043 26985
rect 4985 26976 4997 26979
rect 4709 26939 4767 26945
rect 4908 26948 4997 26976
rect 4798 26908 4804 26920
rect 4264 26880 4804 26908
rect 4798 26868 4804 26880
rect 4856 26868 4862 26920
rect 4908 26917 4936 26948
rect 4985 26945 4997 26948
rect 5031 26945 5043 26979
rect 4985 26939 5043 26945
rect 5169 26979 5227 26985
rect 5169 26945 5181 26979
rect 5215 26976 5227 26979
rect 5442 26976 5448 26988
rect 5215 26948 5448 26976
rect 5215 26945 5227 26948
rect 5169 26939 5227 26945
rect 5442 26936 5448 26948
rect 5500 26936 5506 26988
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26976 9275 26979
rect 9674 26976 9680 26988
rect 9263 26948 9680 26976
rect 9263 26945 9275 26948
rect 9217 26939 9275 26945
rect 9674 26936 9680 26948
rect 9732 26936 9738 26988
rect 10042 26936 10048 26988
rect 10100 26936 10106 26988
rect 10134 26936 10140 26988
rect 10192 26936 10198 26988
rect 10229 26979 10287 26985
rect 10229 26945 10241 26979
rect 10275 26976 10287 26979
rect 10502 26976 10508 26988
rect 10275 26948 10508 26976
rect 10275 26945 10287 26948
rect 10229 26939 10287 26945
rect 4893 26911 4951 26917
rect 4893 26877 4905 26911
rect 4939 26877 4951 26911
rect 5994 26908 6000 26920
rect 4893 26871 4951 26877
rect 5184 26880 6000 26908
rect 4706 26840 4712 26852
rect 4080 26812 4712 26840
rect 4706 26800 4712 26812
rect 4764 26840 4770 26852
rect 4908 26840 4936 26871
rect 5184 26840 5212 26880
rect 5994 26868 6000 26880
rect 6052 26868 6058 26920
rect 7190 26868 7196 26920
rect 7248 26908 7254 26920
rect 8202 26908 8208 26920
rect 7248 26880 8208 26908
rect 7248 26868 7254 26880
rect 8202 26868 8208 26880
rect 8260 26868 8266 26920
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8941 26911 8999 26917
rect 8941 26908 8953 26911
rect 8628 26880 8953 26908
rect 8628 26868 8634 26880
rect 8941 26877 8953 26880
rect 8987 26877 8999 26911
rect 8941 26871 8999 26877
rect 9861 26911 9919 26917
rect 9861 26877 9873 26911
rect 9907 26908 9919 26911
rect 10244 26908 10272 26939
rect 10502 26936 10508 26948
rect 10560 26936 10566 26988
rect 10781 26979 10839 26985
rect 10781 26945 10793 26979
rect 10827 26976 10839 26979
rect 11793 26979 11851 26985
rect 11793 26976 11805 26979
rect 10827 26948 11805 26976
rect 10827 26945 10839 26948
rect 10781 26939 10839 26945
rect 11793 26945 11805 26948
rect 11839 26976 11851 26979
rect 12342 26976 12348 26988
rect 11839 26948 12348 26976
rect 11839 26945 11851 26948
rect 11793 26939 11851 26945
rect 12342 26936 12348 26948
rect 12400 26936 12406 26988
rect 12698 26985 12726 27016
rect 13096 27016 13553 27044
rect 13096 26988 13124 27016
rect 13541 27013 13553 27016
rect 13587 27013 13599 27047
rect 13541 27007 13599 27013
rect 13906 27004 13912 27056
rect 13964 27004 13970 27056
rect 14642 27044 14648 27056
rect 14016 27016 14648 27044
rect 12529 26979 12587 26985
rect 12529 26945 12541 26979
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 12683 26979 12741 26985
rect 12683 26945 12695 26979
rect 12729 26976 12741 26979
rect 13078 26976 13084 26988
rect 12729 26948 13084 26976
rect 12729 26945 12741 26948
rect 12683 26939 12741 26945
rect 9907 26880 10272 26908
rect 9907 26877 9919 26880
rect 9861 26871 9919 26877
rect 10962 26868 10968 26920
rect 11020 26868 11026 26920
rect 11514 26868 11520 26920
rect 11572 26868 11578 26920
rect 4764 26812 4936 26840
rect 5000 26812 5212 26840
rect 4764 26800 4770 26812
rect 842 26732 848 26784
rect 900 26772 906 26784
rect 1489 26775 1547 26781
rect 1489 26772 1501 26775
rect 900 26744 1501 26772
rect 900 26732 906 26744
rect 1489 26741 1501 26744
rect 1535 26741 1547 26775
rect 1489 26735 1547 26741
rect 2866 26732 2872 26784
rect 2924 26732 2930 26784
rect 3786 26732 3792 26784
rect 3844 26732 3850 26784
rect 4525 26775 4583 26781
rect 4525 26741 4537 26775
rect 4571 26772 4583 26775
rect 5000 26772 5028 26812
rect 5258 26800 5264 26852
rect 5316 26840 5322 26852
rect 5718 26840 5724 26852
rect 5316 26812 5724 26840
rect 5316 26800 5322 26812
rect 5718 26800 5724 26812
rect 5776 26800 5782 26852
rect 10226 26800 10232 26852
rect 10284 26840 10290 26852
rect 12544 26840 12572 26939
rect 13078 26936 13084 26948
rect 13136 26936 13142 26988
rect 13354 26936 13360 26988
rect 13412 26936 13418 26988
rect 13817 26979 13875 26985
rect 13817 26945 13829 26979
rect 13863 26945 13875 26979
rect 13817 26939 13875 26945
rect 12989 26911 13047 26917
rect 12989 26877 13001 26911
rect 13035 26908 13047 26911
rect 13170 26908 13176 26920
rect 13035 26880 13176 26908
rect 13035 26877 13047 26880
rect 12989 26871 13047 26877
rect 13170 26868 13176 26880
rect 13228 26868 13234 26920
rect 12618 26840 12624 26852
rect 10284 26812 12624 26840
rect 10284 26800 10290 26812
rect 12618 26800 12624 26812
rect 12676 26840 12682 26852
rect 13725 26843 13783 26849
rect 13725 26840 13737 26843
rect 12676 26812 13737 26840
rect 12676 26800 12682 26812
rect 13725 26809 13737 26812
rect 13771 26809 13783 26843
rect 13832 26840 13860 26939
rect 14016 26917 14044 27016
rect 14642 27004 14648 27016
rect 14700 27004 14706 27056
rect 14752 27053 14780 27084
rect 16666 27072 16672 27124
rect 16724 27112 16730 27124
rect 17494 27112 17500 27124
rect 16724 27084 17500 27112
rect 16724 27072 16730 27084
rect 17494 27072 17500 27084
rect 17552 27112 17558 27124
rect 17770 27112 17776 27124
rect 17552 27084 17776 27112
rect 17552 27072 17558 27084
rect 17770 27072 17776 27084
rect 17828 27072 17834 27124
rect 19978 27112 19984 27124
rect 19720 27084 19984 27112
rect 14737 27047 14795 27053
rect 14737 27013 14749 27047
rect 14783 27013 14795 27047
rect 14737 27007 14795 27013
rect 15194 27004 15200 27056
rect 15252 27004 15258 27056
rect 16298 27004 16304 27056
rect 16356 27044 16362 27056
rect 16485 27047 16543 27053
rect 16485 27044 16497 27047
rect 16356 27016 16497 27044
rect 16356 27004 16362 27016
rect 16485 27013 16497 27016
rect 16531 27013 16543 27047
rect 16485 27007 16543 27013
rect 17402 27004 17408 27056
rect 17460 27044 17466 27056
rect 17957 27047 18015 27053
rect 17957 27044 17969 27047
rect 17460 27016 17969 27044
rect 17460 27004 17466 27016
rect 17957 27013 17969 27016
rect 18003 27013 18015 27047
rect 17957 27007 18015 27013
rect 18138 27004 18144 27056
rect 18196 27004 18202 27056
rect 19720 27044 19748 27084
rect 19978 27072 19984 27084
rect 20036 27112 20042 27124
rect 20036 27084 20668 27112
rect 20036 27072 20042 27084
rect 20640 27044 20668 27084
rect 24946 27072 24952 27124
rect 25004 27112 25010 27124
rect 25777 27115 25835 27121
rect 25777 27112 25789 27115
rect 25004 27084 25789 27112
rect 25004 27072 25010 27084
rect 25777 27081 25789 27084
rect 25823 27112 25835 27115
rect 25866 27112 25872 27124
rect 25823 27084 25872 27112
rect 25823 27081 25835 27084
rect 25777 27075 25835 27081
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 26694 27072 26700 27124
rect 26752 27112 26758 27124
rect 26973 27115 27031 27121
rect 26973 27112 26985 27115
rect 26752 27084 26985 27112
rect 26752 27072 26758 27084
rect 26973 27081 26985 27084
rect 27019 27081 27031 27115
rect 26973 27075 27031 27081
rect 27062 27072 27068 27124
rect 27120 27112 27126 27124
rect 27430 27112 27436 27124
rect 27120 27084 27436 27112
rect 27120 27072 27126 27084
rect 27430 27072 27436 27084
rect 27488 27072 27494 27124
rect 28074 27072 28080 27124
rect 28132 27112 28138 27124
rect 35158 27112 35164 27124
rect 28132 27084 35164 27112
rect 28132 27072 28138 27084
rect 35158 27072 35164 27084
rect 35216 27112 35222 27124
rect 36262 27112 36268 27124
rect 35216 27084 36268 27112
rect 35216 27072 35222 27084
rect 36262 27072 36268 27084
rect 36320 27072 36326 27124
rect 36998 27072 37004 27124
rect 37056 27112 37062 27124
rect 38105 27115 38163 27121
rect 38105 27112 38117 27115
rect 37056 27084 38117 27112
rect 37056 27072 37062 27084
rect 38105 27081 38117 27084
rect 38151 27081 38163 27115
rect 38105 27075 38163 27081
rect 38565 27115 38623 27121
rect 38565 27081 38577 27115
rect 38611 27112 38623 27115
rect 40034 27112 40040 27124
rect 38611 27084 40040 27112
rect 38611 27081 38623 27084
rect 38565 27075 38623 27081
rect 40034 27072 40040 27084
rect 40092 27072 40098 27124
rect 21361 27047 21419 27053
rect 21361 27044 21373 27047
rect 18616 27016 19826 27044
rect 20640 27016 21373 27044
rect 14182 26936 14188 26988
rect 14240 26936 14246 26988
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 18616 26976 18644 27016
rect 21361 27013 21373 27016
rect 21407 27013 21419 27047
rect 21361 27007 21419 27013
rect 21450 27004 21456 27056
rect 21508 27044 21514 27056
rect 21545 27047 21603 27053
rect 21545 27044 21557 27047
rect 21508 27016 21557 27044
rect 21508 27004 21514 27016
rect 21545 27013 21557 27016
rect 21591 27013 21603 27047
rect 21545 27007 21603 27013
rect 22922 27004 22928 27056
rect 22980 27044 22986 27056
rect 24578 27044 24584 27056
rect 22980 27016 24584 27044
rect 22980 27004 22986 27016
rect 24578 27004 24584 27016
rect 24636 27044 24642 27056
rect 24636 27016 24794 27044
rect 24636 27004 24642 27016
rect 26510 27004 26516 27056
rect 26568 27044 26574 27056
rect 26568 27016 27568 27044
rect 26568 27004 26574 27016
rect 18104 26948 18644 26976
rect 18104 26936 18110 26948
rect 18690 26936 18696 26988
rect 18748 26936 18754 26988
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 25700 26948 27169 26976
rect 14001 26911 14059 26917
rect 14001 26877 14013 26911
rect 14047 26877 14059 26911
rect 14001 26871 14059 26877
rect 14090 26868 14096 26920
rect 14148 26908 14154 26920
rect 14461 26911 14519 26917
rect 14461 26908 14473 26911
rect 14148 26880 14473 26908
rect 14148 26868 14154 26880
rect 14461 26877 14473 26880
rect 14507 26877 14519 26911
rect 14461 26871 14519 26877
rect 17770 26868 17776 26920
rect 17828 26908 17834 26920
rect 19426 26908 19432 26920
rect 17828 26880 19432 26908
rect 17828 26868 17834 26880
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 19518 26868 19524 26920
rect 19576 26908 19582 26920
rect 20438 26908 20444 26920
rect 19576 26880 20444 26908
rect 19576 26868 19582 26880
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 20990 26868 20996 26920
rect 21048 26868 21054 26920
rect 21269 26911 21327 26917
rect 21269 26877 21281 26911
rect 21315 26908 21327 26911
rect 21358 26908 21364 26920
rect 21315 26880 21364 26908
rect 21315 26877 21327 26880
rect 21269 26871 21327 26877
rect 21358 26868 21364 26880
rect 21416 26908 21422 26920
rect 24029 26911 24087 26917
rect 24029 26908 24041 26911
rect 21416 26880 24041 26908
rect 21416 26868 21422 26880
rect 24029 26877 24041 26880
rect 24075 26877 24087 26911
rect 24029 26871 24087 26877
rect 24302 26868 24308 26920
rect 24360 26868 24366 26920
rect 18325 26843 18383 26849
rect 13832 26812 14596 26840
rect 13725 26803 13783 26809
rect 4571 26744 5028 26772
rect 5077 26775 5135 26781
rect 4571 26741 4583 26744
rect 4525 26735 4583 26741
rect 5077 26741 5089 26775
rect 5123 26772 5135 26775
rect 6546 26772 6552 26784
rect 5123 26744 6552 26772
rect 5123 26741 5135 26744
rect 5077 26735 5135 26741
rect 6546 26732 6552 26744
rect 6604 26732 6610 26784
rect 8386 26732 8392 26784
rect 8444 26772 8450 26784
rect 9309 26775 9367 26781
rect 9309 26772 9321 26775
rect 8444 26744 9321 26772
rect 8444 26732 8450 26744
rect 9309 26741 9321 26744
rect 9355 26741 9367 26775
rect 9309 26735 9367 26741
rect 11238 26732 11244 26784
rect 11296 26772 11302 26784
rect 11609 26775 11667 26781
rect 11609 26772 11621 26775
rect 11296 26744 11621 26772
rect 11296 26732 11302 26744
rect 11609 26741 11621 26744
rect 11655 26741 11667 26775
rect 11609 26735 11667 26741
rect 11698 26732 11704 26784
rect 11756 26732 11762 26784
rect 13817 26775 13875 26781
rect 13817 26741 13829 26775
rect 13863 26772 13875 26775
rect 13909 26775 13967 26781
rect 13909 26772 13921 26775
rect 13863 26744 13921 26772
rect 13863 26741 13875 26744
rect 13817 26735 13875 26741
rect 13909 26741 13921 26744
rect 13955 26741 13967 26775
rect 14568 26772 14596 26812
rect 18325 26809 18337 26843
rect 18371 26840 18383 26843
rect 18598 26840 18604 26852
rect 18371 26812 18604 26840
rect 18371 26809 18383 26812
rect 18325 26803 18383 26809
rect 18598 26800 18604 26812
rect 18656 26840 18662 26852
rect 23290 26840 23296 26852
rect 18656 26812 19334 26840
rect 18656 26800 18662 26812
rect 14918 26772 14924 26784
rect 14568 26744 14924 26772
rect 13909 26735 13967 26741
rect 14918 26732 14924 26744
rect 14976 26732 14982 26784
rect 16758 26732 16764 26784
rect 16816 26772 16822 26784
rect 18877 26775 18935 26781
rect 18877 26772 18889 26775
rect 16816 26744 18889 26772
rect 16816 26732 16822 26744
rect 18877 26741 18889 26744
rect 18923 26772 18935 26775
rect 19150 26772 19156 26784
rect 18923 26744 19156 26772
rect 18923 26741 18935 26744
rect 18877 26735 18935 26741
rect 19150 26732 19156 26744
rect 19208 26732 19214 26784
rect 19306 26772 19334 26812
rect 21468 26812 23296 26840
rect 21468 26772 21496 26812
rect 23290 26800 23296 26812
rect 23348 26800 23354 26852
rect 19306 26744 21496 26772
rect 21542 26732 21548 26784
rect 21600 26772 21606 26784
rect 25700 26772 25728 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27246 26936 27252 26988
rect 27304 26936 27310 26988
rect 27540 26985 27568 27016
rect 29822 27004 29828 27056
rect 29880 27004 29886 27056
rect 30742 27004 30748 27056
rect 30800 27044 30806 27056
rect 36446 27044 36452 27056
rect 30800 27016 36452 27044
rect 30800 27004 30806 27016
rect 36446 27004 36452 27016
rect 36504 27004 36510 27056
rect 36630 27004 36636 27056
rect 36688 27044 36694 27056
rect 38197 27047 38255 27053
rect 38197 27044 38209 27047
rect 36688 27016 38209 27044
rect 36688 27004 36694 27016
rect 38197 27013 38209 27016
rect 38243 27044 38255 27047
rect 38654 27044 38660 27056
rect 38243 27016 38660 27044
rect 38243 27013 38255 27016
rect 38197 27007 38255 27013
rect 38654 27004 38660 27016
rect 38712 27004 38718 27056
rect 39117 27047 39175 27053
rect 39117 27013 39129 27047
rect 39163 27044 39175 27047
rect 39390 27044 39396 27056
rect 39163 27016 39396 27044
rect 39163 27013 39175 27016
rect 39117 27007 39175 27013
rect 39390 27004 39396 27016
rect 39448 27004 39454 27056
rect 39574 27004 39580 27056
rect 39632 27004 39638 27056
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 25866 26868 25872 26920
rect 25924 26908 25930 26920
rect 26513 26911 26571 26917
rect 26513 26908 26525 26911
rect 25924 26880 26525 26908
rect 25924 26868 25930 26880
rect 26513 26877 26525 26880
rect 26559 26877 26571 26911
rect 26513 26871 26571 26877
rect 26602 26868 26608 26920
rect 26660 26908 26666 26920
rect 27356 26908 27384 26939
rect 29270 26936 29276 26988
rect 29328 26976 29334 26988
rect 29549 26979 29607 26985
rect 29549 26976 29561 26979
rect 29328 26948 29561 26976
rect 29328 26936 29334 26948
rect 29549 26945 29561 26948
rect 29595 26945 29607 26979
rect 29549 26939 29607 26945
rect 29733 26979 29791 26985
rect 29733 26945 29745 26979
rect 29779 26945 29791 26979
rect 29733 26939 29791 26945
rect 26660 26880 27384 26908
rect 26660 26868 26666 26880
rect 27982 26868 27988 26920
rect 28040 26908 28046 26920
rect 29748 26908 29776 26939
rect 29914 26936 29920 26988
rect 29972 26936 29978 26988
rect 32306 26976 32312 26988
rect 31726 26948 32312 26976
rect 31726 26908 31754 26948
rect 32306 26936 32312 26948
rect 32364 26936 32370 26988
rect 41230 26936 41236 26988
rect 41288 26936 41294 26988
rect 28040 26880 31754 26908
rect 28040 26868 28046 26880
rect 34422 26868 34428 26920
rect 34480 26908 34486 26920
rect 38013 26911 38071 26917
rect 38013 26908 38025 26911
rect 34480 26880 38025 26908
rect 34480 26868 34486 26880
rect 38013 26877 38025 26880
rect 38059 26908 38071 26911
rect 38286 26908 38292 26920
rect 38059 26880 38292 26908
rect 38059 26877 38071 26880
rect 38013 26871 38071 26877
rect 38286 26868 38292 26880
rect 38344 26868 38350 26920
rect 38841 26911 38899 26917
rect 38841 26877 38853 26911
rect 38887 26908 38899 26911
rect 40402 26908 40408 26920
rect 38887 26880 40408 26908
rect 38887 26877 38899 26880
rect 38841 26871 38899 26877
rect 40402 26868 40408 26880
rect 40460 26868 40466 26920
rect 42150 26868 42156 26920
rect 42208 26868 42214 26920
rect 40218 26800 40224 26852
rect 40276 26840 40282 26852
rect 40589 26843 40647 26849
rect 40589 26840 40601 26843
rect 40276 26812 40601 26840
rect 40276 26800 40282 26812
rect 40589 26809 40601 26812
rect 40635 26840 40647 26843
rect 41046 26840 41052 26852
rect 40635 26812 41052 26840
rect 40635 26809 40647 26812
rect 40589 26803 40647 26809
rect 41046 26800 41052 26812
rect 41104 26800 41110 26852
rect 41417 26843 41475 26849
rect 41417 26809 41429 26843
rect 41463 26840 41475 26843
rect 41690 26840 41696 26852
rect 41463 26812 41696 26840
rect 41463 26809 41475 26812
rect 41417 26803 41475 26809
rect 41690 26800 41696 26812
rect 41748 26800 41754 26852
rect 21600 26744 25728 26772
rect 21600 26732 21606 26744
rect 25958 26732 25964 26784
rect 26016 26732 26022 26784
rect 30101 26775 30159 26781
rect 30101 26741 30113 26775
rect 30147 26772 30159 26775
rect 40770 26772 40776 26784
rect 30147 26744 40776 26772
rect 30147 26741 30159 26744
rect 30101 26735 30159 26741
rect 40770 26732 40776 26744
rect 40828 26732 40834 26784
rect 41506 26732 41512 26784
rect 41564 26732 41570 26784
rect 1104 26682 42504 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 42504 26682
rect 1104 26608 42504 26630
rect 4798 26528 4804 26580
rect 4856 26568 4862 26580
rect 4893 26571 4951 26577
rect 4893 26568 4905 26571
rect 4856 26540 4905 26568
rect 4856 26528 4862 26540
rect 4893 26537 4905 26540
rect 4939 26537 4951 26571
rect 6178 26568 6184 26580
rect 4893 26531 4951 26537
rect 5092 26540 6184 26568
rect 2961 26435 3019 26441
rect 2961 26401 2973 26435
rect 3007 26432 3019 26435
rect 3786 26432 3792 26444
rect 3007 26404 3792 26432
rect 3007 26401 3019 26404
rect 2961 26395 3019 26401
rect 3786 26392 3792 26404
rect 3844 26392 3850 26444
rect 5092 26432 5120 26540
rect 6178 26528 6184 26540
rect 6236 26528 6242 26580
rect 8570 26528 8576 26580
rect 8628 26528 8634 26580
rect 10226 26568 10232 26580
rect 8680 26540 10232 26568
rect 7558 26460 7564 26512
rect 7616 26500 7622 26512
rect 8680 26500 8708 26540
rect 10226 26528 10232 26540
rect 10284 26528 10290 26580
rect 10321 26571 10379 26577
rect 10321 26537 10333 26571
rect 10367 26568 10379 26571
rect 10502 26568 10508 26580
rect 10367 26540 10508 26568
rect 10367 26537 10379 26540
rect 10321 26531 10379 26537
rect 10502 26528 10508 26540
rect 10560 26528 10566 26580
rect 10870 26528 10876 26580
rect 10928 26568 10934 26580
rect 11330 26568 11336 26580
rect 10928 26540 11336 26568
rect 10928 26528 10934 26540
rect 7616 26472 8708 26500
rect 7616 26460 7622 26472
rect 5718 26432 5724 26444
rect 3896 26404 5120 26432
rect 5368 26404 5724 26432
rect 3896 26373 3924 26404
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26333 3295 26367
rect 3237 26327 3295 26333
rect 3881 26367 3939 26373
rect 3881 26333 3893 26367
rect 3927 26333 3939 26367
rect 3881 26327 3939 26333
rect 3050 26296 3056 26308
rect 2530 26268 3056 26296
rect 3050 26256 3056 26268
rect 3108 26256 3114 26308
rect 3252 26296 3280 26327
rect 4614 26324 4620 26376
rect 4672 26324 4678 26376
rect 4706 26324 4712 26376
rect 4764 26364 4770 26376
rect 4985 26367 5043 26373
rect 4985 26364 4997 26367
rect 4764 26336 4997 26364
rect 4764 26324 4770 26336
rect 4985 26333 4997 26336
rect 5031 26333 5043 26367
rect 4985 26327 5043 26333
rect 5074 26324 5080 26376
rect 5132 26324 5138 26376
rect 5166 26324 5172 26376
rect 5224 26364 5230 26376
rect 5368 26373 5396 26404
rect 5718 26392 5724 26404
rect 5776 26392 5782 26444
rect 10980 26441 11008 26540
rect 11330 26528 11336 26540
rect 11388 26568 11394 26580
rect 12250 26568 12256 26580
rect 11388 26540 12256 26568
rect 11388 26528 11394 26540
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 12618 26528 12624 26580
rect 12676 26568 12682 26580
rect 12989 26571 13047 26577
rect 12989 26568 13001 26571
rect 12676 26540 13001 26568
rect 12676 26528 12682 26540
rect 12989 26537 13001 26540
rect 13035 26537 13047 26571
rect 12989 26531 13047 26537
rect 13722 26528 13728 26580
rect 13780 26528 13786 26580
rect 14182 26528 14188 26580
rect 14240 26568 14246 26580
rect 14829 26571 14887 26577
rect 14829 26568 14841 26571
rect 14240 26540 14841 26568
rect 14240 26528 14246 26540
rect 14829 26537 14841 26540
rect 14875 26568 14887 26571
rect 14875 26540 19012 26568
rect 14875 26537 14887 26540
rect 14829 26531 14887 26537
rect 12713 26503 12771 26509
rect 12713 26469 12725 26503
rect 12759 26500 12771 26503
rect 12802 26500 12808 26512
rect 12759 26472 12808 26500
rect 12759 26469 12771 26472
rect 12713 26463 12771 26469
rect 12802 26460 12808 26472
rect 12860 26460 12866 26512
rect 16942 26500 16948 26512
rect 13188 26472 15056 26500
rect 7193 26435 7251 26441
rect 7193 26401 7205 26435
rect 7239 26432 7251 26435
rect 7837 26435 7895 26441
rect 7837 26432 7849 26435
rect 7239 26404 7849 26432
rect 7239 26401 7251 26404
rect 7193 26395 7251 26401
rect 7837 26401 7849 26404
rect 7883 26401 7895 26435
rect 7837 26395 7895 26401
rect 10965 26435 11023 26441
rect 10965 26401 10977 26435
rect 11011 26401 11023 26435
rect 10965 26395 11023 26401
rect 5261 26367 5319 26373
rect 5261 26364 5273 26367
rect 5224 26336 5273 26364
rect 5224 26324 5230 26336
rect 5261 26333 5273 26336
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26333 5411 26367
rect 5353 26327 5411 26333
rect 5445 26367 5503 26373
rect 5445 26333 5457 26367
rect 5491 26333 5503 26367
rect 5445 26327 5503 26333
rect 4632 26296 4660 26324
rect 5460 26296 5488 26327
rect 8018 26324 8024 26376
rect 8076 26324 8082 26376
rect 8110 26324 8116 26376
rect 8168 26364 8174 26376
rect 8297 26367 8355 26373
rect 8297 26364 8309 26367
rect 8168 26336 8309 26364
rect 8168 26324 8174 26336
rect 8297 26333 8309 26336
rect 8343 26333 8355 26367
rect 8297 26327 8355 26333
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 8570 26364 8576 26376
rect 8435 26336 8576 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 8941 26367 8999 26373
rect 8941 26333 8953 26367
rect 8987 26364 8999 26367
rect 9674 26364 9680 26376
rect 8987 26336 9680 26364
rect 8987 26333 8999 26336
rect 8941 26327 8999 26333
rect 9674 26324 9680 26336
rect 9732 26364 9738 26376
rect 10980 26364 11008 26395
rect 11238 26392 11244 26444
rect 11296 26392 11302 26444
rect 12434 26392 12440 26444
rect 12492 26392 12498 26444
rect 12897 26435 12955 26441
rect 12897 26401 12909 26435
rect 12943 26432 12955 26435
rect 13078 26432 13084 26444
rect 12943 26404 13084 26432
rect 12943 26401 12955 26404
rect 12897 26395 12955 26401
rect 13078 26392 13084 26404
rect 13136 26392 13142 26444
rect 9732 26336 11008 26364
rect 12452 26364 12480 26392
rect 13188 26373 13216 26472
rect 13630 26392 13636 26444
rect 13688 26432 13694 26444
rect 13725 26435 13783 26441
rect 13725 26432 13737 26435
rect 13688 26404 13737 26432
rect 13688 26392 13694 26404
rect 13725 26401 13737 26404
rect 13771 26432 13783 26435
rect 13771 26404 14688 26432
rect 13771 26401 13783 26404
rect 13725 26395 13783 26401
rect 13173 26367 13231 26373
rect 13173 26364 13185 26367
rect 12452 26336 13185 26364
rect 9732 26324 9738 26336
rect 13173 26333 13185 26336
rect 13219 26333 13231 26367
rect 13173 26327 13231 26333
rect 13817 26367 13875 26373
rect 13817 26333 13829 26367
rect 13863 26333 13875 26367
rect 13817 26327 13875 26333
rect 3252 26268 5488 26296
rect 5718 26256 5724 26308
rect 5776 26256 5782 26308
rect 6454 26256 6460 26308
rect 6512 26256 6518 26308
rect 7098 26256 7104 26308
rect 7156 26296 7162 26308
rect 8205 26299 8263 26305
rect 8205 26296 8217 26299
rect 7156 26268 8217 26296
rect 7156 26256 7162 26268
rect 8205 26265 8217 26268
rect 8251 26265 8263 26299
rect 8205 26259 8263 26265
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 9186 26299 9244 26305
rect 9186 26296 9198 26299
rect 8536 26268 9198 26296
rect 8536 26256 8542 26268
rect 9186 26265 9198 26268
rect 9232 26265 9244 26299
rect 13078 26296 13084 26308
rect 12466 26268 13084 26296
rect 9186 26259 9244 26265
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 13357 26299 13415 26305
rect 13357 26265 13369 26299
rect 13403 26296 13415 26299
rect 13832 26296 13860 26327
rect 14550 26324 14556 26376
rect 14608 26324 14614 26376
rect 14660 26373 14688 26404
rect 14645 26367 14703 26373
rect 14645 26333 14657 26367
rect 14691 26364 14703 26367
rect 14734 26364 14740 26376
rect 14691 26336 14740 26364
rect 14691 26333 14703 26336
rect 14645 26327 14703 26333
rect 14734 26324 14740 26336
rect 14792 26324 14798 26376
rect 15028 26364 15056 26472
rect 15120 26472 16948 26500
rect 15120 26441 15148 26472
rect 16942 26460 16948 26472
rect 17000 26500 17006 26512
rect 17770 26500 17776 26512
rect 17000 26472 17776 26500
rect 17000 26460 17006 26472
rect 17770 26460 17776 26472
rect 17828 26500 17834 26512
rect 17865 26503 17923 26509
rect 17865 26500 17877 26503
rect 17828 26472 17877 26500
rect 17828 26460 17834 26472
rect 17865 26469 17877 26472
rect 17911 26469 17923 26503
rect 17865 26463 17923 26469
rect 18138 26460 18144 26512
rect 18196 26500 18202 26512
rect 18325 26503 18383 26509
rect 18325 26500 18337 26503
rect 18196 26472 18337 26500
rect 18196 26460 18202 26472
rect 18325 26469 18337 26472
rect 18371 26469 18383 26503
rect 18325 26463 18383 26469
rect 18693 26503 18751 26509
rect 18693 26469 18705 26503
rect 18739 26500 18751 26503
rect 18782 26500 18788 26512
rect 18739 26472 18788 26500
rect 18739 26469 18751 26472
rect 18693 26463 18751 26469
rect 18782 26460 18788 26472
rect 18840 26460 18846 26512
rect 18984 26500 19012 26540
rect 19150 26528 19156 26580
rect 19208 26568 19214 26580
rect 19245 26571 19303 26577
rect 19245 26568 19257 26571
rect 19208 26540 19257 26568
rect 19208 26528 19214 26540
rect 19245 26537 19257 26540
rect 19291 26537 19303 26571
rect 19245 26531 19303 26537
rect 19610 26528 19616 26580
rect 19668 26528 19674 26580
rect 20809 26571 20867 26577
rect 20809 26537 20821 26571
rect 20855 26568 20867 26571
rect 20990 26568 20996 26580
rect 20855 26540 20996 26568
rect 20855 26537 20867 26540
rect 20809 26531 20867 26537
rect 20990 26528 20996 26540
rect 21048 26528 21054 26580
rect 21450 26568 21456 26580
rect 21192 26540 21456 26568
rect 19628 26500 19656 26528
rect 21192 26500 21220 26540
rect 21450 26528 21456 26540
rect 21508 26528 21514 26580
rect 21542 26528 21548 26580
rect 21600 26568 21606 26580
rect 21600 26540 24256 26568
rect 21600 26528 21606 26540
rect 18984 26472 19288 26500
rect 19628 26472 21220 26500
rect 22833 26503 22891 26509
rect 15105 26435 15163 26441
rect 15105 26401 15117 26435
rect 15151 26401 15163 26435
rect 15105 26395 15163 26401
rect 15194 26392 15200 26444
rect 15252 26392 15258 26444
rect 15565 26435 15623 26441
rect 15565 26401 15577 26435
rect 15611 26432 15623 26435
rect 15654 26432 15660 26444
rect 15611 26404 15660 26432
rect 15611 26401 15623 26404
rect 15565 26395 15623 26401
rect 15654 26392 15660 26404
rect 15712 26392 15718 26444
rect 18230 26432 18236 26444
rect 17972 26404 18236 26432
rect 15473 26367 15531 26373
rect 15473 26364 15485 26367
rect 15028 26336 15485 26364
rect 15473 26333 15485 26336
rect 15519 26333 15531 26367
rect 15473 26327 15531 26333
rect 13403 26268 13860 26296
rect 15488 26296 15516 26327
rect 17586 26324 17592 26376
rect 17644 26324 17650 26376
rect 17678 26324 17684 26376
rect 17736 26324 17742 26376
rect 17972 26373 18000 26404
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 18506 26432 18512 26444
rect 18340 26404 18512 26432
rect 17957 26367 18015 26373
rect 17957 26333 17969 26367
rect 18003 26333 18015 26367
rect 17957 26327 18015 26333
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26364 18107 26367
rect 18340 26364 18368 26404
rect 18506 26392 18512 26404
rect 18564 26392 18570 26444
rect 18984 26441 19012 26472
rect 18969 26435 19027 26441
rect 18969 26401 18981 26435
rect 19015 26401 19027 26435
rect 19260 26432 19288 26472
rect 22833 26469 22845 26503
rect 22879 26500 22891 26503
rect 23198 26500 23204 26512
rect 22879 26472 23204 26500
rect 22879 26469 22891 26472
rect 22833 26463 22891 26469
rect 23198 26460 23204 26472
rect 23256 26460 23262 26512
rect 24228 26500 24256 26540
rect 24302 26528 24308 26580
rect 24360 26568 24366 26580
rect 24581 26571 24639 26577
rect 24581 26568 24593 26571
rect 24360 26540 24593 26568
rect 24360 26528 24366 26540
rect 24581 26537 24593 26540
rect 24627 26537 24639 26571
rect 24581 26531 24639 26537
rect 24670 26528 24676 26580
rect 24728 26568 24734 26580
rect 33318 26568 33324 26580
rect 24728 26540 33324 26568
rect 24728 26528 24734 26540
rect 33318 26528 33324 26540
rect 33376 26528 33382 26580
rect 35434 26528 35440 26580
rect 35492 26528 35498 26580
rect 36357 26571 36415 26577
rect 36357 26537 36369 26571
rect 36403 26568 36415 26571
rect 36630 26568 36636 26580
rect 36403 26540 36636 26568
rect 36403 26537 36415 26540
rect 36357 26531 36415 26537
rect 36630 26528 36636 26540
rect 36688 26528 36694 26580
rect 38473 26571 38531 26577
rect 38473 26537 38485 26571
rect 38519 26568 38531 26571
rect 38930 26568 38936 26580
rect 38519 26540 38936 26568
rect 38519 26537 38531 26540
rect 38473 26531 38531 26537
rect 38930 26528 38936 26540
rect 38988 26528 38994 26580
rect 24857 26503 24915 26509
rect 24228 26472 24808 26500
rect 19337 26435 19395 26441
rect 19337 26432 19349 26435
rect 19260 26404 19349 26432
rect 18969 26395 19027 26401
rect 19337 26401 19349 26404
rect 19383 26401 19395 26435
rect 19337 26395 19395 26401
rect 19426 26392 19432 26444
rect 19484 26432 19490 26444
rect 20257 26435 20315 26441
rect 20257 26432 20269 26435
rect 19484 26404 20269 26432
rect 19484 26392 19490 26404
rect 20257 26401 20269 26404
rect 20303 26432 20315 26435
rect 20346 26432 20352 26444
rect 20303 26404 20352 26432
rect 20303 26401 20315 26404
rect 20257 26395 20315 26401
rect 20346 26392 20352 26404
rect 20404 26392 20410 26444
rect 21085 26435 21143 26441
rect 21085 26401 21097 26435
rect 21131 26432 21143 26435
rect 21358 26432 21364 26444
rect 21131 26404 21364 26432
rect 21131 26401 21143 26404
rect 21085 26395 21143 26401
rect 21358 26392 21364 26404
rect 21416 26392 21422 26444
rect 21450 26392 21456 26444
rect 21508 26432 21514 26444
rect 21508 26404 24532 26432
rect 21508 26392 21514 26404
rect 18598 26364 18604 26376
rect 18095 26336 18368 26364
rect 18432 26336 18604 26364
rect 18095 26333 18107 26336
rect 18049 26327 18107 26333
rect 17862 26296 17868 26308
rect 15488 26268 17868 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 17862 26256 17868 26268
rect 17920 26256 17926 26308
rect 17972 26296 18000 26327
rect 18141 26299 18199 26305
rect 18141 26296 18153 26299
rect 17972 26268 18153 26296
rect 18141 26265 18153 26268
rect 18187 26265 18199 26299
rect 18141 26259 18199 26265
rect 18325 26299 18383 26305
rect 18325 26265 18337 26299
rect 18371 26296 18383 26299
rect 18432 26296 18460 26336
rect 18598 26324 18604 26336
rect 18656 26324 18662 26376
rect 19242 26324 19248 26376
rect 19300 26324 19306 26376
rect 23109 26367 23167 26373
rect 19352 26336 20852 26364
rect 19352 26296 19380 26336
rect 18371 26268 18460 26296
rect 19306 26268 19380 26296
rect 20349 26299 20407 26305
rect 18371 26265 18383 26268
rect 18325 26259 18383 26265
rect 1489 26231 1547 26237
rect 1489 26197 1501 26231
rect 1535 26228 1547 26231
rect 2038 26228 2044 26240
rect 1535 26200 2044 26228
rect 1535 26197 1547 26200
rect 1489 26191 1547 26197
rect 2038 26188 2044 26200
rect 2096 26228 2102 26240
rect 2866 26228 2872 26240
rect 2096 26200 2872 26228
rect 2096 26188 2102 26200
rect 2866 26188 2872 26200
rect 2924 26188 2930 26240
rect 5074 26188 5080 26240
rect 5132 26228 5138 26240
rect 5810 26228 5816 26240
rect 5132 26200 5816 26228
rect 5132 26188 5138 26200
rect 5810 26188 5816 26200
rect 5868 26188 5874 26240
rect 7006 26188 7012 26240
rect 7064 26228 7070 26240
rect 7285 26231 7343 26237
rect 7285 26228 7297 26231
rect 7064 26200 7297 26228
rect 7064 26188 7070 26200
rect 7285 26197 7297 26200
rect 7331 26197 7343 26231
rect 7285 26191 7343 26197
rect 13446 26188 13452 26240
rect 13504 26188 13510 26240
rect 14921 26231 14979 26237
rect 14921 26197 14933 26231
rect 14967 26228 14979 26231
rect 15102 26228 15108 26240
rect 14967 26200 15108 26228
rect 14967 26197 14979 26200
rect 14921 26191 14979 26197
rect 15102 26188 15108 26200
rect 15160 26188 15166 26240
rect 15378 26188 15384 26240
rect 15436 26188 15442 26240
rect 17402 26188 17408 26240
rect 17460 26188 17466 26240
rect 18230 26188 18236 26240
rect 18288 26228 18294 26240
rect 18509 26231 18567 26237
rect 18509 26228 18521 26231
rect 18288 26200 18521 26228
rect 18288 26188 18294 26200
rect 18509 26197 18521 26200
rect 18555 26228 18567 26231
rect 19306 26228 19334 26268
rect 20349 26265 20361 26299
rect 20395 26296 20407 26299
rect 20714 26296 20720 26308
rect 20395 26268 20720 26296
rect 20395 26265 20407 26268
rect 20349 26259 20407 26265
rect 20714 26256 20720 26268
rect 20772 26256 20778 26308
rect 20824 26296 20852 26336
rect 23109 26333 23121 26367
rect 23155 26333 23167 26367
rect 23109 26327 23167 26333
rect 23293 26367 23351 26373
rect 23293 26333 23305 26367
rect 23339 26364 23351 26367
rect 24118 26364 24124 26376
rect 23339 26336 24124 26364
rect 23339 26333 23351 26336
rect 23293 26327 23351 26333
rect 20824 26268 21312 26296
rect 18555 26200 19334 26228
rect 18555 26197 18567 26200
rect 18509 26191 18567 26197
rect 20438 26188 20444 26240
rect 20496 26188 20502 26240
rect 21284 26228 21312 26268
rect 21358 26256 21364 26308
rect 21416 26256 21422 26308
rect 21450 26256 21456 26308
rect 21508 26256 21514 26308
rect 22922 26296 22928 26308
rect 22586 26268 22928 26296
rect 22922 26256 22928 26268
rect 22980 26256 22986 26308
rect 21468 26228 21496 26256
rect 21284 26200 21496 26228
rect 23014 26188 23020 26240
rect 23072 26228 23078 26240
rect 23124 26228 23152 26327
rect 24118 26324 24124 26336
rect 24176 26324 24182 26376
rect 23201 26299 23259 26305
rect 23201 26265 23213 26299
rect 23247 26296 23259 26299
rect 24394 26296 24400 26308
rect 23247 26268 24400 26296
rect 23247 26265 23259 26268
rect 23201 26259 23259 26265
rect 24394 26256 24400 26268
rect 24452 26256 24458 26308
rect 24504 26296 24532 26404
rect 24780 26376 24808 26472
rect 24857 26469 24869 26503
rect 24903 26500 24915 26503
rect 25498 26500 25504 26512
rect 24903 26472 25504 26500
rect 24903 26469 24915 26472
rect 24857 26463 24915 26469
rect 25498 26460 25504 26472
rect 25556 26460 25562 26512
rect 35452 26500 35480 26528
rect 41046 26500 41052 26512
rect 35452 26472 41052 26500
rect 41046 26460 41052 26472
rect 41104 26460 41110 26512
rect 25041 26435 25099 26441
rect 25041 26401 25053 26435
rect 25087 26432 25099 26435
rect 25958 26432 25964 26444
rect 25087 26404 25964 26432
rect 25087 26401 25099 26404
rect 25041 26395 25099 26401
rect 25958 26392 25964 26404
rect 26016 26392 26022 26444
rect 31754 26392 31760 26444
rect 31812 26432 31818 26444
rect 33505 26435 33563 26441
rect 33505 26432 33517 26435
rect 31812 26404 33517 26432
rect 31812 26392 31818 26404
rect 33505 26401 33517 26404
rect 33551 26432 33563 26435
rect 35250 26432 35256 26444
rect 33551 26404 35256 26432
rect 33551 26401 33563 26404
rect 33505 26395 33563 26401
rect 35250 26392 35256 26404
rect 35308 26392 35314 26444
rect 35434 26392 35440 26444
rect 35492 26432 35498 26444
rect 35621 26435 35679 26441
rect 35621 26432 35633 26435
rect 35492 26404 35633 26432
rect 35492 26392 35498 26404
rect 35621 26401 35633 26404
rect 35667 26401 35679 26435
rect 35621 26395 35679 26401
rect 35805 26435 35863 26441
rect 35805 26401 35817 26435
rect 35851 26432 35863 26435
rect 36722 26432 36728 26444
rect 35851 26404 36728 26432
rect 35851 26401 35863 26404
rect 35805 26395 35863 26401
rect 36722 26392 36728 26404
rect 36780 26392 36786 26444
rect 37826 26392 37832 26444
rect 37884 26432 37890 26444
rect 41322 26432 41328 26444
rect 37884 26404 41328 26432
rect 37884 26392 37890 26404
rect 41322 26392 41328 26404
rect 41380 26392 41386 26444
rect 24762 26324 24768 26376
rect 24820 26324 24826 26376
rect 24946 26324 24952 26376
rect 25004 26324 25010 26376
rect 25222 26324 25228 26376
rect 25280 26324 25286 26376
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26364 25743 26367
rect 25774 26364 25780 26376
rect 25731 26336 25780 26364
rect 25731 26333 25743 26336
rect 25685 26327 25743 26333
rect 25774 26324 25780 26336
rect 25832 26324 25838 26376
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26364 25927 26367
rect 26326 26364 26332 26376
rect 25915 26336 26332 26364
rect 25915 26333 25927 26336
rect 25869 26327 25927 26333
rect 26326 26324 26332 26336
rect 26384 26364 26390 26376
rect 27062 26364 27068 26376
rect 26384 26336 27068 26364
rect 26384 26324 26390 26336
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 29546 26324 29552 26376
rect 29604 26364 29610 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 29604 26336 29745 26364
rect 29604 26324 29610 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 33321 26367 33379 26373
rect 33321 26333 33333 26367
rect 33367 26364 33379 26367
rect 33594 26364 33600 26376
rect 33367 26336 33600 26364
rect 33367 26333 33379 26336
rect 33321 26327 33379 26333
rect 33594 26324 33600 26336
rect 33652 26324 33658 26376
rect 35342 26324 35348 26376
rect 35400 26324 35406 26376
rect 35529 26367 35587 26373
rect 35529 26333 35541 26367
rect 35575 26364 35587 26367
rect 36078 26364 36084 26376
rect 35575 26336 36084 26364
rect 35575 26333 35587 26336
rect 35529 26327 35587 26333
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 37458 26324 37464 26376
rect 37516 26364 37522 26376
rect 37921 26367 37979 26373
rect 37921 26364 37933 26367
rect 37516 26336 37933 26364
rect 37516 26324 37522 26336
rect 37921 26333 37933 26336
rect 37967 26333 37979 26367
rect 37921 26327 37979 26333
rect 38010 26324 38016 26376
rect 38068 26364 38074 26376
rect 38289 26367 38347 26373
rect 38289 26364 38301 26367
rect 38068 26336 38301 26364
rect 38068 26324 38074 26336
rect 38289 26333 38301 26336
rect 38335 26333 38347 26367
rect 38289 26327 38347 26333
rect 38746 26324 38752 26376
rect 38804 26324 38810 26376
rect 39853 26367 39911 26373
rect 39853 26333 39865 26367
rect 39899 26364 39911 26367
rect 39899 26336 39933 26364
rect 39899 26333 39911 26336
rect 39853 26327 39911 26333
rect 26970 26296 26976 26308
rect 24504 26268 26976 26296
rect 26970 26256 26976 26268
rect 27028 26256 27034 26308
rect 28718 26256 28724 26308
rect 28776 26296 28782 26308
rect 29641 26299 29699 26305
rect 29641 26296 29653 26299
rect 28776 26268 29653 26296
rect 28776 26256 28782 26268
rect 29641 26265 29653 26268
rect 29687 26265 29699 26299
rect 29641 26259 29699 26265
rect 35805 26299 35863 26305
rect 35805 26265 35817 26299
rect 35851 26296 35863 26299
rect 35986 26296 35992 26308
rect 35851 26268 35992 26296
rect 35851 26265 35863 26268
rect 35805 26259 35863 26265
rect 35986 26256 35992 26268
rect 36044 26256 36050 26308
rect 36096 26296 36124 26324
rect 36538 26296 36544 26308
rect 36096 26268 36544 26296
rect 36538 26256 36544 26268
rect 36596 26256 36602 26308
rect 38102 26256 38108 26308
rect 38160 26256 38166 26308
rect 38197 26299 38255 26305
rect 38197 26265 38209 26299
rect 38243 26296 38255 26299
rect 38378 26296 38384 26308
rect 38243 26268 38384 26296
rect 38243 26265 38255 26268
rect 38197 26259 38255 26265
rect 38378 26256 38384 26268
rect 38436 26256 38442 26308
rect 39577 26299 39635 26305
rect 39577 26265 39589 26299
rect 39623 26296 39635 26299
rect 39868 26296 39896 26327
rect 40402 26296 40408 26308
rect 39623 26268 40408 26296
rect 39623 26265 39635 26268
rect 39577 26259 39635 26265
rect 40402 26256 40408 26268
rect 40460 26256 40466 26308
rect 26602 26228 26608 26240
rect 23072 26200 26608 26228
rect 23072 26188 23078 26200
rect 26602 26188 26608 26200
rect 26660 26188 26666 26240
rect 27154 26188 27160 26240
rect 27212 26228 27218 26240
rect 31754 26228 31760 26240
rect 27212 26200 31760 26228
rect 27212 26188 27218 26200
rect 31754 26188 31760 26200
rect 31812 26188 31818 26240
rect 32950 26188 32956 26240
rect 33008 26188 33014 26240
rect 33410 26188 33416 26240
rect 33468 26188 33474 26240
rect 36170 26188 36176 26240
rect 36228 26188 36234 26240
rect 36341 26231 36399 26237
rect 36341 26197 36353 26231
rect 36387 26228 36399 26231
rect 36906 26228 36912 26240
rect 36387 26200 36912 26228
rect 36387 26197 36399 26200
rect 36341 26191 36399 26197
rect 36906 26188 36912 26200
rect 36964 26188 36970 26240
rect 1104 26138 42504 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 42504 26138
rect 1104 26064 42504 26086
rect 3605 26027 3663 26033
rect 3605 25993 3617 26027
rect 3651 26024 3663 26027
rect 3878 26024 3884 26036
rect 3651 25996 3884 26024
rect 3651 25993 3663 25996
rect 3605 25987 3663 25993
rect 3878 25984 3884 25996
rect 3936 25984 3942 26036
rect 5718 25984 5724 26036
rect 5776 26024 5782 26036
rect 6365 26027 6423 26033
rect 6365 26024 6377 26027
rect 5776 25996 6377 26024
rect 5776 25984 5782 25996
rect 6365 25993 6377 25996
rect 6411 25993 6423 26027
rect 6365 25987 6423 25993
rect 7101 26027 7159 26033
rect 7101 25993 7113 26027
rect 7147 26024 7159 26027
rect 8018 26024 8024 26036
rect 7147 25996 8024 26024
rect 7147 25993 7159 25996
rect 7101 25987 7159 25993
rect 8018 25984 8024 25996
rect 8076 25984 8082 26036
rect 8205 26027 8263 26033
rect 8205 25993 8217 26027
rect 8251 26024 8263 26027
rect 8478 26024 8484 26036
rect 8251 25996 8484 26024
rect 8251 25993 8263 25996
rect 8205 25987 8263 25993
rect 8478 25984 8484 25996
rect 8536 25984 8542 26036
rect 14921 26027 14979 26033
rect 14921 25993 14933 26027
rect 14967 26024 14979 26027
rect 16666 26024 16672 26036
rect 14967 25996 16672 26024
rect 14967 25993 14979 25996
rect 14921 25987 14979 25993
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 20714 25984 20720 26036
rect 20772 25984 20778 26036
rect 21358 25984 21364 26036
rect 21416 26024 21422 26036
rect 21821 26027 21879 26033
rect 21821 26024 21833 26027
rect 21416 25996 21833 26024
rect 21416 25984 21422 25996
rect 21821 25993 21833 25996
rect 21867 25993 21879 26027
rect 21821 25987 21879 25993
rect 22189 26027 22247 26033
rect 22189 25993 22201 26027
rect 22235 26024 22247 26027
rect 22830 26024 22836 26036
rect 22235 25996 22836 26024
rect 22235 25993 22247 25996
rect 22189 25987 22247 25993
rect 22830 25984 22836 25996
rect 22888 26024 22894 26036
rect 23198 26024 23204 26036
rect 22888 25996 23204 26024
rect 22888 25984 22894 25996
rect 23198 25984 23204 25996
rect 23256 25984 23262 26036
rect 23290 25984 23296 26036
rect 23348 26024 23354 26036
rect 25038 26024 25044 26036
rect 23348 25996 25044 26024
rect 23348 25984 23354 25996
rect 25038 25984 25044 25996
rect 25096 25984 25102 26036
rect 25133 26027 25191 26033
rect 25133 25993 25145 26027
rect 25179 26024 25191 26027
rect 25222 26024 25228 26036
rect 25179 25996 25228 26024
rect 25179 25993 25191 25996
rect 25133 25987 25191 25993
rect 25222 25984 25228 25996
rect 25280 25984 25286 26036
rect 25323 25996 26188 26024
rect 3237 25959 3295 25965
rect 2792 25928 3004 25956
rect 2038 25848 2044 25900
rect 2096 25848 2102 25900
rect 2195 25891 2253 25897
rect 2195 25857 2207 25891
rect 2241 25888 2253 25891
rect 2590 25888 2596 25900
rect 2241 25860 2596 25888
rect 2241 25857 2253 25860
rect 2195 25851 2253 25857
rect 2590 25848 2596 25860
rect 2648 25848 2654 25900
rect 2792 25897 2820 25928
rect 2777 25891 2835 25897
rect 2777 25857 2789 25891
rect 2823 25857 2835 25891
rect 2777 25851 2835 25857
rect 2866 25848 2872 25900
rect 2924 25848 2930 25900
rect 2976 25888 3004 25928
rect 3237 25925 3249 25959
rect 3283 25956 3295 25959
rect 4062 25956 4068 25968
rect 3283 25928 4068 25956
rect 3283 25925 3295 25928
rect 3237 25919 3295 25925
rect 4062 25916 4068 25928
rect 4120 25916 4126 25968
rect 4985 25959 5043 25965
rect 4985 25925 4997 25959
rect 5031 25956 5043 25959
rect 5626 25956 5632 25968
rect 5031 25928 5632 25956
rect 5031 25925 5043 25928
rect 4985 25919 5043 25925
rect 5626 25916 5632 25928
rect 5684 25916 5690 25968
rect 7929 25959 7987 25965
rect 7929 25925 7941 25959
rect 7975 25956 7987 25959
rect 8386 25956 8392 25968
rect 7975 25928 8392 25956
rect 7975 25925 7987 25928
rect 7929 25919 7987 25925
rect 8386 25916 8392 25928
rect 8444 25916 8450 25968
rect 8573 25959 8631 25965
rect 8573 25925 8585 25959
rect 8619 25956 8631 25959
rect 8941 25959 8999 25965
rect 8941 25956 8953 25959
rect 8619 25928 8953 25956
rect 8619 25925 8631 25928
rect 8573 25919 8631 25925
rect 8941 25925 8953 25928
rect 8987 25925 8999 25959
rect 10042 25956 10048 25968
rect 8941 25919 8999 25925
rect 9600 25928 10048 25956
rect 3326 25888 3332 25900
rect 2976 25860 3332 25888
rect 3326 25848 3332 25860
rect 3384 25848 3390 25900
rect 3510 25848 3516 25900
rect 3568 25848 3574 25900
rect 4525 25891 4583 25897
rect 4525 25857 4537 25891
rect 4571 25888 4583 25891
rect 4614 25888 4620 25900
rect 4571 25860 4620 25888
rect 4571 25857 4583 25860
rect 4525 25851 4583 25857
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 4798 25848 4804 25900
rect 4856 25897 4862 25900
rect 4856 25891 4905 25897
rect 4856 25857 4859 25891
rect 4893 25857 4905 25891
rect 4856 25851 4905 25857
rect 5077 25891 5135 25897
rect 5077 25857 5089 25891
rect 5123 25857 5135 25891
rect 5258 25888 5264 25900
rect 5219 25860 5264 25888
rect 5077 25851 5135 25857
rect 4856 25848 4862 25851
rect 2409 25823 2467 25829
rect 2409 25789 2421 25823
rect 2455 25820 2467 25823
rect 3528 25820 3556 25848
rect 2455 25792 3556 25820
rect 5092 25820 5120 25851
rect 5258 25848 5264 25860
rect 5316 25848 5322 25900
rect 5350 25848 5356 25900
rect 5408 25848 5414 25900
rect 6546 25848 6552 25900
rect 6604 25848 6610 25900
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25888 6883 25891
rect 7006 25888 7012 25900
rect 6871 25860 7012 25888
rect 6871 25857 6883 25860
rect 6825 25851 6883 25857
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7650 25848 7656 25900
rect 7708 25848 7714 25900
rect 7834 25848 7840 25900
rect 7892 25848 7898 25900
rect 8021 25891 8079 25897
rect 8021 25857 8033 25891
rect 8067 25857 8079 25891
rect 8021 25851 8079 25857
rect 6733 25823 6791 25829
rect 5092 25792 5212 25820
rect 2455 25789 2467 25792
rect 2409 25783 2467 25789
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 4709 25687 4767 25693
rect 4709 25684 4721 25687
rect 4120 25656 4721 25684
rect 4120 25644 4126 25656
rect 4709 25653 4721 25656
rect 4755 25653 4767 25687
rect 5184 25684 5212 25792
rect 6733 25789 6745 25823
rect 6779 25820 6791 25823
rect 7098 25820 7104 25832
rect 6779 25792 7104 25820
rect 6779 25789 6791 25792
rect 6733 25783 6791 25789
rect 7098 25780 7104 25792
rect 7156 25780 7162 25832
rect 6638 25712 6644 25764
rect 6696 25752 6702 25764
rect 8036 25752 8064 25851
rect 8294 25848 8300 25900
rect 8352 25848 8358 25900
rect 9600 25897 9628 25928
rect 10042 25916 10048 25928
rect 10100 25916 10106 25968
rect 13446 25916 13452 25968
rect 13504 25916 13510 25968
rect 15010 25956 15016 25968
rect 14674 25928 15016 25956
rect 15010 25916 15016 25928
rect 15068 25916 15074 25968
rect 17402 25916 17408 25968
rect 17460 25916 17466 25968
rect 18046 25916 18052 25968
rect 18104 25916 18110 25968
rect 19150 25916 19156 25968
rect 19208 25956 19214 25968
rect 20441 25959 20499 25965
rect 19208 25928 20208 25956
rect 19208 25916 19214 25928
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25857 8539 25891
rect 8665 25891 8723 25897
rect 8665 25888 8677 25891
rect 8481 25851 8539 25857
rect 8588 25860 8677 25888
rect 8202 25780 8208 25832
rect 8260 25820 8266 25832
rect 8496 25820 8524 25851
rect 8260 25792 8524 25820
rect 8260 25780 8266 25792
rect 8588 25752 8616 25860
rect 8665 25857 8677 25860
rect 8711 25857 8723 25891
rect 8665 25851 8723 25857
rect 9585 25891 9643 25897
rect 9585 25857 9597 25891
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 9674 25848 9680 25900
rect 9732 25848 9738 25900
rect 9766 25848 9772 25900
rect 9824 25888 9830 25900
rect 9933 25891 9991 25897
rect 9933 25888 9945 25891
rect 9824 25860 9945 25888
rect 9824 25848 9830 25860
rect 9933 25857 9945 25860
rect 9979 25857 9991 25891
rect 9933 25851 9991 25857
rect 14734 25848 14740 25900
rect 14792 25888 14798 25900
rect 16666 25888 16672 25900
rect 14792 25860 16672 25888
rect 14792 25848 14798 25860
rect 16666 25848 16672 25860
rect 16724 25848 16730 25900
rect 20180 25897 20208 25928
rect 20441 25925 20453 25959
rect 20487 25956 20499 25959
rect 20898 25956 20904 25968
rect 20487 25928 20904 25956
rect 20487 25925 20499 25928
rect 20441 25919 20499 25925
rect 20898 25916 20904 25928
rect 20956 25956 20962 25968
rect 21266 25956 21272 25968
rect 20956 25928 21272 25956
rect 20956 25916 20962 25928
rect 21266 25916 21272 25928
rect 21324 25916 21330 25968
rect 25323 25956 25351 25996
rect 21376 25928 24256 25956
rect 20165 25891 20223 25897
rect 20165 25857 20177 25891
rect 20211 25857 20223 25891
rect 20165 25851 20223 25857
rect 20254 25848 20260 25900
rect 20312 25888 20318 25900
rect 20349 25891 20407 25897
rect 20349 25888 20361 25891
rect 20312 25860 20361 25888
rect 20312 25848 20318 25860
rect 20349 25857 20361 25860
rect 20395 25857 20407 25891
rect 20349 25851 20407 25857
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25888 20591 25891
rect 21376 25888 21404 25928
rect 20579 25860 21404 25888
rect 20579 25857 20591 25860
rect 20533 25851 20591 25857
rect 13173 25823 13231 25829
rect 13173 25789 13185 25823
rect 13219 25820 13231 25823
rect 14090 25820 14096 25832
rect 13219 25792 14096 25820
rect 13219 25789 13231 25792
rect 13173 25783 13231 25789
rect 14090 25780 14096 25792
rect 14148 25780 14154 25832
rect 14458 25780 14464 25832
rect 14516 25820 14522 25832
rect 16390 25820 16396 25832
rect 14516 25792 16396 25820
rect 14516 25780 14522 25792
rect 16390 25780 16396 25792
rect 16448 25780 16454 25832
rect 17126 25780 17132 25832
rect 17184 25780 17190 25832
rect 18414 25780 18420 25832
rect 18472 25820 18478 25832
rect 19153 25823 19211 25829
rect 19153 25820 19165 25823
rect 18472 25792 19165 25820
rect 18472 25780 18478 25792
rect 19153 25789 19165 25792
rect 19199 25789 19211 25823
rect 20548 25820 20576 25851
rect 23382 25848 23388 25900
rect 23440 25888 23446 25900
rect 23937 25891 23995 25897
rect 23937 25888 23949 25891
rect 23440 25860 23949 25888
rect 23440 25848 23446 25860
rect 23937 25857 23949 25860
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 19153 25783 19211 25789
rect 19306 25792 20576 25820
rect 9306 25752 9312 25764
rect 6696 25724 9312 25752
rect 6696 25712 6702 25724
rect 9306 25712 9312 25724
rect 9364 25712 9370 25764
rect 18782 25712 18788 25764
rect 18840 25752 18846 25764
rect 19306 25752 19334 25792
rect 21542 25780 21548 25832
rect 21600 25820 21606 25832
rect 22281 25823 22339 25829
rect 22281 25820 22293 25823
rect 21600 25792 22293 25820
rect 21600 25780 21606 25792
rect 22281 25789 22293 25792
rect 22327 25789 22339 25823
rect 22281 25783 22339 25789
rect 22465 25823 22523 25829
rect 22465 25789 22477 25823
rect 22511 25820 22523 25823
rect 23474 25820 23480 25832
rect 22511 25792 23480 25820
rect 22511 25789 22523 25792
rect 22465 25783 22523 25789
rect 18840 25724 19334 25752
rect 18840 25712 18846 25724
rect 20346 25712 20352 25764
rect 20404 25752 20410 25764
rect 22480 25752 22508 25783
rect 23474 25780 23480 25792
rect 23532 25780 23538 25832
rect 23566 25780 23572 25832
rect 23624 25820 23630 25832
rect 23842 25820 23848 25832
rect 23624 25792 23848 25820
rect 23624 25780 23630 25792
rect 23842 25780 23848 25792
rect 23900 25780 23906 25832
rect 20404 25724 22508 25752
rect 20404 25712 20410 25724
rect 7466 25684 7472 25696
rect 5184 25656 7472 25684
rect 4709 25647 4767 25653
rect 7466 25644 7472 25656
rect 7524 25644 7530 25696
rect 8846 25644 8852 25696
rect 8904 25644 8910 25696
rect 11054 25644 11060 25696
rect 11112 25684 11118 25696
rect 12250 25684 12256 25696
rect 11112 25656 12256 25684
rect 11112 25644 11118 25656
rect 12250 25644 12256 25656
rect 12308 25644 12314 25696
rect 17034 25644 17040 25696
rect 17092 25684 17098 25696
rect 17954 25684 17960 25696
rect 17092 25656 17960 25684
rect 17092 25644 17098 25656
rect 17954 25644 17960 25656
rect 18012 25644 18018 25696
rect 18598 25644 18604 25696
rect 18656 25684 18662 25696
rect 19150 25684 19156 25696
rect 18656 25656 19156 25684
rect 18656 25644 18662 25656
rect 19150 25644 19156 25656
rect 19208 25684 19214 25696
rect 22094 25684 22100 25696
rect 19208 25656 22100 25684
rect 19208 25644 19214 25656
rect 22094 25644 22100 25656
rect 22152 25684 22158 25696
rect 23014 25684 23020 25696
rect 22152 25656 23020 25684
rect 22152 25644 22158 25656
rect 23014 25644 23020 25656
rect 23072 25644 23078 25696
rect 23569 25687 23627 25693
rect 23569 25653 23581 25687
rect 23615 25684 23627 25687
rect 23658 25684 23664 25696
rect 23615 25656 23664 25684
rect 23615 25653 23627 25656
rect 23569 25647 23627 25653
rect 23658 25644 23664 25656
rect 23716 25644 23722 25696
rect 23842 25644 23848 25696
rect 23900 25644 23906 25696
rect 24228 25693 24256 25928
rect 24688 25928 24992 25956
rect 24394 25848 24400 25900
rect 24452 25888 24458 25900
rect 24688 25888 24716 25928
rect 24452 25860 24716 25888
rect 24765 25891 24823 25897
rect 24452 25848 24458 25860
rect 24765 25857 24777 25891
rect 24811 25857 24823 25891
rect 24765 25851 24823 25857
rect 24780 25820 24808 25851
rect 24854 25848 24860 25900
rect 24912 25848 24918 25900
rect 24412 25792 24808 25820
rect 24964 25820 24992 25928
rect 25148 25928 25351 25956
rect 25777 25959 25835 25965
rect 25038 25848 25044 25900
rect 25096 25848 25102 25900
rect 25148 25820 25176 25928
rect 25777 25925 25789 25959
rect 25823 25956 25835 25959
rect 26160 25956 26188 25996
rect 27154 25984 27160 26036
rect 27212 25984 27218 26036
rect 31573 26027 31631 26033
rect 28966 25996 29224 26024
rect 28966 25956 28994 25996
rect 25823 25928 26096 25956
rect 26160 25928 28994 25956
rect 29196 25956 29224 25996
rect 31573 25993 31585 26027
rect 31619 26024 31631 26027
rect 32214 26024 32220 26036
rect 31619 25996 32220 26024
rect 31619 25993 31631 25996
rect 31573 25987 31631 25993
rect 32214 25984 32220 25996
rect 32272 25984 32278 26036
rect 34790 26024 34796 26036
rect 32416 25996 34796 26024
rect 29196 25928 32168 25956
rect 25823 25925 25835 25928
rect 25777 25919 25835 25925
rect 25406 25897 25412 25900
rect 25377 25891 25412 25897
rect 25377 25857 25389 25891
rect 25377 25851 25412 25857
rect 25406 25848 25412 25851
rect 25464 25848 25470 25900
rect 25498 25848 25504 25900
rect 25556 25848 25562 25900
rect 25682 25848 25688 25900
rect 25740 25848 25746 25900
rect 25866 25848 25872 25900
rect 25924 25848 25930 25900
rect 25958 25848 25964 25900
rect 26016 25848 26022 25900
rect 26068 25897 26096 25928
rect 26054 25891 26112 25897
rect 26054 25857 26066 25891
rect 26100 25857 26112 25891
rect 26054 25851 26112 25857
rect 26142 25848 26148 25900
rect 26200 25888 26206 25900
rect 26237 25891 26295 25897
rect 26237 25888 26249 25891
rect 26200 25860 26249 25888
rect 26200 25848 26206 25860
rect 26237 25857 26249 25860
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 26326 25848 26332 25900
rect 26384 25848 26390 25900
rect 26426 25891 26484 25897
rect 26426 25857 26438 25891
rect 26472 25888 26484 25891
rect 26472 25860 26556 25888
rect 26472 25857 26484 25860
rect 26426 25851 26484 25857
rect 24964 25792 25176 25820
rect 24412 25764 24440 25792
rect 25590 25780 25596 25832
rect 25648 25780 25654 25832
rect 25774 25780 25780 25832
rect 25832 25820 25838 25832
rect 26528 25820 26556 25860
rect 26970 25848 26976 25900
rect 27028 25848 27034 25900
rect 28718 25848 28724 25900
rect 28776 25848 28782 25900
rect 28810 25848 28816 25900
rect 28868 25848 28874 25900
rect 28902 25848 28908 25900
rect 28960 25848 28966 25900
rect 29043 25891 29101 25897
rect 29043 25857 29055 25891
rect 29089 25857 29101 25891
rect 29043 25851 29101 25857
rect 29457 25891 29515 25897
rect 29457 25857 29469 25891
rect 29503 25888 29515 25891
rect 30006 25888 30012 25900
rect 29503 25860 30012 25888
rect 29503 25857 29515 25860
rect 29457 25851 29515 25857
rect 25832 25792 26556 25820
rect 25832 25780 25838 25792
rect 24394 25712 24400 25764
rect 24452 25712 24458 25764
rect 24854 25752 24860 25764
rect 24688 25724 24860 25752
rect 24213 25687 24271 25693
rect 24213 25653 24225 25687
rect 24259 25684 24271 25687
rect 24688 25684 24716 25724
rect 24854 25712 24860 25724
rect 24912 25712 24918 25764
rect 24946 25712 24952 25764
rect 25004 25752 25010 25764
rect 25041 25755 25099 25761
rect 25041 25752 25053 25755
rect 25004 25724 25053 25752
rect 25004 25712 25010 25724
rect 25041 25721 25053 25724
rect 25087 25721 25099 25755
rect 25041 25715 25099 25721
rect 25130 25712 25136 25764
rect 25188 25752 25194 25764
rect 25792 25752 25820 25780
rect 25188 25724 25820 25752
rect 26528 25752 26556 25792
rect 26602 25780 26608 25832
rect 26660 25820 26666 25832
rect 28920 25820 28948 25848
rect 26660 25792 28948 25820
rect 26660 25780 26666 25792
rect 29058 25764 29086 25851
rect 30006 25848 30012 25860
rect 30064 25848 30070 25900
rect 30161 25891 30219 25897
rect 30161 25857 30173 25891
rect 30207 25888 30219 25891
rect 30207 25857 30236 25888
rect 30161 25851 30236 25857
rect 29181 25823 29239 25829
rect 29181 25789 29193 25823
rect 29227 25820 29239 25823
rect 29270 25820 29276 25832
rect 29227 25792 29276 25820
rect 29227 25789 29239 25792
rect 29181 25783 29239 25789
rect 29270 25780 29276 25792
rect 29328 25780 29334 25832
rect 29546 25780 29552 25832
rect 29604 25780 29610 25832
rect 29656 25792 30144 25820
rect 29058 25752 29092 25764
rect 26528 25724 29092 25752
rect 25188 25712 25194 25724
rect 29086 25712 29092 25724
rect 29144 25712 29150 25764
rect 24259 25656 24716 25684
rect 24259 25653 24271 25656
rect 24213 25647 24271 25653
rect 24762 25644 24768 25696
rect 24820 25684 24826 25696
rect 25958 25684 25964 25696
rect 24820 25656 25964 25684
rect 24820 25644 24826 25656
rect 25958 25644 25964 25656
rect 26016 25644 26022 25696
rect 26602 25644 26608 25696
rect 26660 25644 26666 25696
rect 28534 25644 28540 25696
rect 28592 25644 28598 25696
rect 28718 25644 28724 25696
rect 28776 25684 28782 25696
rect 29656 25684 29684 25792
rect 29825 25755 29883 25761
rect 29825 25721 29837 25755
rect 29871 25752 29883 25755
rect 30006 25752 30012 25764
rect 29871 25724 30012 25752
rect 29871 25721 29883 25724
rect 29825 25715 29883 25721
rect 30006 25712 30012 25724
rect 30064 25712 30070 25764
rect 28776 25656 29684 25684
rect 28776 25644 28782 25656
rect 29730 25644 29736 25696
rect 29788 25684 29794 25696
rect 29917 25687 29975 25693
rect 29917 25684 29929 25687
rect 29788 25656 29929 25684
rect 29788 25644 29794 25656
rect 29917 25653 29929 25656
rect 29963 25653 29975 25687
rect 30116 25684 30144 25792
rect 30208 25752 30236 25851
rect 30374 25848 30380 25900
rect 30432 25888 30438 25900
rect 31386 25888 31392 25900
rect 30432 25860 31392 25888
rect 30432 25848 30438 25860
rect 31386 25848 31392 25860
rect 31444 25848 31450 25900
rect 31665 25891 31723 25897
rect 31665 25857 31677 25891
rect 31711 25888 31723 25891
rect 32030 25888 32036 25900
rect 31711 25860 32036 25888
rect 31711 25857 31723 25860
rect 31665 25851 31723 25857
rect 32030 25848 32036 25860
rect 32088 25848 32094 25900
rect 32140 25897 32168 25928
rect 32416 25897 32444 25996
rect 32677 25959 32735 25965
rect 32677 25925 32689 25959
rect 32723 25956 32735 25959
rect 32950 25956 32956 25968
rect 32723 25928 32956 25956
rect 32723 25925 32735 25928
rect 32677 25919 32735 25925
rect 32950 25916 32956 25928
rect 33008 25916 33014 25968
rect 34146 25916 34152 25968
rect 34204 25916 34210 25968
rect 34440 25956 34468 25996
rect 34790 25984 34796 25996
rect 34848 26024 34854 26036
rect 35342 26024 35348 26036
rect 34848 25996 35348 26024
rect 34848 25984 34854 25996
rect 35342 25984 35348 25996
rect 35400 25984 35406 26036
rect 36722 25984 36728 26036
rect 36780 26024 36786 26036
rect 38657 26027 38715 26033
rect 36780 25996 37688 26024
rect 36780 25984 36786 25996
rect 34348 25928 34468 25956
rect 32125 25891 32183 25897
rect 32125 25857 32137 25891
rect 32171 25857 32183 25891
rect 32125 25851 32183 25857
rect 32401 25891 32459 25897
rect 32401 25857 32413 25891
rect 32447 25857 32459 25891
rect 34164 25888 34192 25916
rect 34348 25897 34376 25928
rect 34333 25891 34391 25897
rect 33810 25860 34284 25888
rect 32401 25851 32459 25857
rect 31754 25780 31760 25832
rect 31812 25780 31818 25832
rect 33686 25780 33692 25832
rect 33744 25820 33750 25832
rect 34146 25820 34152 25832
rect 33744 25792 34152 25820
rect 33744 25780 33750 25792
rect 34146 25780 34152 25792
rect 34204 25780 34210 25832
rect 30374 25752 30380 25764
rect 30208 25724 30380 25752
rect 30374 25712 30380 25724
rect 30432 25712 30438 25764
rect 30285 25687 30343 25693
rect 30285 25684 30297 25687
rect 30116 25656 30297 25684
rect 29917 25647 29975 25653
rect 30285 25653 30297 25656
rect 30331 25653 30343 25687
rect 30285 25647 30343 25653
rect 31202 25644 31208 25696
rect 31260 25644 31266 25696
rect 32309 25687 32367 25693
rect 32309 25653 32321 25687
rect 32355 25684 32367 25687
rect 32490 25684 32496 25696
rect 32355 25656 32496 25684
rect 32355 25653 32367 25656
rect 32309 25647 32367 25653
rect 32490 25644 32496 25656
rect 32548 25644 32554 25696
rect 32766 25644 32772 25696
rect 32824 25684 32830 25696
rect 34256 25684 34284 25860
rect 34333 25857 34345 25891
rect 34379 25857 34391 25891
rect 36633 25891 36691 25897
rect 35742 25874 36492 25888
rect 34333 25851 34391 25857
rect 35728 25860 36492 25874
rect 34606 25780 34612 25832
rect 34664 25780 34670 25832
rect 35728 25684 35756 25860
rect 36357 25823 36415 25829
rect 36357 25789 36369 25823
rect 36403 25789 36415 25823
rect 36464 25820 36492 25860
rect 36633 25857 36645 25891
rect 36679 25888 36691 25891
rect 36740 25888 36768 25984
rect 37660 25965 37688 25996
rect 38657 25993 38669 26027
rect 38703 26024 38715 26027
rect 39206 26024 39212 26036
rect 38703 25996 39212 26024
rect 38703 25993 38715 25996
rect 38657 25987 38715 25993
rect 39206 25984 39212 25996
rect 39264 25984 39270 26036
rect 41598 25984 41604 26036
rect 41656 26024 41662 26036
rect 42153 26027 42211 26033
rect 42153 26024 42165 26027
rect 41656 25996 42165 26024
rect 41656 25984 41662 25996
rect 42153 25993 42165 25996
rect 42199 25993 42211 26027
rect 42153 25987 42211 25993
rect 37001 25959 37059 25965
rect 37001 25925 37013 25959
rect 37047 25956 37059 25959
rect 37553 25959 37611 25965
rect 37553 25956 37565 25959
rect 37047 25928 37565 25956
rect 37047 25925 37059 25928
rect 37001 25919 37059 25925
rect 37553 25925 37565 25928
rect 37599 25925 37611 25959
rect 37553 25919 37611 25925
rect 37645 25959 37703 25965
rect 37645 25925 37657 25959
rect 37691 25925 37703 25959
rect 37645 25919 37703 25925
rect 38933 25959 38991 25965
rect 38933 25925 38945 25959
rect 38979 25956 38991 25959
rect 39482 25956 39488 25968
rect 38979 25928 39488 25956
rect 38979 25925 38991 25928
rect 38933 25919 38991 25925
rect 39482 25916 39488 25928
rect 39540 25916 39546 25968
rect 41414 25916 41420 25968
rect 41472 25916 41478 25968
rect 36679 25860 36768 25888
rect 36679 25857 36691 25860
rect 36633 25851 36691 25857
rect 36906 25848 36912 25900
rect 36964 25848 36970 25900
rect 37366 25848 37372 25900
rect 37424 25888 37430 25900
rect 37461 25891 37519 25897
rect 37461 25888 37473 25891
rect 37424 25860 37473 25888
rect 37424 25848 37430 25860
rect 37461 25857 37473 25860
rect 37507 25857 37519 25891
rect 37763 25891 37821 25897
rect 37763 25888 37775 25891
rect 37461 25851 37519 25857
rect 37752 25857 37775 25888
rect 37809 25857 37821 25891
rect 37752 25851 37821 25857
rect 38841 25891 38899 25897
rect 38841 25857 38853 25891
rect 38887 25857 38899 25891
rect 38841 25851 38899 25857
rect 36998 25820 37004 25832
rect 36464 25792 37004 25820
rect 36357 25783 36415 25789
rect 36372 25752 36400 25783
rect 36998 25780 37004 25792
rect 37056 25780 37062 25832
rect 37550 25780 37556 25832
rect 37608 25820 37614 25832
rect 37752 25820 37780 25851
rect 37608 25792 37780 25820
rect 37921 25823 37979 25829
rect 37608 25780 37614 25792
rect 37921 25789 37933 25823
rect 37967 25820 37979 25823
rect 38102 25820 38108 25832
rect 37967 25792 38108 25820
rect 37967 25789 37979 25792
rect 37921 25783 37979 25789
rect 38102 25780 38108 25792
rect 38160 25820 38166 25832
rect 38562 25820 38568 25832
rect 38160 25792 38568 25820
rect 38160 25780 38166 25792
rect 38562 25780 38568 25792
rect 38620 25780 38626 25832
rect 38856 25820 38884 25851
rect 39022 25848 39028 25900
rect 39080 25848 39086 25900
rect 39209 25891 39267 25897
rect 39209 25857 39221 25891
rect 39255 25888 39267 25891
rect 40218 25888 40224 25900
rect 39255 25860 40224 25888
rect 39255 25857 39267 25860
rect 39209 25851 39267 25857
rect 40218 25848 40224 25860
rect 40276 25848 40282 25900
rect 40313 25891 40371 25897
rect 40313 25857 40325 25891
rect 40359 25857 40371 25891
rect 40313 25851 40371 25857
rect 40126 25820 40132 25832
rect 38856 25792 40132 25820
rect 40126 25780 40132 25792
rect 40184 25780 40190 25832
rect 38470 25752 38476 25764
rect 36372 25724 38476 25752
rect 38470 25712 38476 25724
rect 38528 25712 38534 25764
rect 32824 25656 35756 25684
rect 32824 25644 32830 25656
rect 36078 25644 36084 25696
rect 36136 25644 36142 25696
rect 36262 25644 36268 25696
rect 36320 25684 36326 25696
rect 36449 25687 36507 25693
rect 36449 25684 36461 25687
rect 36320 25656 36461 25684
rect 36320 25644 36326 25656
rect 36449 25653 36461 25656
rect 36495 25653 36507 25687
rect 36449 25647 36507 25653
rect 36817 25687 36875 25693
rect 36817 25653 36829 25687
rect 36863 25684 36875 25687
rect 37090 25684 37096 25696
rect 36863 25656 37096 25684
rect 36863 25653 36875 25656
rect 36817 25647 36875 25653
rect 37090 25644 37096 25656
rect 37148 25644 37154 25696
rect 37274 25644 37280 25696
rect 37332 25644 37338 25696
rect 40126 25644 40132 25696
rect 40184 25644 40190 25696
rect 40328 25684 40356 25851
rect 40402 25780 40408 25832
rect 40460 25780 40466 25832
rect 40681 25823 40739 25829
rect 40681 25789 40693 25823
rect 40727 25820 40739 25823
rect 41138 25820 41144 25832
rect 40727 25792 41144 25820
rect 40727 25789 40739 25792
rect 40681 25783 40739 25789
rect 41138 25780 41144 25792
rect 41196 25780 41202 25832
rect 42058 25684 42064 25696
rect 40328 25656 42064 25684
rect 42058 25644 42064 25656
rect 42116 25644 42122 25696
rect 1104 25594 42504 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 42504 25594
rect 1104 25520 42504 25542
rect 5258 25480 5264 25492
rect 3252 25452 5264 25480
rect 3252 25344 3280 25452
rect 5258 25440 5264 25452
rect 5316 25440 5322 25492
rect 7558 25440 7564 25492
rect 7616 25440 7622 25492
rect 10042 25440 10048 25492
rect 10100 25480 10106 25492
rect 10321 25483 10379 25489
rect 10321 25480 10333 25483
rect 10100 25452 10333 25480
rect 10100 25440 10106 25452
rect 10321 25449 10333 25452
rect 10367 25449 10379 25483
rect 10321 25443 10379 25449
rect 11422 25440 11428 25492
rect 11480 25480 11486 25492
rect 17494 25480 17500 25492
rect 11480 25452 17500 25480
rect 11480 25440 11486 25452
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 17678 25440 17684 25492
rect 17736 25480 17742 25492
rect 17865 25483 17923 25489
rect 17865 25480 17877 25483
rect 17736 25452 17877 25480
rect 17736 25440 17742 25452
rect 17865 25449 17877 25452
rect 17911 25449 17923 25483
rect 17865 25443 17923 25449
rect 20254 25440 20260 25492
rect 20312 25440 20318 25492
rect 21542 25440 21548 25492
rect 21600 25440 21606 25492
rect 22094 25480 22100 25492
rect 22020 25452 22100 25480
rect 14366 25372 14372 25424
rect 14424 25412 14430 25424
rect 16758 25412 16764 25424
rect 14424 25384 16764 25412
rect 14424 25372 14430 25384
rect 16758 25372 16764 25384
rect 16816 25372 16822 25424
rect 17402 25412 17408 25424
rect 17328 25384 17408 25412
rect 3160 25316 3280 25344
rect 3789 25347 3847 25353
rect 3160 25285 3188 25316
rect 3789 25313 3801 25347
rect 3835 25344 3847 25347
rect 4154 25344 4160 25356
rect 3835 25316 4160 25344
rect 3835 25313 3847 25316
rect 3789 25307 3847 25313
rect 4154 25304 4160 25316
rect 4212 25344 4218 25356
rect 4614 25344 4620 25356
rect 4212 25316 4620 25344
rect 4212 25304 4218 25316
rect 4614 25304 4620 25316
rect 4672 25344 4678 25356
rect 6181 25347 6239 25353
rect 6181 25344 6193 25347
rect 4672 25316 6193 25344
rect 4672 25304 4678 25316
rect 6181 25313 6193 25316
rect 6227 25313 6239 25347
rect 6181 25307 6239 25313
rect 11698 25304 11704 25356
rect 11756 25344 11762 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 11756 25316 12265 25344
rect 11756 25304 11762 25316
rect 12253 25313 12265 25316
rect 12299 25344 12311 25347
rect 12434 25344 12440 25356
rect 12299 25316 12440 25344
rect 12299 25313 12311 25316
rect 12253 25307 12311 25313
rect 12434 25304 12440 25316
rect 12492 25344 12498 25356
rect 13170 25344 13176 25356
rect 12492 25316 13176 25344
rect 12492 25304 12498 25316
rect 13170 25304 13176 25316
rect 13228 25304 13234 25356
rect 15381 25347 15439 25353
rect 15381 25313 15393 25347
rect 15427 25344 15439 25347
rect 16393 25347 16451 25353
rect 16393 25344 16405 25347
rect 15427 25316 16405 25344
rect 15427 25313 15439 25316
rect 15381 25307 15439 25313
rect 16393 25313 16405 25316
rect 16439 25313 16451 25347
rect 16393 25307 16451 25313
rect 16666 25304 16672 25356
rect 16724 25344 16730 25356
rect 16724 25316 16804 25344
rect 16724 25304 16730 25316
rect 3145 25279 3203 25285
rect 3145 25245 3157 25279
rect 3191 25245 3203 25279
rect 3145 25239 3203 25245
rect 3237 25279 3295 25285
rect 3237 25245 3249 25279
rect 3283 25245 3295 25279
rect 3237 25239 3295 25245
rect 3329 25279 3387 25285
rect 3329 25245 3341 25279
rect 3375 25276 3387 25279
rect 3418 25276 3424 25288
rect 3375 25248 3424 25276
rect 3375 25245 3387 25248
rect 3329 25239 3387 25245
rect 2866 25100 2872 25152
rect 2924 25100 2930 25152
rect 3252 25140 3280 25239
rect 3418 25236 3424 25248
rect 3476 25236 3482 25288
rect 3510 25236 3516 25288
rect 3568 25236 3574 25288
rect 5350 25276 5356 25288
rect 5198 25248 5356 25276
rect 5350 25236 5356 25248
rect 5408 25276 5414 25288
rect 6270 25276 6276 25288
rect 5408 25248 6276 25276
rect 5408 25236 5414 25248
rect 6270 25236 6276 25248
rect 6328 25236 6334 25288
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25276 8999 25279
rect 9674 25276 9680 25288
rect 8987 25248 9680 25276
rect 8987 25245 8999 25248
rect 8941 25239 8999 25245
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 15102 25236 15108 25288
rect 15160 25236 15166 25288
rect 15197 25279 15255 25285
rect 15197 25245 15209 25279
rect 15243 25245 15255 25279
rect 15197 25239 15255 25245
rect 4062 25168 4068 25220
rect 4120 25168 4126 25220
rect 6454 25217 6460 25220
rect 6448 25171 6460 25217
rect 6454 25168 6460 25171
rect 6512 25168 6518 25220
rect 8846 25168 8852 25220
rect 8904 25208 8910 25220
rect 9186 25211 9244 25217
rect 9186 25208 9198 25211
rect 8904 25180 9198 25208
rect 8904 25168 8910 25180
rect 9186 25177 9198 25180
rect 9232 25177 9244 25211
rect 9186 25171 9244 25177
rect 11422 25168 11428 25220
rect 11480 25208 11486 25220
rect 11977 25211 12035 25217
rect 11977 25208 11989 25211
rect 11480 25180 11989 25208
rect 11480 25168 11486 25180
rect 11977 25177 11989 25180
rect 12023 25177 12035 25211
rect 15212 25208 15240 25239
rect 15470 25236 15476 25288
rect 15528 25236 15534 25288
rect 15562 25236 15568 25288
rect 15620 25276 15626 25288
rect 16022 25276 16028 25288
rect 15620 25248 16028 25276
rect 15620 25236 15626 25248
rect 16022 25236 16028 25248
rect 16080 25276 16086 25288
rect 16209 25279 16267 25285
rect 16209 25276 16221 25279
rect 16080 25248 16221 25276
rect 16080 25236 16086 25248
rect 16209 25245 16221 25248
rect 16255 25245 16267 25279
rect 16209 25239 16267 25245
rect 16574 25236 16580 25288
rect 16632 25236 16638 25288
rect 16776 25276 16804 25316
rect 17034 25304 17040 25356
rect 17092 25304 17098 25356
rect 17221 25347 17279 25353
rect 17221 25313 17233 25347
rect 17267 25344 17279 25347
rect 17328 25344 17356 25384
rect 17402 25372 17408 25384
rect 17460 25372 17466 25424
rect 17586 25372 17592 25424
rect 17644 25412 17650 25424
rect 17773 25415 17831 25421
rect 17773 25412 17785 25415
rect 17644 25384 17785 25412
rect 17644 25372 17650 25384
rect 17773 25381 17785 25384
rect 17819 25381 17831 25415
rect 17773 25375 17831 25381
rect 17267 25316 17356 25344
rect 17267 25313 17279 25316
rect 17221 25307 17279 25313
rect 17954 25304 17960 25356
rect 18012 25344 18018 25356
rect 18230 25344 18236 25356
rect 18012 25316 18236 25344
rect 18012 25304 18018 25316
rect 16879 25279 16937 25285
rect 16879 25278 16891 25279
rect 16868 25276 16891 25278
rect 16776 25248 16891 25276
rect 16879 25245 16891 25248
rect 16925 25245 16937 25279
rect 16879 25239 16937 25245
rect 17129 25279 17187 25285
rect 17129 25245 17141 25279
rect 17175 25276 17187 25279
rect 17313 25279 17371 25285
rect 17175 25248 17264 25276
rect 17175 25245 17187 25248
rect 17129 25239 17187 25245
rect 15657 25211 15715 25217
rect 15657 25208 15669 25211
rect 15212 25180 15669 25208
rect 11977 25171 12035 25177
rect 15657 25177 15669 25180
rect 15703 25177 15715 25211
rect 15657 25171 15715 25177
rect 16666 25168 16672 25220
rect 16724 25168 16730 25220
rect 16758 25168 16764 25220
rect 16816 25168 16822 25220
rect 3418 25140 3424 25152
rect 3252 25112 3424 25140
rect 3418 25100 3424 25112
rect 3476 25140 3482 25152
rect 3970 25140 3976 25152
rect 3476 25112 3976 25140
rect 3476 25100 3482 25112
rect 3970 25100 3976 25112
rect 4028 25100 4034 25152
rect 5537 25143 5595 25149
rect 5537 25109 5549 25143
rect 5583 25140 5595 25143
rect 5626 25140 5632 25152
rect 5583 25112 5632 25140
rect 5583 25109 5595 25112
rect 5537 25103 5595 25109
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 11609 25143 11667 25149
rect 11609 25109 11621 25143
rect 11655 25140 11667 25143
rect 11790 25140 11796 25152
rect 11655 25112 11796 25140
rect 11655 25109 11667 25112
rect 11609 25103 11667 25109
rect 11790 25100 11796 25112
rect 11848 25100 11854 25152
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 13354 25140 13360 25152
rect 12115 25112 13360 25140
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 13354 25100 13360 25112
rect 13412 25100 13418 25152
rect 14550 25100 14556 25152
rect 14608 25140 14614 25152
rect 14921 25143 14979 25149
rect 14921 25140 14933 25143
rect 14608 25112 14933 25140
rect 14608 25100 14614 25112
rect 14921 25109 14933 25112
rect 14967 25109 14979 25143
rect 17236 25140 17264 25248
rect 17313 25245 17325 25279
rect 17359 25245 17371 25279
rect 17313 25239 17371 25245
rect 17328 25208 17356 25239
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 18064 25285 18092 25316
rect 18230 25304 18236 25316
rect 18288 25304 18294 25356
rect 18322 25304 18328 25356
rect 18380 25344 18386 25356
rect 18506 25344 18512 25356
rect 18380 25316 18512 25344
rect 18380 25304 18386 25316
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 17589 25279 17647 25285
rect 17589 25245 17601 25279
rect 17635 25276 17647 25279
rect 18049 25279 18107 25285
rect 17635 25248 18000 25276
rect 17635 25245 17647 25248
rect 17589 25239 17647 25245
rect 17678 25208 17684 25220
rect 17328 25180 17684 25208
rect 17678 25168 17684 25180
rect 17736 25168 17742 25220
rect 17972 25208 18000 25248
rect 18049 25245 18061 25279
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 18138 25236 18144 25288
rect 18196 25236 18202 25288
rect 18414 25236 18420 25288
rect 18472 25236 18478 25288
rect 20254 25236 20260 25288
rect 20312 25236 20318 25288
rect 20441 25279 20499 25285
rect 20441 25245 20453 25279
rect 20487 25276 20499 25279
rect 20990 25276 20996 25288
rect 20487 25248 20996 25276
rect 20487 25245 20499 25248
rect 20441 25239 20499 25245
rect 20990 25236 20996 25248
rect 21048 25236 21054 25288
rect 21726 25236 21732 25288
rect 21784 25236 21790 25288
rect 21913 25279 21971 25285
rect 21913 25245 21925 25279
rect 21959 25276 21971 25279
rect 22020 25276 22048 25452
rect 22094 25440 22100 25452
rect 22152 25440 22158 25492
rect 23201 25483 23259 25489
rect 23201 25449 23213 25483
rect 23247 25480 23259 25483
rect 23842 25480 23848 25492
rect 23247 25452 23848 25480
rect 23247 25449 23259 25452
rect 23201 25443 23259 25449
rect 23842 25440 23848 25452
rect 23900 25440 23906 25492
rect 25317 25483 25375 25489
rect 25317 25449 25329 25483
rect 25363 25480 25375 25483
rect 25866 25480 25872 25492
rect 25363 25452 25872 25480
rect 25363 25449 25375 25452
rect 25317 25443 25375 25449
rect 25866 25440 25872 25452
rect 25924 25440 25930 25492
rect 25961 25483 26019 25489
rect 25961 25449 25973 25483
rect 26007 25480 26019 25483
rect 26142 25480 26148 25492
rect 26007 25452 26148 25480
rect 26007 25449 26019 25452
rect 25961 25443 26019 25449
rect 26142 25440 26148 25452
rect 26200 25440 26206 25492
rect 26252 25452 28764 25480
rect 23385 25415 23443 25421
rect 23385 25381 23397 25415
rect 23431 25412 23443 25415
rect 24394 25412 24400 25424
rect 23431 25384 24400 25412
rect 23431 25381 23443 25384
rect 23385 25375 23443 25381
rect 24394 25372 24400 25384
rect 24452 25412 24458 25424
rect 25590 25412 25596 25424
rect 24452 25384 25596 25412
rect 24452 25372 24458 25384
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 22704 25316 23060 25344
rect 22704 25304 22710 25316
rect 23032 25288 23060 25316
rect 23474 25304 23480 25356
rect 23532 25344 23538 25356
rect 23569 25347 23627 25353
rect 23569 25344 23581 25347
rect 23532 25316 23581 25344
rect 23532 25304 23538 25316
rect 23569 25313 23581 25316
rect 23615 25313 23627 25347
rect 23569 25307 23627 25313
rect 23842 25304 23848 25356
rect 23900 25344 23906 25356
rect 24581 25347 24639 25353
rect 24581 25344 24593 25347
rect 23900 25316 24593 25344
rect 23900 25304 23906 25316
rect 24581 25313 24593 25316
rect 24627 25313 24639 25347
rect 24581 25307 24639 25313
rect 21959 25248 22048 25276
rect 22189 25279 22247 25285
rect 21959 25245 21971 25248
rect 21913 25239 21971 25245
rect 22189 25245 22201 25279
rect 22235 25276 22247 25279
rect 22278 25276 22284 25288
rect 22235 25248 22284 25276
rect 22235 25245 22247 25248
rect 22189 25239 22247 25245
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 22462 25236 22468 25288
rect 22520 25236 22526 25288
rect 22830 25236 22836 25288
rect 22888 25236 22894 25288
rect 23014 25236 23020 25288
rect 23072 25236 23078 25288
rect 23290 25236 23296 25288
rect 23348 25236 23354 25288
rect 23658 25236 23664 25288
rect 23716 25236 23722 25288
rect 23934 25236 23940 25288
rect 23992 25236 23998 25288
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25245 24087 25279
rect 24029 25239 24087 25245
rect 18782 25208 18788 25220
rect 17972 25180 18788 25208
rect 18782 25168 18788 25180
rect 18840 25168 18846 25220
rect 21821 25211 21879 25217
rect 21821 25177 21833 25211
rect 21867 25177 21879 25211
rect 21821 25171 21879 25177
rect 22051 25211 22109 25217
rect 22051 25177 22063 25211
rect 22097 25208 22109 25211
rect 23569 25211 23627 25217
rect 22097 25180 23520 25208
rect 22097 25177 22109 25180
rect 22051 25171 22109 25177
rect 17586 25140 17592 25152
rect 17236 25112 17592 25140
rect 14921 25103 14979 25109
rect 17586 25100 17592 25112
rect 17644 25100 17650 25152
rect 21836 25140 21864 25171
rect 22373 25143 22431 25149
rect 22373 25140 22385 25143
rect 21836 25112 22385 25140
rect 22373 25109 22385 25112
rect 22419 25109 22431 25143
rect 23492 25140 23520 25180
rect 23569 25177 23581 25211
rect 23615 25208 23627 25211
rect 23845 25211 23903 25217
rect 23845 25208 23857 25211
rect 23615 25180 23857 25208
rect 23615 25177 23627 25180
rect 23569 25171 23627 25177
rect 23845 25177 23857 25180
rect 23891 25177 23903 25211
rect 24044 25208 24072 25239
rect 24670 25236 24676 25288
rect 24728 25236 24734 25288
rect 24854 25236 24860 25288
rect 24912 25236 24918 25288
rect 25038 25236 25044 25288
rect 25096 25236 25102 25288
rect 25516 25285 25544 25384
rect 25590 25372 25596 25384
rect 25648 25372 25654 25424
rect 25884 25412 25912 25440
rect 26252 25412 26280 25452
rect 25884 25384 26280 25412
rect 28736 25412 28764 25452
rect 28810 25440 28816 25492
rect 28868 25480 28874 25492
rect 28905 25483 28963 25489
rect 28905 25480 28917 25483
rect 28868 25452 28917 25480
rect 28868 25440 28874 25452
rect 28905 25449 28917 25452
rect 28951 25449 28963 25483
rect 28905 25443 28963 25449
rect 30374 25440 30380 25492
rect 30432 25440 30438 25492
rect 31846 25440 31852 25492
rect 31904 25480 31910 25492
rect 32214 25480 32220 25492
rect 31904 25452 32220 25480
rect 31904 25440 31910 25452
rect 32214 25440 32220 25452
rect 32272 25480 32278 25492
rect 32585 25483 32643 25489
rect 32585 25480 32597 25483
rect 32272 25452 32597 25480
rect 32272 25440 32278 25452
rect 32585 25449 32597 25452
rect 32631 25480 32643 25483
rect 32858 25480 32864 25492
rect 32631 25452 32864 25480
rect 32631 25449 32643 25452
rect 32585 25443 32643 25449
rect 32858 25440 32864 25452
rect 32916 25440 32922 25492
rect 33410 25440 33416 25492
rect 33468 25480 33474 25492
rect 33597 25483 33655 25489
rect 33597 25480 33609 25483
rect 33468 25452 33609 25480
rect 33468 25440 33474 25452
rect 33597 25449 33609 25452
rect 33643 25449 33655 25483
rect 33597 25443 33655 25449
rect 35158 25440 35164 25492
rect 35216 25480 35222 25492
rect 36078 25480 36084 25492
rect 35216 25452 36084 25480
rect 35216 25440 35222 25452
rect 36078 25440 36084 25452
rect 36136 25440 36142 25492
rect 36446 25440 36452 25492
rect 36504 25480 36510 25492
rect 36814 25480 36820 25492
rect 36504 25452 36820 25480
rect 36504 25440 36510 25452
rect 36814 25440 36820 25452
rect 36872 25480 36878 25492
rect 39206 25480 39212 25492
rect 36872 25452 39212 25480
rect 36872 25440 36878 25452
rect 39206 25440 39212 25452
rect 39264 25440 39270 25492
rect 39485 25483 39543 25489
rect 39485 25449 39497 25483
rect 39531 25480 39543 25483
rect 40494 25480 40500 25492
rect 39531 25452 40500 25480
rect 39531 25449 39543 25452
rect 39485 25443 39543 25449
rect 28994 25412 29000 25424
rect 28736 25384 29000 25412
rect 28994 25372 29000 25384
rect 29052 25372 29058 25424
rect 29086 25372 29092 25424
rect 29144 25412 29150 25424
rect 29144 25384 30241 25412
rect 29144 25372 29150 25384
rect 25958 25304 25964 25356
rect 26016 25344 26022 25356
rect 26016 25316 28028 25344
rect 26016 25304 26022 25316
rect 25501 25279 25559 25285
rect 25501 25245 25513 25279
rect 25547 25245 25559 25279
rect 25501 25239 25559 25245
rect 25774 25236 25780 25288
rect 25832 25236 25838 25288
rect 26145 25279 26203 25285
rect 26145 25245 26157 25279
rect 26191 25245 26203 25279
rect 27890 25276 27896 25288
rect 27554 25248 27896 25276
rect 26145 25239 26203 25245
rect 24872 25208 24900 25236
rect 23845 25171 23903 25177
rect 23952 25180 24900 25208
rect 24949 25211 25007 25217
rect 23952 25140 23980 25180
rect 24949 25177 24961 25211
rect 24995 25208 25007 25211
rect 25222 25208 25228 25220
rect 24995 25180 25228 25208
rect 24995 25177 25007 25180
rect 24949 25171 25007 25177
rect 25222 25168 25228 25180
rect 25280 25208 25286 25220
rect 25593 25211 25651 25217
rect 25593 25208 25605 25211
rect 25280 25180 25605 25208
rect 25280 25168 25286 25180
rect 25593 25177 25605 25180
rect 25639 25177 25651 25211
rect 26160 25208 26188 25239
rect 27890 25236 27896 25248
rect 27948 25236 27954 25288
rect 28000 25276 28028 25316
rect 28534 25304 28540 25356
rect 28592 25304 28598 25356
rect 28718 25304 28724 25356
rect 28776 25304 28782 25356
rect 28902 25304 28908 25356
rect 28960 25344 28966 25356
rect 28960 25316 29859 25344
rect 28960 25304 28966 25316
rect 29831 25285 29859 25316
rect 29733 25279 29791 25285
rect 29733 25276 29745 25279
rect 28000 25248 29745 25276
rect 29733 25245 29745 25248
rect 29779 25245 29791 25279
rect 29733 25239 29791 25245
rect 29826 25279 29884 25285
rect 29826 25245 29838 25279
rect 29872 25245 29884 25279
rect 29826 25239 29884 25245
rect 30006 25236 30012 25288
rect 30064 25236 30070 25288
rect 30213 25285 30241 25384
rect 35342 25372 35348 25424
rect 35400 25412 35406 25424
rect 37642 25412 37648 25424
rect 35400 25384 37648 25412
rect 35400 25372 35406 25384
rect 30837 25347 30895 25353
rect 30837 25313 30849 25347
rect 30883 25344 30895 25347
rect 31110 25344 31116 25356
rect 30883 25316 31116 25344
rect 30883 25313 30895 25316
rect 30837 25307 30895 25313
rect 31110 25304 31116 25316
rect 31168 25344 31174 25356
rect 31662 25344 31668 25356
rect 31168 25316 31668 25344
rect 31168 25304 31174 25316
rect 31662 25304 31668 25316
rect 31720 25304 31726 25356
rect 32674 25304 32680 25356
rect 32732 25304 32738 25356
rect 34790 25304 34796 25356
rect 34848 25304 34854 25356
rect 35897 25347 35955 25353
rect 35897 25313 35909 25347
rect 35943 25344 35955 25347
rect 36170 25344 36176 25356
rect 35943 25316 36176 25344
rect 35943 25313 35955 25316
rect 35897 25307 35955 25313
rect 36170 25304 36176 25316
rect 36228 25304 36234 25356
rect 36357 25347 36415 25353
rect 36357 25313 36369 25347
rect 36403 25344 36415 25347
rect 36446 25344 36452 25356
rect 36403 25316 36452 25344
rect 36403 25313 36415 25316
rect 36357 25307 36415 25313
rect 36446 25304 36452 25316
rect 36504 25304 36510 25356
rect 37016 25353 37044 25384
rect 37642 25372 37648 25384
rect 37700 25372 37706 25424
rect 37734 25372 37740 25424
rect 37792 25412 37798 25424
rect 37792 25384 37872 25412
rect 37792 25372 37798 25384
rect 37001 25347 37059 25353
rect 37001 25313 37013 25347
rect 37047 25313 37059 25347
rect 37001 25307 37059 25313
rect 37185 25347 37243 25353
rect 37185 25313 37197 25347
rect 37231 25344 37243 25347
rect 37274 25344 37280 25356
rect 37231 25316 37280 25344
rect 37231 25313 37243 25316
rect 37185 25307 37243 25313
rect 37274 25304 37280 25316
rect 37332 25304 37338 25356
rect 37844 25344 37872 25384
rect 38013 25347 38071 25353
rect 38013 25344 38025 25347
rect 37844 25316 38025 25344
rect 38013 25313 38025 25316
rect 38059 25313 38071 25347
rect 38013 25307 38071 25313
rect 38378 25304 38384 25356
rect 38436 25344 38442 25356
rect 39500 25344 39528 25443
rect 40494 25440 40500 25452
rect 40552 25440 40558 25492
rect 42150 25440 42156 25492
rect 42208 25440 42214 25492
rect 38436 25316 39528 25344
rect 38436 25304 38442 25316
rect 30198 25279 30256 25285
rect 30198 25245 30210 25279
rect 30244 25245 30256 25279
rect 30198 25239 30256 25245
rect 30742 25236 30748 25288
rect 30800 25236 30806 25288
rect 32766 25276 32772 25288
rect 32246 25248 32772 25276
rect 32766 25236 32772 25248
rect 32824 25236 32830 25288
rect 32953 25279 33011 25285
rect 32953 25245 32965 25279
rect 32999 25276 33011 25279
rect 33410 25276 33416 25288
rect 32999 25248 33416 25276
rect 32999 25245 33011 25248
rect 32953 25239 33011 25245
rect 33410 25236 33416 25248
rect 33468 25236 33474 25288
rect 33778 25236 33784 25288
rect 33836 25236 33842 25288
rect 33870 25236 33876 25288
rect 33928 25236 33934 25288
rect 33962 25236 33968 25288
rect 34020 25276 34026 25288
rect 34241 25279 34299 25285
rect 34241 25276 34253 25279
rect 34020 25248 34253 25276
rect 34020 25236 34026 25248
rect 34241 25245 34253 25248
rect 34287 25245 34299 25279
rect 34241 25239 34299 25245
rect 34514 25236 34520 25288
rect 34572 25276 34578 25288
rect 35621 25279 35679 25285
rect 35621 25276 35633 25279
rect 34572 25248 35633 25276
rect 34572 25236 34578 25248
rect 35621 25245 35633 25248
rect 35667 25245 35679 25279
rect 35621 25239 35679 25245
rect 35986 25236 35992 25288
rect 36044 25236 36050 25288
rect 37550 25276 37556 25288
rect 36280 25248 37556 25276
rect 26160 25180 26280 25208
rect 25593 25171 25651 25177
rect 23492 25112 23980 25140
rect 22373 25103 22431 25109
rect 24026 25100 24032 25152
rect 24084 25140 24090 25152
rect 24213 25143 24271 25149
rect 24213 25140 24225 25143
rect 24084 25112 24225 25140
rect 24084 25100 24090 25112
rect 24213 25109 24225 25112
rect 24259 25109 24271 25143
rect 24213 25103 24271 25109
rect 24857 25143 24915 25149
rect 24857 25109 24869 25143
rect 24903 25140 24915 25143
rect 25774 25140 25780 25152
rect 24903 25112 25780 25140
rect 24903 25109 24915 25112
rect 24857 25103 24915 25109
rect 25774 25100 25780 25112
rect 25832 25100 25838 25152
rect 26252 25140 26280 25180
rect 26418 25168 26424 25220
rect 26476 25168 26482 25220
rect 28445 25211 28503 25217
rect 28445 25177 28457 25211
rect 28491 25208 28503 25211
rect 29089 25211 29147 25217
rect 29089 25208 29101 25211
rect 28491 25180 29101 25208
rect 28491 25177 28503 25180
rect 28445 25171 28503 25177
rect 29089 25177 29101 25180
rect 29135 25208 29147 25211
rect 29178 25208 29184 25220
rect 29135 25180 29184 25208
rect 29135 25177 29147 25180
rect 29089 25171 29147 25177
rect 29178 25168 29184 25180
rect 29236 25168 29242 25220
rect 29273 25211 29331 25217
rect 29273 25177 29285 25211
rect 29319 25177 29331 25211
rect 29273 25171 29331 25177
rect 30101 25211 30159 25217
rect 30101 25177 30113 25211
rect 30147 25208 30159 25211
rect 30834 25208 30840 25220
rect 30147 25180 30840 25208
rect 30147 25177 30159 25180
rect 30101 25171 30159 25177
rect 27338 25140 27344 25152
rect 26252 25112 27344 25140
rect 27338 25100 27344 25112
rect 27396 25100 27402 25152
rect 27798 25100 27804 25152
rect 27856 25140 27862 25152
rect 27893 25143 27951 25149
rect 27893 25140 27905 25143
rect 27856 25112 27905 25140
rect 27856 25100 27862 25112
rect 27893 25109 27905 25112
rect 27939 25109 27951 25143
rect 27893 25103 27951 25109
rect 28074 25100 28080 25152
rect 28132 25100 28138 25152
rect 28994 25100 29000 25152
rect 29052 25140 29058 25152
rect 29288 25140 29316 25171
rect 30208 25152 30236 25180
rect 30834 25168 30840 25180
rect 30892 25168 30898 25220
rect 31113 25211 31171 25217
rect 31113 25177 31125 25211
rect 31159 25208 31171 25211
rect 31202 25208 31208 25220
rect 31159 25180 31208 25208
rect 31159 25177 31171 25180
rect 31113 25171 31171 25177
rect 31202 25168 31208 25180
rect 31260 25168 31266 25220
rect 32490 25168 32496 25220
rect 32548 25208 32554 25220
rect 34149 25211 34207 25217
rect 34149 25208 34161 25211
rect 32548 25180 34161 25208
rect 32548 25168 32554 25180
rect 34149 25177 34161 25180
rect 34195 25208 34207 25211
rect 36078 25208 36084 25220
rect 34195 25180 36084 25208
rect 34195 25177 34207 25180
rect 34149 25171 34207 25177
rect 36078 25168 36084 25180
rect 36136 25208 36142 25220
rect 36280 25217 36308 25248
rect 37550 25236 37556 25248
rect 37608 25236 37614 25288
rect 37737 25279 37795 25285
rect 37737 25245 37749 25279
rect 37783 25245 37795 25279
rect 39298 25276 39304 25288
rect 39146 25248 39304 25276
rect 37737 25239 37795 25245
rect 36265 25211 36323 25217
rect 36265 25208 36277 25211
rect 36136 25180 36277 25208
rect 36136 25168 36142 25180
rect 36265 25177 36277 25180
rect 36311 25177 36323 25211
rect 37752 25208 37780 25239
rect 39298 25236 39304 25248
rect 39356 25276 39362 25288
rect 39574 25276 39580 25288
rect 39356 25248 39580 25276
rect 39356 25236 39362 25248
rect 39574 25236 39580 25248
rect 39632 25236 39638 25288
rect 39942 25236 39948 25288
rect 40000 25276 40006 25288
rect 40402 25276 40408 25288
rect 40000 25248 40408 25276
rect 40000 25236 40006 25248
rect 40402 25236 40408 25248
rect 40460 25236 40466 25288
rect 38286 25208 38292 25220
rect 37752 25180 38292 25208
rect 36265 25171 36323 25177
rect 38286 25168 38292 25180
rect 38344 25168 38350 25220
rect 40678 25168 40684 25220
rect 40736 25168 40742 25220
rect 41414 25168 41420 25220
rect 41472 25168 41478 25220
rect 29052 25112 29316 25140
rect 29052 25100 29058 25112
rect 30190 25100 30196 25152
rect 30248 25100 30254 25152
rect 30558 25100 30564 25152
rect 30616 25140 30622 25152
rect 31018 25140 31024 25152
rect 30616 25112 31024 25140
rect 30616 25100 30622 25112
rect 31018 25100 31024 25112
rect 31076 25100 31082 25152
rect 35250 25100 35256 25152
rect 35308 25140 35314 25152
rect 35713 25143 35771 25149
rect 35713 25140 35725 25143
rect 35308 25112 35725 25140
rect 35308 25100 35314 25112
rect 35713 25109 35725 25112
rect 35759 25109 35771 25143
rect 35713 25103 35771 25109
rect 36814 25100 36820 25152
rect 36872 25140 36878 25152
rect 37274 25140 37280 25152
rect 36872 25112 37280 25140
rect 36872 25100 36878 25112
rect 37274 25100 37280 25112
rect 37332 25100 37338 25152
rect 37645 25143 37703 25149
rect 37645 25109 37657 25143
rect 37691 25140 37703 25143
rect 37734 25140 37740 25152
rect 37691 25112 37740 25140
rect 37691 25109 37703 25112
rect 37645 25103 37703 25109
rect 37734 25100 37740 25112
rect 37792 25100 37798 25152
rect 39574 25100 39580 25152
rect 39632 25140 39638 25152
rect 41598 25140 41604 25152
rect 39632 25112 41604 25140
rect 39632 25100 39638 25112
rect 41598 25100 41604 25112
rect 41656 25100 41662 25152
rect 1104 25050 42504 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 42504 25050
rect 1104 24976 42504 24998
rect 2590 24896 2596 24948
rect 2648 24936 2654 24948
rect 3145 24939 3203 24945
rect 3145 24936 3157 24939
rect 2648 24908 3157 24936
rect 2648 24896 2654 24908
rect 3145 24905 3157 24908
rect 3191 24936 3203 24939
rect 3234 24936 3240 24948
rect 3191 24908 3240 24936
rect 3191 24905 3203 24908
rect 3145 24899 3203 24905
rect 3234 24896 3240 24908
rect 3292 24896 3298 24948
rect 3418 24896 3424 24948
rect 3476 24936 3482 24948
rect 3513 24939 3571 24945
rect 3513 24936 3525 24939
rect 3476 24908 3525 24936
rect 3476 24896 3482 24908
rect 3513 24905 3525 24908
rect 3559 24905 3571 24939
rect 5350 24936 5356 24948
rect 3513 24899 3571 24905
rect 4172 24908 5356 24936
rect 4172 24868 4200 24908
rect 5350 24896 5356 24908
rect 5408 24896 5414 24948
rect 6365 24939 6423 24945
rect 6365 24905 6377 24939
rect 6411 24936 6423 24939
rect 6454 24936 6460 24948
rect 6411 24908 6460 24936
rect 6411 24905 6423 24908
rect 6365 24899 6423 24905
rect 6454 24896 6460 24908
rect 6512 24896 6518 24948
rect 7558 24896 7564 24948
rect 7616 24896 7622 24948
rect 7650 24896 7656 24948
rect 7708 24936 7714 24948
rect 8202 24936 8208 24948
rect 7708 24908 8208 24936
rect 7708 24896 7714 24908
rect 8202 24896 8208 24908
rect 8260 24936 8266 24948
rect 8260 24908 8984 24936
rect 8260 24896 8266 24908
rect 4798 24868 4804 24880
rect 3252 24840 4200 24868
rect 4264 24840 4804 24868
rect 3050 24800 3056 24812
rect 2806 24772 3056 24800
rect 3050 24760 3056 24772
rect 3108 24800 3114 24812
rect 3252 24800 3280 24840
rect 3108 24772 3280 24800
rect 3329 24803 3387 24809
rect 3108 24760 3114 24772
rect 3329 24769 3341 24803
rect 3375 24800 3387 24803
rect 3694 24800 3700 24812
rect 3375 24772 3700 24800
rect 3375 24769 3387 24772
rect 3329 24763 3387 24769
rect 3694 24760 3700 24772
rect 3752 24760 3758 24812
rect 3881 24803 3939 24809
rect 3881 24769 3893 24803
rect 3927 24800 3939 24803
rect 4264 24800 4292 24840
rect 4798 24828 4804 24840
rect 4856 24828 4862 24880
rect 6546 24828 6552 24880
rect 6604 24868 6610 24880
rect 7576 24868 7604 24896
rect 7929 24871 7987 24877
rect 7929 24868 7941 24871
rect 6604 24840 6776 24868
rect 6604 24828 6610 24840
rect 3927 24772 4292 24800
rect 4525 24803 4583 24809
rect 3927 24769 3939 24772
rect 3881 24763 3939 24769
rect 4525 24769 4537 24803
rect 4571 24800 4583 24803
rect 4706 24800 4712 24812
rect 4571 24772 4712 24800
rect 4571 24769 4583 24772
rect 4525 24763 4583 24769
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24800 4951 24803
rect 5626 24800 5632 24812
rect 4939 24772 5632 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5626 24760 5632 24772
rect 5684 24760 5690 24812
rect 6638 24760 6644 24812
rect 6696 24760 6702 24812
rect 6748 24809 6776 24840
rect 7300 24840 7604 24868
rect 7760 24840 7941 24868
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24769 6791 24803
rect 6733 24763 6791 24769
rect 6822 24760 6828 24812
rect 6880 24760 6886 24812
rect 7300 24809 7328 24840
rect 7009 24803 7067 24809
rect 7009 24769 7021 24803
rect 7055 24800 7067 24803
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 7055 24772 7113 24800
rect 7055 24769 7067 24772
rect 7009 24763 7067 24769
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 7285 24803 7343 24809
rect 7285 24769 7297 24803
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 7469 24803 7527 24809
rect 7469 24800 7481 24803
rect 7432 24772 7481 24800
rect 7432 24760 7438 24772
rect 7469 24769 7481 24772
rect 7515 24769 7527 24803
rect 7469 24763 7527 24769
rect 7558 24760 7564 24812
rect 7616 24760 7622 24812
rect 7650 24760 7656 24812
rect 7708 24760 7714 24812
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24701 1455 24735
rect 1397 24695 1455 24701
rect 1412 24596 1440 24695
rect 1670 24692 1676 24744
rect 1728 24692 1734 24744
rect 3418 24692 3424 24744
rect 3476 24732 3482 24744
rect 4249 24735 4307 24741
rect 4249 24732 4261 24735
rect 3476 24704 4261 24732
rect 3476 24692 3482 24704
rect 4249 24701 4261 24704
rect 4295 24701 4307 24735
rect 4249 24695 4307 24701
rect 4341 24735 4399 24741
rect 4341 24701 4353 24735
rect 4387 24732 4399 24735
rect 5350 24732 5356 24744
rect 4387 24704 5356 24732
rect 4387 24701 4399 24704
rect 4341 24695 4399 24701
rect 4154 24664 4160 24676
rect 2746 24636 4160 24664
rect 2746 24596 2774 24636
rect 4154 24624 4160 24636
rect 4212 24624 4218 24676
rect 4264 24664 4292 24695
rect 5350 24692 5356 24704
rect 5408 24692 5414 24744
rect 7760 24732 7788 24840
rect 7929 24837 7941 24840
rect 7975 24868 7987 24871
rect 7975 24840 8340 24868
rect 7975 24837 7987 24840
rect 7929 24831 7987 24837
rect 7834 24760 7840 24812
rect 7892 24800 7898 24812
rect 8021 24803 8079 24809
rect 8021 24800 8033 24803
rect 7892 24772 8033 24800
rect 7892 24760 7898 24772
rect 8021 24769 8033 24772
rect 8067 24769 8079 24803
rect 8205 24803 8263 24809
rect 8205 24800 8217 24803
rect 8021 24763 8079 24769
rect 8128 24772 8217 24800
rect 6656 24704 7788 24732
rect 8128 24732 8156 24772
rect 8205 24769 8217 24772
rect 8251 24769 8263 24803
rect 8312 24800 8340 24840
rect 8754 24800 8760 24812
rect 8312 24772 8760 24800
rect 8205 24763 8263 24769
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 8956 24809 8984 24908
rect 14384 24908 14688 24936
rect 9232 24840 9720 24868
rect 9232 24809 9260 24840
rect 8941 24803 8999 24809
rect 8941 24769 8953 24803
rect 8987 24769 8999 24803
rect 8941 24763 8999 24769
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24769 9183 24803
rect 9125 24763 9183 24769
rect 9217 24803 9275 24809
rect 9217 24769 9229 24803
rect 9263 24769 9275 24803
rect 9217 24763 9275 24769
rect 9140 24732 9168 24763
rect 9306 24760 9312 24812
rect 9364 24760 9370 24812
rect 9582 24760 9588 24812
rect 9640 24760 9646 24812
rect 8128 24704 9168 24732
rect 9692 24732 9720 24840
rect 11790 24828 11796 24880
rect 11848 24828 11854 24880
rect 13078 24868 13084 24880
rect 13018 24840 13084 24868
rect 13078 24828 13084 24840
rect 13136 24868 13142 24880
rect 14384 24868 14412 24908
rect 13136 24840 14412 24868
rect 13136 24828 13142 24840
rect 14550 24828 14556 24880
rect 14608 24828 14614 24880
rect 14660 24868 14688 24908
rect 16022 24896 16028 24948
rect 16080 24896 16086 24948
rect 16666 24896 16672 24948
rect 16724 24896 16730 24948
rect 17034 24896 17040 24948
rect 17092 24936 17098 24948
rect 17402 24936 17408 24948
rect 17092 24908 17408 24936
rect 17092 24896 17098 24908
rect 17402 24896 17408 24908
rect 17460 24896 17466 24948
rect 18322 24896 18328 24948
rect 18380 24896 18386 24948
rect 18414 24896 18420 24948
rect 18472 24896 18478 24948
rect 18874 24936 18880 24948
rect 18616 24908 18880 24936
rect 15010 24868 15016 24880
rect 14660 24840 15016 24868
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 16040 24868 16068 24896
rect 16853 24871 16911 24877
rect 16853 24868 16865 24871
rect 16040 24840 16865 24868
rect 16853 24837 16865 24840
rect 16899 24868 16911 24871
rect 17586 24868 17592 24880
rect 16899 24840 17592 24868
rect 16899 24837 16911 24840
rect 16853 24831 16911 24837
rect 17586 24828 17592 24840
rect 17644 24828 17650 24880
rect 18432 24868 18460 24896
rect 18156 24840 18460 24868
rect 9769 24803 9827 24809
rect 9769 24769 9781 24803
rect 9815 24800 9827 24803
rect 10686 24800 10692 24812
rect 9815 24772 10692 24800
rect 9815 24769 9827 24772
rect 9769 24763 9827 24769
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 11330 24760 11336 24812
rect 11388 24800 11394 24812
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 11388 24772 11529 24800
rect 11388 24760 11394 24772
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 13817 24803 13875 24809
rect 13817 24800 13829 24803
rect 11517 24763 11575 24769
rect 13648 24772 13829 24800
rect 11054 24732 11060 24744
rect 9692 24704 11060 24732
rect 6656 24676 6684 24704
rect 4709 24667 4767 24673
rect 4709 24664 4721 24667
rect 4264 24636 4721 24664
rect 4709 24633 4721 24636
rect 4755 24633 4767 24667
rect 4709 24627 4767 24633
rect 6638 24624 6644 24676
rect 6696 24624 6702 24676
rect 7745 24667 7803 24673
rect 7745 24664 7757 24667
rect 6748 24636 7757 24664
rect 1412 24568 2774 24596
rect 5994 24556 6000 24608
rect 6052 24596 6058 24608
rect 6748 24596 6776 24636
rect 7745 24633 7757 24636
rect 7791 24633 7803 24667
rect 7745 24627 7803 24633
rect 6052 24568 6776 24596
rect 6052 24556 6058 24568
rect 7374 24556 7380 24608
rect 7432 24596 7438 24608
rect 8128 24596 8156 24704
rect 11054 24692 11060 24704
rect 11112 24692 11118 24744
rect 8205 24667 8263 24673
rect 8205 24633 8217 24667
rect 8251 24664 8263 24667
rect 8294 24664 8300 24676
rect 8251 24636 8300 24664
rect 8251 24633 8263 24636
rect 8205 24627 8263 24633
rect 8294 24624 8300 24636
rect 8352 24624 8358 24676
rect 9582 24624 9588 24676
rect 9640 24664 9646 24676
rect 9953 24667 10011 24673
rect 9953 24664 9965 24667
rect 9640 24636 9965 24664
rect 9640 24624 9646 24636
rect 9953 24633 9965 24636
rect 9999 24633 10011 24667
rect 13648 24664 13676 24772
rect 13817 24769 13829 24772
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 16206 24760 16212 24812
rect 16264 24760 16270 24812
rect 17034 24760 17040 24812
rect 17092 24760 17098 24812
rect 18156 24809 18184 24840
rect 18616 24809 18644 24908
rect 18874 24896 18880 24908
rect 18932 24896 18938 24948
rect 19613 24939 19671 24945
rect 19613 24905 19625 24939
rect 19659 24936 19671 24939
rect 20070 24936 20076 24948
rect 19659 24908 20076 24936
rect 19659 24905 19671 24908
rect 19613 24899 19671 24905
rect 20070 24896 20076 24908
rect 20128 24896 20134 24948
rect 20254 24896 20260 24948
rect 20312 24936 20318 24948
rect 20441 24939 20499 24945
rect 20441 24936 20453 24939
rect 20312 24908 20453 24936
rect 20312 24896 20318 24908
rect 20441 24905 20453 24908
rect 20487 24905 20499 24939
rect 20441 24899 20499 24905
rect 21637 24939 21695 24945
rect 21637 24905 21649 24939
rect 21683 24936 21695 24939
rect 21726 24936 21732 24948
rect 21683 24908 21732 24936
rect 21683 24905 21695 24908
rect 21637 24899 21695 24905
rect 21726 24896 21732 24908
rect 21784 24896 21790 24948
rect 22462 24896 22468 24948
rect 22520 24896 22526 24948
rect 23934 24896 23940 24948
rect 23992 24936 23998 24948
rect 24762 24936 24768 24948
rect 23992 24908 24768 24936
rect 23992 24896 23998 24908
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 26418 24896 26424 24948
rect 26476 24936 26482 24948
rect 26973 24939 27031 24945
rect 26973 24936 26985 24939
rect 26476 24908 26985 24936
rect 26476 24896 26482 24908
rect 26973 24905 26985 24908
rect 27019 24905 27031 24939
rect 26973 24899 27031 24905
rect 27614 24896 27620 24948
rect 27672 24896 27678 24948
rect 27890 24896 27896 24948
rect 27948 24936 27954 24948
rect 30558 24936 30564 24948
rect 27948 24908 30564 24936
rect 27948 24896 27954 24908
rect 19904 24840 20300 24868
rect 18141 24803 18199 24809
rect 18141 24769 18153 24803
rect 18187 24769 18199 24803
rect 18417 24803 18475 24809
rect 18417 24800 18429 24803
rect 18141 24763 18199 24769
rect 18340 24772 18429 24800
rect 13722 24692 13728 24744
rect 13780 24732 13786 24744
rect 14277 24735 14335 24741
rect 14277 24732 14289 24735
rect 13780 24704 14289 24732
rect 13780 24692 13786 24704
rect 14277 24701 14289 24704
rect 14323 24701 14335 24735
rect 14277 24695 14335 24701
rect 14384 24704 16436 24732
rect 14384 24664 14412 24704
rect 13648 24636 14412 24664
rect 9953 24627 10011 24633
rect 7432 24568 8156 24596
rect 9493 24599 9551 24605
rect 7432 24556 7438 24568
rect 9493 24565 9505 24599
rect 9539 24596 9551 24599
rect 9766 24596 9772 24608
rect 9539 24568 9772 24596
rect 9539 24565 9551 24568
rect 9493 24559 9551 24565
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 13265 24599 13323 24605
rect 13265 24565 13277 24599
rect 13311 24596 13323 24599
rect 13354 24596 13360 24608
rect 13311 24568 13360 24596
rect 13311 24565 13323 24568
rect 13265 24559 13323 24565
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 15746 24596 15752 24608
rect 13596 24568 15752 24596
rect 13596 24556 13602 24568
rect 15746 24556 15752 24568
rect 15804 24556 15810 24608
rect 16408 24605 16436 24704
rect 16393 24599 16451 24605
rect 16393 24565 16405 24599
rect 16439 24596 16451 24599
rect 17954 24596 17960 24608
rect 16439 24568 17960 24596
rect 16439 24565 16451 24568
rect 16393 24559 16451 24565
rect 17954 24556 17960 24568
rect 18012 24556 18018 24608
rect 18340 24596 18368 24772
rect 18417 24769 18429 24772
rect 18463 24769 18475 24803
rect 18417 24763 18475 24769
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24769 18567 24803
rect 18509 24763 18567 24769
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24769 18659 24803
rect 18601 24763 18659 24769
rect 18524 24732 18552 24763
rect 18690 24760 18696 24812
rect 18748 24800 18754 24812
rect 18785 24803 18843 24809
rect 18785 24800 18797 24803
rect 18748 24772 18797 24800
rect 18748 24760 18754 24772
rect 18785 24769 18797 24772
rect 18831 24769 18843 24803
rect 18785 24763 18843 24769
rect 19518 24760 19524 24812
rect 19576 24760 19582 24812
rect 19702 24760 19708 24812
rect 19760 24760 19766 24812
rect 19797 24803 19855 24809
rect 19797 24769 19809 24803
rect 19843 24800 19855 24803
rect 19904 24800 19932 24840
rect 19843 24772 19932 24800
rect 19981 24803 20039 24809
rect 19843 24769 19855 24772
rect 19797 24763 19855 24769
rect 19981 24769 19993 24803
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 18966 24732 18972 24744
rect 18524 24704 18972 24732
rect 18966 24692 18972 24704
rect 19024 24692 19030 24744
rect 18417 24667 18475 24673
rect 18417 24633 18429 24667
rect 18463 24664 18475 24667
rect 18506 24664 18512 24676
rect 18463 24636 18512 24664
rect 18463 24633 18475 24636
rect 18417 24627 18475 24633
rect 18506 24624 18512 24636
rect 18564 24664 18570 24676
rect 19812 24664 19840 24763
rect 18564 24636 19840 24664
rect 19996 24664 20024 24763
rect 20070 24760 20076 24812
rect 20128 24760 20134 24812
rect 20162 24760 20168 24812
rect 20220 24760 20226 24812
rect 20272 24800 20300 24840
rect 20990 24828 20996 24880
rect 21048 24868 21054 24880
rect 22480 24868 22508 24896
rect 23382 24868 23388 24880
rect 21048 24840 22140 24868
rect 22480 24840 23388 24868
rect 21048 24828 21054 24840
rect 21100 24809 21128 24840
rect 20533 24803 20591 24809
rect 20533 24800 20545 24803
rect 20272 24772 20545 24800
rect 20533 24769 20545 24772
rect 20579 24769 20591 24803
rect 20533 24763 20591 24769
rect 20717 24803 20775 24809
rect 20717 24769 20729 24803
rect 20763 24800 20775 24803
rect 21085 24803 21143 24809
rect 20763 24772 21036 24800
rect 20763 24769 20775 24772
rect 20717 24763 20775 24769
rect 20088 24732 20116 24760
rect 20901 24735 20959 24741
rect 20901 24732 20913 24735
rect 20088 24704 20913 24732
rect 20901 24701 20913 24704
rect 20947 24701 20959 24735
rect 20901 24695 20959 24701
rect 21008 24664 21036 24772
rect 21085 24769 21097 24803
rect 21131 24769 21143 24803
rect 21085 24763 21143 24769
rect 21177 24803 21235 24809
rect 21177 24769 21189 24803
rect 21223 24800 21235 24803
rect 21361 24803 21419 24809
rect 21223 24772 21312 24800
rect 21223 24769 21235 24772
rect 21177 24763 21235 24769
rect 19996 24636 21036 24664
rect 21284 24664 21312 24772
rect 21361 24769 21373 24803
rect 21407 24769 21419 24803
rect 21361 24763 21419 24769
rect 21376 24732 21404 24763
rect 21450 24760 21456 24812
rect 21508 24800 21514 24812
rect 22112 24809 22140 24840
rect 23382 24828 23388 24840
rect 23440 24868 23446 24880
rect 24670 24868 24676 24880
rect 23440 24840 24676 24868
rect 23440 24828 23446 24840
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21508 24772 21833 24800
rect 21508 24760 21514 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 22097 24803 22155 24809
rect 22097 24769 22109 24803
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 22189 24803 22247 24809
rect 22189 24769 22201 24803
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 21726 24732 21732 24744
rect 21376 24704 21732 24732
rect 21726 24692 21732 24704
rect 21784 24732 21790 24744
rect 22020 24732 22048 24763
rect 21784 24704 22048 24732
rect 21784 24692 21790 24704
rect 22204 24664 22232 24763
rect 23566 24760 23572 24812
rect 23624 24800 23630 24812
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23624 24772 23673 24800
rect 23624 24760 23630 24772
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 23661 24763 23719 24769
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24800 23995 24803
rect 24026 24800 24032 24812
rect 23983 24772 24032 24800
rect 23983 24769 23995 24772
rect 23937 24763 23995 24769
rect 24026 24760 24032 24772
rect 24084 24760 24090 24812
rect 24320 24809 24348 24840
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 27632 24868 27660 24896
rect 27540 24840 27660 24868
rect 27801 24871 27859 24877
rect 24305 24803 24363 24809
rect 24305 24769 24317 24803
rect 24351 24769 24363 24803
rect 24305 24763 24363 24769
rect 24486 24760 24492 24812
rect 24544 24760 24550 24812
rect 25498 24760 25504 24812
rect 25556 24760 25562 24812
rect 26602 24760 26608 24812
rect 26660 24800 26666 24812
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 26660 24772 27169 24800
rect 26660 24760 26666 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27540 24800 27568 24840
rect 27801 24837 27813 24871
rect 27847 24868 27859 24871
rect 28074 24868 28080 24880
rect 27847 24840 28080 24868
rect 27847 24837 27859 24840
rect 27801 24831 27859 24837
rect 28074 24828 28080 24840
rect 28132 24828 28138 24880
rect 28184 24868 28212 24908
rect 28184 24840 28290 24868
rect 29730 24828 29736 24880
rect 29788 24828 29794 24880
rect 30116 24868 30144 24908
rect 30558 24896 30564 24908
rect 30616 24896 30622 24948
rect 33870 24896 33876 24948
rect 33928 24896 33934 24948
rect 34606 24896 34612 24948
rect 34664 24936 34670 24948
rect 34793 24939 34851 24945
rect 34793 24936 34805 24939
rect 34664 24908 34805 24936
rect 34664 24896 34670 24908
rect 34793 24905 34805 24908
rect 34839 24905 34851 24939
rect 34793 24899 34851 24905
rect 35158 24896 35164 24948
rect 35216 24896 35222 24948
rect 35250 24896 35256 24948
rect 35308 24896 35314 24948
rect 35713 24939 35771 24945
rect 35713 24905 35725 24939
rect 35759 24905 35771 24939
rect 35713 24899 35771 24905
rect 30116 24840 30222 24868
rect 31018 24828 31024 24880
rect 31076 24868 31082 24880
rect 31938 24868 31944 24880
rect 31076 24840 31944 24868
rect 31076 24828 31082 24840
rect 31938 24828 31944 24840
rect 31996 24828 32002 24880
rect 32582 24828 32588 24880
rect 32640 24877 32646 24880
rect 32640 24871 32669 24877
rect 32657 24837 32669 24871
rect 33410 24868 33416 24880
rect 32640 24831 32669 24837
rect 32968 24840 33416 24868
rect 32640 24828 32646 24831
rect 27157 24763 27215 24769
rect 27448 24772 27568 24800
rect 31481 24803 31539 24809
rect 23474 24692 23480 24744
rect 23532 24732 23538 24744
rect 23753 24735 23811 24741
rect 23753 24732 23765 24735
rect 23532 24704 23765 24732
rect 23532 24692 23538 24704
rect 23753 24701 23765 24704
rect 23799 24701 23811 24735
rect 23753 24695 23811 24701
rect 23842 24692 23848 24744
rect 23900 24732 23906 24744
rect 24213 24735 24271 24741
rect 24213 24732 24225 24735
rect 23900 24704 24225 24732
rect 23900 24692 23906 24704
rect 24213 24701 24225 24704
rect 24259 24701 24271 24735
rect 24213 24695 24271 24701
rect 24394 24692 24400 24744
rect 24452 24732 24458 24744
rect 24673 24735 24731 24741
rect 24673 24732 24685 24735
rect 24452 24704 24685 24732
rect 24452 24692 24458 24704
rect 24673 24701 24685 24704
rect 24719 24701 24731 24735
rect 24673 24695 24731 24701
rect 25774 24692 25780 24744
rect 25832 24732 25838 24744
rect 26050 24732 26056 24744
rect 25832 24704 26056 24732
rect 25832 24692 25838 24704
rect 26050 24692 26056 24704
rect 26108 24732 26114 24744
rect 27448 24741 27476 24772
rect 31481 24769 31493 24803
rect 31527 24800 31539 24803
rect 31846 24800 31852 24812
rect 31527 24772 31852 24800
rect 31527 24769 31539 24772
rect 31481 24763 31539 24769
rect 31846 24760 31852 24772
rect 31904 24760 31910 24812
rect 32030 24760 32036 24812
rect 32088 24800 32094 24812
rect 32125 24803 32183 24809
rect 32125 24800 32137 24803
rect 32088 24772 32137 24800
rect 32088 24760 32094 24772
rect 32125 24769 32137 24772
rect 32171 24769 32183 24803
rect 32125 24763 32183 24769
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32401 24803 32459 24809
rect 32401 24769 32413 24803
rect 32447 24769 32459 24803
rect 32401 24763 32459 24769
rect 32493 24803 32551 24809
rect 32493 24769 32505 24803
rect 32539 24800 32551 24803
rect 32968 24800 32996 24840
rect 33410 24828 33416 24840
rect 33468 24828 33474 24880
rect 33686 24868 33692 24880
rect 33520 24840 33692 24868
rect 32539 24772 32996 24800
rect 32539 24769 32551 24772
rect 32493 24763 32551 24769
rect 27433 24735 27491 24741
rect 27433 24732 27445 24735
rect 26108 24704 27445 24732
rect 26108 24692 26114 24704
rect 27433 24701 27445 24704
rect 27479 24701 27491 24735
rect 27433 24695 27491 24701
rect 27522 24692 27528 24744
rect 27580 24732 27586 24744
rect 29457 24735 29515 24741
rect 29457 24732 29469 24735
rect 27580 24704 29469 24732
rect 27580 24692 27586 24704
rect 29457 24701 29469 24704
rect 29503 24701 29515 24735
rect 29457 24695 29515 24701
rect 31205 24735 31263 24741
rect 31205 24701 31217 24735
rect 31251 24732 31263 24735
rect 31386 24732 31392 24744
rect 31251 24704 31392 24732
rect 31251 24701 31263 24704
rect 31205 24695 31263 24701
rect 31386 24692 31392 24704
rect 31444 24732 31450 24744
rect 31573 24735 31631 24741
rect 31573 24732 31585 24735
rect 31444 24704 31585 24732
rect 31444 24692 31450 24704
rect 31573 24701 31585 24704
rect 31619 24701 31631 24735
rect 31573 24695 31631 24701
rect 31665 24735 31723 24741
rect 31665 24701 31677 24735
rect 31711 24701 31723 24735
rect 31665 24695 31723 24701
rect 21284 24636 22232 24664
rect 24121 24667 24179 24673
rect 18564 24624 18570 24636
rect 18693 24599 18751 24605
rect 18693 24596 18705 24599
rect 18340 24568 18705 24596
rect 18693 24565 18705 24568
rect 18739 24596 18751 24599
rect 19610 24596 19616 24608
rect 18739 24568 19616 24596
rect 18739 24565 18751 24568
rect 18693 24559 18751 24565
rect 19610 24556 19616 24568
rect 19668 24596 19674 24608
rect 19996 24596 20024 24636
rect 19668 24568 20024 24596
rect 19668 24556 19674 24568
rect 20162 24556 20168 24608
rect 20220 24596 20226 24608
rect 20438 24596 20444 24608
rect 20220 24568 20444 24596
rect 20220 24556 20226 24568
rect 20438 24556 20444 24568
rect 20496 24596 20502 24608
rect 20809 24599 20867 24605
rect 20809 24596 20821 24599
rect 20496 24568 20821 24596
rect 20496 24556 20502 24568
rect 20809 24565 20821 24568
rect 20855 24596 20867 24599
rect 21284 24596 21312 24636
rect 24121 24633 24133 24667
rect 24167 24664 24179 24667
rect 24578 24664 24584 24676
rect 24167 24636 24584 24664
rect 24167 24633 24179 24636
rect 24121 24627 24179 24633
rect 24578 24624 24584 24636
rect 24636 24624 24642 24676
rect 27154 24624 27160 24676
rect 27212 24664 27218 24676
rect 27341 24667 27399 24673
rect 27341 24664 27353 24667
rect 27212 24636 27353 24664
rect 27212 24624 27218 24636
rect 27341 24633 27353 24636
rect 27387 24633 27399 24667
rect 27341 24627 27399 24633
rect 29178 24624 29184 24676
rect 29236 24664 29242 24676
rect 29273 24667 29331 24673
rect 29273 24664 29285 24667
rect 29236 24636 29285 24664
rect 29236 24624 29242 24636
rect 29273 24633 29285 24636
rect 29319 24633 29331 24667
rect 29273 24627 29331 24633
rect 20855 24568 21312 24596
rect 20855 24565 20867 24568
rect 20809 24559 20867 24565
rect 25314 24556 25320 24608
rect 25372 24596 25378 24608
rect 25593 24599 25651 24605
rect 25593 24596 25605 24599
rect 25372 24568 25605 24596
rect 25372 24556 25378 24568
rect 25593 24565 25605 24568
rect 25639 24565 25651 24599
rect 29288 24596 29316 24627
rect 29822 24596 29828 24608
rect 29288 24568 29828 24596
rect 25593 24559 25651 24565
rect 29822 24556 29828 24568
rect 29880 24596 29886 24608
rect 31680 24596 31708 24695
rect 31754 24692 31760 24744
rect 31812 24692 31818 24744
rect 31941 24735 31999 24741
rect 31941 24701 31953 24735
rect 31987 24732 31999 24735
rect 32324 24732 32352 24763
rect 31987 24704 32352 24732
rect 31987 24701 31999 24704
rect 31941 24695 31999 24701
rect 32416 24664 32444 24763
rect 33042 24760 33048 24812
rect 33100 24760 33106 24812
rect 33520 24809 33548 24840
rect 33686 24828 33692 24840
rect 33744 24828 33750 24880
rect 34698 24828 34704 24880
rect 34756 24868 34762 24880
rect 35176 24868 35204 24896
rect 34756 24840 35204 24868
rect 34756 24828 34762 24840
rect 35618 24828 35624 24880
rect 35676 24868 35682 24880
rect 35728 24868 35756 24899
rect 35986 24896 35992 24948
rect 36044 24936 36050 24948
rect 39574 24936 39580 24948
rect 36044 24908 39580 24936
rect 36044 24896 36050 24908
rect 39574 24896 39580 24908
rect 39632 24896 39638 24948
rect 40678 24896 40684 24948
rect 40736 24936 40742 24948
rect 40865 24939 40923 24945
rect 40865 24936 40877 24939
rect 40736 24908 40877 24936
rect 40736 24896 40742 24908
rect 40865 24905 40877 24908
rect 40911 24905 40923 24939
rect 40865 24899 40923 24905
rect 41046 24896 41052 24948
rect 41104 24936 41110 24948
rect 41233 24939 41291 24945
rect 41233 24936 41245 24939
rect 41104 24908 41245 24936
rect 41104 24896 41110 24908
rect 41233 24905 41245 24908
rect 41279 24905 41291 24939
rect 41233 24899 41291 24905
rect 35676 24840 35756 24868
rect 35676 24828 35682 24840
rect 36262 24828 36268 24880
rect 36320 24868 36326 24880
rect 37734 24868 37740 24880
rect 36320 24840 37044 24868
rect 36320 24828 36326 24840
rect 33505 24803 33563 24809
rect 33505 24769 33517 24803
rect 33551 24769 33563 24803
rect 33505 24763 33563 24769
rect 33597 24803 33655 24809
rect 33597 24769 33609 24803
rect 33643 24800 33655 24803
rect 33643 24772 34100 24800
rect 33643 24769 33655 24772
rect 33597 24763 33655 24769
rect 32674 24692 32680 24744
rect 32732 24732 32738 24744
rect 32769 24735 32827 24741
rect 32769 24732 32781 24735
rect 32732 24704 32781 24732
rect 32732 24692 32738 24704
rect 32769 24701 32781 24704
rect 32815 24732 32827 24735
rect 33226 24732 33232 24744
rect 32815 24704 33232 24732
rect 32815 24701 32827 24704
rect 32769 24695 32827 24701
rect 33226 24692 33232 24704
rect 33284 24692 33290 24744
rect 33410 24692 33416 24744
rect 33468 24732 33474 24744
rect 33873 24735 33931 24741
rect 33873 24732 33885 24735
rect 33468 24704 33885 24732
rect 33468 24692 33474 24704
rect 33873 24701 33885 24704
rect 33919 24701 33931 24735
rect 33873 24695 33931 24701
rect 32953 24667 33011 24673
rect 32953 24664 32965 24667
rect 32416 24636 32965 24664
rect 32953 24633 32965 24636
rect 32999 24633 33011 24667
rect 32953 24627 33011 24633
rect 29880 24568 31708 24596
rect 29880 24556 29886 24568
rect 33778 24556 33784 24608
rect 33836 24556 33842 24608
rect 33888 24596 33916 24695
rect 34072 24673 34100 24772
rect 34146 24760 34152 24812
rect 34204 24760 34210 24812
rect 34514 24760 34520 24812
rect 34572 24760 34578 24812
rect 35158 24800 35164 24812
rect 34624 24772 35164 24800
rect 34333 24735 34391 24741
rect 34333 24701 34345 24735
rect 34379 24732 34391 24735
rect 34624 24732 34652 24772
rect 35158 24760 35164 24772
rect 35216 24760 35222 24812
rect 35434 24760 35440 24812
rect 35492 24800 35498 24812
rect 35897 24803 35955 24809
rect 35897 24800 35909 24803
rect 35492 24772 35909 24800
rect 35492 24760 35498 24772
rect 35897 24769 35909 24772
rect 35943 24769 35955 24803
rect 35897 24763 35955 24769
rect 35989 24803 36047 24809
rect 35989 24769 36001 24803
rect 36035 24800 36047 24803
rect 36538 24800 36544 24812
rect 36035 24772 36544 24800
rect 36035 24769 36047 24772
rect 35989 24763 36047 24769
rect 36538 24760 36544 24772
rect 36596 24760 36602 24812
rect 36648 24809 36676 24840
rect 36633 24803 36691 24809
rect 36633 24769 36645 24803
rect 36679 24769 36691 24803
rect 36633 24763 36691 24769
rect 36725 24803 36783 24809
rect 36725 24769 36737 24803
rect 36771 24769 36783 24803
rect 36725 24763 36783 24769
rect 34379 24704 34652 24732
rect 34701 24735 34759 24741
rect 34379 24701 34391 24704
rect 34333 24695 34391 24701
rect 34701 24701 34713 24735
rect 34747 24732 34759 24735
rect 34882 24732 34888 24744
rect 34747 24704 34888 24732
rect 34747 24701 34759 24704
rect 34701 24695 34759 24701
rect 34882 24692 34888 24704
rect 34940 24692 34946 24744
rect 35342 24692 35348 24744
rect 35400 24692 35406 24744
rect 36078 24692 36084 24744
rect 36136 24732 36142 24744
rect 36265 24735 36323 24741
rect 36265 24732 36277 24735
rect 36136 24704 36277 24732
rect 36136 24692 36142 24704
rect 36265 24701 36277 24704
rect 36311 24701 36323 24735
rect 36265 24695 36323 24701
rect 36354 24692 36360 24744
rect 36412 24692 36418 24744
rect 34057 24667 34115 24673
rect 34057 24633 34069 24667
rect 34103 24664 34115 24667
rect 36170 24664 36176 24676
rect 34103 24636 36176 24664
rect 34103 24633 34115 24636
rect 34057 24627 34115 24633
rect 36170 24624 36176 24636
rect 36228 24624 36234 24676
rect 36372 24664 36400 24692
rect 36630 24664 36636 24676
rect 36372 24636 36636 24664
rect 36630 24624 36636 24636
rect 36688 24624 36694 24676
rect 36740 24664 36768 24763
rect 36814 24760 36820 24812
rect 36872 24800 36878 24812
rect 36909 24803 36967 24809
rect 36909 24800 36921 24803
rect 36872 24772 36921 24800
rect 36872 24760 36878 24772
rect 36909 24769 36921 24772
rect 36955 24769 36967 24803
rect 37016 24800 37044 24840
rect 37476 24840 37740 24868
rect 37476 24809 37504 24840
rect 37734 24828 37740 24840
rect 37792 24868 37798 24880
rect 37921 24871 37979 24877
rect 37921 24868 37933 24871
rect 37792 24840 37933 24868
rect 37792 24828 37798 24840
rect 37921 24837 37933 24840
rect 37967 24868 37979 24871
rect 38562 24868 38568 24880
rect 37967 24840 38568 24868
rect 37967 24837 37979 24840
rect 37921 24831 37979 24837
rect 38562 24828 38568 24840
rect 38620 24828 38626 24880
rect 39298 24828 39304 24880
rect 39356 24828 39362 24880
rect 40696 24840 40908 24868
rect 37277 24803 37335 24809
rect 37277 24800 37289 24803
rect 37016 24772 37289 24800
rect 36909 24763 36967 24769
rect 37277 24769 37289 24772
rect 37323 24769 37335 24803
rect 37277 24763 37335 24769
rect 37461 24803 37519 24809
rect 37461 24769 37473 24803
rect 37507 24769 37519 24803
rect 37461 24763 37519 24769
rect 37093 24735 37151 24741
rect 37093 24701 37105 24735
rect 37139 24732 37151 24735
rect 37366 24732 37372 24744
rect 37139 24704 37372 24732
rect 37139 24701 37151 24704
rect 37093 24695 37151 24701
rect 37366 24692 37372 24704
rect 37424 24692 37430 24744
rect 37476 24664 37504 24763
rect 38286 24760 38292 24812
rect 38344 24800 38350 24812
rect 38381 24803 38439 24809
rect 38381 24800 38393 24803
rect 38344 24772 38393 24800
rect 38344 24760 38350 24772
rect 38381 24769 38393 24772
rect 38427 24769 38439 24803
rect 40696 24800 40724 24840
rect 38381 24763 38439 24769
rect 39868 24772 40724 24800
rect 40773 24803 40831 24809
rect 37642 24692 37648 24744
rect 37700 24692 37706 24744
rect 37826 24692 37832 24744
rect 37884 24692 37890 24744
rect 38657 24735 38715 24741
rect 38657 24732 38669 24735
rect 38304 24704 38669 24732
rect 38304 24673 38332 24704
rect 38657 24701 38669 24704
rect 38703 24701 38715 24735
rect 38657 24695 38715 24701
rect 39022 24692 39028 24744
rect 39080 24732 39086 24744
rect 39868 24732 39896 24772
rect 40773 24769 40785 24803
rect 40819 24769 40831 24803
rect 40773 24763 40831 24769
rect 39080 24704 39896 24732
rect 40405 24735 40463 24741
rect 39080 24692 39086 24704
rect 40405 24701 40417 24735
rect 40451 24701 40463 24735
rect 40405 24695 40463 24701
rect 36740 24636 37504 24664
rect 38289 24667 38347 24673
rect 38289 24633 38301 24667
rect 38335 24633 38347 24667
rect 38289 24627 38347 24633
rect 36722 24596 36728 24608
rect 33888 24568 36728 24596
rect 36722 24556 36728 24568
rect 36780 24556 36786 24608
rect 37274 24556 37280 24608
rect 37332 24596 37338 24608
rect 37369 24599 37427 24605
rect 37369 24596 37381 24599
rect 37332 24568 37381 24596
rect 37332 24556 37338 24568
rect 37369 24565 37381 24568
rect 37415 24565 37427 24599
rect 37369 24559 37427 24565
rect 38470 24556 38476 24608
rect 38528 24596 38534 24608
rect 40420 24596 40448 24695
rect 40788 24664 40816 24763
rect 40880 24732 40908 24840
rect 41414 24828 41420 24880
rect 41472 24868 41478 24880
rect 41472 24840 41736 24868
rect 41472 24828 41478 24840
rect 41325 24803 41383 24809
rect 41325 24769 41337 24803
rect 41371 24800 41383 24803
rect 41506 24800 41512 24812
rect 41371 24772 41512 24800
rect 41371 24769 41383 24772
rect 41325 24763 41383 24769
rect 41506 24760 41512 24772
rect 41564 24760 41570 24812
rect 41708 24809 41736 24840
rect 41693 24803 41751 24809
rect 41693 24769 41705 24803
rect 41739 24769 41751 24803
rect 41693 24763 41751 24769
rect 41966 24760 41972 24812
rect 42024 24800 42030 24812
rect 42061 24803 42119 24809
rect 42061 24800 42073 24803
rect 42024 24772 42073 24800
rect 42024 24760 42030 24772
rect 42061 24769 42073 24772
rect 42107 24769 42119 24803
rect 42061 24763 42119 24769
rect 41417 24735 41475 24741
rect 41417 24732 41429 24735
rect 40880 24704 41429 24732
rect 41417 24701 41429 24704
rect 41463 24732 41475 24735
rect 41463 24704 41552 24732
rect 41463 24701 41475 24704
rect 41417 24695 41475 24701
rect 41524 24676 41552 24704
rect 40788 24636 41414 24664
rect 38528 24568 40448 24596
rect 38528 24556 38534 24568
rect 40586 24556 40592 24608
rect 40644 24556 40650 24608
rect 41386 24596 41414 24636
rect 41506 24624 41512 24676
rect 41564 24624 41570 24676
rect 41690 24596 41696 24608
rect 41386 24568 41696 24596
rect 41690 24556 41696 24568
rect 41748 24556 41754 24608
rect 1104 24506 42504 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 42504 24506
rect 1104 24432 42504 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 1857 24395 1915 24401
rect 1857 24392 1869 24395
rect 1728 24364 1869 24392
rect 1728 24352 1734 24364
rect 1857 24361 1869 24364
rect 1903 24361 1915 24395
rect 1857 24355 1915 24361
rect 3053 24395 3111 24401
rect 3053 24361 3065 24395
rect 3099 24392 3111 24395
rect 3510 24392 3516 24404
rect 3099 24364 3516 24392
rect 3099 24361 3111 24364
rect 3053 24355 3111 24361
rect 3510 24352 3516 24364
rect 3568 24352 3574 24404
rect 6914 24352 6920 24404
rect 6972 24392 6978 24404
rect 7561 24395 7619 24401
rect 7561 24392 7573 24395
rect 6972 24364 7573 24392
rect 6972 24352 6978 24364
rect 7561 24361 7573 24364
rect 7607 24361 7619 24395
rect 9674 24392 9680 24404
rect 7561 24355 7619 24361
rect 9324 24364 9680 24392
rect 1762 24284 1768 24336
rect 1820 24324 1826 24336
rect 1820 24296 3188 24324
rect 1820 24284 1826 24296
rect 2866 24256 2872 24268
rect 1872 24228 2872 24256
rect 1872 24197 1900 24228
rect 2866 24216 2872 24228
rect 2924 24216 2930 24268
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 1857 24151 1915 24157
rect 2133 24191 2191 24197
rect 2133 24157 2145 24191
rect 2179 24157 2191 24191
rect 2133 24151 2191 24157
rect 2317 24191 2375 24197
rect 2317 24157 2329 24191
rect 2363 24188 2375 24191
rect 2774 24188 2780 24200
rect 2363 24160 2780 24188
rect 2363 24157 2375 24160
rect 2317 24151 2375 24157
rect 2148 24120 2176 24151
rect 2774 24148 2780 24160
rect 2832 24148 2838 24200
rect 2958 24148 2964 24200
rect 3016 24148 3022 24200
rect 3160 24197 3188 24296
rect 7098 24284 7104 24336
rect 7156 24324 7162 24336
rect 7745 24327 7803 24333
rect 7745 24324 7757 24327
rect 7156 24296 7757 24324
rect 7156 24284 7162 24296
rect 7745 24293 7757 24296
rect 7791 24293 7803 24327
rect 7745 24287 7803 24293
rect 3329 24259 3387 24265
rect 3329 24225 3341 24259
rect 3375 24256 3387 24259
rect 3375 24228 4844 24256
rect 3375 24225 3387 24228
rect 3329 24219 3387 24225
rect 4816 24200 4844 24228
rect 5994 24216 6000 24268
rect 6052 24216 6058 24268
rect 6270 24216 6276 24268
rect 6328 24256 6334 24268
rect 7193 24259 7251 24265
rect 7193 24256 7205 24259
rect 6328 24228 7205 24256
rect 6328 24216 6334 24228
rect 7193 24225 7205 24228
rect 7239 24256 7251 24259
rect 7282 24256 7288 24268
rect 7239 24228 7288 24256
rect 7239 24225 7251 24228
rect 7193 24219 7251 24225
rect 7282 24216 7288 24228
rect 7340 24216 7346 24268
rect 7650 24216 7656 24268
rect 7708 24256 7714 24268
rect 8113 24259 8171 24265
rect 8113 24256 8125 24259
rect 7708 24228 8125 24256
rect 7708 24216 7714 24228
rect 8113 24225 8125 24228
rect 8159 24225 8171 24259
rect 8113 24219 8171 24225
rect 8202 24216 8208 24268
rect 8260 24216 8266 24268
rect 8294 24216 8300 24268
rect 8352 24216 8358 24268
rect 9324 24265 9352 24364
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 10686 24352 10692 24404
rect 10744 24352 10750 24404
rect 15010 24352 15016 24404
rect 15068 24392 15074 24404
rect 16117 24395 16175 24401
rect 16117 24392 16129 24395
rect 15068 24364 16129 24392
rect 15068 24352 15074 24364
rect 16117 24361 16129 24364
rect 16163 24361 16175 24395
rect 16117 24355 16175 24361
rect 18598 24352 18604 24404
rect 18656 24392 18662 24404
rect 19058 24392 19064 24404
rect 18656 24364 18736 24392
rect 18656 24352 18662 24364
rect 9309 24259 9367 24265
rect 9309 24225 9321 24259
rect 9355 24225 9367 24259
rect 10704 24256 10732 24352
rect 10781 24259 10839 24265
rect 10781 24256 10793 24259
rect 10704 24228 10793 24256
rect 9309 24219 9367 24225
rect 10781 24225 10793 24228
rect 10827 24225 10839 24259
rect 10781 24219 10839 24225
rect 11330 24216 11336 24268
rect 11388 24256 11394 24268
rect 11517 24259 11575 24265
rect 11517 24256 11529 24259
rect 11388 24228 11529 24256
rect 11388 24216 11394 24228
rect 11517 24225 11529 24228
rect 11563 24225 11575 24259
rect 14553 24259 14611 24265
rect 14553 24256 14565 24259
rect 11517 24219 11575 24225
rect 13372 24228 14565 24256
rect 3145 24191 3203 24197
rect 3145 24157 3157 24191
rect 3191 24157 3203 24191
rect 3145 24151 3203 24157
rect 3050 24120 3056 24132
rect 2148 24092 3056 24120
rect 3050 24080 3056 24092
rect 3108 24080 3114 24132
rect 3160 24120 3188 24151
rect 3234 24148 3240 24200
rect 3292 24148 3298 24200
rect 3418 24148 3424 24200
rect 3476 24148 3482 24200
rect 4798 24148 4804 24200
rect 4856 24188 4862 24200
rect 4893 24191 4951 24197
rect 4893 24188 4905 24191
rect 4856 24160 4905 24188
rect 4856 24148 4862 24160
rect 4893 24157 4905 24160
rect 4939 24157 4951 24191
rect 4893 24151 4951 24157
rect 5534 24148 5540 24200
rect 5592 24148 5598 24200
rect 5626 24148 5632 24200
rect 5684 24148 5690 24200
rect 6638 24148 6644 24200
rect 6696 24148 6702 24200
rect 8021 24191 8079 24197
rect 6748 24160 7328 24188
rect 5350 24120 5356 24132
rect 3160 24092 5356 24120
rect 5350 24080 5356 24092
rect 5408 24080 5414 24132
rect 2041 24055 2099 24061
rect 2041 24021 2053 24055
rect 2087 24052 2099 24055
rect 2682 24052 2688 24064
rect 2087 24024 2688 24052
rect 2087 24021 2099 24024
rect 2041 24015 2099 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 2866 24012 2872 24064
rect 2924 24012 2930 24064
rect 6748 24061 6776 24160
rect 7300 24132 7328 24160
rect 7607 24157 7665 24163
rect 7607 24154 7619 24157
rect 6917 24123 6975 24129
rect 6917 24089 6929 24123
rect 6963 24120 6975 24123
rect 7006 24120 7012 24132
rect 6963 24092 7012 24120
rect 6963 24089 6975 24092
rect 6917 24083 6975 24089
rect 7006 24080 7012 24092
rect 7064 24120 7070 24132
rect 7190 24120 7196 24132
rect 7064 24092 7196 24120
rect 7064 24080 7070 24092
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 7282 24080 7288 24132
rect 7340 24080 7346 24132
rect 7377 24123 7435 24129
rect 7377 24089 7389 24123
rect 7423 24120 7435 24123
rect 7466 24120 7472 24132
rect 7423 24092 7472 24120
rect 7423 24089 7435 24092
rect 7377 24083 7435 24089
rect 6733 24055 6791 24061
rect 6733 24021 6745 24055
rect 6779 24021 6791 24055
rect 6733 24015 6791 24021
rect 7098 24012 7104 24064
rect 7156 24052 7162 24064
rect 7392 24052 7420 24083
rect 7466 24080 7472 24092
rect 7524 24080 7530 24132
rect 7592 24123 7619 24154
rect 7653 24132 7665 24157
rect 8021 24157 8033 24191
rect 8067 24188 8079 24191
rect 8570 24188 8576 24200
rect 8067 24160 8576 24188
rect 8067 24157 8079 24160
rect 8021 24151 8079 24157
rect 8570 24148 8576 24160
rect 8628 24148 8634 24200
rect 13372 24197 13400 24228
rect 14553 24225 14565 24228
rect 14599 24225 14611 24259
rect 14553 24219 14611 24225
rect 15933 24259 15991 24265
rect 15933 24225 15945 24259
rect 15979 24256 15991 24259
rect 16022 24256 16028 24268
rect 15979 24228 16028 24256
rect 15979 24225 15991 24228
rect 15933 24219 15991 24225
rect 16022 24216 16028 24228
rect 16080 24216 16086 24268
rect 16942 24216 16948 24268
rect 17000 24256 17006 24268
rect 17221 24259 17279 24265
rect 17221 24256 17233 24259
rect 17000 24228 17233 24256
rect 17000 24216 17006 24228
rect 17221 24225 17233 24228
rect 17267 24225 17279 24259
rect 17221 24219 17279 24225
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24157 13415 24191
rect 13357 24151 13415 24157
rect 13538 24148 13544 24200
rect 13596 24148 13602 24200
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24188 13783 24191
rect 15010 24188 15016 24200
rect 13771 24160 15016 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 15010 24148 15016 24160
rect 15068 24148 15074 24200
rect 15102 24148 15108 24200
rect 15160 24148 15166 24200
rect 16666 24148 16672 24200
rect 16724 24188 16730 24200
rect 17126 24188 17132 24200
rect 16724 24160 17132 24188
rect 16724 24148 16730 24160
rect 17126 24148 17132 24160
rect 17184 24188 17190 24200
rect 17586 24188 17592 24200
rect 17184 24160 17592 24188
rect 17184 24148 17190 24160
rect 17586 24148 17592 24160
rect 17644 24148 17650 24200
rect 18325 24191 18383 24197
rect 18325 24188 18337 24191
rect 17880 24160 18337 24188
rect 7653 24123 7656 24132
rect 7592 24092 7656 24123
rect 7650 24080 7656 24092
rect 7708 24080 7714 24132
rect 9582 24129 9588 24132
rect 9576 24083 9588 24129
rect 9582 24080 9588 24083
rect 9640 24080 9646 24132
rect 11790 24080 11796 24132
rect 11848 24080 11854 24132
rect 13078 24120 13084 24132
rect 13018 24092 13084 24120
rect 13078 24080 13084 24092
rect 13136 24080 13142 24132
rect 13633 24123 13691 24129
rect 13633 24089 13645 24123
rect 13679 24120 13691 24123
rect 15289 24123 15347 24129
rect 15289 24120 15301 24123
rect 13679 24092 15301 24120
rect 13679 24089 13691 24092
rect 13633 24083 13691 24089
rect 15289 24089 15301 24092
rect 15335 24089 15347 24123
rect 15289 24083 15347 24089
rect 16393 24123 16451 24129
rect 16393 24089 16405 24123
rect 16439 24120 16451 24123
rect 16574 24120 16580 24132
rect 16439 24092 16580 24120
rect 16439 24089 16451 24092
rect 16393 24083 16451 24089
rect 16574 24080 16580 24092
rect 16632 24080 16638 24132
rect 17037 24123 17095 24129
rect 17037 24089 17049 24123
rect 17083 24120 17095 24123
rect 17770 24120 17776 24132
rect 17083 24092 17776 24120
rect 17083 24089 17095 24092
rect 17037 24083 17095 24089
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 7156 24024 7420 24052
rect 8481 24055 8539 24061
rect 7156 24012 7162 24024
rect 8481 24021 8493 24055
rect 8527 24052 8539 24055
rect 9306 24052 9312 24064
rect 8527 24024 9312 24052
rect 8527 24021 8539 24024
rect 8481 24015 8539 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 11422 24012 11428 24064
rect 11480 24012 11486 24064
rect 13262 24012 13268 24064
rect 13320 24012 13326 24064
rect 13909 24055 13967 24061
rect 13909 24021 13921 24055
rect 13955 24052 13967 24055
rect 13998 24052 14004 24064
rect 13955 24024 14004 24052
rect 13955 24021 13967 24024
rect 13909 24015 13967 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 16669 24055 16727 24061
rect 16669 24021 16681 24055
rect 16715 24052 16727 24055
rect 16942 24052 16948 24064
rect 16715 24024 16948 24052
rect 16715 24021 16727 24024
rect 16669 24015 16727 24021
rect 16942 24012 16948 24024
rect 17000 24012 17006 24064
rect 17129 24055 17187 24061
rect 17129 24021 17141 24055
rect 17175 24052 17187 24055
rect 17880 24052 17908 24160
rect 18325 24157 18337 24160
rect 18371 24157 18383 24191
rect 18506 24188 18512 24200
rect 18468 24160 18512 24188
rect 18325 24151 18383 24157
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 18708 24197 18736 24364
rect 18892 24364 19064 24392
rect 18892 24256 18920 24364
rect 19058 24352 19064 24364
rect 19116 24352 19122 24404
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 20438 24352 20444 24404
rect 20496 24352 20502 24404
rect 21450 24352 21456 24404
rect 21508 24392 21514 24404
rect 21545 24395 21603 24401
rect 21545 24392 21557 24395
rect 21508 24364 21557 24392
rect 21508 24352 21514 24364
rect 21545 24361 21557 24364
rect 21591 24361 21603 24395
rect 21545 24355 21603 24361
rect 21726 24352 21732 24404
rect 21784 24352 21790 24404
rect 29546 24352 29552 24404
rect 29604 24352 29610 24404
rect 31849 24395 31907 24401
rect 31849 24361 31861 24395
rect 31895 24392 31907 24395
rect 33042 24392 33048 24404
rect 31895 24364 33048 24392
rect 31895 24361 31907 24364
rect 31849 24355 31907 24361
rect 33042 24352 33048 24364
rect 33100 24392 33106 24404
rect 33100 24364 34468 24392
rect 33100 24352 33106 24364
rect 18966 24284 18972 24336
rect 19024 24284 19030 24336
rect 25501 24327 25559 24333
rect 25501 24293 25513 24327
rect 25547 24324 25559 24327
rect 26878 24324 26884 24336
rect 25547 24296 26884 24324
rect 25547 24293 25559 24296
rect 25501 24287 25559 24293
rect 26878 24284 26884 24296
rect 26936 24284 26942 24336
rect 31297 24327 31355 24333
rect 31297 24293 31309 24327
rect 31343 24324 31355 24327
rect 31938 24324 31944 24336
rect 31343 24296 31944 24324
rect 31343 24293 31355 24296
rect 31297 24287 31355 24293
rect 31938 24284 31944 24296
rect 31996 24324 32002 24336
rect 32398 24324 32404 24336
rect 31996 24296 32404 24324
rect 31996 24284 32002 24296
rect 32398 24284 32404 24296
rect 32456 24284 32462 24336
rect 18800 24228 18920 24256
rect 18984 24256 19012 24284
rect 18984 24228 19840 24256
rect 18800 24198 18828 24228
rect 19058 24198 19064 24200
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18800 24191 19064 24198
rect 18800 24170 18981 24191
rect 18693 24151 18751 24157
rect 18969 24157 18981 24170
rect 19015 24170 19064 24191
rect 19015 24157 19027 24170
rect 18969 24151 19027 24157
rect 19058 24148 19064 24170
rect 19116 24148 19122 24200
rect 19150 24148 19156 24200
rect 19208 24182 19214 24200
rect 19429 24191 19487 24197
rect 19429 24188 19441 24191
rect 19260 24182 19441 24188
rect 19208 24160 19441 24182
rect 19208 24154 19288 24160
rect 19429 24157 19441 24160
rect 19475 24157 19487 24191
rect 19208 24148 19214 24154
rect 19429 24151 19487 24157
rect 19610 24148 19616 24200
rect 19668 24148 19674 24200
rect 19812 24197 19840 24228
rect 19886 24216 19892 24268
rect 19944 24256 19950 24268
rect 22830 24256 22836 24268
rect 19944 24228 20300 24256
rect 19944 24216 19950 24228
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24157 19855 24191
rect 20070 24188 20076 24200
rect 19797 24151 19855 24157
rect 19996 24160 20076 24188
rect 18230 24080 18236 24132
rect 18288 24120 18294 24132
rect 18602 24123 18660 24129
rect 18288 24092 18368 24120
rect 18288 24080 18294 24092
rect 17175 24024 17908 24052
rect 18340 24052 18368 24092
rect 18602 24089 18614 24123
rect 18648 24089 18660 24123
rect 18602 24083 18660 24089
rect 18616 24052 18644 24083
rect 18782 24080 18788 24132
rect 18840 24129 18846 24132
rect 18840 24123 18889 24129
rect 18840 24089 18843 24123
rect 18877 24089 18889 24123
rect 18840 24083 18889 24089
rect 19260 24092 19472 24120
rect 18840 24080 18846 24083
rect 19260 24064 19288 24092
rect 18340 24024 18644 24052
rect 17175 24021 17187 24024
rect 17129 24015 17187 24021
rect 19242 24012 19248 24064
rect 19300 24012 19306 24064
rect 19444 24052 19472 24092
rect 19518 24080 19524 24132
rect 19576 24080 19582 24132
rect 19702 24080 19708 24132
rect 19760 24120 19766 24132
rect 19996 24120 20024 24160
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20272 24197 20300 24228
rect 21652 24228 22836 24256
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20990 24148 20996 24200
rect 21048 24188 21054 24200
rect 21652 24197 21680 24228
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 23198 24216 23204 24268
rect 23256 24256 23262 24268
rect 33778 24256 33784 24268
rect 23256 24228 33784 24256
rect 23256 24216 23262 24228
rect 33778 24216 33784 24228
rect 33836 24216 33842 24268
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21048 24160 21373 24188
rect 21048 24148 21054 24160
rect 21361 24157 21373 24160
rect 21407 24188 21419 24191
rect 21637 24191 21695 24197
rect 21637 24188 21649 24191
rect 21407 24160 21649 24188
rect 21407 24157 21419 24160
rect 21361 24151 21419 24157
rect 21637 24157 21649 24160
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 21821 24191 21879 24197
rect 21821 24157 21833 24191
rect 21867 24188 21879 24191
rect 23014 24188 23020 24200
rect 21867 24160 23020 24188
rect 21867 24157 21879 24160
rect 21821 24151 21879 24157
rect 19760 24092 20024 24120
rect 21177 24123 21235 24129
rect 19760 24080 19766 24092
rect 21177 24089 21189 24123
rect 21223 24120 21235 24123
rect 21836 24120 21864 24151
rect 23014 24148 23020 24160
rect 23072 24148 23078 24200
rect 24946 24148 24952 24200
rect 25004 24148 25010 24200
rect 25222 24148 25228 24200
rect 25280 24148 25286 24200
rect 25314 24148 25320 24200
rect 25372 24148 25378 24200
rect 25958 24148 25964 24200
rect 26016 24148 26022 24200
rect 26050 24148 26056 24200
rect 26108 24148 26114 24200
rect 26329 24191 26387 24197
rect 26329 24157 26341 24191
rect 26375 24188 26387 24191
rect 26694 24188 26700 24200
rect 26375 24160 26700 24188
rect 26375 24157 26387 24160
rect 26329 24151 26387 24157
rect 26694 24148 26700 24160
rect 26752 24148 26758 24200
rect 28718 24148 28724 24200
rect 28776 24148 28782 24200
rect 28994 24148 29000 24200
rect 29052 24188 29058 24200
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 29052 24160 29745 24188
rect 29052 24148 29058 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 21223 24092 21864 24120
rect 21223 24089 21235 24092
rect 21177 24083 21235 24089
rect 21192 24052 21220 24083
rect 24394 24080 24400 24132
rect 24452 24120 24458 24132
rect 25133 24123 25191 24129
rect 25133 24120 25145 24123
rect 24452 24092 25145 24120
rect 24452 24080 24458 24092
rect 25133 24089 25145 24092
rect 25179 24120 25191 24123
rect 26145 24123 26203 24129
rect 26145 24120 26157 24123
rect 25179 24092 26157 24120
rect 25179 24089 25191 24092
rect 25133 24083 25191 24089
rect 26145 24089 26157 24092
rect 26191 24089 26203 24123
rect 29748 24120 29776 24151
rect 29822 24148 29828 24200
rect 29880 24148 29886 24200
rect 31386 24148 31392 24200
rect 31444 24188 31450 24200
rect 31481 24191 31539 24197
rect 31481 24188 31493 24191
rect 31444 24160 31493 24188
rect 31444 24148 31450 24160
rect 31481 24157 31493 24160
rect 31527 24157 31539 24191
rect 31481 24151 31539 24157
rect 31665 24123 31723 24129
rect 31665 24120 31677 24123
rect 29748 24092 31677 24120
rect 26145 24083 26203 24089
rect 31665 24089 31677 24092
rect 31711 24120 31723 24123
rect 31754 24120 31760 24132
rect 31711 24092 31760 24120
rect 31711 24089 31723 24092
rect 31665 24083 31723 24089
rect 31754 24080 31760 24092
rect 31812 24080 31818 24132
rect 34440 24120 34468 24364
rect 35250 24352 35256 24404
rect 35308 24392 35314 24404
rect 35345 24395 35403 24401
rect 35345 24392 35357 24395
rect 35308 24364 35357 24392
rect 35308 24352 35314 24364
rect 35345 24361 35357 24364
rect 35391 24361 35403 24395
rect 35345 24355 35403 24361
rect 35434 24352 35440 24404
rect 35492 24392 35498 24404
rect 36446 24392 36452 24404
rect 35492 24364 36452 24392
rect 35492 24352 35498 24364
rect 36446 24352 36452 24364
rect 36504 24352 36510 24404
rect 36538 24352 36544 24404
rect 36596 24352 36602 24404
rect 36633 24395 36691 24401
rect 36633 24361 36645 24395
rect 36679 24392 36691 24395
rect 36906 24392 36912 24404
rect 36679 24364 36912 24392
rect 36679 24361 36691 24364
rect 36633 24355 36691 24361
rect 34514 24284 34520 24336
rect 34572 24324 34578 24336
rect 35161 24327 35219 24333
rect 35161 24324 35173 24327
rect 34572 24296 35173 24324
rect 34572 24284 34578 24296
rect 35161 24293 35173 24296
rect 35207 24324 35219 24327
rect 36648 24324 36676 24355
rect 36906 24352 36912 24364
rect 36964 24352 36970 24404
rect 37645 24395 37703 24401
rect 37645 24361 37657 24395
rect 37691 24392 37703 24395
rect 37826 24392 37832 24404
rect 37691 24364 37832 24392
rect 37691 24361 37703 24364
rect 37645 24355 37703 24361
rect 37826 24352 37832 24364
rect 37884 24352 37890 24404
rect 41690 24352 41696 24404
rect 41748 24392 41754 24404
rect 42058 24392 42064 24404
rect 41748 24364 42064 24392
rect 41748 24352 41754 24364
rect 42058 24352 42064 24364
rect 42116 24392 42122 24404
rect 42153 24395 42211 24401
rect 42153 24392 42165 24395
rect 42116 24364 42165 24392
rect 42116 24352 42122 24364
rect 42153 24361 42165 24364
rect 42199 24361 42211 24395
rect 42153 24355 42211 24361
rect 35207 24296 36676 24324
rect 35207 24293 35219 24296
rect 35161 24287 35219 24293
rect 36722 24284 36728 24336
rect 36780 24284 36786 24336
rect 35618 24216 35624 24268
rect 35676 24256 35682 24268
rect 36081 24259 36139 24265
rect 36081 24256 36093 24259
rect 35676 24228 36093 24256
rect 35676 24216 35682 24228
rect 36081 24225 36093 24228
rect 36127 24225 36139 24259
rect 36081 24219 36139 24225
rect 36170 24216 36176 24268
rect 36228 24216 36234 24268
rect 36449 24259 36507 24265
rect 36449 24225 36461 24259
rect 36495 24256 36507 24259
rect 36740 24256 36768 24284
rect 36495 24228 36768 24256
rect 36495 24225 36507 24228
rect 36449 24219 36507 24225
rect 36262 24188 36268 24200
rect 35452 24160 36268 24188
rect 35313 24123 35371 24129
rect 35313 24120 35325 24123
rect 34440 24092 35325 24120
rect 35313 24089 35325 24092
rect 35359 24120 35371 24123
rect 35452 24120 35480 24160
rect 36262 24148 36268 24160
rect 36320 24148 36326 24200
rect 36538 24148 36544 24200
rect 36596 24188 36602 24200
rect 36725 24191 36783 24197
rect 36725 24188 36737 24191
rect 36596 24160 36737 24188
rect 36596 24148 36602 24160
rect 36725 24157 36737 24160
rect 36771 24157 36783 24191
rect 36725 24151 36783 24157
rect 37090 24148 37096 24200
rect 37148 24148 37154 24200
rect 37274 24148 37280 24200
rect 37332 24148 37338 24200
rect 37461 24191 37519 24197
rect 37461 24157 37473 24191
rect 37507 24188 37519 24191
rect 37550 24188 37556 24200
rect 37507 24160 37556 24188
rect 37507 24157 37519 24160
rect 37461 24151 37519 24157
rect 37550 24148 37556 24160
rect 37608 24148 37614 24200
rect 39390 24148 39396 24200
rect 39448 24188 39454 24200
rect 39942 24188 39948 24200
rect 39448 24160 39948 24188
rect 39448 24148 39454 24160
rect 39942 24148 39948 24160
rect 40000 24188 40006 24200
rect 40405 24191 40463 24197
rect 40405 24188 40417 24191
rect 40000 24160 40417 24188
rect 40000 24148 40006 24160
rect 40405 24157 40417 24160
rect 40451 24157 40463 24191
rect 40405 24151 40463 24157
rect 35359 24092 35480 24120
rect 35359 24089 35371 24092
rect 35313 24083 35371 24089
rect 35526 24080 35532 24132
rect 35584 24120 35590 24132
rect 36814 24120 36820 24132
rect 35584 24092 36820 24120
rect 35584 24080 35590 24092
rect 36814 24080 36820 24092
rect 36872 24080 36878 24132
rect 37369 24123 37427 24129
rect 37369 24089 37381 24123
rect 37415 24089 37427 24123
rect 37369 24083 37427 24089
rect 40681 24123 40739 24129
rect 40681 24089 40693 24123
rect 40727 24120 40739 24123
rect 40954 24120 40960 24132
rect 40727 24092 40960 24120
rect 40727 24089 40739 24092
rect 40681 24083 40739 24089
rect 19444 24024 21220 24052
rect 25777 24055 25835 24061
rect 25777 24021 25789 24055
rect 25823 24052 25835 24055
rect 26970 24052 26976 24064
rect 25823 24024 26976 24052
rect 25823 24021 25835 24024
rect 25777 24015 25835 24021
rect 26970 24012 26976 24024
rect 27028 24012 27034 24064
rect 28537 24055 28595 24061
rect 28537 24021 28549 24055
rect 28583 24052 28595 24055
rect 28810 24052 28816 24064
rect 28583 24024 28816 24052
rect 28583 24021 28595 24024
rect 28537 24015 28595 24021
rect 28810 24012 28816 24024
rect 28868 24012 28874 24064
rect 29822 24012 29828 24064
rect 29880 24052 29886 24064
rect 31573 24055 31631 24061
rect 31573 24052 31585 24055
rect 29880 24024 31585 24052
rect 29880 24012 29886 24024
rect 31573 24021 31585 24024
rect 31619 24021 31631 24055
rect 31573 24015 31631 24021
rect 35434 24012 35440 24064
rect 35492 24052 35498 24064
rect 35621 24055 35679 24061
rect 35621 24052 35633 24055
rect 35492 24024 35633 24052
rect 35492 24012 35498 24024
rect 35621 24021 35633 24024
rect 35667 24021 35679 24055
rect 35621 24015 35679 24021
rect 35989 24055 36047 24061
rect 35989 24021 36001 24055
rect 36035 24052 36047 24055
rect 36446 24052 36452 24064
rect 36035 24024 36452 24052
rect 36035 24021 36047 24024
rect 35989 24015 36047 24021
rect 36446 24012 36452 24024
rect 36504 24012 36510 24064
rect 37384 24052 37412 24083
rect 40954 24080 40960 24092
rect 41012 24080 41018 24132
rect 41414 24080 41420 24132
rect 41472 24080 41478 24132
rect 37458 24052 37464 24064
rect 37384 24024 37464 24052
rect 37458 24012 37464 24024
rect 37516 24012 37522 24064
rect 1104 23962 42504 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 42504 23962
rect 1104 23888 42504 23910
rect 2774 23848 2780 23860
rect 2746 23808 2780 23848
rect 2832 23808 2838 23860
rect 3050 23808 3056 23860
rect 3108 23808 3114 23860
rect 6457 23851 6515 23857
rect 6457 23817 6469 23851
rect 6503 23848 6515 23851
rect 6822 23848 6828 23860
rect 6503 23820 6828 23848
rect 6503 23817 6515 23820
rect 6457 23811 6515 23817
rect 6822 23808 6828 23820
rect 6880 23808 6886 23860
rect 6914 23808 6920 23860
rect 6972 23808 6978 23860
rect 7653 23851 7711 23857
rect 7653 23817 7665 23851
rect 7699 23848 7711 23851
rect 7834 23848 7840 23860
rect 7699 23820 7840 23848
rect 7699 23817 7711 23820
rect 7653 23811 7711 23817
rect 7834 23808 7840 23820
rect 7892 23808 7898 23860
rect 9232 23820 9536 23848
rect 2746 23780 2774 23808
rect 3418 23780 3424 23792
rect 2608 23752 3424 23780
rect 2608 23721 2636 23752
rect 3418 23740 3424 23752
rect 3476 23740 3482 23792
rect 6546 23780 6552 23792
rect 4908 23752 6552 23780
rect 2593 23715 2651 23721
rect 2593 23681 2605 23715
rect 2639 23681 2651 23715
rect 2593 23675 2651 23681
rect 2682 23672 2688 23724
rect 2740 23672 2746 23724
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23712 2835 23715
rect 3234 23712 3240 23724
rect 2823 23684 3240 23712
rect 2823 23681 2835 23684
rect 2777 23675 2835 23681
rect 3234 23672 3240 23684
rect 3292 23712 3298 23724
rect 4908 23721 4936 23752
rect 6546 23740 6552 23752
rect 6604 23740 6610 23792
rect 6932 23780 6960 23808
rect 6748 23752 6960 23780
rect 3605 23715 3663 23721
rect 3605 23712 3617 23715
rect 3292 23684 3617 23712
rect 3292 23672 3298 23684
rect 3605 23681 3617 23684
rect 3651 23681 3663 23715
rect 3605 23675 3663 23681
rect 4893 23715 4951 23721
rect 4893 23681 4905 23715
rect 4939 23681 4951 23715
rect 4893 23675 4951 23681
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5258 23712 5264 23724
rect 5123 23684 5264 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 6270 23672 6276 23724
rect 6328 23712 6334 23724
rect 6748 23721 6776 23752
rect 7282 23740 7288 23792
rect 7340 23780 7346 23792
rect 9099 23783 9157 23789
rect 7340 23752 8616 23780
rect 7340 23740 7346 23752
rect 6457 23715 6515 23721
rect 6457 23712 6469 23715
rect 6328 23684 6469 23712
rect 6328 23672 6334 23684
rect 6457 23681 6469 23684
rect 6503 23681 6515 23715
rect 6457 23675 6515 23681
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23681 6791 23715
rect 6733 23675 6791 23681
rect 6822 23672 6828 23724
rect 6880 23672 6886 23724
rect 7374 23672 7380 23724
rect 7432 23712 7438 23724
rect 7469 23715 7527 23721
rect 7469 23712 7481 23715
rect 7432 23684 7481 23712
rect 7432 23672 7438 23684
rect 7469 23681 7481 23684
rect 7515 23681 7527 23715
rect 7469 23675 7527 23681
rect 7745 23715 7803 23721
rect 7745 23681 7757 23715
rect 7791 23712 7803 23715
rect 7926 23712 7932 23724
rect 7791 23684 7932 23712
rect 7791 23681 7803 23684
rect 7745 23675 7803 23681
rect 7926 23672 7932 23684
rect 7984 23672 7990 23724
rect 8588 23712 8616 23752
rect 9099 23749 9111 23783
rect 9145 23780 9157 23783
rect 9232 23780 9260 23820
rect 9145 23752 9260 23780
rect 9145 23749 9157 23752
rect 9099 23743 9157 23749
rect 9306 23740 9312 23792
rect 9364 23740 9370 23792
rect 9508 23780 9536 23820
rect 9582 23808 9588 23860
rect 9640 23808 9646 23860
rect 11790 23808 11796 23860
rect 11848 23808 11854 23860
rect 12253 23851 12311 23857
rect 12253 23817 12265 23851
rect 12299 23848 12311 23851
rect 13262 23848 13268 23860
rect 12299 23820 13268 23848
rect 12299 23817 12311 23820
rect 12253 23811 12311 23817
rect 13262 23808 13268 23820
rect 13320 23848 13326 23860
rect 13320 23820 14964 23848
rect 13320 23808 13326 23820
rect 11422 23780 11428 23792
rect 9508 23752 11428 23780
rect 11422 23740 11428 23752
rect 11480 23740 11486 23792
rect 14936 23780 14964 23820
rect 15010 23808 15016 23860
rect 15068 23848 15074 23860
rect 16301 23851 16359 23857
rect 16301 23848 16313 23851
rect 15068 23820 16313 23848
rect 15068 23808 15074 23820
rect 16301 23817 16313 23820
rect 16347 23848 16359 23851
rect 16347 23820 18276 23848
rect 16347 23817 16359 23820
rect 16301 23811 16359 23817
rect 18248 23792 18276 23820
rect 18414 23808 18420 23860
rect 18472 23848 18478 23860
rect 18690 23848 18696 23860
rect 18472 23820 18696 23848
rect 18472 23808 18478 23820
rect 18690 23808 18696 23820
rect 18748 23808 18754 23860
rect 18966 23808 18972 23860
rect 19024 23808 19030 23860
rect 19996 23820 22324 23848
rect 14936 23752 15424 23780
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 8588 23684 9229 23712
rect 9217 23681 9229 23684
rect 9263 23681 9275 23715
rect 9217 23675 9275 23681
rect 9401 23715 9459 23721
rect 9401 23681 9413 23715
rect 9447 23712 9459 23715
rect 9490 23712 9496 23724
rect 9447 23684 9496 23712
rect 9447 23681 9459 23684
rect 9401 23675 9459 23681
rect 2700 23644 2728 23672
rect 3142 23644 3148 23656
rect 2700 23616 3148 23644
rect 3142 23604 3148 23616
rect 3200 23644 3206 23656
rect 3326 23644 3332 23656
rect 3200 23616 3332 23644
rect 3200 23604 3206 23616
rect 3326 23604 3332 23616
rect 3384 23604 3390 23656
rect 3694 23604 3700 23656
rect 3752 23644 3758 23656
rect 3752 23616 3924 23644
rect 3752 23604 3758 23616
rect 2958 23536 2964 23588
rect 3016 23576 3022 23588
rect 3786 23576 3792 23588
rect 3016 23548 3792 23576
rect 3016 23536 3022 23548
rect 3786 23536 3792 23548
rect 3844 23536 3850 23588
rect 3896 23576 3924 23616
rect 5166 23604 5172 23656
rect 5224 23644 5230 23656
rect 6288 23644 6316 23672
rect 5224 23616 6316 23644
rect 5224 23604 5230 23616
rect 6546 23604 6552 23656
rect 6604 23644 6610 23656
rect 7098 23644 7104 23656
rect 6604 23616 7104 23644
rect 6604 23604 6610 23616
rect 7098 23604 7104 23616
rect 7156 23604 7162 23656
rect 7190 23604 7196 23656
rect 7248 23604 7254 23656
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9122 23644 9128 23656
rect 8987 23616 9128 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 9232 23644 9260 23675
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 9674 23672 9680 23724
rect 9732 23712 9738 23724
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 9732 23684 9781 23712
rect 9732 23672 9738 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9858 23672 9864 23724
rect 9916 23712 9922 23724
rect 10025 23715 10083 23721
rect 10025 23712 10037 23715
rect 9916 23684 10037 23712
rect 9916 23672 9922 23684
rect 10025 23681 10037 23684
rect 10071 23681 10083 23715
rect 10025 23675 10083 23681
rect 11054 23672 11060 23724
rect 11112 23712 11118 23724
rect 12161 23715 12219 23721
rect 12161 23712 12173 23715
rect 11112 23684 12173 23712
rect 11112 23672 11118 23684
rect 12161 23681 12173 23684
rect 12207 23681 12219 23715
rect 12161 23675 12219 23681
rect 13722 23672 13728 23724
rect 13780 23672 13786 23724
rect 13998 23721 14004 23724
rect 13992 23712 14004 23721
rect 13959 23684 14004 23712
rect 13992 23675 14004 23684
rect 13998 23672 14004 23675
rect 14056 23672 14062 23724
rect 9306 23644 9312 23656
rect 9232 23616 9312 23644
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 12434 23604 12440 23656
rect 12492 23604 12498 23656
rect 15396 23644 15424 23752
rect 16942 23740 16948 23792
rect 17000 23740 17006 23792
rect 18230 23740 18236 23792
rect 18288 23780 18294 23792
rect 19996 23780 20024 23820
rect 18288 23752 20024 23780
rect 18288 23740 18294 23752
rect 15562 23672 15568 23724
rect 15620 23672 15626 23724
rect 16390 23672 16396 23724
rect 16448 23672 16454 23724
rect 16666 23712 16672 23724
rect 16724 23721 16730 23724
rect 16500 23684 16672 23712
rect 15396 23616 15608 23644
rect 8570 23576 8576 23588
rect 3896 23548 8576 23576
rect 8570 23536 8576 23548
rect 8628 23536 8634 23588
rect 4982 23468 4988 23520
rect 5040 23468 5046 23520
rect 7377 23511 7435 23517
rect 7377 23477 7389 23511
rect 7423 23508 7435 23511
rect 7834 23508 7840 23520
rect 7423 23480 7840 23508
rect 7423 23477 7435 23480
rect 7377 23471 7435 23477
rect 7834 23468 7840 23480
rect 7892 23468 7898 23520
rect 10502 23468 10508 23520
rect 10560 23508 10566 23520
rect 11149 23511 11207 23517
rect 11149 23508 11161 23511
rect 10560 23480 11161 23508
rect 10560 23468 10566 23480
rect 11149 23477 11161 23480
rect 11195 23477 11207 23511
rect 11149 23471 11207 23477
rect 14734 23468 14740 23520
rect 14792 23508 14798 23520
rect 15102 23508 15108 23520
rect 14792 23480 15108 23508
rect 14792 23468 14798 23480
rect 15102 23468 15108 23480
rect 15160 23468 15166 23520
rect 15194 23468 15200 23520
rect 15252 23468 15258 23520
rect 15580 23508 15608 23616
rect 15654 23604 15660 23656
rect 15712 23604 15718 23656
rect 15746 23604 15752 23656
rect 15804 23604 15810 23656
rect 15930 23604 15936 23656
rect 15988 23644 15994 23656
rect 16500 23644 16528 23684
rect 16666 23672 16672 23684
rect 16724 23675 16734 23721
rect 16724 23672 16730 23675
rect 18046 23672 18052 23724
rect 18104 23672 18110 23724
rect 18598 23672 18604 23724
rect 18656 23672 18662 23724
rect 18690 23672 18696 23724
rect 18748 23712 18754 23724
rect 19996 23721 20024 23752
rect 20070 23740 20076 23792
rect 20128 23740 20134 23792
rect 22296 23780 22324 23820
rect 22370 23808 22376 23860
rect 22428 23808 22434 23860
rect 24486 23848 24492 23860
rect 22848 23820 24492 23848
rect 22848 23780 22876 23820
rect 24486 23808 24492 23820
rect 24544 23848 24550 23860
rect 25958 23848 25964 23860
rect 24544 23820 25964 23848
rect 24544 23808 24550 23820
rect 25958 23808 25964 23820
rect 26016 23808 26022 23860
rect 26786 23808 26792 23860
rect 26844 23848 26850 23860
rect 26973 23851 27031 23857
rect 26973 23848 26985 23851
rect 26844 23820 26985 23848
rect 26844 23808 26850 23820
rect 26973 23817 26985 23820
rect 27019 23848 27031 23851
rect 28994 23848 29000 23860
rect 27019 23820 29000 23848
rect 27019 23817 27031 23820
rect 26973 23811 27031 23817
rect 28994 23808 29000 23820
rect 29052 23808 29058 23860
rect 29641 23851 29699 23857
rect 29641 23817 29653 23851
rect 29687 23848 29699 23851
rect 29914 23848 29920 23860
rect 29687 23820 29920 23848
rect 29687 23817 29699 23820
rect 29641 23811 29699 23817
rect 29914 23808 29920 23820
rect 29972 23808 29978 23860
rect 32306 23808 32312 23860
rect 32364 23848 32370 23860
rect 32364 23820 35112 23848
rect 32364 23808 32370 23820
rect 22296 23752 22876 23780
rect 22922 23740 22928 23792
rect 22980 23780 22986 23792
rect 22980 23752 23506 23780
rect 22980 23740 22986 23752
rect 24578 23740 24584 23792
rect 24636 23780 24642 23792
rect 24673 23783 24731 23789
rect 24673 23780 24685 23783
rect 24636 23752 24685 23780
rect 24636 23740 24642 23752
rect 24673 23749 24685 23752
rect 24719 23749 24731 23783
rect 24673 23743 24731 23749
rect 25314 23740 25320 23792
rect 25372 23780 25378 23792
rect 33778 23780 33784 23792
rect 25372 23752 33784 23780
rect 25372 23740 25378 23752
rect 33778 23740 33784 23752
rect 33836 23740 33842 23792
rect 35084 23789 35112 23820
rect 38194 23808 38200 23860
rect 38252 23848 38258 23860
rect 38381 23851 38439 23857
rect 38381 23848 38393 23851
rect 38252 23820 38393 23848
rect 38252 23808 38258 23820
rect 38381 23817 38393 23820
rect 38427 23817 38439 23851
rect 38381 23811 38439 23817
rect 40954 23808 40960 23860
rect 41012 23808 41018 23860
rect 41322 23808 41328 23860
rect 41380 23808 41386 23860
rect 35069 23783 35127 23789
rect 35069 23749 35081 23783
rect 35115 23749 35127 23783
rect 35069 23743 35127 23749
rect 35158 23740 35164 23792
rect 35216 23780 35222 23792
rect 37734 23780 37740 23792
rect 35216 23752 37740 23780
rect 35216 23740 35222 23752
rect 37734 23740 37740 23752
rect 37792 23740 37798 23792
rect 18785 23715 18843 23721
rect 18785 23712 18797 23715
rect 18748 23684 18797 23712
rect 18748 23672 18754 23684
rect 18785 23681 18797 23684
rect 18831 23681 18843 23715
rect 18785 23675 18843 23681
rect 19981 23715 20039 23721
rect 19981 23681 19993 23715
rect 20027 23681 20039 23715
rect 19981 23675 20039 23681
rect 20162 23672 20168 23724
rect 20220 23672 20226 23724
rect 20349 23715 20407 23721
rect 20349 23681 20361 23715
rect 20395 23712 20407 23715
rect 21082 23712 21088 23724
rect 20395 23684 21088 23712
rect 20395 23681 20407 23684
rect 20349 23675 20407 23681
rect 21082 23672 21088 23684
rect 21140 23672 21146 23724
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23712 25007 23715
rect 26418 23712 26424 23724
rect 24995 23684 26424 23712
rect 24995 23681 25007 23684
rect 24949 23675 25007 23681
rect 26418 23672 26424 23684
rect 26476 23672 26482 23724
rect 28097 23715 28155 23721
rect 28097 23681 28109 23715
rect 28143 23712 28155 23715
rect 28258 23712 28264 23724
rect 28143 23684 28264 23712
rect 28143 23681 28155 23684
rect 28097 23675 28155 23681
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 28994 23672 29000 23724
rect 29052 23672 29058 23724
rect 32125 23715 32183 23721
rect 32125 23681 32137 23715
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 15988 23616 16528 23644
rect 15988 23604 15994 23616
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 20530 23644 20536 23656
rect 16632 23616 20536 23644
rect 16632 23604 16638 23616
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 21358 23604 21364 23656
rect 21416 23604 21422 23656
rect 22462 23604 22468 23656
rect 22520 23604 22526 23656
rect 22557 23647 22615 23653
rect 22557 23613 22569 23647
rect 22603 23613 22615 23647
rect 22557 23607 22615 23613
rect 25685 23647 25743 23653
rect 25685 23613 25697 23647
rect 25731 23644 25743 23647
rect 25774 23644 25780 23656
rect 25731 23616 25780 23644
rect 25731 23613 25743 23616
rect 25685 23607 25743 23613
rect 15764 23576 15792 23604
rect 16666 23576 16672 23588
rect 15764 23548 16672 23576
rect 16666 23536 16672 23548
rect 16724 23536 16730 23588
rect 17954 23536 17960 23588
rect 18012 23576 18018 23588
rect 21910 23576 21916 23588
rect 18012 23548 21916 23576
rect 18012 23536 18018 23548
rect 21910 23536 21916 23548
rect 21968 23576 21974 23588
rect 22572 23576 22600 23607
rect 25774 23604 25780 23616
rect 25832 23604 25838 23656
rect 25866 23604 25872 23656
rect 25924 23604 25930 23656
rect 28353 23647 28411 23653
rect 28353 23613 28365 23647
rect 28399 23613 28411 23647
rect 28353 23607 28411 23613
rect 21968 23548 22600 23576
rect 23201 23579 23259 23585
rect 21968 23536 21974 23548
rect 23201 23545 23213 23579
rect 23247 23576 23259 23579
rect 23566 23576 23572 23588
rect 23247 23548 23572 23576
rect 23247 23545 23259 23548
rect 23201 23539 23259 23545
rect 23566 23536 23572 23548
rect 23624 23536 23630 23588
rect 28368 23576 28396 23607
rect 28810 23604 28816 23656
rect 28868 23644 28874 23656
rect 29365 23647 29423 23653
rect 29365 23644 29377 23647
rect 28868 23616 29377 23644
rect 28868 23604 28874 23616
rect 29365 23613 29377 23616
rect 29411 23613 29423 23647
rect 29365 23607 29423 23613
rect 29549 23647 29607 23653
rect 29549 23613 29561 23647
rect 29595 23613 29607 23647
rect 29549 23607 29607 23613
rect 28994 23576 29000 23588
rect 28368 23548 29000 23576
rect 19702 23508 19708 23520
rect 15580 23480 19708 23508
rect 19702 23468 19708 23480
rect 19760 23468 19766 23520
rect 19797 23511 19855 23517
rect 19797 23477 19809 23511
rect 19843 23508 19855 23511
rect 20070 23508 20076 23520
rect 19843 23480 20076 23508
rect 19843 23477 19855 23480
rect 19797 23471 19855 23477
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 21082 23508 21088 23520
rect 20855 23480 21088 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 21082 23468 21088 23480
rect 21140 23468 21146 23520
rect 22002 23468 22008 23520
rect 22060 23468 22066 23520
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 25041 23511 25099 23517
rect 25041 23508 25053 23511
rect 24912 23480 25053 23508
rect 24912 23468 24918 23480
rect 25041 23477 25053 23480
rect 25087 23477 25099 23511
rect 25041 23471 25099 23477
rect 26513 23511 26571 23517
rect 26513 23477 26525 23511
rect 26559 23508 26571 23511
rect 26694 23508 26700 23520
rect 26559 23480 26700 23508
rect 26559 23477 26571 23480
rect 26513 23471 26571 23477
rect 26694 23468 26700 23480
rect 26752 23468 26758 23520
rect 27430 23468 27436 23520
rect 27488 23508 27494 23520
rect 28368 23508 28396 23548
rect 28994 23536 29000 23548
rect 29052 23536 29058 23588
rect 29564 23576 29592 23607
rect 30926 23604 30932 23656
rect 30984 23604 30990 23656
rect 32140 23644 32168 23675
rect 32306 23672 32312 23724
rect 32364 23672 32370 23724
rect 32398 23672 32404 23724
rect 32456 23672 32462 23724
rect 32490 23672 32496 23724
rect 32548 23712 32554 23724
rect 34885 23715 34943 23721
rect 34885 23712 34897 23715
rect 32548 23684 34897 23712
rect 32548 23672 32554 23684
rect 34885 23681 34897 23684
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 34977 23715 35035 23721
rect 34977 23681 34989 23715
rect 35023 23712 35035 23715
rect 35176 23712 35204 23740
rect 35023 23684 35204 23712
rect 35253 23715 35311 23721
rect 35023 23681 35035 23684
rect 34977 23675 35035 23681
rect 35253 23681 35265 23715
rect 35299 23712 35311 23715
rect 35342 23712 35348 23724
rect 35299 23684 35348 23712
rect 35299 23681 35311 23684
rect 35253 23675 35311 23681
rect 35342 23672 35348 23684
rect 35400 23672 35406 23724
rect 38286 23672 38292 23724
rect 38344 23712 38350 23724
rect 39390 23712 39396 23724
rect 38344 23684 39396 23712
rect 38344 23672 38350 23684
rect 39390 23672 39396 23684
rect 39448 23672 39454 23724
rect 39666 23721 39672 23724
rect 39660 23675 39672 23721
rect 39666 23672 39672 23675
rect 39724 23672 39730 23724
rect 33413 23647 33471 23653
rect 33413 23644 33425 23647
rect 32140 23616 33425 23644
rect 32416 23588 32444 23616
rect 33413 23613 33425 23616
rect 33459 23613 33471 23647
rect 33413 23607 33471 23613
rect 34057 23647 34115 23653
rect 34057 23613 34069 23647
rect 34103 23644 34115 23647
rect 34514 23644 34520 23656
rect 34103 23616 34520 23644
rect 34103 23613 34115 23616
rect 34057 23607 34115 23613
rect 34514 23604 34520 23616
rect 34572 23604 34578 23656
rect 38473 23647 38531 23653
rect 38473 23644 38485 23647
rect 38396 23616 38485 23644
rect 38396 23588 38424 23616
rect 38473 23613 38485 23616
rect 38519 23613 38531 23647
rect 38473 23607 38531 23613
rect 38562 23604 38568 23656
rect 38620 23604 38626 23656
rect 41414 23604 41420 23656
rect 41472 23604 41478 23656
rect 41506 23604 41512 23656
rect 41564 23604 41570 23656
rect 29914 23576 29920 23588
rect 29564 23548 29920 23576
rect 29914 23536 29920 23548
rect 29972 23576 29978 23588
rect 30285 23579 30343 23585
rect 30285 23576 30297 23579
rect 29972 23548 30297 23576
rect 29972 23536 29978 23548
rect 30285 23545 30297 23548
rect 30331 23545 30343 23579
rect 30285 23539 30343 23545
rect 32398 23536 32404 23588
rect 32456 23536 32462 23588
rect 38378 23536 38384 23588
rect 38436 23536 38442 23588
rect 27488 23480 28396 23508
rect 28445 23511 28503 23517
rect 27488 23468 27494 23480
rect 28445 23477 28457 23511
rect 28491 23508 28503 23511
rect 28902 23508 28908 23520
rect 28491 23480 28908 23508
rect 28491 23477 28503 23480
rect 28445 23471 28503 23477
rect 28902 23468 28908 23480
rect 28960 23468 28966 23520
rect 30006 23468 30012 23520
rect 30064 23468 30070 23520
rect 32677 23511 32735 23517
rect 32677 23477 32689 23511
rect 32723 23508 32735 23511
rect 33318 23508 33324 23520
rect 32723 23480 33324 23508
rect 32723 23477 32735 23480
rect 32677 23471 32735 23477
rect 33318 23468 33324 23480
rect 33376 23468 33382 23520
rect 34698 23468 34704 23520
rect 34756 23468 34762 23520
rect 37918 23468 37924 23520
rect 37976 23508 37982 23520
rect 38013 23511 38071 23517
rect 38013 23508 38025 23511
rect 37976 23480 38025 23508
rect 37976 23468 37982 23480
rect 38013 23477 38025 23480
rect 38059 23477 38071 23511
rect 38013 23471 38071 23477
rect 40770 23468 40776 23520
rect 40828 23468 40834 23520
rect 1104 23418 42504 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 42504 23418
rect 1104 23344 42504 23366
rect 3234 23264 3240 23316
rect 3292 23304 3298 23316
rect 3329 23307 3387 23313
rect 3329 23304 3341 23307
rect 3292 23276 3341 23304
rect 3292 23264 3298 23276
rect 3329 23273 3341 23276
rect 3375 23273 3387 23307
rect 3329 23267 3387 23273
rect 6454 23264 6460 23316
rect 6512 23304 6518 23316
rect 7190 23304 7196 23316
rect 6512 23276 7196 23304
rect 6512 23264 6518 23276
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 7469 23307 7527 23313
rect 7469 23273 7481 23307
rect 7515 23304 7527 23307
rect 7742 23304 7748 23316
rect 7515 23276 7748 23304
rect 7515 23273 7527 23276
rect 7469 23267 7527 23273
rect 7742 23264 7748 23276
rect 7800 23304 7806 23316
rect 8202 23304 8208 23316
rect 7800 23276 8208 23304
rect 7800 23264 7806 23276
rect 8202 23264 8208 23276
rect 8260 23264 8266 23316
rect 9769 23307 9827 23313
rect 9769 23273 9781 23307
rect 9815 23304 9827 23307
rect 9858 23304 9864 23316
rect 9815 23276 9864 23304
rect 9815 23273 9827 23276
rect 9769 23267 9827 23273
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 11054 23264 11060 23316
rect 11112 23264 11118 23316
rect 13722 23264 13728 23316
rect 13780 23304 13786 23316
rect 15565 23307 15623 23313
rect 13780 23276 15516 23304
rect 13780 23264 13786 23276
rect 2869 23239 2927 23245
rect 2869 23205 2881 23239
rect 2915 23236 2927 23239
rect 3694 23236 3700 23248
rect 2915 23208 3700 23236
rect 2915 23205 2927 23208
rect 2869 23199 2927 23205
rect 3694 23196 3700 23208
rect 3752 23196 3758 23248
rect 8294 23196 8300 23248
rect 8352 23236 8358 23248
rect 12710 23236 12716 23248
rect 8352 23208 12716 23236
rect 8352 23196 8358 23208
rect 12710 23196 12716 23208
rect 12768 23196 12774 23248
rect 15488 23236 15516 23276
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 15654 23304 15660 23316
rect 15611 23276 15660 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 18598 23304 18604 23316
rect 16040 23276 18604 23304
rect 15930 23236 15936 23248
rect 15488 23208 15936 23236
rect 2774 23168 2780 23180
rect 2608 23140 2780 23168
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 2608 23109 2636 23140
rect 2774 23128 2780 23140
rect 2832 23168 2838 23180
rect 4341 23171 4399 23177
rect 2832 23140 3372 23168
rect 2832 23128 2838 23140
rect 2501 23103 2559 23109
rect 2501 23069 2513 23103
rect 2547 23069 2559 23103
rect 2501 23063 2559 23069
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 3234 23100 3240 23112
rect 2731 23072 3240 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 2516 23032 2544 23063
rect 3234 23060 3240 23072
rect 3292 23060 3298 23112
rect 2961 23035 3019 23041
rect 2961 23032 2973 23035
rect 2516 23004 2973 23032
rect 2961 23001 2973 23004
rect 3007 23032 3019 23035
rect 3142 23032 3148 23044
rect 3007 23004 3148 23032
rect 3007 23001 3019 23004
rect 2961 22995 3019 23001
rect 3142 22992 3148 23004
rect 3200 22992 3206 23044
rect 3344 23041 3372 23140
rect 4341 23137 4353 23171
rect 4387 23168 4399 23171
rect 4614 23168 4620 23180
rect 4387 23140 4620 23168
rect 4387 23137 4399 23140
rect 4341 23131 4399 23137
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 4709 23171 4767 23177
rect 4709 23137 4721 23171
rect 4755 23168 4767 23171
rect 4982 23168 4988 23180
rect 4755 23140 4988 23168
rect 4755 23137 4767 23140
rect 4709 23131 4767 23137
rect 4982 23128 4988 23140
rect 5040 23128 5046 23180
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23168 6423 23171
rect 10502 23168 10508 23180
rect 6411 23140 7696 23168
rect 6411 23137 6423 23140
rect 6365 23131 6423 23137
rect 7668 23112 7696 23140
rect 8496 23140 10508 23168
rect 3602 23060 3608 23112
rect 3660 23060 3666 23112
rect 3786 23060 3792 23112
rect 3844 23060 3850 23112
rect 6273 23103 6331 23109
rect 6273 23069 6285 23103
rect 6319 23069 6331 23103
rect 6273 23063 6331 23069
rect 3338 23035 3396 23041
rect 3338 23001 3350 23035
rect 3384 23001 3396 23035
rect 3338 22995 3396 23001
rect 5074 22992 5080 23044
rect 5132 22992 5138 23044
rect 5902 22992 5908 23044
rect 5960 23032 5966 23044
rect 6135 23035 6193 23041
rect 6135 23032 6147 23035
rect 5960 23004 6147 23032
rect 5960 22992 5966 23004
rect 6135 23001 6147 23004
rect 6181 23032 6193 23035
rect 6288 23032 6316 23063
rect 6454 23060 6460 23112
rect 6512 23060 6518 23112
rect 6822 23060 6828 23112
rect 6880 23060 6886 23112
rect 7006 23060 7012 23112
rect 7064 23100 7070 23112
rect 7064 23072 7620 23100
rect 7064 23060 7070 23072
rect 6730 23032 6736 23044
rect 6181 23004 6736 23032
rect 6181 23001 6193 23004
rect 6135 22995 6193 23001
rect 6730 22992 6736 23004
rect 6788 23032 6794 23044
rect 7098 23032 7104 23044
rect 6788 23004 7104 23032
rect 6788 22992 6794 23004
rect 7098 22992 7104 23004
rect 7156 22992 7162 23044
rect 7190 22992 7196 23044
rect 7248 23032 7254 23044
rect 7285 23035 7343 23041
rect 7285 23032 7297 23035
rect 7248 23004 7297 23032
rect 7248 22992 7254 23004
rect 7285 23001 7297 23004
rect 7331 23001 7343 23035
rect 7592 23032 7620 23072
rect 7650 23060 7656 23112
rect 7708 23060 7714 23112
rect 7926 23060 7932 23112
rect 7984 23060 7990 23112
rect 8496 23109 8524 23140
rect 10502 23128 10508 23140
rect 10560 23128 10566 23180
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12529 23171 12587 23177
rect 12529 23168 12541 23171
rect 12492 23140 12541 23168
rect 12492 23128 12498 23140
rect 12529 23137 12541 23140
rect 12575 23168 12587 23171
rect 12986 23168 12992 23180
rect 12575 23140 12992 23168
rect 12575 23137 12587 23140
rect 12529 23131 12587 23137
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 15488 23177 15516 23208
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23137 15531 23171
rect 15473 23131 15531 23137
rect 8113 23103 8171 23109
rect 8113 23069 8125 23103
rect 8159 23100 8171 23103
rect 8205 23103 8263 23109
rect 8205 23100 8217 23103
rect 8159 23072 8217 23100
rect 8159 23069 8171 23072
rect 8113 23063 8171 23069
rect 8205 23069 8217 23072
rect 8251 23069 8263 23103
rect 8205 23063 8263 23069
rect 8481 23103 8539 23109
rect 8481 23069 8493 23103
rect 8527 23069 8539 23103
rect 8481 23063 8539 23069
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23069 8631 23103
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 8573 23063 8631 23069
rect 8772 23072 9229 23100
rect 7592 23004 8340 23032
rect 7285 22995 7343 23001
rect 842 22924 848 22976
rect 900 22964 906 22976
rect 1581 22967 1639 22973
rect 1581 22964 1593 22967
rect 900 22936 1593 22964
rect 900 22924 906 22936
rect 1581 22933 1593 22936
rect 1627 22933 1639 22967
rect 1581 22927 1639 22933
rect 3973 22967 4031 22973
rect 3973 22933 3985 22967
rect 4019 22964 4031 22967
rect 5626 22964 5632 22976
rect 4019 22936 5632 22964
rect 4019 22933 4031 22936
rect 3973 22927 4031 22933
rect 5626 22924 5632 22936
rect 5684 22924 5690 22976
rect 6641 22967 6699 22973
rect 6641 22933 6653 22967
rect 6687 22964 6699 22967
rect 6914 22964 6920 22976
rect 6687 22936 6920 22964
rect 6687 22933 6699 22936
rect 6641 22927 6699 22933
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 7374 22924 7380 22976
rect 7432 22964 7438 22976
rect 7745 22967 7803 22973
rect 7745 22964 7757 22967
rect 7432 22936 7757 22964
rect 7432 22924 7438 22936
rect 7745 22933 7757 22936
rect 7791 22933 7803 22967
rect 8312 22964 8340 23004
rect 8386 22992 8392 23044
rect 8444 22992 8450 23044
rect 8588 22964 8616 23063
rect 8662 22964 8668 22976
rect 8312 22936 8668 22964
rect 7745 22927 7803 22933
rect 8662 22924 8668 22936
rect 8720 22924 8726 22976
rect 8772 22973 8800 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 9364 23072 9413 23100
rect 9364 23060 9370 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 11054 23100 11060 23112
rect 9631 23072 11060 23100
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 15194 23060 15200 23112
rect 15252 23109 15258 23112
rect 15252 23100 15264 23109
rect 15252 23072 15297 23100
rect 15252 23063 15264 23072
rect 15252 23060 15258 23063
rect 9122 22992 9128 23044
rect 9180 23032 9186 23044
rect 9493 23035 9551 23041
rect 9493 23032 9505 23035
rect 9180 23004 9505 23032
rect 9180 22992 9186 23004
rect 9493 23001 9505 23004
rect 9539 23001 9551 23035
rect 12253 23035 12311 23041
rect 12253 23032 12265 23035
rect 9493 22995 9551 23001
rect 11808 23004 12265 23032
rect 8757 22967 8815 22973
rect 8757 22933 8769 22967
rect 8803 22933 8815 22967
rect 8757 22927 8815 22933
rect 11422 22924 11428 22976
rect 11480 22964 11486 22976
rect 11808 22973 11836 23004
rect 12253 23001 12265 23004
rect 12299 23001 12311 23035
rect 16040 23032 16068 23276
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 23106 23264 23112 23316
rect 23164 23304 23170 23316
rect 23201 23307 23259 23313
rect 23201 23304 23213 23307
rect 23164 23276 23213 23304
rect 23164 23264 23170 23276
rect 23201 23273 23213 23276
rect 23247 23304 23259 23307
rect 23290 23304 23296 23316
rect 23247 23276 23296 23304
rect 23247 23273 23259 23276
rect 23201 23267 23259 23273
rect 23290 23264 23296 23276
rect 23348 23264 23354 23316
rect 28258 23264 28264 23316
rect 28316 23304 28322 23316
rect 28353 23307 28411 23313
rect 28353 23304 28365 23307
rect 28316 23276 28365 23304
rect 28316 23264 28322 23276
rect 28353 23273 28365 23276
rect 28399 23273 28411 23307
rect 28353 23267 28411 23273
rect 28552 23276 30604 23304
rect 17218 23196 17224 23248
rect 17276 23236 17282 23248
rect 17276 23208 18368 23236
rect 17276 23196 17282 23208
rect 17586 23128 17592 23180
rect 17644 23168 17650 23180
rect 18233 23171 18291 23177
rect 18233 23168 18245 23171
rect 17644 23140 18245 23168
rect 17644 23128 17650 23140
rect 18233 23137 18245 23140
rect 18279 23137 18291 23171
rect 18340 23168 18368 23208
rect 27249 23171 27307 23177
rect 18340 23140 20576 23168
rect 18233 23131 18291 23137
rect 16117 23103 16175 23109
rect 16117 23069 16129 23103
rect 16163 23069 16175 23103
rect 16117 23063 16175 23069
rect 12253 22995 12311 23001
rect 13280 23004 16068 23032
rect 13280 22976 13308 23004
rect 11793 22967 11851 22973
rect 11793 22964 11805 22967
rect 11480 22936 11805 22964
rect 11480 22924 11486 22936
rect 11793 22933 11805 22936
rect 11839 22933 11851 22967
rect 11793 22927 11851 22933
rect 11882 22924 11888 22976
rect 11940 22924 11946 22976
rect 12345 22967 12403 22973
rect 12345 22933 12357 22967
rect 12391 22964 12403 22967
rect 13262 22964 13268 22976
rect 12391 22936 13268 22964
rect 12391 22933 12403 22936
rect 12345 22927 12403 22933
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 14093 22967 14151 22973
rect 14093 22933 14105 22967
rect 14139 22964 14151 22967
rect 14826 22964 14832 22976
rect 14139 22936 14832 22964
rect 14139 22933 14151 22936
rect 14093 22927 14151 22933
rect 14826 22924 14832 22936
rect 14884 22964 14890 22976
rect 16132 22964 16160 23063
rect 17494 23060 17500 23112
rect 17552 23060 17558 23112
rect 19794 23060 19800 23112
rect 19852 23060 19858 23112
rect 19886 23060 19892 23112
rect 19944 23100 19950 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 19944 23072 20453 23100
rect 19944 23060 19950 23072
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20548 23100 20576 23140
rect 27249 23137 27261 23171
rect 27295 23168 27307 23171
rect 27430 23168 27436 23180
rect 27295 23140 27436 23168
rect 27295 23137 27307 23140
rect 27249 23131 27307 23137
rect 27430 23128 27436 23140
rect 27488 23128 27494 23180
rect 21913 23103 21971 23109
rect 21913 23100 21925 23103
rect 20548 23072 21925 23100
rect 20441 23063 20499 23069
rect 21913 23069 21925 23072
rect 21959 23069 21971 23103
rect 21913 23063 21971 23069
rect 24397 23103 24455 23109
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 26418 23100 26424 23112
rect 24443 23072 26424 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 26970 23060 26976 23112
rect 27028 23109 27034 23112
rect 28552 23109 28580 23276
rect 27028 23100 27040 23109
rect 28537 23103 28595 23109
rect 28537 23100 28549 23103
rect 27028 23072 27073 23100
rect 27172 23072 28549 23100
rect 27028 23063 27040 23072
rect 27028 23060 27034 23063
rect 20708 23035 20766 23041
rect 20708 23001 20720 23035
rect 20754 23032 20766 23035
rect 22002 23032 22008 23044
rect 20754 23004 22008 23032
rect 20754 23001 20766 23004
rect 20708 22995 20766 23001
rect 22002 22992 22008 23004
rect 22060 22992 22066 23044
rect 24486 22992 24492 23044
rect 24544 23032 24550 23044
rect 24642 23035 24700 23041
rect 24642 23032 24654 23035
rect 24544 23004 24654 23032
rect 24544 22992 24550 23004
rect 24642 23001 24654 23004
rect 24688 23001 24700 23035
rect 24642 22995 24700 23001
rect 25958 22992 25964 23044
rect 26016 23032 26022 23044
rect 27172 23032 27200 23072
rect 28537 23069 28549 23072
rect 28583 23069 28595 23103
rect 28537 23063 28595 23069
rect 28629 23103 28687 23109
rect 28629 23069 28641 23103
rect 28675 23100 28687 23103
rect 28675 23072 28856 23100
rect 28675 23069 28687 23072
rect 28629 23063 28687 23069
rect 26016 23004 27200 23032
rect 26016 22992 26022 23004
rect 28258 22992 28264 23044
rect 28316 22992 28322 23044
rect 28721 23035 28779 23041
rect 28721 23001 28733 23035
rect 28767 23001 28779 23035
rect 28828 23032 28856 23072
rect 28902 23060 28908 23112
rect 28960 23060 28966 23112
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29549 23103 29607 23109
rect 29549 23100 29561 23103
rect 29052 23072 29561 23100
rect 29052 23060 29058 23072
rect 29549 23069 29561 23072
rect 29595 23100 29607 23103
rect 30098 23100 30104 23112
rect 29595 23072 30104 23100
rect 29595 23069 29607 23072
rect 29549 23063 29607 23069
rect 30098 23060 30104 23072
rect 30156 23060 30162 23112
rect 29178 23032 29184 23044
rect 28828 23004 29184 23032
rect 28721 22995 28779 23001
rect 14884 22936 16160 22964
rect 14884 22924 14890 22936
rect 17678 22924 17684 22976
rect 17736 22964 17742 22976
rect 19245 22967 19303 22973
rect 19245 22964 19257 22967
rect 17736 22936 19257 22964
rect 17736 22924 17742 22936
rect 19245 22933 19257 22936
rect 19291 22933 19303 22967
rect 19245 22927 19303 22933
rect 21821 22967 21879 22973
rect 21821 22933 21833 22967
rect 21867 22964 21879 22967
rect 22830 22964 22836 22976
rect 21867 22936 22836 22964
rect 21867 22933 21879 22936
rect 21821 22927 21879 22933
rect 22830 22924 22836 22936
rect 22888 22924 22894 22976
rect 25774 22924 25780 22976
rect 25832 22924 25838 22976
rect 25866 22924 25872 22976
rect 25924 22924 25930 22976
rect 28736 22964 28764 22995
rect 29178 22992 29184 23004
rect 29236 22992 29242 23044
rect 29816 23035 29874 23041
rect 29816 23001 29828 23035
rect 29862 23032 29874 23035
rect 30006 23032 30012 23044
rect 29862 23004 30012 23032
rect 29862 23001 29874 23004
rect 29816 22995 29874 23001
rect 30006 22992 30012 23004
rect 30064 22992 30070 23044
rect 30576 23032 30604 23276
rect 30926 23264 30932 23316
rect 30984 23264 30990 23316
rect 32030 23304 32036 23316
rect 31036 23276 32036 23304
rect 31036 23109 31064 23276
rect 32030 23264 32036 23276
rect 32088 23264 32094 23316
rect 34790 23304 34796 23316
rect 33152 23276 34796 23304
rect 31662 23128 31668 23180
rect 31720 23128 31726 23180
rect 33152 23177 33180 23276
rect 34790 23264 34796 23276
rect 34848 23264 34854 23316
rect 36078 23264 36084 23316
rect 36136 23304 36142 23316
rect 36446 23304 36452 23316
rect 36136 23276 36452 23304
rect 36136 23264 36142 23276
rect 36446 23264 36452 23276
rect 36504 23304 36510 23316
rect 37185 23307 37243 23313
rect 37185 23304 37197 23307
rect 36504 23276 37197 23304
rect 36504 23264 36510 23276
rect 37185 23273 37197 23276
rect 37231 23273 37243 23307
rect 38286 23304 38292 23316
rect 37185 23267 37243 23273
rect 37660 23276 38292 23304
rect 33137 23171 33195 23177
rect 33137 23137 33149 23171
rect 33183 23137 33195 23171
rect 34808 23168 34836 23264
rect 37660 23177 37688 23276
rect 38286 23264 38292 23276
rect 38344 23264 38350 23316
rect 39666 23264 39672 23316
rect 39724 23304 39730 23316
rect 39853 23307 39911 23313
rect 39853 23304 39865 23307
rect 39724 23276 39865 23304
rect 39724 23264 39730 23276
rect 39853 23273 39865 23276
rect 39899 23273 39911 23307
rect 39853 23267 39911 23273
rect 41414 23264 41420 23316
rect 41472 23304 41478 23316
rect 41509 23307 41567 23313
rect 41509 23304 41521 23307
rect 41472 23276 41521 23304
rect 41472 23264 41478 23276
rect 41509 23273 41521 23276
rect 41555 23273 41567 23307
rect 41509 23267 41567 23273
rect 35437 23171 35495 23177
rect 35437 23168 35449 23171
rect 34808 23140 35449 23168
rect 33137 23131 33195 23137
rect 35437 23137 35449 23140
rect 35483 23137 35495 23171
rect 35437 23131 35495 23137
rect 37645 23171 37703 23177
rect 37645 23137 37657 23171
rect 37691 23137 37703 23171
rect 37645 23131 37703 23137
rect 38654 23128 38660 23180
rect 38712 23168 38718 23180
rect 40405 23171 40463 23177
rect 40405 23168 40417 23171
rect 38712 23140 40417 23168
rect 38712 23128 38718 23140
rect 40405 23137 40417 23140
rect 40451 23137 40463 23171
rect 40405 23131 40463 23137
rect 40770 23128 40776 23180
rect 40828 23128 40834 23180
rect 42058 23128 42064 23180
rect 42116 23128 42122 23180
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23069 31079 23103
rect 31389 23103 31447 23109
rect 31389 23100 31401 23103
rect 31021 23063 31079 23069
rect 31128 23072 31401 23100
rect 31128 23032 31156 23072
rect 31389 23069 31401 23072
rect 31435 23100 31447 23103
rect 32490 23100 32496 23112
rect 31435 23072 32496 23100
rect 31435 23069 31447 23072
rect 31389 23063 31447 23069
rect 32490 23060 32496 23072
rect 32548 23060 32554 23112
rect 33404 23103 33462 23109
rect 33404 23069 33416 23103
rect 33450 23069 33462 23103
rect 33404 23063 33462 23069
rect 34701 23103 34759 23109
rect 34701 23069 34713 23103
rect 34747 23100 34759 23103
rect 34882 23100 34888 23112
rect 34747 23072 34888 23100
rect 34747 23069 34759 23072
rect 34701 23063 34759 23069
rect 30576 23004 31156 23032
rect 31202 22992 31208 23044
rect 31260 22992 31266 23044
rect 31297 23035 31355 23041
rect 31297 23001 31309 23035
rect 31343 23032 31355 23035
rect 31910 23035 31968 23041
rect 31910 23032 31922 23035
rect 31343 23004 31432 23032
rect 31343 23001 31355 23004
rect 31297 22995 31355 23001
rect 28810 22964 28816 22976
rect 28736 22936 28816 22964
rect 28810 22924 28816 22936
rect 28868 22964 28874 22976
rect 31220 22964 31248 22992
rect 31404 22976 31432 23004
rect 31726 23004 31922 23032
rect 28868 22936 31248 22964
rect 28868 22924 28874 22936
rect 31386 22924 31392 22976
rect 31444 22924 31450 22976
rect 31573 22967 31631 22973
rect 31573 22933 31585 22967
rect 31619 22964 31631 22967
rect 31726 22964 31754 23004
rect 31910 23001 31922 23004
rect 31956 23001 31968 23035
rect 31910 22995 31968 23001
rect 33318 22992 33324 23044
rect 33376 23032 33382 23044
rect 33428 23032 33456 23063
rect 34882 23060 34888 23072
rect 34940 23060 34946 23112
rect 37918 23109 37924 23112
rect 37912 23100 37924 23109
rect 37879 23072 37924 23100
rect 37912 23063 37924 23072
rect 37918 23060 37924 23063
rect 37976 23060 37982 23112
rect 40034 23060 40040 23112
rect 40092 23100 40098 23112
rect 40221 23103 40279 23109
rect 40221 23100 40233 23103
rect 40092 23072 40233 23100
rect 40092 23060 40098 23072
rect 40221 23069 40233 23072
rect 40267 23069 40279 23103
rect 40221 23063 40279 23069
rect 33376 23004 33456 23032
rect 33376 22992 33382 23004
rect 35434 22992 35440 23044
rect 35492 23032 35498 23044
rect 35713 23035 35771 23041
rect 35713 23032 35725 23035
rect 35492 23004 35725 23032
rect 35492 22992 35498 23004
rect 35713 23001 35725 23004
rect 35759 23001 35771 23035
rect 36998 23032 37004 23044
rect 36938 23004 37004 23032
rect 35713 22995 35771 23001
rect 36998 22992 37004 23004
rect 37056 23032 37062 23044
rect 41966 23032 41972 23044
rect 37056 23004 41972 23032
rect 37056 22992 37062 23004
rect 41966 22992 41972 23004
rect 42024 22992 42030 23044
rect 31619 22936 31754 22964
rect 31619 22933 31631 22936
rect 31573 22927 31631 22933
rect 32766 22924 32772 22976
rect 32824 22964 32830 22976
rect 33045 22967 33103 22973
rect 33045 22964 33057 22967
rect 32824 22936 33057 22964
rect 32824 22924 32830 22936
rect 33045 22933 33057 22936
rect 33091 22933 33103 22967
rect 33045 22927 33103 22933
rect 34514 22924 34520 22976
rect 34572 22924 34578 22976
rect 35342 22924 35348 22976
rect 35400 22924 35406 22976
rect 39022 22924 39028 22976
rect 39080 22924 39086 22976
rect 40313 22967 40371 22973
rect 40313 22933 40325 22967
rect 40359 22964 40371 22967
rect 41046 22964 41052 22976
rect 40359 22936 41052 22964
rect 40359 22933 40371 22936
rect 40313 22927 40371 22933
rect 41046 22924 41052 22936
rect 41104 22964 41110 22976
rect 41417 22967 41475 22973
rect 41417 22964 41429 22967
rect 41104 22936 41429 22964
rect 41104 22924 41110 22936
rect 41417 22933 41429 22936
rect 41463 22933 41475 22967
rect 41417 22927 41475 22933
rect 1104 22874 42504 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 42504 22874
rect 1104 22800 42504 22822
rect 1394 22720 1400 22772
rect 1452 22720 1458 22772
rect 5169 22763 5227 22769
rect 5169 22729 5181 22763
rect 5215 22760 5227 22763
rect 5258 22760 5264 22772
rect 5215 22732 5264 22760
rect 5215 22729 5227 22732
rect 5169 22723 5227 22729
rect 5258 22720 5264 22732
rect 5316 22720 5322 22772
rect 6914 22720 6920 22772
rect 6972 22760 6978 22772
rect 7374 22760 7380 22772
rect 6972 22732 7380 22760
rect 6972 22720 6978 22732
rect 7374 22720 7380 22732
rect 7432 22720 7438 22772
rect 8478 22720 8484 22772
rect 8536 22760 8542 22772
rect 9122 22760 9128 22772
rect 8536 22732 9128 22760
rect 8536 22720 8542 22732
rect 9122 22720 9128 22732
rect 9180 22760 9186 22772
rect 9677 22763 9735 22769
rect 9180 22732 9444 22760
rect 9180 22720 9186 22732
rect 2869 22695 2927 22701
rect 2869 22661 2881 22695
rect 2915 22692 2927 22695
rect 3142 22692 3148 22704
rect 2915 22664 3148 22692
rect 2915 22661 2927 22664
rect 2869 22655 2927 22661
rect 3142 22652 3148 22664
rect 3200 22652 3206 22704
rect 3970 22652 3976 22704
rect 4028 22692 4034 22704
rect 5902 22692 5908 22704
rect 4028 22664 4844 22692
rect 4028 22652 4034 22664
rect 1762 22584 1768 22636
rect 1820 22584 1826 22636
rect 4525 22627 4583 22633
rect 4525 22593 4537 22627
rect 4571 22624 4583 22627
rect 4614 22624 4620 22636
rect 4571 22596 4620 22624
rect 4571 22593 4583 22596
rect 4525 22587 4583 22593
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 4706 22584 4712 22636
rect 4764 22584 4770 22636
rect 4816 22633 4844 22664
rect 4908 22664 5908 22692
rect 4908 22633 4936 22664
rect 5902 22652 5908 22664
rect 5960 22652 5966 22704
rect 6733 22695 6791 22701
rect 6733 22661 6745 22695
rect 6779 22692 6791 22695
rect 8386 22692 8392 22704
rect 6779 22664 8392 22692
rect 6779 22661 6791 22664
rect 6733 22655 6791 22661
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22593 4859 22627
rect 4801 22587 4859 22593
rect 4893 22627 4951 22633
rect 4893 22593 4905 22627
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 5261 22627 5319 22633
rect 5261 22593 5273 22627
rect 5307 22624 5319 22627
rect 5534 22624 5540 22636
rect 5307 22596 5540 22624
rect 5307 22593 5319 22596
rect 5261 22587 5319 22593
rect 3142 22516 3148 22568
rect 3200 22516 3206 22568
rect 4816 22488 4844 22587
rect 5534 22584 5540 22596
rect 5592 22624 5598 22636
rect 5718 22624 5724 22636
rect 5592 22596 5724 22624
rect 5592 22584 5598 22596
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 6825 22627 6883 22633
rect 6825 22593 6837 22627
rect 6871 22624 6883 22627
rect 6917 22627 6975 22633
rect 6917 22624 6929 22627
rect 6871 22596 6929 22624
rect 6871 22593 6883 22596
rect 6825 22587 6883 22593
rect 6917 22593 6929 22596
rect 6963 22593 6975 22627
rect 6917 22587 6975 22593
rect 7101 22627 7159 22633
rect 7101 22593 7113 22627
rect 7147 22624 7159 22627
rect 7282 22624 7288 22636
rect 7147 22596 7288 22624
rect 7147 22593 7159 22596
rect 7101 22587 7159 22593
rect 5166 22516 5172 22568
rect 5224 22516 5230 22568
rect 6656 22556 6684 22587
rect 7282 22584 7288 22596
rect 7340 22584 7346 22636
rect 7374 22584 7380 22636
rect 7432 22584 7438 22636
rect 7466 22584 7472 22636
rect 7524 22624 7530 22636
rect 8312 22633 8340 22664
rect 8386 22652 8392 22664
rect 8444 22652 8450 22704
rect 9306 22652 9312 22704
rect 9364 22652 9370 22704
rect 9416 22701 9444 22732
rect 9677 22729 9689 22763
rect 9723 22729 9735 22763
rect 9677 22723 9735 22729
rect 9401 22695 9459 22701
rect 9401 22661 9413 22695
rect 9447 22661 9459 22695
rect 9692 22692 9720 22723
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 9824 22732 11560 22760
rect 9824 22720 9830 22732
rect 10014 22695 10072 22701
rect 10014 22692 10026 22695
rect 9692 22664 10026 22692
rect 9401 22655 9459 22661
rect 10014 22661 10026 22664
rect 10060 22661 10072 22695
rect 10014 22655 10072 22661
rect 11532 22636 11560 22732
rect 13262 22720 13268 22772
rect 13320 22720 13326 22772
rect 18233 22763 18291 22769
rect 18233 22729 18245 22763
rect 18279 22760 18291 22763
rect 18279 22732 18460 22760
rect 18279 22729 18291 22732
rect 18233 22723 18291 22729
rect 11793 22695 11851 22701
rect 11793 22661 11805 22695
rect 11839 22692 11851 22695
rect 11882 22692 11888 22704
rect 11839 22664 11888 22692
rect 11839 22661 11851 22664
rect 11793 22655 11851 22661
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 16666 22652 16672 22704
rect 16724 22692 16730 22704
rect 17494 22692 17500 22704
rect 16724 22664 17500 22692
rect 16724 22652 16730 22664
rect 17494 22652 17500 22664
rect 17552 22692 17558 22704
rect 17865 22695 17923 22701
rect 17865 22692 17877 22695
rect 17552 22664 17877 22692
rect 17552 22652 17558 22664
rect 17865 22661 17877 22664
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 17957 22695 18015 22701
rect 17957 22661 17969 22695
rect 18003 22692 18015 22695
rect 18138 22692 18144 22704
rect 18003 22664 18144 22692
rect 18003 22661 18015 22664
rect 17957 22655 18015 22661
rect 18138 22652 18144 22664
rect 18196 22652 18202 22704
rect 7837 22627 7895 22633
rect 7837 22624 7849 22627
rect 7524 22596 7849 22624
rect 7524 22584 7530 22596
rect 7837 22593 7849 22596
rect 7883 22593 7895 22627
rect 7837 22587 7895 22593
rect 8297 22627 8355 22633
rect 8297 22593 8309 22627
rect 8343 22593 8355 22627
rect 8297 22587 8355 22593
rect 8481 22627 8539 22633
rect 8481 22593 8493 22627
rect 8527 22593 8539 22627
rect 8481 22587 8539 22593
rect 8573 22627 8631 22633
rect 8573 22593 8585 22627
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 7006 22556 7012 22568
rect 6656 22528 7012 22556
rect 6656 22488 6684 22528
rect 7006 22516 7012 22528
rect 7064 22516 7070 22568
rect 4816 22460 6684 22488
rect 7300 22488 7328 22584
rect 7561 22559 7619 22565
rect 7561 22525 7573 22559
rect 7607 22525 7619 22559
rect 7561 22519 7619 22525
rect 7576 22488 7604 22519
rect 7650 22516 7656 22568
rect 7708 22516 7714 22568
rect 7742 22516 7748 22568
rect 7800 22516 7806 22568
rect 8021 22559 8079 22565
rect 8021 22525 8033 22559
rect 8067 22556 8079 22559
rect 8496 22556 8524 22587
rect 8067 22528 8524 22556
rect 8067 22525 8079 22528
rect 8021 22519 8079 22525
rect 7926 22488 7932 22500
rect 7300 22460 7932 22488
rect 7926 22448 7932 22460
rect 7984 22448 7990 22500
rect 4525 22423 4583 22429
rect 4525 22389 4537 22423
rect 4571 22420 4583 22423
rect 4798 22420 4804 22432
rect 4571 22392 4804 22420
rect 4571 22389 4583 22392
rect 4525 22383 4583 22389
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 4982 22380 4988 22432
rect 5040 22380 5046 22432
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 5350 22420 5356 22432
rect 5132 22392 5356 22420
rect 5132 22380 5138 22392
rect 5350 22380 5356 22392
rect 5408 22380 5414 22432
rect 7006 22380 7012 22432
rect 7064 22420 7070 22432
rect 7190 22420 7196 22432
rect 7064 22392 7196 22420
rect 7064 22380 7070 22392
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 7285 22423 7343 22429
rect 7285 22389 7297 22423
rect 7331 22420 7343 22423
rect 7742 22420 7748 22432
rect 7331 22392 7748 22420
rect 7331 22389 7343 22392
rect 7285 22383 7343 22389
rect 7742 22380 7748 22392
rect 7800 22380 7806 22432
rect 8588 22420 8616 22587
rect 8662 22584 8668 22636
rect 8720 22584 8726 22636
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 8864 22596 9137 22624
rect 8864 22497 8892 22596
rect 9125 22593 9137 22596
rect 9171 22593 9183 22627
rect 9125 22587 9183 22593
rect 9493 22627 9551 22633
rect 9493 22593 9505 22627
rect 9539 22624 9551 22627
rect 11422 22624 11428 22636
rect 9539 22596 11428 22624
rect 9539 22593 9551 22596
rect 9493 22587 9551 22593
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 11514 22584 11520 22636
rect 11572 22584 11578 22636
rect 12894 22584 12900 22636
rect 12952 22584 12958 22636
rect 14734 22584 14740 22636
rect 14792 22584 14798 22636
rect 17313 22627 17371 22633
rect 17313 22593 17325 22627
rect 17359 22624 17371 22627
rect 17402 22624 17408 22636
rect 17359 22596 17408 22624
rect 17359 22593 17371 22596
rect 17313 22587 17371 22593
rect 17402 22584 17408 22596
rect 17460 22584 17466 22636
rect 17678 22584 17684 22636
rect 17736 22584 17742 22636
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22624 18107 22627
rect 18230 22624 18236 22636
rect 18095 22596 18236 22624
rect 18095 22593 18107 22596
rect 18049 22587 18107 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18432 22624 18460 22732
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19668 22732 19717 22760
rect 19668 22720 19674 22732
rect 19705 22729 19717 22732
rect 19751 22760 19763 22763
rect 19794 22760 19800 22772
rect 19751 22732 19800 22760
rect 19751 22729 19763 22732
rect 19705 22723 19763 22729
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 20772 22732 21189 22760
rect 20772 22720 20778 22732
rect 21177 22729 21189 22732
rect 21223 22760 21235 22763
rect 21358 22760 21364 22772
rect 21223 22732 21364 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 21358 22720 21364 22732
rect 21416 22720 21422 22772
rect 32030 22720 32036 22772
rect 32088 22760 32094 22772
rect 32125 22763 32183 22769
rect 32125 22760 32137 22763
rect 32088 22732 32137 22760
rect 32088 22720 32094 22732
rect 32125 22729 32137 22732
rect 32171 22729 32183 22763
rect 32125 22723 32183 22729
rect 33413 22763 33471 22769
rect 33413 22729 33425 22763
rect 33459 22760 33471 22763
rect 34882 22760 34888 22772
rect 33459 22732 34888 22760
rect 33459 22729 33471 22732
rect 33413 22723 33471 22729
rect 34882 22720 34888 22732
rect 34940 22760 34946 22772
rect 35434 22760 35440 22772
rect 34940 22732 35440 22760
rect 34940 22720 34946 22732
rect 35434 22720 35440 22732
rect 35492 22720 35498 22772
rect 41046 22720 41052 22772
rect 41104 22720 41110 22772
rect 41877 22763 41935 22769
rect 41877 22729 41889 22763
rect 41923 22760 41935 22763
rect 41966 22760 41972 22772
rect 41923 22732 41972 22760
rect 41923 22729 41935 22732
rect 41877 22723 41935 22729
rect 41966 22720 41972 22732
rect 42024 22720 42030 22772
rect 23293 22695 23351 22701
rect 23293 22661 23305 22695
rect 23339 22692 23351 22695
rect 23661 22695 23719 22701
rect 23661 22692 23673 22695
rect 23339 22664 23673 22692
rect 23339 22661 23351 22664
rect 23293 22655 23351 22661
rect 23661 22661 23673 22664
rect 23707 22661 23719 22695
rect 23661 22655 23719 22661
rect 25992 22695 26050 22701
rect 25992 22661 26004 22695
rect 26038 22692 26050 22695
rect 26326 22692 26332 22704
rect 26038 22664 26332 22692
rect 26038 22661 26050 22664
rect 25992 22655 26050 22661
rect 26326 22652 26332 22664
rect 26384 22652 26390 22704
rect 27430 22692 27436 22704
rect 26988 22664 27436 22692
rect 20070 22633 20076 22636
rect 18581 22627 18639 22633
rect 18581 22624 18593 22627
rect 18432 22596 18593 22624
rect 18581 22593 18593 22596
rect 18627 22593 18639 22627
rect 20064 22624 20076 22633
rect 20031 22596 20076 22624
rect 18581 22587 18639 22593
rect 20064 22587 20076 22596
rect 20070 22584 20076 22587
rect 20128 22584 20134 22636
rect 26237 22627 26295 22633
rect 22112 22596 22218 22624
rect 22112 22568 22140 22596
rect 26237 22593 26249 22627
rect 26283 22624 26295 22627
rect 26418 22624 26424 22636
rect 26283 22596 26424 22624
rect 26283 22593 26295 22596
rect 26237 22587 26295 22593
rect 26418 22584 26424 22596
rect 26476 22624 26482 22636
rect 26988 22633 27016 22664
rect 27430 22652 27436 22664
rect 27488 22652 27494 22704
rect 30834 22692 30840 22704
rect 29946 22664 30840 22692
rect 30834 22652 30840 22664
rect 30892 22652 30898 22704
rect 34548 22695 34606 22701
rect 34548 22661 34560 22695
rect 34594 22692 34606 22695
rect 34698 22692 34704 22704
rect 34594 22664 34704 22692
rect 34594 22661 34606 22664
rect 34548 22655 34606 22661
rect 34698 22652 34704 22664
rect 34756 22652 34762 22704
rect 35526 22692 35532 22704
rect 34808 22664 35532 22692
rect 27246 22633 27252 22636
rect 26973 22627 27031 22633
rect 26973 22624 26985 22627
rect 26476 22596 26985 22624
rect 26476 22584 26482 22596
rect 26973 22593 26985 22596
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 27240 22587 27252 22633
rect 27246 22584 27252 22587
rect 27304 22584 27310 22636
rect 30552 22627 30610 22633
rect 30552 22593 30564 22627
rect 30598 22624 30610 22627
rect 30926 22624 30932 22636
rect 30598 22596 30932 22624
rect 30598 22593 30610 22596
rect 30552 22587 30610 22593
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 34808 22633 34836 22664
rect 35526 22652 35532 22664
rect 35584 22692 35590 22704
rect 39850 22692 39856 22704
rect 35584 22664 36308 22692
rect 35584 22652 35590 22664
rect 36280 22633 36308 22664
rect 37292 22664 39856 22692
rect 37292 22636 37320 22664
rect 34793 22627 34851 22633
rect 34793 22593 34805 22627
rect 34839 22593 34851 22627
rect 34793 22587 34851 22593
rect 36009 22627 36067 22633
rect 36009 22593 36021 22627
rect 36055 22624 36067 22627
rect 36265 22627 36323 22633
rect 36055 22596 36216 22624
rect 36055 22593 36067 22596
rect 36009 22587 36067 22593
rect 9766 22516 9772 22568
rect 9824 22516 9830 22568
rect 14826 22516 14832 22568
rect 14884 22516 14890 22568
rect 17586 22516 17592 22568
rect 17644 22556 17650 22568
rect 18325 22559 18383 22565
rect 18325 22556 18337 22559
rect 17644 22528 18337 22556
rect 17644 22516 17650 22528
rect 18325 22525 18337 22528
rect 18371 22525 18383 22559
rect 18325 22519 18383 22525
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22525 19855 22559
rect 19797 22519 19855 22525
rect 8849 22491 8907 22497
rect 8849 22457 8861 22491
rect 8895 22457 8907 22491
rect 8849 22451 8907 22457
rect 11146 22420 11152 22432
rect 8588 22392 11152 22420
rect 11146 22380 11152 22392
rect 11204 22380 11210 22432
rect 15102 22380 15108 22432
rect 15160 22380 15166 22432
rect 16666 22380 16672 22432
rect 16724 22380 16730 22432
rect 18340 22420 18368 22519
rect 19812 22432 19840 22519
rect 22094 22516 22100 22568
rect 22152 22516 22158 22568
rect 23569 22559 23627 22565
rect 23569 22525 23581 22559
rect 23615 22525 23627 22559
rect 23569 22519 23627 22525
rect 19794 22420 19800 22432
rect 18340 22392 19800 22420
rect 19794 22380 19800 22392
rect 19852 22380 19858 22432
rect 21821 22423 21879 22429
rect 21821 22389 21833 22423
rect 21867 22420 21879 22423
rect 22554 22420 22560 22432
rect 21867 22392 22560 22420
rect 21867 22389 21879 22392
rect 21821 22383 21879 22389
rect 22554 22380 22560 22392
rect 22612 22380 22618 22432
rect 22922 22380 22928 22432
rect 22980 22420 22986 22432
rect 23584 22420 23612 22519
rect 24210 22516 24216 22568
rect 24268 22516 24274 22568
rect 26510 22516 26516 22568
rect 26568 22556 26574 22568
rect 26786 22556 26792 22568
rect 26568 22528 26792 22556
rect 26568 22516 26574 22528
rect 26786 22516 26792 22528
rect 26844 22516 26850 22568
rect 28445 22559 28503 22565
rect 28445 22525 28457 22559
rect 28491 22556 28503 22559
rect 28721 22559 28779 22565
rect 28491 22528 28580 22556
rect 28491 22525 28503 22528
rect 28445 22519 28503 22525
rect 22980 22392 23612 22420
rect 24857 22423 24915 22429
rect 22980 22380 22986 22392
rect 24857 22389 24869 22423
rect 24903 22420 24915 22423
rect 25958 22420 25964 22432
rect 24903 22392 25964 22420
rect 24903 22389 24915 22392
rect 24857 22383 24915 22389
rect 25958 22380 25964 22392
rect 26016 22380 26022 22432
rect 28350 22380 28356 22432
rect 28408 22380 28414 22432
rect 28552 22420 28580 22528
rect 28721 22525 28733 22559
rect 28767 22556 28779 22559
rect 29454 22556 29460 22568
rect 28767 22528 29460 22556
rect 28767 22525 28779 22528
rect 28721 22519 28779 22525
rect 29454 22516 29460 22528
rect 29512 22516 29518 22568
rect 30098 22516 30104 22568
rect 30156 22556 30162 22568
rect 30285 22559 30343 22565
rect 30285 22556 30297 22559
rect 30156 22528 30297 22556
rect 30156 22516 30162 22528
rect 30285 22525 30297 22528
rect 30331 22525 30343 22559
rect 30285 22519 30343 22525
rect 32766 22516 32772 22568
rect 32824 22516 32830 22568
rect 36188 22556 36216 22596
rect 36265 22593 36277 22627
rect 36311 22624 36323 22627
rect 37274 22624 37280 22636
rect 36311 22596 37280 22624
rect 36311 22593 36323 22596
rect 36265 22587 36323 22593
rect 37274 22584 37280 22596
rect 37332 22584 37338 22636
rect 37550 22633 37556 22636
rect 37544 22587 37556 22633
rect 37550 22584 37556 22587
rect 37608 22584 37614 22636
rect 39316 22633 39344 22664
rect 39850 22652 39856 22664
rect 39908 22652 39914 22704
rect 41598 22652 41604 22704
rect 41656 22692 41662 22704
rect 41785 22695 41843 22701
rect 41785 22692 41797 22695
rect 41656 22664 41797 22692
rect 41656 22652 41662 22664
rect 41785 22661 41797 22664
rect 41831 22661 41843 22695
rect 41785 22655 41843 22661
rect 39574 22633 39580 22636
rect 39301 22627 39359 22633
rect 39301 22593 39313 22627
rect 39347 22593 39359 22627
rect 39301 22587 39359 22593
rect 39568 22587 39580 22633
rect 39574 22584 39580 22587
rect 39632 22584 39638 22636
rect 41141 22627 41199 22633
rect 41141 22593 41153 22627
rect 41187 22624 41199 22627
rect 41690 22624 41696 22636
rect 41187 22596 41696 22624
rect 41187 22593 41199 22596
rect 41141 22587 41199 22593
rect 41690 22584 41696 22596
rect 41748 22584 41754 22636
rect 36357 22559 36415 22565
rect 36357 22556 36369 22559
rect 36188 22528 36369 22556
rect 36357 22525 36369 22528
rect 36403 22525 36415 22559
rect 36357 22519 36415 22525
rect 36906 22516 36912 22568
rect 36964 22516 36970 22568
rect 40770 22516 40776 22568
rect 40828 22556 40834 22568
rect 40865 22559 40923 22565
rect 40865 22556 40877 22559
rect 40828 22528 40877 22556
rect 40828 22516 40834 22528
rect 40865 22525 40877 22528
rect 40911 22525 40923 22559
rect 40865 22519 40923 22525
rect 30098 22420 30104 22432
rect 28552 22392 30104 22420
rect 30098 22380 30104 22392
rect 30156 22380 30162 22432
rect 30193 22423 30251 22429
rect 30193 22389 30205 22423
rect 30239 22420 30251 22423
rect 30650 22420 30656 22432
rect 30239 22392 30656 22420
rect 30239 22389 30251 22392
rect 30193 22383 30251 22389
rect 30650 22380 30656 22392
rect 30708 22380 30714 22432
rect 31665 22423 31723 22429
rect 31665 22389 31677 22423
rect 31711 22420 31723 22423
rect 32030 22420 32036 22432
rect 31711 22392 32036 22420
rect 31711 22389 31723 22392
rect 31665 22383 31723 22389
rect 32030 22380 32036 22392
rect 32088 22380 32094 22432
rect 34790 22380 34796 22432
rect 34848 22420 34854 22432
rect 34885 22423 34943 22429
rect 34885 22420 34897 22423
rect 34848 22392 34897 22420
rect 34848 22380 34854 22392
rect 34885 22389 34897 22392
rect 34931 22389 34943 22423
rect 34885 22383 34943 22389
rect 38654 22380 38660 22432
rect 38712 22380 38718 22432
rect 40678 22380 40684 22432
rect 40736 22380 40742 22432
rect 41506 22380 41512 22432
rect 41564 22380 41570 22432
rect 1104 22330 42504 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 42504 22330
rect 1104 22256 42504 22278
rect 2887 22219 2945 22225
rect 2887 22185 2899 22219
rect 2933 22216 2945 22219
rect 3050 22216 3056 22228
rect 2933 22188 3056 22216
rect 2933 22185 2945 22188
rect 2887 22179 2945 22185
rect 3050 22176 3056 22188
rect 3108 22176 3114 22228
rect 4706 22176 4712 22228
rect 4764 22216 4770 22228
rect 4764 22188 5304 22216
rect 4764 22176 4770 22188
rect 5276 22148 5304 22188
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 9306 22216 9312 22228
rect 5408 22188 7236 22216
rect 5408 22176 5414 22188
rect 5721 22151 5779 22157
rect 5721 22148 5733 22151
rect 5276 22120 5733 22148
rect 5721 22117 5733 22120
rect 5767 22148 5779 22151
rect 7006 22148 7012 22160
rect 5767 22120 7012 22148
rect 5767 22117 5779 22120
rect 5721 22111 5779 22117
rect 7006 22108 7012 22120
rect 7064 22108 7070 22160
rect 4338 22040 4344 22092
rect 4396 22080 4402 22092
rect 4614 22080 4620 22092
rect 4396 22052 4620 22080
rect 4396 22040 4402 22052
rect 4614 22040 4620 22052
rect 4672 22040 4678 22092
rect 7098 22040 7104 22092
rect 7156 22040 7162 22092
rect 7208 22080 7236 22188
rect 8496 22188 9312 22216
rect 7282 22080 7288 22092
rect 7208 22052 7288 22080
rect 7282 22040 7288 22052
rect 7340 22040 7346 22092
rect 8018 22040 8024 22092
rect 8076 22040 8082 22092
rect 1762 21972 1768 22024
rect 1820 21972 1826 22024
rect 3142 21972 3148 22024
rect 3200 22012 3206 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3200 21984 3985 22012
rect 3200 21972 3206 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 6822 21972 6828 22024
rect 6880 21972 6886 22024
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 7190 22012 7196 22024
rect 7064 21984 7196 22012
rect 7064 21972 7070 21984
rect 7190 21972 7196 21984
rect 7248 21972 7254 22024
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 7300 21984 7389 22012
rect 4246 21904 4252 21956
rect 4304 21904 4310 21956
rect 6917 21947 6975 21953
rect 4356 21916 4738 21944
rect 1394 21836 1400 21888
rect 1452 21836 1458 21888
rect 3694 21836 3700 21888
rect 3752 21876 3758 21888
rect 4356 21876 4384 21916
rect 6917 21913 6929 21947
rect 6963 21944 6975 21947
rect 7300 21944 7328 21984
rect 7377 21981 7389 21984
rect 7423 22012 7435 22015
rect 7466 22012 7472 22024
rect 7423 21984 7472 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 7745 22015 7803 22021
rect 7745 21981 7757 22015
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 7760 21944 7788 21975
rect 7834 21972 7840 22024
rect 7892 21972 7898 22024
rect 8110 21972 8116 22024
rect 8168 21972 8174 22024
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 21981 8263 22015
rect 8205 21975 8263 21981
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 22012 8447 22015
rect 8496 22012 8524 22188
rect 9306 22176 9312 22188
rect 9364 22176 9370 22228
rect 18322 22216 18328 22228
rect 13924 22188 18328 22216
rect 8435 21984 8524 22012
rect 8435 21981 8447 21984
rect 8389 21975 8447 21981
rect 6963 21916 7328 21944
rect 7392 21916 7788 21944
rect 6963 21913 6975 21916
rect 6917 21907 6975 21913
rect 3752 21848 4384 21876
rect 3752 21836 3758 21848
rect 4614 21836 4620 21888
rect 4672 21876 4678 21888
rect 4982 21876 4988 21888
rect 4672 21848 4988 21876
rect 4672 21836 4678 21848
rect 4982 21836 4988 21848
rect 5040 21876 5046 21888
rect 6546 21876 6552 21888
rect 5040 21848 6552 21876
rect 5040 21836 5046 21848
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 7392 21885 7420 21916
rect 7377 21879 7435 21885
rect 7377 21845 7389 21879
rect 7423 21845 7435 21879
rect 7377 21839 7435 21845
rect 7561 21879 7619 21885
rect 7561 21845 7573 21879
rect 7607 21876 7619 21879
rect 8220 21876 8248 21975
rect 8570 21972 8576 22024
rect 8628 21972 8634 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9766 22012 9772 22024
rect 9171 21984 9772 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 11882 21972 11888 22024
rect 11940 21972 11946 22024
rect 13924 21956 13952 22188
rect 18322 22176 18328 22188
rect 18380 22176 18386 22228
rect 20162 22216 20168 22228
rect 18892 22188 20168 22216
rect 15102 22108 15108 22160
rect 15160 22148 15166 22160
rect 15160 22120 15332 22148
rect 15160 22108 15166 22120
rect 15304 22089 15332 22120
rect 17770 22108 17776 22160
rect 17828 22148 17834 22160
rect 18892 22148 18920 22188
rect 20162 22176 20168 22188
rect 20220 22176 20226 22228
rect 27246 22176 27252 22228
rect 27304 22216 27310 22228
rect 27341 22219 27399 22225
rect 27341 22216 27353 22219
rect 27304 22188 27353 22216
rect 27304 22176 27310 22188
rect 27341 22185 27353 22188
rect 27387 22185 27399 22219
rect 27341 22179 27399 22185
rect 29454 22176 29460 22228
rect 29512 22216 29518 22228
rect 29549 22219 29607 22225
rect 29549 22216 29561 22219
rect 29512 22188 29561 22216
rect 29512 22176 29518 22188
rect 29549 22185 29561 22188
rect 29595 22185 29607 22219
rect 29549 22179 29607 22185
rect 30926 22176 30932 22228
rect 30984 22176 30990 22228
rect 34790 22176 34796 22228
rect 34848 22216 34854 22228
rect 35342 22216 35348 22228
rect 34848 22188 35348 22216
rect 34848 22176 34854 22188
rect 35342 22176 35348 22188
rect 35400 22176 35406 22228
rect 37550 22176 37556 22228
rect 37608 22216 37614 22228
rect 37737 22219 37795 22225
rect 37737 22216 37749 22219
rect 37608 22188 37749 22216
rect 37608 22176 37614 22188
rect 37737 22185 37749 22188
rect 37783 22185 37795 22219
rect 37737 22179 37795 22185
rect 24670 22148 24676 22160
rect 17828 22120 18920 22148
rect 17828 22108 17834 22120
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 15335 22052 15369 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 15470 22040 15476 22092
rect 15528 22040 15534 22092
rect 18892 22089 18920 22120
rect 22388 22120 24676 22148
rect 16301 22083 16359 22089
rect 16301 22049 16313 22083
rect 16347 22080 16359 22083
rect 18877 22083 18935 22089
rect 16347 22052 16896 22080
rect 16347 22049 16359 22052
rect 16301 22043 16359 22049
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 22012 16083 22015
rect 16666 22012 16672 22024
rect 16071 21984 16672 22012
rect 16071 21981 16083 21984
rect 16025 21975 16083 21981
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 16758 21972 16764 22024
rect 16816 21972 16822 22024
rect 16868 22012 16896 22052
rect 18877 22049 18889 22083
rect 18923 22080 18935 22083
rect 18923 22052 18957 22080
rect 18923 22049 18935 22052
rect 18877 22043 18935 22049
rect 19794 22040 19800 22092
rect 19852 22040 19858 22092
rect 21910 22040 21916 22092
rect 21968 22040 21974 22092
rect 22388 22089 22416 22120
rect 24670 22108 24676 22120
rect 24728 22108 24734 22160
rect 28810 22148 28816 22160
rect 28000 22120 28816 22148
rect 22373 22083 22431 22089
rect 22373 22049 22385 22083
rect 22419 22080 22431 22083
rect 22419 22052 22453 22080
rect 22419 22049 22431 22052
rect 22373 22043 22431 22049
rect 22830 22040 22836 22092
rect 22888 22080 22894 22092
rect 23569 22083 23627 22089
rect 23569 22080 23581 22083
rect 22888 22052 23581 22080
rect 22888 22040 22894 22052
rect 23569 22049 23581 22052
rect 23615 22049 23627 22083
rect 23569 22043 23627 22049
rect 26326 22040 26332 22092
rect 26384 22080 26390 22092
rect 26421 22083 26479 22089
rect 26421 22080 26433 22083
rect 26384 22052 26433 22080
rect 26384 22040 26390 22052
rect 26421 22049 26433 22052
rect 26467 22049 26479 22083
rect 26421 22043 26479 22049
rect 26970 22040 26976 22092
rect 27028 22040 27034 22092
rect 28000 22089 28028 22120
rect 28810 22108 28816 22120
rect 28868 22108 28874 22160
rect 31202 22108 31208 22160
rect 31260 22148 31266 22160
rect 33134 22148 33140 22160
rect 31260 22120 31616 22148
rect 31260 22108 31266 22120
rect 27985 22083 28043 22089
rect 27985 22049 27997 22083
rect 28031 22080 28043 22083
rect 28031 22052 28065 22080
rect 28031 22049 28043 22052
rect 27985 22043 28043 22049
rect 28350 22040 28356 22092
rect 28408 22080 28414 22092
rect 28721 22083 28779 22089
rect 28721 22080 28733 22083
rect 28408 22052 28733 22080
rect 28408 22040 28414 22052
rect 28721 22049 28733 22052
rect 28767 22049 28779 22083
rect 28721 22043 28779 22049
rect 30006 22040 30012 22092
rect 30064 22040 30070 22092
rect 30193 22083 30251 22089
rect 30193 22049 30205 22083
rect 30239 22080 30251 22083
rect 31386 22080 31392 22092
rect 30239 22052 31392 22080
rect 30239 22049 30251 22052
rect 30193 22043 30251 22049
rect 31386 22040 31392 22052
rect 31444 22040 31450 22092
rect 31588 22089 31616 22120
rect 32968 22120 33140 22148
rect 31573 22083 31631 22089
rect 31573 22049 31585 22083
rect 31619 22080 31631 22083
rect 31619 22052 31754 22080
rect 31619 22049 31631 22052
rect 31573 22043 31631 22049
rect 17494 22012 17500 22024
rect 16868 21984 17500 22012
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 18598 21972 18604 22024
rect 18656 21972 18662 22024
rect 21634 21972 21640 22024
rect 21692 21972 21698 22024
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 23017 22015 23075 22021
rect 23017 22012 23029 22015
rect 22520 21984 23029 22012
rect 22520 21972 22526 21984
rect 23017 21981 23029 21984
rect 23063 21981 23075 22015
rect 23017 21975 23075 21981
rect 25593 22015 25651 22021
rect 25593 21981 25605 22015
rect 25639 22012 25651 22015
rect 25774 22012 25780 22024
rect 25639 21984 25780 22012
rect 25639 21981 25651 21984
rect 25593 21975 25651 21981
rect 25774 21972 25780 21984
rect 25832 22012 25838 22024
rect 25958 22012 25964 22024
rect 25832 21984 25964 22012
rect 25832 21972 25838 21984
rect 25958 21972 25964 21984
rect 26016 21972 26022 22024
rect 26237 22015 26295 22021
rect 26237 21981 26249 22015
rect 26283 21981 26295 22015
rect 26237 21975 26295 21981
rect 8478 21904 8484 21956
rect 8536 21904 8542 21956
rect 9370 21947 9428 21953
rect 9370 21944 9382 21947
rect 8772 21916 9382 21944
rect 8772 21885 8800 21916
rect 9370 21913 9382 21916
rect 9416 21913 9428 21947
rect 9370 21907 9428 21913
rect 12158 21904 12164 21956
rect 12216 21904 12222 21956
rect 12894 21904 12900 21956
rect 12952 21904 12958 21956
rect 13906 21904 13912 21956
rect 13964 21904 13970 21956
rect 15197 21947 15255 21953
rect 15197 21913 15209 21947
rect 15243 21944 15255 21947
rect 17028 21947 17086 21953
rect 15243 21916 16160 21944
rect 15243 21913 15255 21916
rect 15197 21907 15255 21913
rect 7607 21848 8248 21876
rect 8757 21879 8815 21885
rect 7607 21845 7619 21848
rect 7561 21839 7619 21845
rect 8757 21845 8769 21879
rect 8803 21845 8815 21879
rect 8757 21839 8815 21845
rect 10502 21836 10508 21888
rect 10560 21836 10566 21888
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 16132 21885 16160 21916
rect 17028 21913 17040 21947
rect 17074 21944 17086 21947
rect 20064 21947 20122 21953
rect 17074 21916 18276 21944
rect 17074 21913 17086 21916
rect 17028 21907 17086 21913
rect 15657 21879 15715 21885
rect 15657 21876 15669 21879
rect 15344 21848 15669 21876
rect 15344 21836 15350 21848
rect 15657 21845 15669 21848
rect 15703 21845 15715 21879
rect 15657 21839 15715 21845
rect 16117 21879 16175 21885
rect 16117 21845 16129 21879
rect 16163 21876 16175 21879
rect 16574 21876 16580 21888
rect 16163 21848 16580 21876
rect 16163 21845 16175 21848
rect 16117 21839 16175 21845
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 18138 21836 18144 21888
rect 18196 21836 18202 21888
rect 18248 21885 18276 21916
rect 20064 21913 20076 21947
rect 20110 21944 20122 21947
rect 20110 21916 21312 21944
rect 20110 21913 20122 21916
rect 20064 21907 20122 21913
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21845 18291 21879
rect 18233 21839 18291 21845
rect 18690 21836 18696 21888
rect 18748 21836 18754 21888
rect 21174 21836 21180 21888
rect 21232 21836 21238 21888
rect 21284 21885 21312 21916
rect 22554 21904 22560 21956
rect 22612 21904 22618 21956
rect 24302 21904 24308 21956
rect 24360 21944 24366 21956
rect 26252 21944 26280 21975
rect 27706 21972 27712 22024
rect 27764 21972 27770 22024
rect 31294 21972 31300 22024
rect 31352 21972 31358 22024
rect 24360 21916 26280 21944
rect 31726 21944 31754 22052
rect 32030 22040 32036 22092
rect 32088 22080 32094 22092
rect 32309 22083 32367 22089
rect 32309 22080 32321 22083
rect 32088 22052 32321 22080
rect 32088 22040 32094 22052
rect 32309 22049 32321 22052
rect 32355 22049 32367 22083
rect 32309 22043 32367 22049
rect 32968 22021 32996 22120
rect 33134 22108 33140 22120
rect 33192 22108 33198 22160
rect 33229 22083 33287 22089
rect 33229 22049 33241 22083
rect 33275 22080 33287 22083
rect 33870 22080 33876 22092
rect 33275 22052 33876 22080
rect 33275 22049 33287 22052
rect 33229 22043 33287 22049
rect 32953 22015 33011 22021
rect 32953 21981 32965 22015
rect 32999 21981 33011 22015
rect 32953 21975 33011 21981
rect 32306 21944 32312 21956
rect 31726 21916 32312 21944
rect 24360 21904 24366 21916
rect 32306 21904 32312 21916
rect 32364 21944 32370 21956
rect 33244 21944 33272 22043
rect 33870 22040 33876 22052
rect 33928 22040 33934 22092
rect 36004 22052 37136 22080
rect 33502 21972 33508 22024
rect 33560 22012 33566 22024
rect 33965 22015 34023 22021
rect 33965 22012 33977 22015
rect 33560 21984 33977 22012
rect 33560 21972 33566 21984
rect 33965 21981 33977 21984
rect 34011 21981 34023 22015
rect 33965 21975 34023 21981
rect 34977 22015 35035 22021
rect 34977 21981 34989 22015
rect 35023 22012 35035 22015
rect 35526 22012 35532 22024
rect 35023 21984 35532 22012
rect 35023 21981 35035 21984
rect 34977 21975 35035 21981
rect 35526 21972 35532 21984
rect 35584 21972 35590 22024
rect 35250 21953 35256 21956
rect 32364 21916 33272 21944
rect 32364 21904 32370 21916
rect 35244 21907 35256 21953
rect 35250 21904 35256 21907
rect 35308 21904 35314 21956
rect 21269 21879 21327 21885
rect 21269 21845 21281 21879
rect 21315 21845 21327 21879
rect 21269 21839 21327 21845
rect 21726 21836 21732 21888
rect 21784 21836 21790 21888
rect 22925 21879 22983 21885
rect 22925 21845 22937 21879
rect 22971 21876 22983 21879
rect 24210 21876 24216 21888
rect 22971 21848 24216 21876
rect 22971 21845 22983 21848
rect 22925 21839 22983 21845
rect 24210 21836 24216 21848
rect 24268 21836 24274 21888
rect 24946 21836 24952 21888
rect 25004 21836 25010 21888
rect 25682 21836 25688 21888
rect 25740 21836 25746 21888
rect 27801 21879 27859 21885
rect 27801 21845 27813 21879
rect 27847 21876 27859 21879
rect 28166 21876 28172 21888
rect 27847 21848 28172 21876
rect 27847 21845 27859 21848
rect 27801 21839 27859 21845
rect 28166 21836 28172 21848
rect 28224 21836 28230 21888
rect 29914 21836 29920 21888
rect 29972 21836 29978 21888
rect 31294 21836 31300 21888
rect 31352 21876 31358 21888
rect 31389 21879 31447 21885
rect 31389 21876 31401 21879
rect 31352 21848 31401 21876
rect 31352 21836 31358 21848
rect 31389 21845 31401 21848
rect 31435 21876 31447 21879
rect 31757 21879 31815 21885
rect 31757 21876 31769 21879
rect 31435 21848 31769 21876
rect 31435 21845 31447 21848
rect 31389 21839 31447 21845
rect 31757 21845 31769 21848
rect 31803 21845 31815 21879
rect 31757 21839 31815 21845
rect 32582 21836 32588 21888
rect 32640 21836 32646 21888
rect 33045 21879 33103 21885
rect 33045 21845 33057 21879
rect 33091 21876 33103 21879
rect 33226 21876 33232 21888
rect 33091 21848 33232 21876
rect 33091 21845 33103 21848
rect 33045 21839 33103 21845
rect 33226 21836 33232 21848
rect 33284 21876 33290 21888
rect 33413 21879 33471 21885
rect 33413 21876 33425 21879
rect 33284 21848 33425 21876
rect 33284 21836 33290 21848
rect 33413 21845 33425 21848
rect 33459 21845 33471 21879
rect 33413 21839 33471 21845
rect 33594 21836 33600 21888
rect 33652 21876 33658 21888
rect 36004 21876 36032 22052
rect 37001 22015 37059 22021
rect 37001 22012 37013 22015
rect 36372 21984 37013 22012
rect 33652 21848 36032 21876
rect 33652 21836 33658 21848
rect 36078 21836 36084 21888
rect 36136 21876 36142 21888
rect 36372 21885 36400 21984
rect 37001 21981 37013 21984
rect 37047 21981 37059 22015
rect 37001 21975 37059 21981
rect 37108 21944 37136 22052
rect 38286 22040 38292 22092
rect 38344 22080 38350 22092
rect 38562 22080 38568 22092
rect 38344 22052 38568 22080
rect 38344 22040 38350 22052
rect 38562 22040 38568 22052
rect 38620 22040 38626 22092
rect 38654 22040 38660 22092
rect 38712 22080 38718 22092
rect 39117 22083 39175 22089
rect 39117 22080 39129 22083
rect 38712 22052 39129 22080
rect 38712 22040 38718 22052
rect 39117 22049 39129 22052
rect 39163 22049 39175 22083
rect 39117 22043 39175 22049
rect 40497 22083 40555 22089
rect 40497 22049 40509 22083
rect 40543 22080 40555 22083
rect 41138 22080 41144 22092
rect 40543 22052 41144 22080
rect 40543 22049 40555 22052
rect 40497 22043 40555 22049
rect 41138 22040 41144 22052
rect 41196 22040 41202 22092
rect 41690 22040 41696 22092
rect 41748 22080 41754 22092
rect 41874 22080 41880 22092
rect 41748 22052 41880 22080
rect 41748 22040 41754 22052
rect 41874 22040 41880 22052
rect 41932 22080 41938 22092
rect 41969 22083 42027 22089
rect 41969 22080 41981 22083
rect 41932 22052 41981 22080
rect 41932 22040 41938 22052
rect 41969 22049 41981 22052
rect 42015 22049 42027 22083
rect 41969 22043 42027 22049
rect 38010 21972 38016 22024
rect 38068 22012 38074 22024
rect 38105 22015 38163 22021
rect 38105 22012 38117 22015
rect 38068 21984 38117 22012
rect 38068 21972 38074 21984
rect 38105 21981 38117 21984
rect 38151 21981 38163 22015
rect 38105 21975 38163 21981
rect 39850 21972 39856 22024
rect 39908 22012 39914 22024
rect 40218 22012 40224 22024
rect 39908 21984 40224 22012
rect 39908 21972 39914 21984
rect 40218 21972 40224 21984
rect 40276 21972 40282 22024
rect 37108 21916 38700 21944
rect 36357 21879 36415 21885
rect 36357 21876 36369 21879
rect 36136 21848 36369 21876
rect 36136 21836 36142 21848
rect 36357 21845 36369 21848
rect 36403 21845 36415 21879
rect 36357 21839 36415 21845
rect 36446 21836 36452 21888
rect 36504 21836 36510 21888
rect 37642 21836 37648 21888
rect 37700 21876 37706 21888
rect 38197 21879 38255 21885
rect 38197 21876 38209 21879
rect 37700 21848 38209 21876
rect 37700 21836 37706 21848
rect 38197 21845 38209 21848
rect 38243 21876 38255 21879
rect 38565 21879 38623 21885
rect 38565 21876 38577 21879
rect 38243 21848 38577 21876
rect 38243 21845 38255 21848
rect 38197 21839 38255 21845
rect 38565 21845 38577 21848
rect 38611 21845 38623 21879
rect 38672 21876 38700 21916
rect 40586 21904 40592 21956
rect 40644 21944 40650 21956
rect 40644 21916 40986 21944
rect 40644 21904 40650 21916
rect 40770 21876 40776 21888
rect 38672 21848 40776 21876
rect 38565 21839 38623 21845
rect 40770 21836 40776 21848
rect 40828 21836 40834 21888
rect 40880 21876 40908 21916
rect 41414 21876 41420 21888
rect 40880 21848 41420 21876
rect 41414 21836 41420 21848
rect 41472 21836 41478 21888
rect 1104 21786 42504 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 42504 21786
rect 1104 21712 42504 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1360 21644 1593 21672
rect 1360 21632 1366 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 1581 21635 1639 21641
rect 4338 21632 4344 21684
rect 4396 21632 4402 21684
rect 7745 21675 7803 21681
rect 7745 21641 7757 21675
rect 7791 21672 7803 21675
rect 7834 21672 7840 21684
rect 7791 21644 7840 21672
rect 7791 21641 7803 21644
rect 7745 21635 7803 21641
rect 7834 21632 7840 21644
rect 7892 21632 7898 21684
rect 12158 21632 12164 21684
rect 12216 21672 12222 21684
rect 12345 21675 12403 21681
rect 12345 21672 12357 21675
rect 12216 21644 12357 21672
rect 12216 21632 12222 21644
rect 12345 21641 12357 21644
rect 12391 21641 12403 21675
rect 12345 21635 12403 21641
rect 12805 21675 12863 21681
rect 12805 21641 12817 21675
rect 12851 21672 12863 21675
rect 13906 21672 13912 21684
rect 12851 21644 13912 21672
rect 12851 21641 12863 21644
rect 12805 21635 12863 21641
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 14918 21672 14924 21684
rect 14016 21644 14924 21672
rect 3602 21564 3608 21616
rect 3660 21604 3666 21616
rect 4509 21607 4567 21613
rect 4509 21604 4521 21607
rect 3660 21576 4521 21604
rect 3660 21564 3666 21576
rect 4509 21573 4521 21576
rect 4555 21604 4567 21607
rect 4614 21604 4620 21616
rect 4555 21576 4620 21604
rect 4555 21573 4567 21576
rect 4509 21567 4567 21573
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 4709 21607 4767 21613
rect 4709 21573 4721 21607
rect 4755 21573 4767 21607
rect 5994 21604 6000 21616
rect 4709 21567 4767 21573
rect 5000 21576 6000 21604
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1762 21496 1768 21548
rect 1820 21496 1826 21548
rect 3970 21496 3976 21548
rect 4028 21536 4034 21548
rect 4724 21536 4752 21567
rect 5000 21548 5028 21576
rect 5994 21564 6000 21576
rect 6052 21564 6058 21616
rect 8570 21564 8576 21616
rect 8628 21604 8634 21616
rect 9585 21607 9643 21613
rect 9585 21604 9597 21607
rect 8628 21576 9597 21604
rect 8628 21564 8634 21576
rect 9585 21573 9597 21576
rect 9631 21604 9643 21607
rect 12713 21607 12771 21613
rect 12713 21604 12725 21607
rect 9631 21576 12725 21604
rect 9631 21573 9643 21576
rect 9585 21567 9643 21573
rect 12713 21573 12725 21576
rect 12759 21573 12771 21607
rect 12713 21567 12771 21573
rect 12894 21564 12900 21616
rect 12952 21604 12958 21616
rect 14016 21604 14044 21644
rect 14918 21632 14924 21644
rect 14976 21672 14982 21684
rect 16485 21675 16543 21681
rect 14976 21644 15415 21672
rect 14976 21632 14982 21644
rect 12952 21576 14044 21604
rect 14093 21607 14151 21613
rect 12952 21564 12958 21576
rect 14093 21573 14105 21607
rect 14139 21604 14151 21607
rect 14182 21604 14188 21616
rect 14139 21576 14188 21604
rect 14139 21573 14151 21576
rect 14093 21567 14151 21573
rect 14182 21564 14188 21576
rect 14240 21604 14246 21616
rect 14369 21607 14427 21613
rect 14369 21604 14381 21607
rect 14240 21576 14381 21604
rect 14240 21564 14246 21576
rect 14369 21573 14381 21576
rect 14415 21573 14427 21607
rect 14369 21567 14427 21573
rect 15013 21607 15071 21613
rect 15013 21573 15025 21607
rect 15059 21604 15071 21607
rect 15286 21604 15292 21616
rect 15059 21576 15292 21604
rect 15059 21573 15071 21576
rect 15013 21567 15071 21573
rect 15286 21564 15292 21576
rect 15344 21564 15350 21616
rect 15387 21604 15415 21644
rect 16485 21641 16497 21675
rect 16531 21672 16543 21675
rect 17402 21672 17408 21684
rect 16531 21644 17408 21672
rect 16531 21641 16543 21644
rect 16485 21635 16543 21641
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 20162 21632 20168 21684
rect 20220 21672 20226 21684
rect 20220 21644 23152 21672
rect 20220 21632 20226 21644
rect 21450 21604 21456 21616
rect 15387 21576 15502 21604
rect 18630 21576 21456 21604
rect 21450 21564 21456 21576
rect 21508 21564 21514 21616
rect 23124 21604 23152 21644
rect 24302 21632 24308 21684
rect 24360 21632 24366 21684
rect 24397 21675 24455 21681
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24486 21672 24492 21684
rect 24443 21644 24492 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 28166 21632 28172 21684
rect 28224 21632 28230 21684
rect 29914 21632 29920 21684
rect 29972 21672 29978 21684
rect 30101 21675 30159 21681
rect 30101 21672 30113 21675
rect 29972 21644 30113 21672
rect 29972 21632 29978 21644
rect 30101 21641 30113 21644
rect 30147 21641 30159 21675
rect 30101 21635 30159 21641
rect 31294 21632 31300 21684
rect 31352 21632 31358 21684
rect 33502 21632 33508 21684
rect 33560 21632 33566 21684
rect 33870 21632 33876 21684
rect 33928 21672 33934 21684
rect 33928 21644 34100 21672
rect 33928 21632 33934 21644
rect 25038 21604 25044 21616
rect 23124 21576 23612 21604
rect 4028 21508 4752 21536
rect 4028 21496 4034 21508
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 4982 21496 4988 21548
rect 5040 21496 5046 21548
rect 7006 21496 7012 21548
rect 7064 21536 7070 21548
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 7064 21508 7481 21536
rect 7064 21496 7070 21508
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 8110 21496 8116 21548
rect 8168 21536 8174 21548
rect 10137 21539 10195 21545
rect 10137 21536 10149 21539
rect 8168 21508 10149 21536
rect 8168 21496 8174 21508
rect 10137 21505 10149 21508
rect 10183 21536 10195 21539
rect 10502 21536 10508 21548
rect 10183 21508 10508 21536
rect 10183 21505 10195 21508
rect 10137 21499 10195 21505
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 14550 21496 14556 21548
rect 14608 21496 14614 21548
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 21232 21508 22094 21536
rect 21232 21496 21238 21508
rect 6546 21428 6552 21480
rect 6604 21468 6610 21480
rect 7745 21471 7803 21477
rect 7745 21468 7757 21471
rect 6604 21440 7757 21468
rect 6604 21428 6610 21440
rect 7745 21437 7757 21440
rect 7791 21468 7803 21471
rect 8018 21468 8024 21480
rect 7791 21440 8024 21468
rect 7791 21437 7803 21440
rect 7745 21431 7803 21437
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 12986 21428 12992 21480
rect 13044 21428 13050 21480
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 13872 21440 14749 21468
rect 13872 21428 13878 21440
rect 14737 21437 14749 21440
rect 14783 21468 14795 21471
rect 16758 21468 16764 21480
rect 14783 21440 16764 21468
rect 14783 21437 14795 21440
rect 14737 21431 14795 21437
rect 16758 21428 16764 21440
rect 16816 21468 16822 21480
rect 17129 21471 17187 21477
rect 17129 21468 17141 21471
rect 16816 21440 17141 21468
rect 16816 21428 16822 21440
rect 17129 21437 17141 21440
rect 17175 21437 17187 21471
rect 17129 21431 17187 21437
rect 17402 21428 17408 21480
rect 17460 21428 17466 21480
rect 18138 21428 18144 21480
rect 18196 21468 18202 21480
rect 19521 21471 19579 21477
rect 19521 21468 19533 21471
rect 18196 21440 19533 21468
rect 18196 21428 18202 21440
rect 19521 21437 19533 21440
rect 19567 21437 19579 21471
rect 19521 21431 19579 21437
rect 20257 21471 20315 21477
rect 20257 21437 20269 21471
rect 20303 21437 20315 21471
rect 20257 21431 20315 21437
rect 1026 21360 1032 21412
rect 1084 21400 1090 21412
rect 1949 21403 2007 21409
rect 1949 21400 1961 21403
rect 1084 21372 1961 21400
rect 1084 21360 1090 21372
rect 1949 21369 1961 21372
rect 1995 21369 2007 21403
rect 1949 21363 2007 21369
rect 4246 21360 4252 21412
rect 4304 21400 4310 21412
rect 4801 21403 4859 21409
rect 4801 21400 4813 21403
rect 4304 21372 4813 21400
rect 4304 21360 4310 21372
rect 4801 21369 4813 21372
rect 4847 21369 4859 21403
rect 4801 21363 4859 21369
rect 18877 21403 18935 21409
rect 18877 21369 18889 21403
rect 18923 21400 18935 21403
rect 19886 21400 19892 21412
rect 18923 21372 19892 21400
rect 18923 21369 18935 21372
rect 18877 21363 18935 21369
rect 19886 21360 19892 21372
rect 19944 21400 19950 21412
rect 20272 21400 20300 21431
rect 21634 21428 21640 21480
rect 21692 21428 21698 21480
rect 22066 21468 22094 21508
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22922 21536 22928 21548
rect 22244 21508 22928 21536
rect 22244 21496 22250 21508
rect 22922 21496 22928 21508
rect 22980 21496 22986 21548
rect 23192 21539 23250 21545
rect 23192 21505 23204 21539
rect 23238 21536 23250 21539
rect 23474 21536 23480 21548
rect 23238 21508 23480 21536
rect 23238 21505 23250 21508
rect 23192 21499 23250 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 23584 21536 23612 21576
rect 24688 21576 25044 21604
rect 24394 21536 24400 21548
rect 23584 21508 24400 21536
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 24578 21496 24584 21548
rect 24636 21496 24642 21548
rect 24688 21545 24716 21576
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 26418 21604 26424 21616
rect 25240 21576 26424 21604
rect 24673 21539 24731 21545
rect 24673 21505 24685 21539
rect 24719 21505 24731 21539
rect 24673 21499 24731 21505
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 22373 21471 22431 21477
rect 22373 21468 22385 21471
rect 22066 21440 22385 21468
rect 22373 21437 22385 21440
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 19944 21372 20300 21400
rect 24412 21400 24440 21496
rect 24780 21400 24808 21499
rect 24946 21496 24952 21548
rect 25004 21496 25010 21548
rect 25240 21536 25268 21576
rect 26418 21564 26424 21576
rect 26476 21564 26482 21616
rect 32392 21607 32450 21613
rect 32392 21573 32404 21607
rect 32438 21604 32450 21607
rect 32582 21604 32588 21616
rect 32438 21576 32588 21604
rect 32438 21573 32450 21576
rect 32392 21567 32450 21573
rect 32582 21564 32588 21576
rect 32640 21564 32646 21616
rect 33778 21564 33784 21616
rect 33836 21604 33842 21616
rect 34072 21613 34100 21644
rect 35250 21632 35256 21684
rect 35308 21632 35314 21684
rect 39485 21675 39543 21681
rect 39485 21641 39497 21675
rect 39531 21672 39543 21675
rect 39574 21672 39580 21684
rect 39531 21644 39580 21672
rect 39531 21641 39543 21644
rect 39485 21635 39543 21641
rect 39574 21632 39580 21644
rect 39632 21632 39638 21684
rect 39758 21632 39764 21684
rect 39816 21672 39822 21684
rect 39853 21675 39911 21681
rect 39853 21672 39865 21675
rect 39816 21644 39865 21672
rect 39816 21632 39822 21644
rect 39853 21641 39865 21644
rect 39899 21641 39911 21675
rect 39853 21635 39911 21641
rect 34057 21607 34115 21613
rect 33836 21576 34008 21604
rect 33836 21564 33842 21576
rect 25056 21508 25268 21536
rect 25308 21539 25366 21545
rect 25056 21480 25084 21508
rect 25308 21505 25320 21539
rect 25354 21536 25366 21539
rect 25590 21536 25596 21548
rect 25354 21508 25596 21536
rect 25354 21505 25366 21508
rect 25308 21499 25366 21505
rect 25590 21496 25596 21508
rect 25648 21496 25654 21548
rect 28077 21539 28135 21545
rect 28077 21505 28089 21539
rect 28123 21536 28135 21539
rect 28537 21539 28595 21545
rect 28537 21536 28549 21539
rect 28123 21508 28549 21536
rect 28123 21505 28135 21508
rect 28077 21499 28135 21505
rect 28537 21505 28549 21508
rect 28583 21505 28595 21539
rect 28537 21499 28595 21505
rect 30650 21496 30656 21548
rect 30708 21496 30714 21548
rect 31205 21539 31263 21545
rect 31205 21505 31217 21539
rect 31251 21536 31263 21539
rect 31938 21536 31944 21548
rect 31251 21508 31944 21536
rect 31251 21505 31263 21508
rect 31205 21499 31263 21505
rect 31938 21496 31944 21508
rect 31996 21496 32002 21548
rect 33873 21539 33931 21545
rect 33873 21505 33885 21539
rect 33919 21505 33931 21539
rect 33980 21536 34008 21576
rect 34057 21573 34069 21607
rect 34103 21573 34115 21607
rect 34057 21567 34115 21573
rect 34149 21607 34207 21613
rect 34149 21573 34161 21607
rect 34195 21604 34207 21607
rect 34330 21604 34336 21616
rect 34195 21576 34336 21604
rect 34195 21573 34207 21576
rect 34149 21567 34207 21573
rect 34330 21564 34336 21576
rect 34388 21564 34394 21616
rect 35529 21607 35587 21613
rect 35529 21573 35541 21607
rect 35575 21604 35587 21607
rect 35986 21604 35992 21616
rect 35575 21576 35992 21604
rect 35575 21573 35587 21576
rect 35529 21567 35587 21573
rect 35986 21564 35992 21576
rect 36044 21564 36050 21616
rect 40586 21604 40592 21616
rect 38778 21576 40592 21604
rect 40586 21564 40592 21576
rect 40644 21564 40650 21616
rect 41322 21564 41328 21616
rect 41380 21564 41386 21616
rect 34241 21539 34299 21545
rect 34241 21536 34253 21539
rect 33980 21508 34253 21536
rect 33873 21499 33931 21505
rect 34241 21505 34253 21508
rect 34287 21536 34299 21539
rect 35342 21536 35348 21548
rect 34287 21508 35348 21536
rect 34287 21505 34299 21508
rect 34241 21499 34299 21505
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 26973 21471 27031 21477
rect 26973 21437 26985 21471
rect 27019 21437 27031 21471
rect 26973 21431 27031 21437
rect 24412 21372 24808 21400
rect 26421 21403 26479 21409
rect 19944 21360 19950 21372
rect 26421 21369 26433 21403
rect 26467 21400 26479 21403
rect 26988 21400 27016 21431
rect 27246 21428 27252 21480
rect 27304 21468 27310 21480
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 27304 21440 28273 21468
rect 27304 21428 27310 21440
rect 28261 21437 28273 21440
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 28902 21428 28908 21480
rect 28960 21468 28966 21480
rect 29089 21471 29147 21477
rect 29089 21468 29101 21471
rect 28960 21440 29101 21468
rect 28960 21428 28966 21440
rect 29089 21437 29101 21440
rect 29135 21437 29147 21471
rect 29089 21431 29147 21437
rect 31386 21428 31392 21480
rect 31444 21428 31450 21480
rect 32122 21428 32128 21480
rect 32180 21428 32186 21480
rect 26467 21372 27016 21400
rect 26467 21369 26479 21372
rect 26421 21363 26479 21369
rect 4522 21292 4528 21344
rect 4580 21292 4586 21344
rect 6914 21292 6920 21344
rect 6972 21332 6978 21344
rect 7558 21332 7564 21344
rect 6972 21304 7564 21332
rect 6972 21292 6978 21304
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 14090 21292 14096 21344
rect 14148 21332 14154 21344
rect 14185 21335 14243 21341
rect 14185 21332 14197 21335
rect 14148 21304 14197 21332
rect 14148 21292 14154 21304
rect 14185 21301 14197 21304
rect 14231 21301 14243 21335
rect 14185 21295 14243 21301
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 18690 21332 18696 21344
rect 18196 21304 18696 21332
rect 18196 21292 18202 21304
rect 18690 21292 18696 21304
rect 18748 21332 18754 21344
rect 18969 21335 19027 21341
rect 18969 21332 18981 21335
rect 18748 21304 18981 21332
rect 18748 21292 18754 21304
rect 18969 21301 18981 21304
rect 19015 21301 19027 21335
rect 18969 21295 19027 21301
rect 19702 21292 19708 21344
rect 19760 21292 19766 21344
rect 20806 21292 20812 21344
rect 20864 21332 20870 21344
rect 20993 21335 21051 21341
rect 20993 21332 21005 21335
rect 20864 21304 21005 21332
rect 20864 21292 20870 21304
rect 20993 21301 21005 21304
rect 21039 21301 21051 21335
rect 20993 21295 21051 21301
rect 21174 21292 21180 21344
rect 21232 21332 21238 21344
rect 21726 21332 21732 21344
rect 21232 21304 21732 21332
rect 21232 21292 21238 21304
rect 21726 21292 21732 21304
rect 21784 21332 21790 21344
rect 21821 21335 21879 21341
rect 21821 21332 21833 21335
rect 21784 21304 21833 21332
rect 21784 21292 21790 21304
rect 21821 21301 21833 21304
rect 21867 21301 21879 21335
rect 21821 21295 21879 21301
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 23198 21332 23204 21344
rect 22152 21304 23204 21332
rect 22152 21292 22158 21304
rect 23198 21292 23204 21304
rect 23256 21292 23262 21344
rect 24670 21292 24676 21344
rect 24728 21332 24734 21344
rect 25222 21332 25228 21344
rect 24728 21304 25228 21332
rect 24728 21292 24734 21304
rect 25222 21292 25228 21304
rect 25280 21332 25286 21344
rect 27246 21332 27252 21344
rect 25280 21304 27252 21332
rect 25280 21292 25286 21304
rect 27246 21292 27252 21304
rect 27304 21292 27310 21344
rect 27522 21292 27528 21344
rect 27580 21332 27586 21344
rect 27617 21335 27675 21341
rect 27617 21332 27629 21335
rect 27580 21304 27629 21332
rect 27580 21292 27586 21304
rect 27617 21301 27629 21304
rect 27663 21301 27675 21335
rect 27617 21295 27675 21301
rect 27706 21292 27712 21344
rect 27764 21292 27770 21344
rect 30374 21292 30380 21344
rect 30432 21332 30438 21344
rect 30837 21335 30895 21341
rect 30837 21332 30849 21335
rect 30432 21304 30849 21332
rect 30432 21292 30438 21304
rect 30837 21301 30849 21304
rect 30883 21301 30895 21335
rect 33888 21332 33916 21499
rect 35342 21496 35348 21508
rect 35400 21536 35406 21548
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 35400 21508 35449 21536
rect 35400 21496 35406 21508
rect 35437 21505 35449 21508
rect 35483 21505 35495 21539
rect 35437 21499 35495 21505
rect 35618 21496 35624 21548
rect 35676 21496 35682 21548
rect 35805 21539 35863 21545
rect 35805 21505 35817 21539
rect 35851 21536 35863 21539
rect 36446 21536 36452 21548
rect 35851 21508 36452 21536
rect 35851 21505 35863 21508
rect 35805 21499 35863 21505
rect 36446 21496 36452 21508
rect 36504 21496 36510 21548
rect 39945 21539 40003 21545
rect 39945 21505 39957 21539
rect 39991 21536 40003 21539
rect 40126 21536 40132 21548
rect 39991 21508 40132 21536
rect 39991 21505 40003 21508
rect 39945 21499 40003 21505
rect 40126 21496 40132 21508
rect 40184 21496 40190 21548
rect 34698 21428 34704 21480
rect 34756 21468 34762 21480
rect 35069 21471 35127 21477
rect 35069 21468 35081 21471
rect 34756 21440 35081 21468
rect 34756 21428 34762 21440
rect 35069 21437 35081 21440
rect 35115 21437 35127 21471
rect 35069 21431 35127 21437
rect 37274 21428 37280 21480
rect 37332 21428 37338 21480
rect 37550 21428 37556 21480
rect 37608 21428 37614 21480
rect 37918 21428 37924 21480
rect 37976 21468 37982 21480
rect 38286 21468 38292 21480
rect 37976 21440 38292 21468
rect 37976 21428 37982 21440
rect 38286 21428 38292 21440
rect 38344 21468 38350 21480
rect 40037 21471 40095 21477
rect 40037 21468 40049 21471
rect 38344 21440 40049 21468
rect 38344 21428 38350 21440
rect 40037 21437 40049 21440
rect 40083 21437 40095 21471
rect 40037 21431 40095 21437
rect 40218 21428 40224 21480
rect 40276 21468 40282 21480
rect 40313 21471 40371 21477
rect 40313 21468 40325 21471
rect 40276 21440 40325 21468
rect 40276 21428 40282 21440
rect 40313 21437 40325 21440
rect 40359 21437 40371 21471
rect 40313 21431 40371 21437
rect 34425 21403 34483 21409
rect 34425 21369 34437 21403
rect 34471 21400 34483 21403
rect 36906 21400 36912 21412
rect 34471 21372 36912 21400
rect 34471 21369 34483 21372
rect 34425 21363 34483 21369
rect 36906 21360 36912 21372
rect 36964 21360 36970 21412
rect 39206 21360 39212 21412
rect 39264 21400 39270 21412
rect 40328 21400 40356 21431
rect 40586 21428 40592 21480
rect 40644 21428 40650 21480
rect 39264 21372 40356 21400
rect 39264 21360 39270 21372
rect 34330 21332 34336 21344
rect 33888 21304 34336 21332
rect 30837 21295 30895 21301
rect 34330 21292 34336 21304
rect 34388 21332 34394 21344
rect 34517 21335 34575 21341
rect 34517 21332 34529 21335
rect 34388 21304 34529 21332
rect 34388 21292 34394 21304
rect 34517 21301 34529 21304
rect 34563 21301 34575 21335
rect 34517 21295 34575 21301
rect 35618 21292 35624 21344
rect 35676 21332 35682 21344
rect 37918 21332 37924 21344
rect 35676 21304 37924 21332
rect 35676 21292 35682 21304
rect 37918 21292 37924 21304
rect 37976 21292 37982 21344
rect 38562 21292 38568 21344
rect 38620 21332 38626 21344
rect 39025 21335 39083 21341
rect 39025 21332 39037 21335
rect 38620 21304 39037 21332
rect 38620 21292 38626 21304
rect 39025 21301 39037 21304
rect 39071 21301 39083 21335
rect 39025 21295 39083 21301
rect 42058 21292 42064 21344
rect 42116 21292 42122 21344
rect 1104 21242 42504 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 42504 21242
rect 1104 21168 42504 21190
rect 1397 21131 1455 21137
rect 1397 21097 1409 21131
rect 1443 21128 1455 21131
rect 1762 21128 1768 21140
rect 1443 21100 1768 21128
rect 1443 21097 1455 21100
rect 1397 21091 1455 21097
rect 1762 21088 1768 21100
rect 1820 21088 1826 21140
rect 4890 21088 4896 21140
rect 4948 21128 4954 21140
rect 4948 21100 5396 21128
rect 4948 21088 4954 21100
rect 2866 20952 2872 21004
rect 2924 20952 2930 21004
rect 4706 20992 4712 21004
rect 3988 20964 4712 20992
rect 3142 20884 3148 20936
rect 3200 20884 3206 20936
rect 3878 20884 3884 20936
rect 3936 20924 3942 20936
rect 3988 20933 4016 20964
rect 4706 20952 4712 20964
rect 4764 20992 4770 21004
rect 4764 20964 5304 20992
rect 4764 20952 4770 20964
rect 3973 20927 4031 20933
rect 3973 20924 3985 20927
rect 3936 20896 3985 20924
rect 3936 20884 3942 20896
rect 3973 20893 3985 20896
rect 4019 20893 4031 20927
rect 3973 20887 4031 20893
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 4154 20924 4160 20936
rect 4111 20896 4160 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 4154 20884 4160 20896
rect 4212 20884 4218 20936
rect 4249 20927 4307 20933
rect 4249 20893 4261 20927
rect 4295 20893 4307 20927
rect 4249 20887 4307 20893
rect 4341 20927 4399 20933
rect 4341 20893 4353 20927
rect 4387 20924 4399 20927
rect 4798 20924 4804 20936
rect 4387 20896 4804 20924
rect 4387 20893 4399 20896
rect 4341 20887 4399 20893
rect 1854 20816 1860 20868
rect 1912 20816 1918 20868
rect 4264 20856 4292 20887
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 4890 20884 4896 20936
rect 4948 20884 4954 20936
rect 4982 20884 4988 20936
rect 5040 20884 5046 20936
rect 5276 20933 5304 20964
rect 5368 20936 5396 21100
rect 11146 21088 11152 21140
rect 11204 21088 11210 21140
rect 16574 21088 16580 21140
rect 16632 21088 16638 21140
rect 17402 21088 17408 21140
rect 17460 21128 17466 21140
rect 17681 21131 17739 21137
rect 17681 21128 17693 21131
rect 17460 21100 17693 21128
rect 17460 21088 17466 21100
rect 17681 21097 17693 21100
rect 17727 21097 17739 21131
rect 20990 21128 20996 21140
rect 17681 21091 17739 21097
rect 18524 21100 20996 21128
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 17862 21060 17868 21072
rect 15528 21032 17868 21060
rect 15528 21020 15534 21032
rect 17862 21020 17868 21032
rect 17920 21060 17926 21072
rect 17920 21032 18276 21060
rect 17920 21020 17926 21032
rect 18248 21004 18276 21032
rect 5537 20995 5595 21001
rect 5537 20961 5549 20995
rect 5583 20992 5595 20995
rect 6362 20992 6368 21004
rect 5583 20964 6368 20992
rect 5583 20961 5595 20964
rect 5537 20955 5595 20961
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 11882 20952 11888 21004
rect 11940 20992 11946 21004
rect 13814 20992 13820 21004
rect 11940 20964 13820 20992
rect 11940 20952 11946 20964
rect 13814 20952 13820 20964
rect 13872 20992 13878 21004
rect 14093 20995 14151 21001
rect 14093 20992 14105 20995
rect 13872 20964 14105 20992
rect 13872 20952 13878 20964
rect 14093 20961 14105 20964
rect 14139 20961 14151 20995
rect 14093 20955 14151 20961
rect 14369 20995 14427 21001
rect 14369 20961 14381 20995
rect 14415 20992 14427 20995
rect 14826 20992 14832 21004
rect 14415 20964 14832 20992
rect 14415 20961 14427 20964
rect 14369 20955 14427 20961
rect 14826 20952 14832 20964
rect 14884 20952 14890 21004
rect 15841 20995 15899 21001
rect 15841 20961 15853 20995
rect 15887 20992 15899 20995
rect 15933 20995 15991 21001
rect 15933 20992 15945 20995
rect 15887 20964 15945 20992
rect 15887 20961 15899 20964
rect 15841 20955 15899 20961
rect 15933 20961 15945 20964
rect 15979 20961 15991 20995
rect 15933 20955 15991 20961
rect 18138 20952 18144 21004
rect 18196 20952 18202 21004
rect 18230 20952 18236 21004
rect 18288 20952 18294 21004
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20893 5227 20927
rect 5169 20887 5227 20893
rect 5261 20927 5319 20933
rect 5261 20893 5273 20927
rect 5307 20893 5319 20927
rect 5261 20887 5319 20893
rect 5000 20856 5028 20884
rect 4264 20828 5028 20856
rect 3326 20748 3332 20800
rect 3384 20788 3390 20800
rect 3789 20791 3847 20797
rect 3789 20788 3801 20791
rect 3384 20760 3801 20788
rect 3384 20748 3390 20760
rect 3789 20757 3801 20760
rect 3835 20757 3847 20791
rect 5184 20788 5212 20887
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5445 20927 5503 20933
rect 5445 20893 5457 20927
rect 5491 20924 5503 20927
rect 5905 20927 5963 20933
rect 5905 20924 5917 20927
rect 5491 20896 5917 20924
rect 5491 20893 5503 20896
rect 5445 20887 5503 20893
rect 5905 20893 5917 20896
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 18524 20933 18552 21100
rect 20990 21088 20996 21100
rect 21048 21088 21054 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 23017 21131 23075 21137
rect 23017 21128 23029 21131
rect 22336 21100 23029 21128
rect 22336 21088 22342 21100
rect 23017 21097 23029 21100
rect 23063 21097 23075 21131
rect 23017 21091 23075 21097
rect 23474 21088 23480 21140
rect 23532 21088 23538 21140
rect 26252 21100 28488 21128
rect 21174 21060 21180 21072
rect 20916 21032 21180 21060
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 19150 20992 19156 21004
rect 18800 20964 19156 20992
rect 18800 20933 18828 20964
rect 19150 20952 19156 20964
rect 19208 20952 19214 21004
rect 20916 21001 20944 21032
rect 21174 21020 21180 21032
rect 21232 21020 21238 21072
rect 25682 21060 25688 21072
rect 23952 21032 25688 21060
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 20993 20995 21051 21001
rect 20993 20961 21005 20995
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 21269 20995 21327 21001
rect 21269 20961 21281 20995
rect 21315 20992 21327 20995
rect 22186 20992 22192 21004
rect 21315 20964 22192 20992
rect 21315 20961 21327 20964
rect 21269 20955 21327 20961
rect 16761 20927 16819 20933
rect 16761 20924 16773 20927
rect 16632 20896 16773 20924
rect 16632 20884 16638 20896
rect 16761 20893 16773 20896
rect 16807 20893 16819 20927
rect 16761 20887 16819 20893
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20893 18567 20927
rect 18509 20887 18567 20893
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 18874 20884 18880 20936
rect 18932 20884 18938 20936
rect 19061 20927 19119 20933
rect 19061 20893 19073 20927
rect 19107 20924 19119 20927
rect 19337 20927 19395 20933
rect 19337 20924 19349 20927
rect 19107 20896 19349 20924
rect 19107 20893 19119 20896
rect 19061 20887 19119 20893
rect 19337 20893 19349 20896
rect 19383 20893 19395 20927
rect 19337 20887 19395 20893
rect 20806 20884 20812 20936
rect 20864 20884 20870 20936
rect 6638 20816 6644 20868
rect 6696 20816 6702 20868
rect 7377 20859 7435 20865
rect 7377 20825 7389 20859
rect 7423 20856 7435 20859
rect 7558 20856 7564 20868
rect 7423 20828 7564 20856
rect 7423 20825 7435 20828
rect 7377 20819 7435 20825
rect 7392 20788 7420 20819
rect 7558 20816 7564 20828
rect 7616 20816 7622 20868
rect 10962 20816 10968 20868
rect 11020 20816 11026 20868
rect 11181 20859 11239 20865
rect 11181 20825 11193 20859
rect 11227 20856 11239 20859
rect 12158 20856 12164 20868
rect 11227 20828 12164 20856
rect 11227 20825 11239 20828
rect 11181 20819 11239 20825
rect 12158 20816 12164 20828
rect 12216 20816 12222 20868
rect 14918 20816 14924 20868
rect 14976 20816 14982 20868
rect 18049 20859 18107 20865
rect 18049 20825 18061 20859
rect 18095 20856 18107 20859
rect 19702 20856 19708 20868
rect 18095 20828 19708 20856
rect 18095 20825 18107 20828
rect 18049 20819 18107 20825
rect 19702 20816 19708 20828
rect 19760 20816 19766 20868
rect 21008 20856 21036 20955
rect 22186 20952 22192 20964
rect 22244 20952 22250 21004
rect 23952 21001 23980 21032
rect 24872 21001 24900 21032
rect 25682 21020 25688 21032
rect 25740 21020 25746 21072
rect 23937 20995 23995 21001
rect 23937 20961 23949 20995
rect 23983 20961 23995 20995
rect 23937 20955 23995 20961
rect 24029 20995 24087 21001
rect 24029 20961 24041 20995
rect 24075 20961 24087 20995
rect 24029 20955 24087 20961
rect 24857 20995 24915 21001
rect 24857 20961 24869 20995
rect 24903 20961 24915 20995
rect 24857 20955 24915 20961
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20992 25099 20995
rect 25222 20992 25228 21004
rect 25087 20964 25228 20992
rect 25087 20961 25099 20964
rect 25041 20955 25099 20961
rect 23750 20884 23756 20936
rect 23808 20924 23814 20936
rect 23845 20927 23903 20933
rect 23845 20924 23857 20927
rect 23808 20896 23857 20924
rect 23808 20884 23814 20896
rect 23845 20893 23857 20896
rect 23891 20893 23903 20927
rect 24044 20924 24072 20955
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 26145 20995 26203 21001
rect 26145 20992 26157 20995
rect 25323 20964 26157 20992
rect 25323 20924 25351 20964
rect 26145 20961 26157 20964
rect 26191 20992 26203 20995
rect 26252 20992 26280 21100
rect 28460 21060 28488 21100
rect 28902 21088 28908 21140
rect 28960 21088 28966 21140
rect 29012 21100 31432 21128
rect 28718 21060 28724 21072
rect 28460 21032 28724 21060
rect 28718 21020 28724 21032
rect 28776 21060 28782 21072
rect 29012 21060 29040 21100
rect 28776 21032 29040 21060
rect 28776 21020 28782 21032
rect 26191 20964 26280 20992
rect 27157 20995 27215 21001
rect 26191 20961 26203 20964
rect 26145 20955 26203 20961
rect 27157 20961 27169 20995
rect 27203 20992 27215 20995
rect 27430 20992 27436 21004
rect 27203 20964 27436 20992
rect 27203 20961 27215 20964
rect 27157 20955 27215 20961
rect 27430 20952 27436 20964
rect 27488 20952 27494 21004
rect 30098 20952 30104 21004
rect 30156 20952 30162 21004
rect 30374 20952 30380 21004
rect 30432 20952 30438 21004
rect 31404 20992 31432 21100
rect 31938 21088 31944 21140
rect 31996 21088 32002 21140
rect 35618 21128 35624 21140
rect 34900 21100 35624 21128
rect 34900 21072 34928 21100
rect 35618 21088 35624 21100
rect 35676 21088 35682 21140
rect 37185 21131 37243 21137
rect 37185 21097 37197 21131
rect 37231 21128 37243 21131
rect 37550 21128 37556 21140
rect 37231 21100 37556 21128
rect 37231 21097 37243 21100
rect 37185 21091 37243 21097
rect 37550 21088 37556 21100
rect 37608 21088 37614 21140
rect 40497 21131 40555 21137
rect 40497 21097 40509 21131
rect 40543 21128 40555 21131
rect 40586 21128 40592 21140
rect 40543 21100 40592 21128
rect 40543 21097 40555 21100
rect 40497 21091 40555 21097
rect 40586 21088 40592 21100
rect 40644 21088 40650 21140
rect 41138 21088 41144 21140
rect 41196 21128 41202 21140
rect 41325 21131 41383 21137
rect 41325 21128 41337 21131
rect 41196 21100 41337 21128
rect 41196 21088 41202 21100
rect 41325 21097 41337 21100
rect 41371 21097 41383 21131
rect 41325 21091 41383 21097
rect 31478 21020 31484 21072
rect 31536 21060 31542 21072
rect 33594 21060 33600 21072
rect 31536 21032 33600 21060
rect 31536 21020 31542 21032
rect 33594 21020 33600 21032
rect 33652 21020 33658 21072
rect 34882 21060 34888 21072
rect 33796 21032 34888 21060
rect 31404 20964 33456 20992
rect 23845 20887 23903 20893
rect 23952 20896 25351 20924
rect 25961 20927 26019 20933
rect 19904 20828 21036 20856
rect 5184 20760 7420 20788
rect 3789 20751 3847 20757
rect 11330 20748 11336 20800
rect 11388 20748 11394 20800
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17405 20791 17463 20797
rect 17405 20788 17417 20791
rect 17184 20760 17417 20788
rect 17184 20748 17190 20760
rect 17405 20757 17417 20760
rect 17451 20757 17463 20791
rect 17405 20751 17463 20757
rect 18230 20748 18236 20800
rect 18288 20788 18294 20800
rect 19904 20788 19932 20828
rect 21542 20816 21548 20868
rect 21600 20816 21606 20868
rect 22094 20816 22100 20868
rect 22152 20816 22158 20868
rect 18288 20760 19932 20788
rect 18288 20748 18294 20760
rect 19978 20748 19984 20800
rect 20036 20748 20042 20800
rect 20438 20748 20444 20800
rect 20496 20748 20502 20800
rect 21910 20748 21916 20800
rect 21968 20788 21974 20800
rect 23952 20788 23980 20896
rect 25961 20893 25973 20927
rect 26007 20924 26019 20927
rect 26786 20924 26792 20936
rect 26007 20896 26792 20924
rect 26007 20893 26019 20896
rect 25961 20887 26019 20893
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 26970 20884 26976 20936
rect 27028 20884 27034 20936
rect 33428 20933 33456 20964
rect 33796 20936 33824 21032
rect 34882 21020 34888 21032
rect 34940 21020 34946 21072
rect 35253 21063 35311 21069
rect 35253 21029 35265 21063
rect 35299 21060 35311 21063
rect 36722 21060 36728 21072
rect 35299 21032 36728 21060
rect 35299 21029 35311 21032
rect 35253 21023 35311 21029
rect 36722 21020 36728 21032
rect 36780 21020 36786 21072
rect 37274 21020 37280 21072
rect 37332 21060 37338 21072
rect 37332 21032 41092 21060
rect 37332 21020 37338 21032
rect 37642 20952 37648 21004
rect 37700 20952 37706 21004
rect 37844 21001 37872 21032
rect 37829 20995 37887 21001
rect 37829 20961 37841 20995
rect 37875 20961 37887 20995
rect 37829 20955 37887 20961
rect 38562 20952 38568 21004
rect 38620 20992 38626 21004
rect 41064 21001 41092 21032
rect 39577 20995 39635 21001
rect 39577 20992 39589 20995
rect 38620 20964 39589 20992
rect 38620 20952 38626 20964
rect 39577 20961 39589 20964
rect 39623 20961 39635 20995
rect 39577 20955 39635 20961
rect 41049 20995 41107 21001
rect 41049 20961 41061 20995
rect 41095 20961 41107 20995
rect 41049 20955 41107 20961
rect 41506 20952 41512 21004
rect 41564 20992 41570 21004
rect 41877 20995 41935 21001
rect 41877 20992 41889 20995
rect 41564 20964 41889 20992
rect 41564 20952 41570 20964
rect 41877 20961 41889 20964
rect 41923 20961 41935 20995
rect 41877 20955 41935 20961
rect 32493 20927 32551 20933
rect 32493 20924 32505 20927
rect 31864 20896 32505 20924
rect 24210 20816 24216 20868
rect 24268 20856 24274 20868
rect 24765 20859 24823 20865
rect 24268 20828 24716 20856
rect 24268 20816 24274 20828
rect 21968 20760 23980 20788
rect 21968 20748 21974 20760
rect 24026 20748 24032 20800
rect 24084 20788 24090 20800
rect 24397 20791 24455 20797
rect 24397 20788 24409 20791
rect 24084 20760 24409 20788
rect 24084 20748 24090 20760
rect 24397 20757 24409 20760
rect 24443 20757 24455 20791
rect 24688 20788 24716 20828
rect 24765 20825 24777 20859
rect 24811 20856 24823 20859
rect 26421 20859 26479 20865
rect 26421 20856 26433 20859
rect 24811 20828 26433 20856
rect 24811 20825 24823 20828
rect 24765 20819 24823 20825
rect 26421 20825 26433 20828
rect 26467 20825 26479 20859
rect 26421 20819 26479 20825
rect 27433 20859 27491 20865
rect 27433 20825 27445 20859
rect 27479 20856 27491 20859
rect 27706 20856 27712 20868
rect 27479 20828 27712 20856
rect 27479 20825 27491 20828
rect 27433 20819 27491 20825
rect 27706 20816 27712 20828
rect 27764 20816 27770 20868
rect 29454 20856 29460 20868
rect 28658 20828 29460 20856
rect 29454 20816 29460 20828
rect 29512 20816 29518 20868
rect 30374 20816 30380 20868
rect 30432 20856 30438 20868
rect 30834 20856 30840 20868
rect 30432 20828 30840 20856
rect 30432 20816 30438 20828
rect 30834 20816 30840 20828
rect 30892 20816 30898 20868
rect 24946 20788 24952 20800
rect 24688 20760 24952 20788
rect 24397 20751 24455 20757
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 25590 20748 25596 20800
rect 25648 20748 25654 20800
rect 26053 20791 26111 20797
rect 26053 20757 26065 20791
rect 26099 20788 26111 20791
rect 27522 20788 27528 20800
rect 26099 20760 27528 20788
rect 26099 20757 26111 20760
rect 26053 20751 26111 20757
rect 27522 20748 27528 20760
rect 27580 20748 27586 20800
rect 31754 20748 31760 20800
rect 31812 20788 31818 20800
rect 31864 20797 31892 20896
rect 32493 20893 32505 20896
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 33413 20927 33471 20933
rect 33413 20893 33425 20927
rect 33459 20893 33471 20927
rect 33413 20887 33471 20893
rect 33597 20927 33655 20933
rect 33597 20893 33609 20927
rect 33643 20924 33655 20927
rect 33778 20924 33784 20936
rect 33643 20896 33784 20924
rect 33643 20893 33655 20896
rect 33597 20887 33655 20893
rect 33778 20884 33784 20896
rect 33836 20884 33842 20936
rect 34054 20884 34060 20936
rect 34112 20924 34118 20936
rect 34241 20927 34299 20933
rect 34241 20924 34253 20927
rect 34112 20896 34253 20924
rect 34112 20884 34118 20896
rect 34241 20893 34253 20896
rect 34287 20893 34299 20927
rect 34241 20887 34299 20893
rect 34701 20927 34759 20933
rect 34701 20893 34713 20927
rect 34747 20893 34759 20927
rect 34701 20887 34759 20893
rect 31849 20791 31907 20797
rect 31849 20788 31861 20791
rect 31812 20760 31861 20788
rect 31812 20748 31818 20760
rect 31849 20757 31861 20760
rect 31895 20757 31907 20791
rect 31849 20751 31907 20757
rect 33594 20748 33600 20800
rect 33652 20788 33658 20800
rect 33689 20791 33747 20797
rect 33689 20788 33701 20791
rect 33652 20760 33701 20788
rect 33652 20748 33658 20760
rect 33689 20757 33701 20760
rect 33735 20757 33747 20791
rect 34716 20788 34744 20887
rect 34974 20884 34980 20936
rect 35032 20884 35038 20936
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20924 35127 20927
rect 35250 20924 35256 20936
rect 35115 20896 35256 20924
rect 35115 20893 35127 20896
rect 35069 20887 35127 20893
rect 35250 20884 35256 20896
rect 35308 20884 35314 20936
rect 35342 20884 35348 20936
rect 35400 20884 35406 20936
rect 37553 20927 37611 20933
rect 37553 20893 37565 20927
rect 37599 20924 37611 20927
rect 39025 20927 39083 20933
rect 39025 20924 39037 20927
rect 37599 20896 39037 20924
rect 37599 20893 37611 20896
rect 37553 20887 37611 20893
rect 39025 20893 39037 20896
rect 39071 20893 39083 20927
rect 39025 20887 39083 20893
rect 34882 20816 34888 20868
rect 34940 20816 34946 20868
rect 38010 20816 38016 20868
rect 38068 20816 38074 20868
rect 38841 20859 38899 20865
rect 38841 20825 38853 20859
rect 38887 20856 38899 20859
rect 39206 20856 39212 20868
rect 38887 20828 39212 20856
rect 38887 20825 38899 20828
rect 38841 20819 38899 20825
rect 39206 20816 39212 20828
rect 39264 20856 39270 20868
rect 39853 20859 39911 20865
rect 39853 20856 39865 20859
rect 39264 20828 39865 20856
rect 39264 20816 39270 20828
rect 39853 20825 39865 20828
rect 39899 20825 39911 20859
rect 39853 20819 39911 20825
rect 40865 20859 40923 20865
rect 40865 20825 40877 20859
rect 40911 20856 40923 20859
rect 41506 20856 41512 20868
rect 40911 20828 41512 20856
rect 40911 20825 40923 20828
rect 40865 20819 40923 20825
rect 41506 20816 41512 20828
rect 41564 20816 41570 20868
rect 35989 20791 36047 20797
rect 35989 20788 36001 20791
rect 34716 20760 36001 20788
rect 33689 20751 33747 20757
rect 35989 20757 36001 20760
rect 36035 20788 36047 20791
rect 36262 20788 36268 20800
rect 36035 20760 36268 20788
rect 36035 20757 36047 20760
rect 35989 20751 36047 20757
rect 36262 20748 36268 20760
rect 36320 20748 36326 20800
rect 40126 20748 40132 20800
rect 40184 20788 40190 20800
rect 40957 20791 41015 20797
rect 40957 20788 40969 20791
rect 40184 20760 40969 20788
rect 40184 20748 40190 20760
rect 40957 20757 40969 20760
rect 41003 20757 41015 20791
rect 40957 20751 41015 20757
rect 1104 20698 42504 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 42504 20698
rect 1104 20624 42504 20646
rect 1854 20544 1860 20596
rect 1912 20584 1918 20596
rect 1912 20556 3648 20584
rect 1912 20544 1918 20556
rect 3620 20516 3648 20556
rect 4614 20544 4620 20596
rect 4672 20584 4678 20596
rect 5166 20584 5172 20596
rect 4672 20556 5172 20584
rect 4672 20544 4678 20556
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 5258 20544 5264 20596
rect 5316 20544 5322 20596
rect 5350 20544 5356 20596
rect 5408 20584 5414 20596
rect 5445 20587 5503 20593
rect 5445 20584 5457 20587
rect 5408 20556 5457 20584
rect 5408 20544 5414 20556
rect 5445 20553 5457 20556
rect 5491 20553 5503 20587
rect 5445 20547 5503 20553
rect 5810 20544 5816 20596
rect 5868 20544 5874 20596
rect 8754 20544 8760 20596
rect 8812 20584 8818 20596
rect 14090 20584 14096 20596
rect 8812 20556 14096 20584
rect 8812 20544 8818 20556
rect 3694 20516 3700 20528
rect 3620 20488 3700 20516
rect 3694 20476 3700 20488
rect 3752 20476 3758 20528
rect 6086 20516 6092 20528
rect 4908 20488 5580 20516
rect 2222 20408 2228 20460
rect 2280 20448 2286 20460
rect 2280 20420 3280 20448
rect 2280 20408 2286 20420
rect 2961 20383 3019 20389
rect 2961 20349 2973 20383
rect 3007 20380 3019 20383
rect 3142 20380 3148 20392
rect 3007 20352 3148 20380
rect 3007 20349 3019 20352
rect 2961 20343 3019 20349
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 3252 20380 3280 20420
rect 3326 20408 3332 20460
rect 3384 20408 3390 20460
rect 4706 20408 4712 20460
rect 4764 20448 4770 20460
rect 4908 20457 4936 20488
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 4764 20420 4905 20448
rect 4764 20408 4770 20420
rect 4893 20417 4905 20420
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 5350 20408 5356 20460
rect 5408 20408 5414 20460
rect 5552 20457 5580 20488
rect 5644 20488 6092 20516
rect 5644 20460 5672 20488
rect 6086 20476 6092 20488
rect 6144 20476 6150 20528
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20417 5595 20451
rect 5537 20411 5595 20417
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 8956 20457 8984 20556
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14608 20556 15025 20584
rect 14608 20544 14614 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 16850 20544 16856 20596
rect 16908 20584 16914 20596
rect 17037 20587 17095 20593
rect 17037 20584 17049 20587
rect 16908 20556 17049 20584
rect 16908 20544 16914 20556
rect 17037 20553 17049 20556
rect 17083 20553 17095 20587
rect 22094 20584 22100 20596
rect 17037 20547 17095 20553
rect 19904 20556 22100 20584
rect 10689 20519 10747 20525
rect 10689 20516 10701 20519
rect 10244 20488 10701 20516
rect 10244 20457 10272 20488
rect 10689 20485 10701 20488
rect 10735 20485 10747 20519
rect 10689 20479 10747 20485
rect 11330 20476 11336 20528
rect 11388 20516 11394 20528
rect 11762 20519 11820 20525
rect 11762 20516 11774 20519
rect 11388 20488 11774 20516
rect 11388 20476 11394 20488
rect 11762 20485 11774 20488
rect 11808 20485 11820 20519
rect 11762 20479 11820 20485
rect 13814 20476 13820 20528
rect 13872 20516 13878 20528
rect 15194 20516 15200 20528
rect 13872 20488 15200 20516
rect 13872 20476 13878 20488
rect 15194 20476 15200 20488
rect 15252 20516 15258 20528
rect 15289 20519 15347 20525
rect 15289 20516 15301 20519
rect 15252 20488 15301 20516
rect 15252 20476 15258 20488
rect 15289 20485 15301 20488
rect 15335 20485 15347 20519
rect 15289 20479 15347 20485
rect 16117 20519 16175 20525
rect 16117 20485 16129 20519
rect 16163 20516 16175 20519
rect 16163 20488 19288 20516
rect 16163 20485 16175 20488
rect 16117 20479 16175 20485
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5776 20420 5825 20448
rect 5776 20408 5782 20420
rect 5813 20417 5825 20420
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 10594 20408 10600 20460
rect 10652 20448 10658 20460
rect 11514 20448 11520 20460
rect 10652 20420 11520 20448
rect 10652 20408 10658 20420
rect 11514 20408 11520 20420
rect 11572 20408 11578 20460
rect 11606 20408 11612 20460
rect 11664 20408 11670 20460
rect 12986 20408 12992 20460
rect 13044 20448 13050 20460
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 13044 20420 14197 20448
rect 13044 20408 13050 20420
rect 14185 20417 14197 20420
rect 14231 20417 14243 20451
rect 14185 20411 14243 20417
rect 14366 20408 14372 20460
rect 14424 20408 14430 20460
rect 14553 20451 14611 20457
rect 14553 20417 14565 20451
rect 14599 20448 14611 20451
rect 14829 20451 14887 20457
rect 14599 20420 14780 20448
rect 14599 20417 14611 20420
rect 14553 20411 14611 20417
rect 4985 20383 5043 20389
rect 4985 20380 4997 20383
rect 3252 20352 4997 20380
rect 4985 20349 4997 20352
rect 5031 20349 5043 20383
rect 4985 20343 5043 20349
rect 9950 20340 9956 20392
rect 10008 20340 10014 20392
rect 10318 20340 10324 20392
rect 10376 20340 10382 20392
rect 11333 20383 11391 20389
rect 11333 20349 11345 20383
rect 11379 20380 11391 20383
rect 11624 20380 11652 20408
rect 11379 20352 11652 20380
rect 11379 20349 11391 20352
rect 11333 20343 11391 20349
rect 14090 20340 14096 20392
rect 14148 20340 14154 20392
rect 14752 20380 14780 20420
rect 14829 20417 14841 20451
rect 14875 20448 14887 20451
rect 15010 20448 15016 20460
rect 14875 20420 15016 20448
rect 14875 20417 14887 20420
rect 14829 20411 14887 20417
rect 15010 20408 15016 20420
rect 15068 20408 15074 20460
rect 15102 20408 15108 20460
rect 15160 20408 15166 20460
rect 16022 20380 16028 20392
rect 14200 20352 14596 20380
rect 14752 20352 16028 20380
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 4755 20315 4813 20321
rect 4755 20312 4767 20315
rect 4212 20284 4767 20312
rect 4212 20272 4218 20284
rect 4755 20281 4767 20284
rect 4801 20312 4813 20315
rect 5442 20312 5448 20324
rect 4801 20284 5448 20312
rect 4801 20281 4813 20284
rect 4755 20275 4813 20281
rect 5442 20272 5448 20284
rect 5500 20272 5506 20324
rect 8202 20272 8208 20324
rect 8260 20312 8266 20324
rect 9309 20315 9367 20321
rect 9309 20312 9321 20315
rect 8260 20284 9321 20312
rect 8260 20272 8266 20284
rect 9309 20281 9321 20284
rect 9355 20281 9367 20315
rect 14200 20312 14228 20352
rect 9309 20275 9367 20281
rect 12820 20284 14228 20312
rect 14568 20312 14596 20352
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 16132 20312 16160 20479
rect 16209 20451 16267 20457
rect 16209 20417 16221 20451
rect 16255 20448 16267 20451
rect 16255 20420 17356 20448
rect 16255 20417 16267 20420
rect 16209 20411 16267 20417
rect 17126 20340 17132 20392
rect 17184 20340 17190 20392
rect 17328 20389 17356 20420
rect 17770 20408 17776 20460
rect 17828 20448 17834 20460
rect 17937 20451 17995 20457
rect 17937 20448 17949 20451
rect 17828 20420 17949 20448
rect 17828 20408 17834 20420
rect 17937 20417 17949 20420
rect 17983 20417 17995 20451
rect 17937 20411 17995 20417
rect 17313 20383 17371 20389
rect 17313 20349 17325 20383
rect 17359 20380 17371 20383
rect 17586 20380 17592 20392
rect 17359 20352 17592 20380
rect 17359 20349 17371 20352
rect 17313 20343 17371 20349
rect 17586 20340 17592 20352
rect 17644 20340 17650 20392
rect 17678 20340 17684 20392
rect 17736 20340 17742 20392
rect 14568 20284 16160 20312
rect 16224 20284 16804 20312
rect 5077 20247 5135 20253
rect 5077 20213 5089 20247
rect 5123 20244 5135 20247
rect 5718 20244 5724 20256
rect 5123 20216 5724 20244
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 9125 20247 9183 20253
rect 9125 20244 9137 20247
rect 8536 20216 9137 20244
rect 8536 20204 8542 20216
rect 9125 20213 9137 20216
rect 9171 20244 9183 20247
rect 9582 20244 9588 20256
rect 9171 20216 9588 20244
rect 9171 20213 9183 20216
rect 9125 20207 9183 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10686 20244 10692 20256
rect 10643 20216 10692 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 10778 20204 10784 20256
rect 10836 20244 10842 20256
rect 12820 20244 12848 20284
rect 10836 20216 12848 20244
rect 10836 20204 10842 20216
rect 12894 20204 12900 20256
rect 12952 20204 12958 20256
rect 14366 20204 14372 20256
rect 14424 20244 14430 20256
rect 14737 20247 14795 20253
rect 14737 20244 14749 20247
rect 14424 20216 14749 20244
rect 14424 20204 14430 20216
rect 14737 20213 14749 20216
rect 14783 20244 14795 20247
rect 16224 20244 16252 20284
rect 14783 20216 16252 20244
rect 14783 20213 14795 20216
rect 14737 20207 14795 20213
rect 16298 20204 16304 20256
rect 16356 20204 16362 20256
rect 16482 20204 16488 20256
rect 16540 20244 16546 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16540 20216 16681 20244
rect 16540 20204 16546 20216
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 16776 20244 16804 20284
rect 18598 20244 18604 20256
rect 16776 20216 18604 20244
rect 16669 20207 16727 20213
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 19024 20216 19073 20244
rect 19024 20204 19030 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 19150 20204 19156 20256
rect 19208 20204 19214 20256
rect 19260 20244 19288 20488
rect 19904 20457 19932 20556
rect 22094 20544 22100 20556
rect 22152 20544 22158 20596
rect 22278 20544 22284 20596
rect 22336 20544 22342 20596
rect 23934 20544 23940 20596
rect 23992 20584 23998 20596
rect 24765 20587 24823 20593
rect 24765 20584 24777 20587
rect 23992 20556 24777 20584
rect 23992 20544 23998 20556
rect 24765 20553 24777 20556
rect 24811 20584 24823 20587
rect 26970 20584 26976 20596
rect 24811 20556 26976 20584
rect 24811 20553 24823 20556
rect 24765 20547 24823 20553
rect 26970 20544 26976 20556
rect 27028 20544 27034 20596
rect 27433 20587 27491 20593
rect 27433 20553 27445 20587
rect 27479 20584 27491 20587
rect 27522 20584 27528 20596
rect 27479 20556 27528 20584
rect 27479 20553 27491 20556
rect 27433 20547 27491 20553
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 29362 20544 29368 20596
rect 29420 20584 29426 20596
rect 29549 20587 29607 20593
rect 29549 20584 29561 20587
rect 29420 20556 29561 20584
rect 29420 20544 29426 20556
rect 29549 20553 29561 20556
rect 29595 20553 29607 20587
rect 29549 20547 29607 20553
rect 31938 20544 31944 20596
rect 31996 20584 32002 20596
rect 32674 20584 32680 20596
rect 31996 20556 32680 20584
rect 31996 20544 32002 20556
rect 32674 20544 32680 20556
rect 32732 20544 32738 20596
rect 33410 20544 33416 20596
rect 33468 20584 33474 20596
rect 34054 20584 34060 20596
rect 33468 20556 34060 20584
rect 33468 20544 33474 20556
rect 34054 20544 34060 20556
rect 34112 20544 34118 20596
rect 36648 20556 41414 20584
rect 20165 20519 20223 20525
rect 20165 20485 20177 20519
rect 20211 20516 20223 20519
rect 20438 20516 20444 20528
rect 20211 20488 20444 20516
rect 20211 20485 20223 20488
rect 20165 20479 20223 20485
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 21450 20516 21456 20528
rect 21390 20488 21456 20516
rect 21450 20476 21456 20488
rect 21508 20516 21514 20528
rect 21726 20516 21732 20528
rect 21508 20488 21732 20516
rect 21508 20476 21514 20488
rect 21726 20476 21732 20488
rect 21784 20476 21790 20528
rect 23198 20476 23204 20528
rect 23256 20516 23262 20528
rect 23750 20516 23756 20528
rect 23256 20488 23756 20516
rect 23256 20476 23262 20488
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 25406 20476 25412 20528
rect 25464 20516 25470 20528
rect 29454 20516 29460 20528
rect 25464 20488 25806 20516
rect 29302 20488 29460 20516
rect 25464 20476 25470 20488
rect 29454 20476 29460 20488
rect 29512 20516 29518 20528
rect 36648 20516 36676 20556
rect 29512 20488 30958 20516
rect 33810 20488 36676 20516
rect 29512 20476 29518 20488
rect 36722 20476 36728 20528
rect 36780 20525 36786 20528
rect 36780 20516 36792 20525
rect 36780 20488 36825 20516
rect 36780 20479 36792 20488
rect 36780 20476 36786 20479
rect 37458 20476 37464 20528
rect 37516 20516 37522 20528
rect 37645 20519 37703 20525
rect 37645 20516 37657 20519
rect 37516 20488 37657 20516
rect 37516 20476 37522 20488
rect 37645 20485 37657 20488
rect 37691 20485 37703 20519
rect 37645 20479 37703 20485
rect 37826 20476 37832 20528
rect 37884 20516 37890 20528
rect 37884 20488 38410 20516
rect 37884 20476 37890 20488
rect 40126 20476 40132 20528
rect 40184 20516 40190 20528
rect 40313 20519 40371 20525
rect 40313 20516 40325 20519
rect 40184 20488 40325 20516
rect 40184 20476 40190 20488
rect 40313 20485 40325 20488
rect 40359 20485 40371 20519
rect 41386 20516 41414 20556
rect 41506 20544 41512 20596
rect 41564 20544 41570 20596
rect 41690 20516 41696 20528
rect 41386 20488 41696 20516
rect 40313 20479 40371 20485
rect 41690 20476 41696 20488
rect 41748 20476 41754 20528
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 22278 20408 22284 20460
rect 22336 20448 22342 20460
rect 22336 20420 22508 20448
rect 22336 20408 22342 20420
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20380 19855 20383
rect 20898 20380 20904 20392
rect 19843 20352 20904 20380
rect 19843 20349 19855 20352
rect 19797 20343 19855 20349
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 21634 20340 21640 20392
rect 21692 20340 21698 20392
rect 22370 20340 22376 20392
rect 22428 20340 22434 20392
rect 22480 20389 22508 20420
rect 26786 20408 26792 20460
rect 26844 20448 26850 20460
rect 26844 20420 27292 20448
rect 26844 20408 26850 20420
rect 27264 20392 27292 20420
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27430 20408 27436 20460
rect 27488 20448 27494 20460
rect 27801 20451 27859 20457
rect 27801 20448 27813 20451
rect 27488 20420 27813 20448
rect 27488 20408 27494 20420
rect 27801 20417 27813 20420
rect 27847 20417 27859 20451
rect 27801 20411 27859 20417
rect 33870 20408 33876 20460
rect 33928 20448 33934 20460
rect 34054 20448 34060 20460
rect 33928 20420 34060 20448
rect 33928 20408 33934 20420
rect 34054 20408 34060 20420
rect 34112 20408 34118 20460
rect 34422 20457 34428 20460
rect 34416 20411 34428 20457
rect 34422 20408 34428 20411
rect 34480 20408 34486 20460
rect 40678 20408 40684 20460
rect 40736 20448 40742 20460
rect 40865 20451 40923 20457
rect 40865 20448 40877 20451
rect 40736 20420 40877 20448
rect 40736 20408 40742 20420
rect 40865 20417 40877 20420
rect 40911 20417 40923 20451
rect 41263 20451 41321 20457
rect 41263 20448 41275 20451
rect 40865 20411 40923 20417
rect 40972 20420 41275 20448
rect 22465 20383 22523 20389
rect 22465 20349 22477 20383
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 23017 20383 23075 20389
rect 23017 20349 23029 20383
rect 23063 20349 23075 20383
rect 23017 20343 23075 20349
rect 23293 20383 23351 20389
rect 23293 20349 23305 20383
rect 23339 20380 23351 20383
rect 24026 20380 24032 20392
rect 23339 20352 24032 20380
rect 23339 20349 23351 20352
rect 23293 20343 23351 20349
rect 21542 20272 21548 20324
rect 21600 20312 21606 20324
rect 21913 20315 21971 20321
rect 21913 20312 21925 20315
rect 21600 20284 21925 20312
rect 21600 20272 21606 20284
rect 21913 20281 21925 20284
rect 21959 20281 21971 20315
rect 21913 20275 21971 20281
rect 22094 20272 22100 20324
rect 22152 20312 22158 20324
rect 23032 20312 23060 20343
rect 24026 20340 24032 20352
rect 24084 20340 24090 20392
rect 25038 20340 25044 20392
rect 25096 20340 25102 20392
rect 25317 20383 25375 20389
rect 25317 20349 25329 20383
rect 25363 20380 25375 20383
rect 25363 20352 27016 20380
rect 25363 20349 25375 20352
rect 25317 20343 25375 20349
rect 26988 20321 27016 20352
rect 27246 20340 27252 20392
rect 27304 20380 27310 20392
rect 27525 20383 27583 20389
rect 27525 20380 27537 20383
rect 27304 20352 27537 20380
rect 27304 20340 27310 20352
rect 27525 20349 27537 20352
rect 27571 20349 27583 20383
rect 27525 20343 27583 20349
rect 28077 20383 28135 20389
rect 28077 20349 28089 20383
rect 28123 20380 28135 20383
rect 28442 20380 28448 20392
rect 28123 20352 28448 20380
rect 28123 20349 28135 20352
rect 28077 20343 28135 20349
rect 28442 20340 28448 20352
rect 28500 20340 28506 20392
rect 30193 20383 30251 20389
rect 30193 20349 30205 20383
rect 30239 20349 30251 20383
rect 30193 20343 30251 20349
rect 30469 20383 30527 20389
rect 30469 20349 30481 20383
rect 30515 20380 30527 20383
rect 31202 20380 31208 20392
rect 30515 20352 31208 20380
rect 30515 20349 30527 20352
rect 30469 20343 30527 20349
rect 22152 20284 23060 20312
rect 26973 20315 27031 20321
rect 22152 20272 22158 20284
rect 26973 20281 26985 20315
rect 27019 20281 27031 20315
rect 26973 20275 27031 20281
rect 21266 20244 21272 20256
rect 19260 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 23014 20244 23020 20256
rect 21876 20216 23020 20244
rect 21876 20204 21882 20216
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 26789 20247 26847 20253
rect 26789 20213 26801 20247
rect 26835 20244 26847 20247
rect 27154 20244 27160 20256
rect 26835 20216 27160 20244
rect 26835 20213 26847 20216
rect 26789 20207 26847 20213
rect 27154 20204 27160 20216
rect 27212 20204 27218 20256
rect 30208 20244 30236 20343
rect 31202 20340 31208 20352
rect 31260 20340 31266 20392
rect 32309 20383 32367 20389
rect 32309 20349 32321 20383
rect 32355 20349 32367 20383
rect 32309 20343 32367 20349
rect 32122 20244 32128 20256
rect 30208 20216 32128 20244
rect 32122 20204 32128 20216
rect 32180 20244 32186 20256
rect 32324 20244 32352 20343
rect 32582 20340 32588 20392
rect 32640 20340 32646 20392
rect 34149 20383 34207 20389
rect 34149 20349 34161 20383
rect 34195 20349 34207 20383
rect 34149 20343 34207 20349
rect 37001 20383 37059 20389
rect 37001 20349 37013 20383
rect 37047 20380 37059 20383
rect 37366 20380 37372 20392
rect 37047 20352 37372 20380
rect 37047 20349 37059 20352
rect 37001 20343 37059 20349
rect 32766 20244 32772 20256
rect 32180 20216 32772 20244
rect 32180 20204 32186 20216
rect 32766 20204 32772 20216
rect 32824 20244 32830 20256
rect 34164 20244 34192 20343
rect 37366 20340 37372 20352
rect 37424 20340 37430 20392
rect 37734 20340 37740 20392
rect 37792 20340 37798 20392
rect 37921 20383 37979 20389
rect 37921 20349 37933 20383
rect 37967 20380 37979 20383
rect 37967 20352 38056 20380
rect 37967 20349 37979 20352
rect 37921 20343 37979 20349
rect 35342 20272 35348 20324
rect 35400 20312 35406 20324
rect 35621 20315 35679 20321
rect 35621 20312 35633 20315
rect 35400 20284 35633 20312
rect 35400 20272 35406 20284
rect 35621 20281 35633 20284
rect 35667 20281 35679 20315
rect 35621 20275 35679 20281
rect 32824 20216 34192 20244
rect 32824 20204 32830 20216
rect 35526 20204 35532 20256
rect 35584 20204 35590 20256
rect 36354 20204 36360 20256
rect 36412 20244 36418 20256
rect 37277 20247 37335 20253
rect 37277 20244 37289 20247
rect 36412 20216 37289 20244
rect 36412 20204 36418 20216
rect 37277 20213 37289 20216
rect 37323 20213 37335 20247
rect 38028 20244 38056 20352
rect 38102 20340 38108 20392
rect 38160 20340 38166 20392
rect 39574 20340 39580 20392
rect 39632 20340 39638 20392
rect 39853 20383 39911 20389
rect 39853 20349 39865 20383
rect 39899 20349 39911 20383
rect 39853 20343 39911 20349
rect 38470 20244 38476 20256
rect 38028 20216 38476 20244
rect 37277 20207 37335 20213
rect 38470 20204 38476 20216
rect 38528 20244 38534 20256
rect 39114 20244 39120 20256
rect 38528 20216 39120 20244
rect 38528 20204 38534 20216
rect 39114 20204 39120 20216
rect 39172 20204 39178 20256
rect 39206 20204 39212 20256
rect 39264 20244 39270 20256
rect 39868 20244 39896 20343
rect 40310 20340 40316 20392
rect 40368 20380 40374 20392
rect 40972 20380 41000 20420
rect 41263 20417 41275 20420
rect 41309 20417 41321 20451
rect 41263 20411 41321 20417
rect 41417 20451 41475 20457
rect 41417 20417 41429 20451
rect 41463 20448 41475 20451
rect 41782 20448 41788 20460
rect 41463 20420 41788 20448
rect 41463 20417 41475 20420
rect 41417 20411 41475 20417
rect 41782 20408 41788 20420
rect 41840 20408 41846 20460
rect 42058 20408 42064 20460
rect 42116 20408 42122 20460
rect 40368 20352 41000 20380
rect 40368 20340 40374 20352
rect 40034 20272 40040 20324
rect 40092 20312 40098 20324
rect 41049 20315 41107 20321
rect 41049 20312 41061 20315
rect 40092 20284 41061 20312
rect 40092 20272 40098 20284
rect 41049 20281 41061 20284
rect 41095 20281 41107 20315
rect 41049 20275 41107 20281
rect 39264 20216 39896 20244
rect 39264 20204 39270 20216
rect 1104 20154 42504 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 42504 20154
rect 1104 20080 42504 20102
rect 5810 20000 5816 20052
rect 5868 20040 5874 20052
rect 5868 20012 9904 20040
rect 5868 20000 5874 20012
rect 5718 19932 5724 19984
rect 5776 19932 5782 19984
rect 9876 19972 9904 20012
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10008 20012 10333 20040
rect 10008 20000 10014 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 12158 20000 12164 20052
rect 12216 20000 12222 20052
rect 16301 20043 16359 20049
rect 16301 20009 16313 20043
rect 16347 20040 16359 20043
rect 16574 20040 16580 20052
rect 16347 20012 16580 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17770 20000 17776 20052
rect 17828 20000 17834 20052
rect 18233 20043 18291 20049
rect 18233 20009 18245 20043
rect 18279 20040 18291 20043
rect 18598 20040 18604 20052
rect 18279 20012 18604 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 18598 20000 18604 20012
rect 18656 20000 18662 20052
rect 19150 20000 19156 20052
rect 19208 20040 19214 20052
rect 22462 20040 22468 20052
rect 19208 20012 22468 20040
rect 19208 20000 19214 20012
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 27062 20000 27068 20052
rect 27120 20000 27126 20052
rect 27338 20000 27344 20052
rect 27396 20040 27402 20052
rect 27801 20043 27859 20049
rect 27801 20040 27813 20043
rect 27396 20012 27813 20040
rect 27396 20000 27402 20012
rect 27801 20009 27813 20012
rect 27847 20009 27859 20043
rect 27801 20003 27859 20009
rect 28442 20000 28448 20052
rect 28500 20000 28506 20052
rect 31202 20000 31208 20052
rect 31260 20000 31266 20052
rect 32582 20000 32588 20052
rect 32640 20040 32646 20052
rect 32769 20043 32827 20049
rect 32769 20040 32781 20043
rect 32640 20012 32781 20040
rect 32640 20000 32646 20012
rect 32769 20009 32781 20012
rect 32815 20009 32827 20043
rect 32769 20003 32827 20009
rect 34422 20000 34428 20052
rect 34480 20040 34486 20052
rect 34517 20043 34575 20049
rect 34517 20040 34529 20043
rect 34480 20012 34529 20040
rect 34480 20000 34486 20012
rect 34517 20009 34529 20012
rect 34563 20009 34575 20043
rect 34517 20003 34575 20009
rect 37458 20000 37464 20052
rect 37516 20040 37522 20052
rect 37829 20043 37887 20049
rect 37829 20040 37841 20043
rect 37516 20012 37841 20040
rect 37516 20000 37522 20012
rect 37829 20009 37841 20012
rect 37875 20009 37887 20043
rect 37829 20003 37887 20009
rect 38657 20043 38715 20049
rect 38657 20009 38669 20043
rect 38703 20040 38715 20043
rect 39574 20040 39580 20052
rect 38703 20012 39580 20040
rect 38703 20009 38715 20012
rect 38657 20003 38715 20009
rect 39574 20000 39580 20012
rect 39632 20000 39638 20052
rect 10502 19972 10508 19984
rect 9876 19944 10508 19972
rect 10502 19932 10508 19944
rect 10560 19932 10566 19984
rect 41322 19972 41328 19984
rect 38212 19944 41328 19972
rect 5736 19904 5764 19932
rect 5994 19904 6000 19916
rect 5736 19876 6000 19904
rect 5994 19864 6000 19876
rect 6052 19864 6058 19916
rect 6086 19864 6092 19916
rect 6144 19864 6150 19916
rect 8113 19907 8171 19913
rect 8113 19873 8125 19907
rect 8159 19904 8171 19907
rect 8294 19904 8300 19916
rect 8159 19876 8300 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 14921 19907 14979 19913
rect 14921 19904 14933 19907
rect 13872 19876 14933 19904
rect 13872 19864 13878 19876
rect 14921 19873 14933 19876
rect 14967 19873 14979 19907
rect 14921 19867 14979 19873
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 5813 19839 5871 19845
rect 5813 19836 5825 19839
rect 5776 19808 5825 19836
rect 5776 19796 5782 19808
rect 5813 19805 5825 19808
rect 5859 19805 5871 19839
rect 5813 19799 5871 19805
rect 5902 19796 5908 19848
rect 5960 19836 5966 19848
rect 5960 19808 6500 19836
rect 5960 19796 5966 19808
rect 2406 19728 2412 19780
rect 2464 19768 2470 19780
rect 3142 19768 3148 19780
rect 2464 19740 3148 19768
rect 2464 19728 2470 19740
rect 3142 19728 3148 19740
rect 3200 19768 3206 19780
rect 3789 19771 3847 19777
rect 3789 19768 3801 19771
rect 3200 19740 3801 19768
rect 3200 19728 3206 19740
rect 3789 19737 3801 19740
rect 3835 19768 3847 19771
rect 4614 19768 4620 19780
rect 3835 19740 4620 19768
rect 3835 19737 3847 19740
rect 3789 19731 3847 19737
rect 4614 19728 4620 19740
rect 4672 19768 4678 19780
rect 6362 19768 6368 19780
rect 4672 19740 6368 19768
rect 4672 19728 4678 19740
rect 6362 19728 6368 19740
rect 6420 19728 6426 19780
rect 6270 19660 6276 19712
rect 6328 19660 6334 19712
rect 6472 19709 6500 19808
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 8202 19796 8208 19848
rect 8260 19796 8266 19848
rect 8941 19839 8999 19845
rect 8941 19805 8953 19839
rect 8987 19836 8999 19839
rect 10594 19836 10600 19848
rect 8987 19808 10600 19836
rect 8987 19805 8999 19808
rect 8941 19799 8999 19805
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 10686 19796 10692 19848
rect 10744 19836 10750 19848
rect 10853 19839 10911 19845
rect 10853 19836 10865 19839
rect 10744 19808 10865 19836
rect 10744 19796 10750 19808
rect 10853 19805 10865 19808
rect 10899 19805 10911 19839
rect 10853 19799 10911 19805
rect 12250 19796 12256 19848
rect 12308 19796 12314 19848
rect 14936 19836 14964 19867
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 18874 19904 18880 19916
rect 16356 19876 18880 19904
rect 16356 19864 16362 19876
rect 16393 19839 16451 19845
rect 16393 19836 16405 19839
rect 14936 19808 16405 19836
rect 16393 19805 16405 19808
rect 16439 19836 16451 19839
rect 16666 19836 16672 19848
rect 16439 19808 16672 19836
rect 16439 19805 16451 19808
rect 16393 19799 16451 19805
rect 16666 19796 16672 19808
rect 16724 19836 16730 19848
rect 17678 19836 17684 19848
rect 16724 19808 17684 19836
rect 16724 19796 16730 19808
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 17972 19845 18000 19876
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 25038 19864 25044 19916
rect 25096 19904 25102 19916
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 25096 19876 25329 19904
rect 25096 19864 25102 19876
rect 25317 19873 25329 19876
rect 25363 19904 25375 19907
rect 27430 19904 27436 19916
rect 25363 19876 27436 19904
rect 25363 19873 25375 19876
rect 25317 19867 25375 19873
rect 27430 19864 27436 19876
rect 27488 19864 27494 19916
rect 28074 19864 28080 19916
rect 28132 19904 28138 19916
rect 28997 19907 29055 19913
rect 28997 19904 29009 19907
rect 28132 19876 29009 19904
rect 28132 19864 28138 19876
rect 28997 19873 29009 19876
rect 29043 19904 29055 19907
rect 31757 19907 31815 19913
rect 31757 19904 31769 19907
rect 29043 19876 31769 19904
rect 29043 19873 29055 19876
rect 28997 19867 29055 19873
rect 31757 19873 31769 19876
rect 31803 19873 31815 19907
rect 31757 19867 31815 19873
rect 33226 19864 33232 19916
rect 33284 19864 33290 19916
rect 33413 19907 33471 19913
rect 33413 19873 33425 19907
rect 33459 19904 33471 19907
rect 33502 19904 33508 19916
rect 33459 19876 33508 19904
rect 33459 19873 33471 19876
rect 33413 19867 33471 19873
rect 33502 19864 33508 19876
rect 33560 19864 33566 19916
rect 33778 19864 33784 19916
rect 33836 19904 33842 19916
rect 33873 19907 33931 19913
rect 33873 19904 33885 19907
rect 33836 19876 33885 19904
rect 33836 19864 33842 19876
rect 33873 19873 33885 19876
rect 33919 19873 33931 19907
rect 33873 19867 33931 19873
rect 35526 19864 35532 19916
rect 35584 19864 35590 19916
rect 36081 19907 36139 19913
rect 36081 19873 36093 19907
rect 36127 19904 36139 19907
rect 37366 19904 37372 19916
rect 36127 19876 37372 19904
rect 36127 19873 36139 19876
rect 36081 19867 36139 19873
rect 37366 19864 37372 19876
rect 37424 19864 37430 19916
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 17957 19799 18015 19805
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 18325 19839 18383 19845
rect 18325 19805 18337 19839
rect 18371 19836 18383 19839
rect 18414 19836 18420 19848
rect 18371 19808 18420 19836
rect 18371 19805 18383 19808
rect 18325 19799 18383 19805
rect 9186 19771 9244 19777
rect 9186 19768 9198 19771
rect 8588 19740 9198 19768
rect 8588 19709 8616 19740
rect 9186 19737 9198 19740
rect 9232 19737 9244 19771
rect 9186 19731 9244 19737
rect 13572 19771 13630 19777
rect 13572 19737 13584 19771
rect 13618 19768 13630 19771
rect 13906 19768 13912 19780
rect 13618 19740 13912 19768
rect 13618 19737 13630 19740
rect 13572 19731 13630 19737
rect 13906 19728 13912 19740
rect 13964 19728 13970 19780
rect 15188 19771 15246 19777
rect 15188 19737 15200 19771
rect 15234 19768 15246 19771
rect 16482 19768 16488 19780
rect 15234 19740 16488 19768
rect 15234 19737 15246 19740
rect 15188 19731 15246 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 6457 19703 6515 19709
rect 6457 19669 6469 19703
rect 6503 19669 6515 19703
rect 6457 19663 6515 19669
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19669 8631 19703
rect 8573 19663 8631 19669
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 11664 19672 11989 19700
rect 11664 19660 11670 19672
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 11977 19663 12035 19669
rect 12342 19660 12348 19712
rect 12400 19700 12406 19712
rect 12437 19703 12495 19709
rect 12437 19700 12449 19703
rect 12400 19672 12449 19700
rect 12400 19660 12406 19672
rect 12437 19669 12449 19672
rect 12483 19669 12495 19703
rect 12437 19663 12495 19669
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 15746 19700 15752 19712
rect 14148 19672 15752 19700
rect 14148 19660 14154 19672
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 18064 19700 18092 19799
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19061 19839 19119 19845
rect 19061 19836 19073 19839
rect 19024 19808 19073 19836
rect 19024 19796 19030 19808
rect 19061 19805 19073 19808
rect 19107 19836 19119 19839
rect 19150 19836 19156 19848
rect 19107 19808 19156 19836
rect 19107 19805 19119 19808
rect 19061 19799 19119 19805
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 19242 19796 19248 19848
rect 19300 19796 19306 19848
rect 19512 19839 19570 19845
rect 19512 19805 19524 19839
rect 19558 19836 19570 19839
rect 19978 19836 19984 19848
rect 19558 19808 19984 19836
rect 19558 19805 19570 19808
rect 19512 19799 19570 19805
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 27154 19796 27160 19848
rect 27212 19796 27218 19848
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 29270 19836 29276 19848
rect 28859 19808 29276 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 29270 19796 29276 19808
rect 29328 19796 29334 19848
rect 31573 19839 31631 19845
rect 31573 19805 31585 19839
rect 31619 19836 31631 19839
rect 31938 19836 31944 19848
rect 31619 19808 31944 19836
rect 31619 19805 31631 19808
rect 31573 19799 31631 19805
rect 31938 19796 31944 19808
rect 31996 19796 32002 19848
rect 33137 19839 33195 19845
rect 33137 19805 33149 19839
rect 33183 19836 33195 19839
rect 33594 19836 33600 19848
rect 33183 19808 33600 19836
rect 33183 19805 33195 19808
rect 33137 19799 33195 19805
rect 33594 19796 33600 19808
rect 33652 19796 33658 19848
rect 34146 19796 34152 19848
rect 34204 19796 34210 19848
rect 38102 19796 38108 19848
rect 38160 19796 38166 19848
rect 38212 19845 38240 19944
rect 41322 19932 41328 19944
rect 41380 19932 41386 19984
rect 38286 19864 38292 19916
rect 38344 19904 38350 19916
rect 38344 19876 39068 19904
rect 38344 19864 38350 19876
rect 38197 19839 38255 19845
rect 38197 19805 38209 19839
rect 38243 19805 38255 19839
rect 38197 19799 38255 19805
rect 38473 19839 38531 19845
rect 38473 19805 38485 19839
rect 38519 19836 38531 19839
rect 38930 19836 38936 19848
rect 38519 19808 38936 19836
rect 38519 19805 38531 19808
rect 38473 19799 38531 19805
rect 38930 19796 38936 19808
rect 38988 19796 38994 19848
rect 39040 19845 39068 19876
rect 39114 19864 39120 19916
rect 39172 19904 39178 19916
rect 39209 19907 39267 19913
rect 39209 19904 39221 19907
rect 39172 19876 39221 19904
rect 39172 19864 39178 19876
rect 39209 19873 39221 19876
rect 39255 19873 39267 19907
rect 39209 19867 39267 19873
rect 39316 19876 40172 19904
rect 39025 19839 39083 19845
rect 39025 19805 39037 19839
rect 39071 19805 39083 19839
rect 39316 19836 39344 19876
rect 39025 19799 39083 19805
rect 39132 19808 39344 19836
rect 25590 19728 25596 19780
rect 25648 19728 25654 19780
rect 25700 19740 26082 19768
rect 18417 19703 18475 19709
rect 18417 19700 18429 19703
rect 18064 19672 18429 19700
rect 18417 19669 18429 19672
rect 18463 19700 18475 19703
rect 18506 19700 18512 19712
rect 18463 19672 18512 19700
rect 18463 19669 18475 19672
rect 18417 19663 18475 19669
rect 18506 19660 18512 19672
rect 18564 19660 18570 19712
rect 20625 19703 20683 19709
rect 20625 19669 20637 19703
rect 20671 19700 20683 19703
rect 20898 19700 20904 19712
rect 20671 19672 20904 19700
rect 20671 19669 20683 19672
rect 20625 19663 20683 19669
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 25700 19700 25728 19740
rect 28718 19728 28724 19780
rect 28776 19768 28782 19780
rect 28905 19771 28963 19777
rect 28905 19768 28917 19771
rect 28776 19740 28917 19768
rect 28776 19728 28782 19740
rect 28905 19737 28917 19740
rect 28951 19737 28963 19771
rect 28905 19731 28963 19737
rect 36354 19728 36360 19780
rect 36412 19728 36418 19780
rect 37826 19768 37832 19780
rect 37582 19740 37832 19768
rect 37826 19728 37832 19740
rect 37884 19728 37890 19780
rect 38286 19728 38292 19780
rect 38344 19728 38350 19780
rect 39132 19777 39160 19808
rect 39390 19796 39396 19848
rect 39448 19836 39454 19848
rect 40144 19845 40172 19876
rect 40037 19839 40095 19845
rect 40037 19836 40049 19839
rect 39448 19808 40049 19836
rect 39448 19796 39454 19808
rect 40037 19805 40049 19808
rect 40083 19805 40095 19839
rect 40037 19799 40095 19805
rect 40129 19839 40187 19845
rect 40129 19805 40141 19839
rect 40175 19805 40187 19839
rect 40129 19799 40187 19805
rect 40405 19839 40463 19845
rect 40405 19805 40417 19839
rect 40451 19836 40463 19839
rect 40586 19836 40592 19848
rect 40451 19808 40592 19836
rect 40451 19805 40463 19808
rect 40405 19799 40463 19805
rect 39117 19771 39175 19777
rect 39117 19737 39129 19771
rect 39163 19737 39175 19771
rect 39117 19731 39175 19737
rect 23808 19672 25728 19700
rect 23808 19660 23814 19672
rect 28166 19660 28172 19712
rect 28224 19700 28230 19712
rect 30374 19700 30380 19712
rect 28224 19672 30380 19700
rect 28224 19660 28230 19672
rect 30374 19660 30380 19672
rect 30432 19660 30438 19712
rect 31662 19660 31668 19712
rect 31720 19660 31726 19712
rect 34057 19703 34115 19709
rect 34057 19669 34069 19703
rect 34103 19700 34115 19703
rect 34790 19700 34796 19712
rect 34103 19672 34796 19700
rect 34103 19669 34115 19672
rect 34057 19663 34115 19669
rect 34790 19660 34796 19672
rect 34848 19700 34854 19712
rect 34885 19703 34943 19709
rect 34885 19700 34897 19703
rect 34848 19672 34897 19700
rect 34848 19660 34854 19672
rect 34885 19669 34897 19672
rect 34931 19669 34943 19703
rect 34885 19663 34943 19669
rect 37918 19660 37924 19712
rect 37976 19660 37982 19712
rect 38010 19660 38016 19712
rect 38068 19700 38074 19712
rect 39390 19700 39396 19712
rect 38068 19672 39396 19700
rect 38068 19660 38074 19672
rect 39390 19660 39396 19672
rect 39448 19660 39454 19712
rect 39482 19660 39488 19712
rect 39540 19700 39546 19712
rect 39853 19703 39911 19709
rect 39853 19700 39865 19703
rect 39540 19672 39865 19700
rect 39540 19660 39546 19672
rect 39853 19669 39865 19672
rect 39899 19669 39911 19703
rect 40144 19700 40172 19799
rect 40586 19796 40592 19808
rect 40644 19796 40650 19848
rect 41138 19796 41144 19848
rect 41196 19796 41202 19848
rect 42150 19796 42156 19848
rect 42208 19796 42214 19848
rect 40218 19728 40224 19780
rect 40276 19728 40282 19780
rect 40589 19703 40647 19709
rect 40589 19700 40601 19703
rect 40144 19672 40601 19700
rect 39853 19663 39911 19669
rect 40589 19669 40601 19672
rect 40635 19669 40647 19703
rect 40589 19663 40647 19669
rect 41506 19660 41512 19712
rect 41564 19660 41570 19712
rect 1104 19610 42504 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 42504 19610
rect 1104 19536 42504 19558
rect 5810 19496 5816 19508
rect 3896 19468 5816 19496
rect 3786 19388 3792 19440
rect 3844 19428 3850 19440
rect 3896 19428 3924 19468
rect 5810 19456 5816 19468
rect 5868 19456 5874 19508
rect 5997 19499 6055 19505
rect 5997 19465 6009 19499
rect 6043 19496 6055 19499
rect 6086 19496 6092 19508
rect 6043 19468 6092 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 8205 19499 8263 19505
rect 8205 19465 8217 19499
rect 8251 19496 8263 19499
rect 8294 19496 8300 19508
rect 8251 19468 8300 19496
rect 8251 19465 8263 19468
rect 8205 19459 8263 19465
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 12069 19499 12127 19505
rect 12069 19465 12081 19499
rect 12115 19496 12127 19499
rect 12434 19496 12440 19508
rect 12115 19468 12440 19496
rect 12115 19465 12127 19468
rect 12069 19459 12127 19465
rect 12434 19456 12440 19468
rect 12492 19496 12498 19508
rect 12894 19496 12900 19508
rect 12492 19468 12900 19496
rect 12492 19456 12498 19468
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 15102 19456 15108 19508
rect 15160 19496 15166 19508
rect 16390 19496 16396 19508
rect 15160 19468 16396 19496
rect 15160 19456 15166 19468
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 16485 19499 16543 19505
rect 16485 19465 16497 19499
rect 16531 19496 16543 19499
rect 16574 19496 16580 19508
rect 16531 19468 16580 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 18414 19456 18420 19508
rect 18472 19496 18478 19508
rect 19058 19496 19064 19508
rect 18472 19468 19064 19496
rect 18472 19456 18478 19468
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 19536 19468 21864 19496
rect 3844 19400 3924 19428
rect 9432 19431 9490 19437
rect 3844 19388 3850 19400
rect 9432 19397 9444 19431
rect 9478 19428 9490 19431
rect 9674 19428 9680 19440
rect 9478 19400 9680 19428
rect 9478 19397 9490 19400
rect 9432 19391 9490 19397
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 10134 19388 10140 19440
rect 10192 19428 10198 19440
rect 10778 19428 10784 19440
rect 10192 19400 10784 19428
rect 10192 19388 10198 19400
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 11164 19400 12173 19428
rect 2406 19320 2412 19372
rect 2464 19320 2470 19372
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 4341 19363 4399 19369
rect 4341 19360 4353 19363
rect 2823 19332 2930 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 2902 19292 2930 19332
rect 3528 19332 4353 19360
rect 3528 19292 3556 19332
rect 4341 19329 4353 19332
rect 4387 19329 4399 19363
rect 4341 19323 4399 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5905 19363 5963 19369
rect 5905 19360 5917 19363
rect 4764 19332 5917 19360
rect 4764 19320 4770 19332
rect 5905 19329 5917 19332
rect 5951 19360 5963 19363
rect 5994 19360 6000 19372
rect 5951 19332 6000 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 6362 19320 6368 19372
rect 6420 19320 6426 19372
rect 6638 19369 6644 19372
rect 6632 19323 6644 19369
rect 6638 19320 6644 19323
rect 6696 19320 6702 19372
rect 8018 19320 8024 19372
rect 8076 19320 8082 19372
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19360 8263 19363
rect 8251 19332 8340 19360
rect 8251 19329 8263 19332
rect 8205 19323 8263 19329
rect 2902 19264 3556 19292
rect 3602 19252 3608 19304
rect 3660 19292 3666 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 3660 19264 4905 19292
rect 3660 19252 3666 19264
rect 4893 19261 4905 19264
rect 4939 19261 4951 19295
rect 4893 19255 4951 19261
rect 5074 19184 5080 19236
rect 5132 19224 5138 19236
rect 5442 19224 5448 19236
rect 5132 19196 5448 19224
rect 5132 19184 5138 19196
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 5629 19227 5687 19233
rect 5629 19193 5641 19227
rect 5675 19224 5687 19227
rect 5718 19224 5724 19236
rect 5675 19196 5724 19224
rect 5675 19193 5687 19196
rect 5629 19187 5687 19193
rect 5718 19184 5724 19196
rect 5776 19224 5782 19236
rect 8312 19233 8340 19332
rect 10318 19320 10324 19372
rect 10376 19360 10382 19372
rect 11164 19369 11192 19400
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 13817 19431 13875 19437
rect 13817 19397 13829 19431
rect 13863 19428 13875 19431
rect 13863 19400 13952 19428
rect 13863 19397 13875 19400
rect 13817 19391 13875 19397
rect 13924 19369 13952 19400
rect 17678 19388 17684 19440
rect 17736 19388 17742 19440
rect 11149 19363 11207 19369
rect 11149 19360 11161 19363
rect 10376 19332 11161 19360
rect 10376 19320 10382 19332
rect 11149 19329 11161 19332
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 11977 19323 12035 19329
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 13541 19363 13599 19369
rect 13541 19360 13553 19363
rect 13495 19332 13553 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 13541 19329 13553 19332
rect 13587 19329 13599 19363
rect 13541 19323 13599 19329
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19329 13967 19363
rect 13909 19323 13967 19329
rect 14093 19363 14151 19369
rect 14093 19329 14105 19363
rect 14139 19329 14151 19363
rect 14093 19323 14151 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19360 15163 19363
rect 15194 19360 15200 19372
rect 15151 19332 15200 19360
rect 15151 19329 15163 19332
rect 15105 19323 15163 19329
rect 9677 19295 9735 19301
rect 9677 19261 9689 19295
rect 9723 19292 9735 19295
rect 10686 19292 10692 19304
rect 9723 19264 10692 19292
rect 9723 19261 9735 19264
rect 9677 19255 9735 19261
rect 10686 19252 10692 19264
rect 10744 19292 10750 19304
rect 10873 19295 10931 19301
rect 10873 19292 10885 19295
rect 10744 19264 10885 19292
rect 10744 19252 10750 19264
rect 10873 19261 10885 19264
rect 10919 19292 10931 19295
rect 11422 19292 11428 19304
rect 10919 19264 11428 19292
rect 10919 19261 10931 19264
rect 10873 19255 10931 19261
rect 11422 19252 11428 19264
rect 11480 19252 11486 19304
rect 11992 19292 12020 19323
rect 12342 19292 12348 19304
rect 11992 19264 12348 19292
rect 12342 19252 12348 19264
rect 12400 19292 12406 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12400 19264 12817 19292
rect 12400 19252 12406 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13814 19252 13820 19304
rect 13872 19252 13878 19304
rect 8297 19227 8355 19233
rect 5776 19196 6408 19224
rect 5776 19184 5782 19196
rect 4203 19159 4261 19165
rect 4203 19125 4215 19159
rect 4249 19156 4261 19159
rect 4982 19156 4988 19168
rect 4249 19128 4988 19156
rect 4249 19125 4261 19128
rect 4203 19119 4261 19125
rect 4982 19116 4988 19128
rect 5040 19156 5046 19168
rect 5810 19156 5816 19168
rect 5040 19128 5816 19156
rect 5040 19116 5046 19128
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 6178 19116 6184 19168
rect 6236 19116 6242 19168
rect 6380 19156 6408 19196
rect 8297 19193 8309 19227
rect 8343 19224 8355 19227
rect 8662 19224 8668 19236
rect 8343 19196 8668 19224
rect 8343 19193 8355 19196
rect 8297 19187 8355 19193
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 11606 19184 11612 19236
rect 11664 19224 11670 19236
rect 11793 19227 11851 19233
rect 11793 19224 11805 19227
rect 11664 19196 11805 19224
rect 11664 19184 11670 19196
rect 11793 19193 11805 19196
rect 11839 19193 11851 19227
rect 11793 19187 11851 19193
rect 11882 19184 11888 19236
rect 11940 19224 11946 19236
rect 12250 19224 12256 19236
rect 11940 19196 12256 19224
rect 11940 19184 11946 19196
rect 12250 19184 12256 19196
rect 12308 19224 12314 19236
rect 13633 19227 13691 19233
rect 13633 19224 13645 19227
rect 12308 19196 13645 19224
rect 12308 19184 12314 19196
rect 13633 19193 13645 19196
rect 13679 19193 13691 19227
rect 13633 19187 13691 19193
rect 13906 19184 13912 19236
rect 13964 19184 13970 19236
rect 7742 19156 7748 19168
rect 6380 19128 7748 19156
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 11241 19159 11299 19165
rect 11241 19125 11253 19159
rect 11287 19156 11299 19159
rect 12066 19156 12072 19168
rect 11287 19128 12072 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 12345 19159 12403 19165
rect 12345 19125 12357 19159
rect 12391 19156 12403 19159
rect 13078 19156 13084 19168
rect 12391 19128 13084 19156
rect 12391 19125 12403 19128
rect 12345 19119 12403 19125
rect 13078 19116 13084 19128
rect 13136 19156 13142 19168
rect 14108 19156 14136 19323
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15378 19369 15384 19372
rect 15372 19323 15384 19369
rect 15378 19320 15384 19323
rect 15436 19320 15442 19372
rect 16666 19320 16672 19372
rect 16724 19320 16730 19372
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 19536 19369 19564 19468
rect 21174 19428 21180 19440
rect 21022 19400 21180 19428
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 21836 19428 21864 19468
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 23661 19499 23719 19505
rect 23661 19496 23673 19499
rect 22428 19468 23673 19496
rect 22428 19456 22434 19468
rect 23661 19465 23673 19468
rect 23707 19465 23719 19499
rect 23661 19459 23719 19465
rect 25590 19456 25596 19508
rect 25648 19456 25654 19508
rect 25961 19499 26019 19505
rect 25961 19465 25973 19499
rect 26007 19496 26019 19499
rect 27062 19496 27068 19508
rect 26007 19468 27068 19496
rect 26007 19465 26019 19468
rect 25961 19459 26019 19465
rect 27062 19456 27068 19468
rect 27120 19456 27126 19508
rect 28718 19456 28724 19508
rect 28776 19496 28782 19508
rect 29273 19499 29331 19505
rect 29273 19496 29285 19499
rect 28776 19468 29285 19496
rect 28776 19456 28782 19468
rect 29273 19465 29285 19468
rect 29319 19465 29331 19499
rect 33042 19496 33048 19508
rect 29273 19459 29331 19465
rect 32692 19468 33048 19496
rect 22094 19428 22100 19440
rect 21836 19400 22100 19428
rect 21836 19369 21864 19400
rect 22094 19388 22100 19400
rect 22152 19388 22158 19440
rect 25038 19428 25044 19440
rect 23322 19400 25044 19428
rect 25038 19388 25044 19400
rect 25096 19428 25102 19440
rect 25406 19428 25412 19440
rect 25096 19400 25412 19428
rect 25096 19388 25102 19400
rect 25406 19388 25412 19400
rect 25464 19428 25470 19440
rect 28166 19428 28172 19440
rect 25464 19400 28172 19428
rect 25464 19388 25470 19400
rect 28166 19388 28172 19400
rect 28224 19388 28230 19440
rect 32692 19437 32720 19468
rect 33042 19456 33048 19468
rect 33100 19496 33106 19508
rect 33229 19499 33287 19505
rect 33229 19496 33241 19499
rect 33100 19468 33241 19496
rect 33100 19456 33106 19468
rect 33229 19465 33241 19468
rect 33275 19465 33287 19499
rect 33229 19459 33287 19465
rect 33686 19456 33692 19508
rect 33744 19496 33750 19508
rect 34330 19496 34336 19508
rect 33744 19468 34336 19496
rect 33744 19456 33750 19468
rect 34330 19456 34336 19468
rect 34388 19456 34394 19508
rect 38286 19456 38292 19508
rect 38344 19496 38350 19508
rect 38473 19499 38531 19505
rect 38473 19496 38485 19499
rect 38344 19468 38485 19496
rect 38344 19456 38350 19468
rect 38473 19465 38485 19468
rect 38519 19465 38531 19499
rect 38473 19459 38531 19465
rect 38930 19456 38936 19508
rect 38988 19496 38994 19508
rect 40770 19496 40776 19508
rect 38988 19468 40776 19496
rect 38988 19456 38994 19468
rect 40770 19456 40776 19468
rect 40828 19456 40834 19508
rect 40957 19499 41015 19505
rect 40957 19465 40969 19499
rect 41003 19496 41015 19499
rect 41138 19496 41144 19508
rect 41003 19468 41144 19496
rect 41003 19465 41015 19468
rect 40957 19459 41015 19465
rect 41138 19456 41144 19468
rect 41196 19456 41202 19508
rect 32677 19431 32735 19437
rect 32677 19397 32689 19431
rect 32723 19397 32735 19431
rect 38562 19428 38568 19440
rect 32677 19391 32735 19397
rect 32876 19400 34652 19428
rect 32876 19372 32904 19400
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19300 19332 19533 19360
rect 19300 19320 19306 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 27430 19320 27436 19372
rect 27488 19320 27494 19372
rect 29914 19320 29920 19372
rect 29972 19360 29978 19372
rect 30193 19363 30251 19369
rect 30193 19360 30205 19363
rect 29972 19332 30205 19360
rect 29972 19320 29978 19332
rect 30193 19329 30205 19332
rect 30239 19329 30251 19363
rect 30193 19323 30251 19329
rect 32122 19320 32128 19372
rect 32180 19360 32186 19372
rect 32493 19363 32551 19369
rect 32493 19360 32505 19363
rect 32180 19332 32505 19360
rect 32180 19320 32186 19332
rect 32493 19329 32505 19332
rect 32539 19329 32551 19363
rect 32493 19323 32551 19329
rect 32769 19363 32827 19369
rect 32769 19329 32781 19363
rect 32815 19329 32827 19363
rect 32769 19323 32827 19329
rect 16942 19252 16948 19304
rect 17000 19252 17006 19304
rect 19797 19295 19855 19301
rect 19797 19261 19809 19295
rect 19843 19292 19855 19295
rect 20254 19292 20260 19304
rect 19843 19264 20260 19292
rect 19843 19261 19855 19264
rect 19797 19255 19855 19261
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 21269 19295 21327 19301
rect 21269 19261 21281 19295
rect 21315 19292 21327 19295
rect 21358 19292 21364 19304
rect 21315 19264 21364 19292
rect 21315 19261 21327 19264
rect 21269 19255 21327 19261
rect 21358 19252 21364 19264
rect 21416 19252 21422 19304
rect 22097 19295 22155 19301
rect 22097 19292 22109 19295
rect 21928 19264 22109 19292
rect 21818 19184 21824 19236
rect 21876 19224 21882 19236
rect 21928 19224 21956 19264
rect 22097 19261 22109 19264
rect 22143 19261 22155 19295
rect 22097 19255 22155 19261
rect 23474 19252 23480 19304
rect 23532 19292 23538 19304
rect 23569 19295 23627 19301
rect 23569 19292 23581 19295
rect 23532 19264 23581 19292
rect 23532 19252 23538 19264
rect 23569 19261 23581 19264
rect 23615 19292 23627 19295
rect 24213 19295 24271 19301
rect 24213 19292 24225 19295
rect 23615 19264 24225 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 24213 19261 24225 19264
rect 24259 19261 24271 19295
rect 24213 19255 24271 19261
rect 26050 19252 26056 19304
rect 26108 19252 26114 19304
rect 26145 19295 26203 19301
rect 26145 19261 26157 19295
rect 26191 19261 26203 19295
rect 26145 19255 26203 19261
rect 27709 19295 27767 19301
rect 27709 19261 27721 19295
rect 27755 19292 27767 19295
rect 28166 19292 28172 19304
rect 27755 19264 28172 19292
rect 27755 19261 27767 19264
rect 27709 19255 27767 19261
rect 26160 19224 26188 19255
rect 28166 19252 28172 19264
rect 28224 19252 28230 19304
rect 29181 19295 29239 19301
rect 29181 19261 29193 19295
rect 29227 19292 29239 19295
rect 29730 19292 29736 19304
rect 29227 19264 29736 19292
rect 29227 19261 29239 19264
rect 29181 19255 29239 19261
rect 29730 19252 29736 19264
rect 29788 19292 29794 19304
rect 29825 19295 29883 19301
rect 29825 19292 29837 19295
rect 29788 19264 29837 19292
rect 29788 19252 29794 19264
rect 29825 19261 29837 19264
rect 29871 19261 29883 19295
rect 29825 19255 29883 19261
rect 30650 19252 30656 19304
rect 30708 19292 30714 19304
rect 30745 19295 30803 19301
rect 30745 19292 30757 19295
rect 30708 19264 30757 19292
rect 30708 19252 30714 19264
rect 30745 19261 30757 19264
rect 30791 19261 30803 19295
rect 30745 19255 30803 19261
rect 21876 19196 21956 19224
rect 26068 19196 26188 19224
rect 21876 19184 21882 19196
rect 15102 19156 15108 19168
rect 13136 19128 15108 19156
rect 13136 19116 13142 19128
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 22278 19116 22284 19168
rect 22336 19156 22342 19168
rect 23198 19156 23204 19168
rect 22336 19128 23204 19156
rect 22336 19116 22342 19128
rect 23198 19116 23204 19128
rect 23256 19156 23262 19168
rect 26068 19156 26096 19196
rect 32674 19184 32680 19236
rect 32732 19224 32738 19236
rect 32784 19224 32812 19323
rect 32858 19320 32864 19372
rect 32916 19320 32922 19372
rect 33229 19363 33287 19369
rect 33229 19329 33241 19363
rect 33275 19329 33287 19363
rect 33229 19323 33287 19329
rect 33244 19292 33272 19323
rect 33410 19320 33416 19372
rect 33468 19320 33474 19372
rect 33965 19363 34023 19369
rect 33965 19329 33977 19363
rect 34011 19329 34023 19363
rect 33965 19323 34023 19329
rect 33686 19292 33692 19304
rect 33244 19264 33692 19292
rect 33686 19252 33692 19264
rect 33744 19252 33750 19304
rect 33980 19292 34008 19323
rect 34054 19320 34060 19372
rect 34112 19360 34118 19372
rect 34149 19363 34207 19369
rect 34149 19360 34161 19363
rect 34112 19332 34161 19360
rect 34112 19320 34118 19332
rect 34149 19329 34161 19332
rect 34195 19329 34207 19363
rect 34149 19323 34207 19329
rect 34238 19320 34244 19372
rect 34296 19320 34302 19372
rect 34330 19320 34336 19372
rect 34388 19320 34394 19372
rect 34624 19369 34652 19400
rect 34808 19400 36768 19428
rect 34609 19363 34667 19369
rect 34609 19329 34621 19363
rect 34655 19329 34667 19363
rect 34808 19360 34836 19400
rect 36740 19372 36768 19400
rect 36924 19400 38568 19428
rect 34609 19323 34667 19329
rect 34716 19332 34836 19360
rect 34876 19363 34934 19369
rect 34716 19292 34744 19332
rect 34876 19329 34888 19363
rect 34922 19360 34934 19363
rect 35618 19360 35624 19372
rect 34922 19332 35624 19360
rect 34922 19329 34934 19332
rect 34876 19323 34934 19329
rect 35618 19320 35624 19332
rect 35676 19320 35682 19372
rect 36722 19320 36728 19372
rect 36780 19320 36786 19372
rect 36924 19369 36952 19400
rect 37476 19369 37504 19400
rect 38562 19388 38568 19400
rect 38620 19388 38626 19440
rect 39482 19388 39488 19440
rect 39540 19388 39546 19440
rect 40126 19388 40132 19440
rect 40184 19388 40190 19440
rect 36909 19363 36967 19369
rect 36909 19329 36921 19363
rect 36955 19329 36967 19363
rect 36909 19323 36967 19329
rect 37093 19363 37151 19369
rect 37093 19329 37105 19363
rect 37139 19360 37151 19363
rect 37277 19363 37335 19369
rect 37277 19360 37289 19363
rect 37139 19332 37289 19360
rect 37139 19329 37151 19332
rect 37093 19323 37151 19329
rect 37277 19329 37289 19332
rect 37323 19329 37335 19363
rect 37277 19323 37335 19329
rect 37461 19363 37519 19369
rect 37461 19329 37473 19363
rect 37507 19329 37519 19363
rect 37461 19323 37519 19329
rect 37645 19363 37703 19369
rect 37645 19329 37657 19363
rect 37691 19360 37703 19363
rect 37918 19360 37924 19372
rect 37691 19332 37924 19360
rect 37691 19329 37703 19332
rect 37645 19323 37703 19329
rect 33980 19264 34744 19292
rect 36081 19295 36139 19301
rect 36081 19261 36093 19295
rect 36127 19261 36139 19295
rect 37292 19292 37320 19323
rect 37918 19320 37924 19332
rect 37976 19320 37982 19372
rect 41690 19320 41696 19372
rect 41748 19360 41754 19372
rect 41785 19363 41843 19369
rect 41785 19360 41797 19363
rect 41748 19332 41797 19360
rect 41748 19320 41754 19332
rect 41785 19329 41797 19332
rect 41831 19329 41843 19363
rect 41785 19323 41843 19329
rect 37550 19292 37556 19304
rect 37292 19264 37556 19292
rect 36081 19255 36139 19261
rect 32732 19196 32812 19224
rect 32732 19184 32738 19196
rect 33502 19184 33508 19236
rect 33560 19224 33566 19236
rect 33560 19196 34652 19224
rect 33560 19184 33566 19196
rect 23256 19128 26096 19156
rect 23256 19116 23262 19128
rect 31478 19116 31484 19168
rect 31536 19156 31542 19168
rect 32585 19159 32643 19165
rect 32585 19156 32597 19159
rect 31536 19128 32597 19156
rect 31536 19116 31542 19128
rect 32585 19125 32597 19128
rect 32631 19125 32643 19159
rect 32585 19119 32643 19125
rect 34514 19116 34520 19168
rect 34572 19116 34578 19168
rect 34624 19156 34652 19196
rect 36096 19168 36124 19255
rect 37550 19252 37556 19264
rect 37608 19292 37614 19304
rect 39025 19295 39083 19301
rect 39025 19292 39037 19295
rect 37608 19264 39037 19292
rect 37608 19252 37614 19264
rect 39025 19261 39037 19264
rect 39071 19261 39083 19295
rect 39025 19255 39083 19261
rect 39206 19252 39212 19304
rect 39264 19252 39270 19304
rect 40126 19252 40132 19304
rect 40184 19292 40190 19304
rect 40184 19264 40540 19292
rect 40184 19252 40190 19264
rect 40512 19224 40540 19264
rect 41598 19252 41604 19304
rect 41656 19252 41662 19304
rect 41414 19224 41420 19236
rect 40512 19196 41420 19224
rect 41414 19184 41420 19196
rect 41472 19224 41478 19236
rect 41969 19227 42027 19233
rect 41969 19224 41981 19227
rect 41472 19196 41981 19224
rect 41472 19184 41478 19196
rect 41969 19193 41981 19196
rect 42015 19193 42027 19227
rect 41969 19187 42027 19193
rect 34882 19156 34888 19168
rect 34624 19128 34888 19156
rect 34882 19116 34888 19128
rect 34940 19116 34946 19168
rect 35989 19159 36047 19165
rect 35989 19125 36001 19159
rect 36035 19156 36047 19159
rect 36078 19156 36084 19168
rect 36035 19128 36084 19156
rect 36035 19125 36047 19128
rect 35989 19119 36047 19125
rect 36078 19116 36084 19128
rect 36136 19116 36142 19168
rect 37001 19159 37059 19165
rect 37001 19125 37013 19159
rect 37047 19156 37059 19159
rect 37182 19156 37188 19168
rect 37047 19128 37188 19156
rect 37047 19125 37059 19128
rect 37001 19119 37059 19125
rect 37182 19116 37188 19128
rect 37240 19116 37246 19168
rect 37274 19116 37280 19168
rect 37332 19156 37338 19168
rect 37461 19159 37519 19165
rect 37461 19156 37473 19159
rect 37332 19128 37473 19156
rect 37332 19116 37338 19128
rect 37461 19125 37473 19128
rect 37507 19156 37519 19159
rect 37918 19156 37924 19168
rect 37507 19128 37924 19156
rect 37507 19125 37519 19128
rect 37461 19119 37519 19125
rect 37918 19116 37924 19128
rect 37976 19116 37982 19168
rect 38194 19116 38200 19168
rect 38252 19116 38258 19168
rect 41046 19116 41052 19168
rect 41104 19116 41110 19168
rect 1104 19066 42504 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 42504 19066
rect 1104 18992 42504 19014
rect 3191 18955 3249 18961
rect 3191 18921 3203 18955
rect 3237 18952 3249 18955
rect 3602 18952 3608 18964
rect 3237 18924 3608 18952
rect 3237 18921 3249 18924
rect 3191 18915 3249 18921
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 4798 18912 4804 18964
rect 4856 18912 4862 18964
rect 4908 18924 5488 18952
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 2314 18816 2320 18828
rect 1452 18788 2320 18816
rect 1452 18776 1458 18788
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 3973 18819 4031 18825
rect 3973 18785 3985 18819
rect 4019 18816 4031 18819
rect 4614 18816 4620 18828
rect 4019 18788 4620 18816
rect 4019 18785 4031 18788
rect 3973 18779 4031 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 1762 18708 1768 18760
rect 1820 18708 1826 18760
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4908 18748 4936 18924
rect 5074 18844 5080 18896
rect 5132 18844 5138 18896
rect 5258 18844 5264 18896
rect 5316 18884 5322 18896
rect 5316 18856 5396 18884
rect 5316 18844 5322 18856
rect 4755 18720 4936 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4982 18708 4988 18760
rect 5040 18708 5046 18760
rect 5166 18708 5172 18760
rect 5224 18708 5230 18760
rect 5258 18708 5264 18760
rect 5316 18708 5322 18760
rect 5368 18748 5396 18856
rect 5460 18816 5488 18924
rect 6270 18912 6276 18964
rect 6328 18952 6334 18964
rect 6549 18955 6607 18961
rect 6549 18952 6561 18955
rect 6328 18924 6561 18952
rect 6328 18912 6334 18924
rect 6549 18921 6561 18924
rect 6595 18921 6607 18955
rect 6549 18915 6607 18921
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 6696 18924 6745 18952
rect 6696 18912 6702 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 9766 18952 9772 18964
rect 6733 18915 6791 18921
rect 6840 18924 9772 18952
rect 6178 18844 6184 18896
rect 6236 18844 6242 18896
rect 6840 18884 6868 18924
rect 9766 18912 9772 18924
rect 9824 18952 9830 18964
rect 10134 18952 10140 18964
rect 9824 18924 10140 18952
rect 9824 18912 9830 18924
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 10318 18912 10324 18964
rect 10376 18912 10382 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11333 18955 11391 18961
rect 11333 18952 11345 18955
rect 11204 18924 11345 18952
rect 11204 18912 11210 18924
rect 11333 18921 11345 18924
rect 11379 18921 11391 18955
rect 11333 18915 11391 18921
rect 11698 18912 11704 18964
rect 11756 18912 11762 18964
rect 11882 18912 11888 18964
rect 11940 18912 11946 18964
rect 12158 18912 12164 18964
rect 12216 18912 12222 18964
rect 12805 18955 12863 18961
rect 12805 18921 12817 18955
rect 12851 18952 12863 18955
rect 13814 18952 13820 18964
rect 12851 18924 13820 18952
rect 12851 18921 12863 18924
rect 12805 18915 12863 18921
rect 6288 18856 6868 18884
rect 8588 18856 11008 18884
rect 6288 18816 6316 18856
rect 5460 18788 6316 18816
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 5368 18720 5457 18748
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 5537 18751 5595 18757
rect 5537 18717 5549 18751
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 5629 18751 5687 18757
rect 5629 18717 5641 18751
rect 5675 18748 5687 18751
rect 5718 18748 5724 18760
rect 5675 18720 5724 18748
rect 5675 18717 5687 18720
rect 5629 18711 5687 18717
rect 3694 18680 3700 18692
rect 2806 18652 3700 18680
rect 3694 18640 3700 18652
rect 3752 18640 3758 18692
rect 4246 18640 4252 18692
rect 4304 18680 4310 18692
rect 5552 18680 5580 18711
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 8588 18748 8616 18856
rect 10980 18828 11008 18856
rect 11238 18844 11244 18896
rect 11296 18884 11302 18896
rect 11716 18884 11744 18912
rect 12434 18884 12440 18896
rect 11296 18856 12440 18884
rect 11296 18844 11302 18856
rect 12434 18844 12440 18856
rect 12492 18844 12498 18896
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 8720 18788 9229 18816
rect 8720 18776 8726 18788
rect 9217 18785 9229 18788
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 6564 18720 8616 18748
rect 8680 18720 8953 18748
rect 6564 18689 6592 18720
rect 4304 18652 5580 18680
rect 6549 18683 6607 18689
rect 4304 18640 4310 18652
rect 6549 18649 6561 18683
rect 6595 18649 6607 18683
rect 6549 18643 6607 18649
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 8680 18680 8708 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 8352 18652 8708 18680
rect 8352 18640 8358 18652
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 5166 18612 5172 18624
rect 4764 18584 5172 18612
rect 4764 18572 4770 18584
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 5997 18615 6055 18621
rect 5997 18612 6009 18615
rect 5684 18584 6009 18612
rect 5684 18572 5690 18584
rect 5997 18581 6009 18584
rect 6043 18581 6055 18615
rect 5997 18575 6055 18581
rect 8018 18572 8024 18624
rect 8076 18612 8082 18624
rect 9140 18612 9168 18711
rect 8076 18584 9168 18612
rect 9232 18612 9260 18779
rect 9674 18776 9680 18828
rect 9732 18776 9738 18828
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10376 18788 10916 18816
rect 10376 18776 10382 18788
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9582 18748 9588 18760
rect 9539 18720 9588 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9324 18680 9352 18711
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9950 18748 9956 18760
rect 9784 18720 9956 18748
rect 9674 18680 9680 18692
rect 9324 18652 9680 18680
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 9784 18689 9812 18720
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 10686 18708 10692 18760
rect 10744 18708 10750 18760
rect 10888 18757 10916 18788
rect 10962 18776 10968 18828
rect 11020 18816 11026 18828
rect 12820 18816 12848 18915
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 15378 18912 15384 18964
rect 15436 18912 15442 18964
rect 16942 18912 16948 18964
rect 17000 18952 17006 18964
rect 17221 18955 17279 18961
rect 17221 18952 17233 18955
rect 17000 18924 17233 18952
rect 17000 18912 17006 18924
rect 17221 18921 17233 18924
rect 17267 18921 17279 18955
rect 17221 18915 17279 18921
rect 20254 18912 20260 18964
rect 20312 18912 20318 18964
rect 23106 18912 23112 18964
rect 23164 18952 23170 18964
rect 23750 18952 23756 18964
rect 23164 18924 23756 18952
rect 23164 18912 23170 18924
rect 23750 18912 23756 18924
rect 23808 18912 23814 18964
rect 28166 18912 28172 18964
rect 28224 18912 28230 18964
rect 35437 18955 35495 18961
rect 35437 18921 35449 18955
rect 35483 18952 35495 18955
rect 35618 18952 35624 18964
rect 35483 18924 35624 18952
rect 35483 18921 35495 18924
rect 35437 18915 35495 18921
rect 35618 18912 35624 18924
rect 35676 18912 35682 18964
rect 37369 18955 37427 18961
rect 37369 18921 37381 18955
rect 37415 18952 37427 18955
rect 41782 18952 41788 18964
rect 37415 18924 39160 18952
rect 37415 18921 37427 18924
rect 37369 18915 37427 18921
rect 22278 18884 22284 18896
rect 20824 18856 22284 18884
rect 16298 18816 16304 18828
rect 11020 18788 12848 18816
rect 15580 18788 16304 18816
rect 11020 18776 11026 18788
rect 10873 18751 10931 18757
rect 10873 18717 10885 18751
rect 10919 18717 10931 18751
rect 10873 18711 10931 18717
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18748 11207 18751
rect 11238 18748 11244 18760
rect 11195 18720 11244 18748
rect 11195 18717 11207 18720
rect 11149 18711 11207 18717
rect 9769 18683 9827 18689
rect 9769 18649 9781 18683
rect 9815 18649 9827 18683
rect 10888 18680 10916 18711
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 11517 18683 11575 18689
rect 10888 18652 11100 18680
rect 9769 18643 9827 18649
rect 9582 18612 9588 18624
rect 9232 18584 9588 18612
rect 8076 18572 8082 18584
rect 9582 18572 9588 18584
rect 9640 18612 9646 18624
rect 9953 18615 10011 18621
rect 9953 18612 9965 18615
rect 9640 18584 9965 18612
rect 9640 18572 9646 18584
rect 9953 18581 9965 18584
rect 9999 18581 10011 18615
rect 9953 18575 10011 18581
rect 10042 18572 10048 18624
rect 10100 18572 10106 18624
rect 10134 18572 10140 18624
rect 10192 18572 10198 18624
rect 10962 18572 10968 18624
rect 11020 18572 11026 18624
rect 11072 18612 11100 18652
rect 11517 18649 11529 18683
rect 11563 18680 11575 18683
rect 11606 18680 11612 18692
rect 11563 18652 11612 18680
rect 11563 18649 11575 18652
rect 11517 18643 11575 18649
rect 11606 18640 11612 18652
rect 11664 18640 11670 18692
rect 12066 18640 12072 18692
rect 12124 18689 12130 18692
rect 12360 18689 12388 18788
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 12621 18751 12679 18757
rect 12621 18748 12633 18751
rect 12584 18720 12633 18748
rect 12584 18708 12590 18720
rect 12621 18717 12633 18720
rect 12667 18717 12679 18751
rect 12621 18711 12679 18717
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 15580 18757 15608 18788
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 16942 18776 16948 18828
rect 17000 18816 17006 18828
rect 17494 18816 17500 18828
rect 17000 18788 17500 18816
rect 17000 18776 17006 18788
rect 17494 18776 17500 18788
rect 17552 18816 17558 18828
rect 20824 18825 20852 18856
rect 22278 18844 22284 18856
rect 22336 18844 22342 18896
rect 30558 18884 30564 18896
rect 29380 18856 30564 18884
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17552 18788 17785 18816
rect 17552 18776 17558 18788
rect 17773 18785 17785 18788
rect 17819 18816 17831 18819
rect 20809 18819 20867 18825
rect 20809 18816 20821 18819
rect 17819 18788 20821 18816
rect 17819 18785 17831 18788
rect 17773 18779 17831 18785
rect 20809 18785 20821 18788
rect 20855 18785 20867 18819
rect 20809 18779 20867 18785
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24949 18819 25007 18825
rect 24949 18816 24961 18819
rect 24176 18788 24961 18816
rect 24176 18776 24182 18788
rect 24949 18785 24961 18788
rect 24995 18785 25007 18819
rect 24949 18779 25007 18785
rect 25130 18776 25136 18828
rect 25188 18816 25194 18828
rect 28813 18819 28871 18825
rect 25188 18788 28580 18816
rect 25188 18776 25194 18788
rect 28552 18760 28580 18788
rect 28813 18785 28825 18819
rect 28859 18816 28871 18819
rect 29270 18816 29276 18828
rect 28859 18788 29276 18816
rect 28859 18785 28871 18788
rect 28813 18779 28871 18785
rect 29270 18776 29276 18788
rect 29328 18776 29334 18828
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14608 18720 14657 18748
rect 14608 18708 14614 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 15565 18751 15623 18757
rect 15565 18717 15577 18751
rect 15611 18717 15623 18751
rect 15565 18711 15623 18717
rect 15746 18708 15752 18760
rect 15804 18708 15810 18760
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 18414 18748 18420 18760
rect 17635 18720 18420 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 12124 18683 12187 18689
rect 12124 18649 12141 18683
rect 12175 18649 12187 18683
rect 12124 18643 12187 18649
rect 12345 18683 12403 18689
rect 12345 18649 12357 18683
rect 12391 18649 12403 18683
rect 12345 18643 12403 18649
rect 12437 18683 12495 18689
rect 12437 18649 12449 18683
rect 12483 18649 12495 18683
rect 15856 18680 15884 18711
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 21266 18708 21272 18760
rect 21324 18708 21330 18760
rect 22373 18751 22431 18757
rect 22373 18717 22385 18751
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 17862 18680 17868 18692
rect 15856 18652 17868 18680
rect 12437 18643 12495 18649
rect 12124 18640 12130 18643
rect 11717 18615 11775 18621
rect 11717 18612 11729 18615
rect 11072 18584 11729 18612
rect 11717 18581 11729 18584
rect 11763 18581 11775 18615
rect 11717 18575 11775 18581
rect 11974 18572 11980 18624
rect 12032 18572 12038 18624
rect 12250 18572 12256 18624
rect 12308 18612 12314 18624
rect 12452 18612 12480 18643
rect 17862 18640 17868 18652
rect 17920 18640 17926 18692
rect 20530 18640 20536 18692
rect 20588 18680 20594 18692
rect 20717 18683 20775 18689
rect 20717 18680 20729 18683
rect 20588 18652 20729 18680
rect 20588 18640 20594 18652
rect 20717 18649 20729 18652
rect 20763 18649 20775 18683
rect 20717 18643 20775 18649
rect 22094 18640 22100 18692
rect 22152 18680 22158 18692
rect 22388 18680 22416 18711
rect 28350 18708 28356 18760
rect 28408 18708 28414 18760
rect 28534 18708 28540 18760
rect 28592 18708 28598 18760
rect 28718 18757 28724 18760
rect 28675 18751 28724 18757
rect 28675 18717 28687 18751
rect 28721 18717 28724 18751
rect 28675 18711 28724 18717
rect 28718 18708 28724 18711
rect 28776 18708 28782 18760
rect 29380 18757 29408 18856
rect 30558 18844 30564 18856
rect 30616 18844 30622 18896
rect 32401 18887 32459 18893
rect 32401 18853 32413 18887
rect 32447 18884 32459 18887
rect 36633 18887 36691 18893
rect 32447 18856 33088 18884
rect 32447 18853 32459 18856
rect 32401 18847 32459 18853
rect 30374 18776 30380 18828
rect 30432 18816 30438 18828
rect 30653 18819 30711 18825
rect 30653 18816 30665 18819
rect 30432 18788 30665 18816
rect 30432 18776 30438 18788
rect 30653 18785 30665 18788
rect 30699 18816 30711 18819
rect 32766 18816 32772 18828
rect 30699 18788 32772 18816
rect 30699 18785 30711 18788
rect 30653 18779 30711 18785
rect 32766 18776 32772 18788
rect 32824 18776 32830 18828
rect 33060 18825 33088 18856
rect 36633 18853 36645 18887
rect 36679 18884 36691 18887
rect 37642 18884 37648 18896
rect 36679 18856 37648 18884
rect 36679 18853 36691 18856
rect 36633 18847 36691 18853
rect 37642 18844 37648 18856
rect 37700 18844 37706 18896
rect 39132 18884 39160 18924
rect 40236 18924 41788 18952
rect 39758 18884 39764 18896
rect 39132 18856 39764 18884
rect 39758 18844 39764 18856
rect 39816 18884 39822 18896
rect 40129 18887 40187 18893
rect 40129 18884 40141 18887
rect 39816 18856 40141 18884
rect 39816 18844 39822 18856
rect 40129 18853 40141 18856
rect 40175 18853 40187 18887
rect 40129 18847 40187 18853
rect 33045 18819 33103 18825
rect 33045 18785 33057 18819
rect 33091 18785 33103 18819
rect 33045 18779 33103 18785
rect 34514 18776 34520 18828
rect 34572 18816 34578 18828
rect 34793 18819 34851 18825
rect 34793 18816 34805 18819
rect 34572 18788 34805 18816
rect 34572 18776 34578 18788
rect 34793 18785 34805 18788
rect 34839 18785 34851 18819
rect 34793 18779 34851 18785
rect 36170 18776 36176 18828
rect 36228 18816 36234 18828
rect 36909 18819 36967 18825
rect 36228 18788 36492 18816
rect 36228 18776 36234 18788
rect 29181 18751 29239 18757
rect 29181 18717 29193 18751
rect 29227 18717 29239 18751
rect 29181 18711 29239 18717
rect 29365 18751 29423 18757
rect 29365 18717 29377 18751
rect 29411 18717 29423 18751
rect 29365 18711 29423 18717
rect 22152 18652 22416 18680
rect 22152 18640 22158 18652
rect 22554 18640 22560 18692
rect 22612 18680 22618 18692
rect 22649 18683 22707 18689
rect 22649 18680 22661 18683
rect 22612 18652 22661 18680
rect 22612 18640 22618 18652
rect 22649 18649 22661 18652
rect 22695 18649 22707 18683
rect 22649 18643 22707 18649
rect 23106 18640 23112 18692
rect 23164 18640 23170 18692
rect 24397 18683 24455 18689
rect 24397 18680 24409 18683
rect 23952 18652 24409 18680
rect 12308 18584 12480 18612
rect 12308 18572 12314 18584
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 13228 18584 14105 18612
rect 13228 18572 13234 18584
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 18874 18612 18880 18624
rect 17727 18584 18880 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 18874 18572 18880 18584
rect 18932 18572 18938 18624
rect 20625 18615 20683 18621
rect 20625 18581 20637 18615
rect 20671 18612 20683 18615
rect 21358 18612 21364 18624
rect 20671 18584 21364 18612
rect 20671 18581 20683 18584
rect 20625 18575 20683 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 23952 18612 23980 18652
rect 24397 18649 24409 18652
rect 24443 18649 24455 18683
rect 24397 18643 24455 18649
rect 28442 18640 28448 18692
rect 28500 18640 28506 18692
rect 29196 18680 29224 18711
rect 29546 18708 29552 18760
rect 29604 18708 29610 18760
rect 33686 18708 33692 18760
rect 33744 18748 33750 18760
rect 33965 18751 34023 18757
rect 33965 18748 33977 18751
rect 33744 18720 33977 18748
rect 33744 18708 33750 18720
rect 33965 18717 33977 18720
rect 34011 18717 34023 18751
rect 33965 18711 34023 18717
rect 36265 18751 36323 18757
rect 36265 18717 36277 18751
rect 36311 18717 36323 18751
rect 36464 18748 36492 18788
rect 36909 18785 36921 18819
rect 36955 18816 36967 18819
rect 37274 18816 37280 18828
rect 36955 18788 37280 18816
rect 36955 18785 36967 18788
rect 36909 18779 36967 18785
rect 37274 18776 37280 18788
rect 37332 18776 37338 18828
rect 37461 18819 37519 18825
rect 37461 18785 37473 18819
rect 37507 18816 37519 18819
rect 37550 18816 37556 18828
rect 37507 18788 37556 18816
rect 37507 18785 37519 18788
rect 37461 18779 37519 18785
rect 37550 18776 37556 18788
rect 37608 18776 37614 18828
rect 38194 18776 38200 18828
rect 38252 18816 38258 18828
rect 38933 18819 38991 18825
rect 38933 18816 38945 18819
rect 38252 18788 38945 18816
rect 38252 18776 38258 18788
rect 38933 18785 38945 18788
rect 38979 18785 38991 18819
rect 40236 18816 40264 18924
rect 41782 18912 41788 18924
rect 41840 18912 41846 18964
rect 42150 18912 42156 18964
rect 42208 18912 42214 18964
rect 38933 18779 38991 18785
rect 40052 18788 40264 18816
rect 37001 18751 37059 18757
rect 37001 18748 37013 18751
rect 36464 18720 37013 18748
rect 36265 18711 36323 18717
rect 37001 18717 37013 18720
rect 37047 18717 37059 18751
rect 37001 18711 37059 18717
rect 30650 18680 30656 18692
rect 28736 18652 30656 18680
rect 23716 18584 23980 18612
rect 23716 18572 23722 18584
rect 28626 18572 28632 18624
rect 28684 18612 28690 18624
rect 28736 18612 28764 18652
rect 30650 18640 30656 18652
rect 30708 18640 30714 18692
rect 30929 18683 30987 18689
rect 30929 18649 30941 18683
rect 30975 18680 30987 18683
rect 31202 18680 31208 18692
rect 30975 18652 31208 18680
rect 30975 18649 30987 18652
rect 30929 18643 30987 18649
rect 31202 18640 31208 18652
rect 31260 18640 31266 18692
rect 36280 18680 36308 18711
rect 37182 18708 37188 18760
rect 37240 18708 37246 18760
rect 39206 18708 39212 18760
rect 39264 18708 39270 18760
rect 40052 18757 40080 18788
rect 40310 18776 40316 18828
rect 40368 18776 40374 18828
rect 40681 18819 40739 18825
rect 40681 18785 40693 18819
rect 40727 18816 40739 18819
rect 41046 18816 41052 18828
rect 40727 18788 41052 18816
rect 40727 18785 40739 18788
rect 40681 18779 40739 18785
rect 41046 18776 41052 18788
rect 41104 18776 41110 18828
rect 40037 18751 40095 18757
rect 40037 18717 40049 18751
rect 40083 18717 40095 18751
rect 40037 18711 40095 18717
rect 40405 18751 40463 18757
rect 40405 18717 40417 18751
rect 40451 18717 40463 18751
rect 40405 18711 40463 18717
rect 37550 18680 37556 18692
rect 31312 18652 31418 18680
rect 36280 18652 37556 18680
rect 28684 18584 28764 18612
rect 28684 18572 28690 18584
rect 29178 18572 29184 18624
rect 29236 18572 29242 18624
rect 30098 18572 30104 18624
rect 30156 18612 30162 18624
rect 30193 18615 30251 18621
rect 30193 18612 30205 18615
rect 30156 18584 30205 18612
rect 30156 18572 30162 18584
rect 30193 18581 30205 18584
rect 30239 18581 30251 18615
rect 30193 18575 30251 18581
rect 30466 18572 30472 18624
rect 30524 18612 30530 18624
rect 31018 18612 31024 18624
rect 30524 18584 31024 18612
rect 30524 18572 30530 18584
rect 31018 18572 31024 18584
rect 31076 18612 31082 18624
rect 31312 18612 31340 18652
rect 37550 18640 37556 18652
rect 37608 18640 37614 18692
rect 39224 18680 39252 18708
rect 40420 18680 40448 18711
rect 37660 18652 37766 18680
rect 39224 18652 40448 18680
rect 31076 18584 31340 18612
rect 31076 18572 31082 18584
rect 31662 18572 31668 18624
rect 31720 18612 31726 18624
rect 32490 18612 32496 18624
rect 31720 18584 32496 18612
rect 31720 18572 31726 18584
rect 32490 18572 32496 18584
rect 32548 18572 32554 18624
rect 32582 18572 32588 18624
rect 32640 18612 32646 18624
rect 33413 18615 33471 18621
rect 33413 18612 33425 18615
rect 32640 18584 33425 18612
rect 32640 18572 32646 18584
rect 33413 18581 33425 18584
rect 33459 18581 33471 18615
rect 33413 18575 33471 18581
rect 34054 18572 34060 18624
rect 34112 18612 34118 18624
rect 35526 18612 35532 18624
rect 34112 18584 35532 18612
rect 34112 18572 34118 18584
rect 35526 18572 35532 18584
rect 35584 18572 35590 18624
rect 37458 18572 37464 18624
rect 37516 18612 37522 18624
rect 37660 18612 37688 18652
rect 41414 18640 41420 18692
rect 41472 18640 41478 18692
rect 40126 18612 40132 18624
rect 37516 18584 40132 18612
rect 37516 18572 37522 18584
rect 40126 18572 40132 18584
rect 40184 18572 40190 18624
rect 40310 18572 40316 18624
rect 40368 18572 40374 18624
rect 1104 18522 42504 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 42504 18522
rect 1104 18448 42504 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 1762 18408 1768 18420
rect 1627 18380 1768 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 4246 18368 4252 18420
rect 4304 18368 4310 18420
rect 4614 18408 4620 18420
rect 4448 18380 4620 18408
rect 3602 18300 3608 18352
rect 3660 18300 3666 18352
rect 4448 18349 4476 18380
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 5258 18368 5264 18420
rect 5316 18368 5322 18420
rect 9953 18411 10011 18417
rect 9953 18377 9965 18411
rect 9999 18408 10011 18411
rect 10042 18408 10048 18420
rect 9999 18380 10048 18408
rect 9999 18377 10011 18380
rect 9953 18371 10011 18377
rect 4433 18343 4491 18349
rect 4433 18309 4445 18343
rect 4479 18309 4491 18343
rect 4433 18303 4491 18309
rect 4798 18300 4804 18352
rect 4856 18300 4862 18352
rect 4893 18343 4951 18349
rect 4893 18309 4905 18343
rect 4939 18340 4951 18343
rect 5718 18340 5724 18352
rect 4939 18312 5724 18340
rect 4939 18309 4951 18312
rect 4893 18303 4951 18309
rect 5718 18300 5724 18312
rect 5776 18340 5782 18352
rect 5902 18340 5908 18352
rect 5776 18312 5908 18340
rect 5776 18300 5782 18312
rect 5902 18300 5908 18312
rect 5960 18300 5966 18352
rect 1397 18275 1455 18281
rect 1397 18241 1409 18275
rect 1443 18272 1455 18275
rect 1486 18272 1492 18284
rect 1443 18244 1492 18272
rect 1443 18241 1455 18244
rect 1397 18235 1455 18241
rect 1486 18232 1492 18244
rect 1544 18232 1550 18284
rect 4019 18275 4077 18281
rect 4019 18241 4031 18275
rect 4065 18272 4077 18275
rect 4157 18275 4215 18281
rect 4157 18272 4169 18275
rect 4065 18244 4169 18272
rect 4065 18241 4077 18244
rect 4019 18235 4077 18241
rect 4157 18241 4169 18244
rect 4203 18272 4215 18275
rect 4614 18272 4620 18284
rect 4203 18244 4620 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 4985 18235 5043 18241
rect 5184 18244 5641 18272
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2406 18204 2412 18216
rect 2271 18176 2412 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2406 18164 2412 18176
rect 2464 18164 2470 18216
rect 2593 18207 2651 18213
rect 2593 18173 2605 18207
rect 2639 18204 2651 18207
rect 3786 18204 3792 18216
rect 2639 18176 3792 18204
rect 2639 18173 2651 18176
rect 2593 18167 2651 18173
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 4798 18164 4804 18216
rect 4856 18204 4862 18216
rect 5000 18204 5028 18235
rect 5184 18216 5212 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 6178 18232 6184 18284
rect 6236 18272 6242 18284
rect 7745 18275 7803 18281
rect 7745 18272 7757 18275
rect 6236 18244 7757 18272
rect 6236 18232 6242 18244
rect 7745 18241 7757 18244
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 7834 18232 7840 18284
rect 7892 18232 7898 18284
rect 7929 18275 7987 18281
rect 7929 18241 7941 18275
rect 7975 18272 7987 18275
rect 8294 18272 8300 18284
rect 7975 18244 8300 18272
rect 7975 18241 7987 18244
rect 7929 18235 7987 18241
rect 8294 18232 8300 18244
rect 8352 18272 8358 18284
rect 8754 18272 8760 18284
rect 8352 18244 8760 18272
rect 8352 18232 8358 18244
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 9309 18275 9367 18281
rect 9309 18241 9321 18275
rect 9355 18241 9367 18275
rect 9309 18235 9367 18241
rect 4856 18176 5028 18204
rect 4856 18164 4862 18176
rect 5166 18164 5172 18216
rect 5224 18164 5230 18216
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5445 18207 5503 18213
rect 5445 18204 5457 18207
rect 5316 18176 5457 18204
rect 5316 18164 5322 18176
rect 5445 18173 5457 18176
rect 5491 18173 5503 18207
rect 5445 18167 5503 18173
rect 5534 18164 5540 18216
rect 5592 18164 5598 18216
rect 5718 18164 5724 18216
rect 5776 18164 5782 18216
rect 9324 18204 9352 18235
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9640 18244 9689 18272
rect 9640 18232 9646 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18272 9827 18275
rect 9858 18272 9864 18284
rect 9815 18244 9864 18272
rect 9815 18241 9827 18244
rect 9769 18235 9827 18241
rect 9858 18232 9864 18244
rect 9916 18272 9922 18284
rect 9968 18272 9996 18371
rect 10042 18368 10048 18380
rect 10100 18408 10106 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 10100 18380 11805 18408
rect 10100 18368 10106 18380
rect 11793 18377 11805 18380
rect 11839 18377 11851 18411
rect 11793 18371 11851 18377
rect 11885 18411 11943 18417
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 12342 18408 12348 18420
rect 11931 18380 12348 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 12342 18368 12348 18380
rect 12400 18408 12406 18420
rect 14090 18408 14096 18420
rect 12400 18380 14096 18408
rect 12400 18368 12406 18380
rect 14090 18368 14096 18380
rect 14148 18368 14154 18420
rect 15102 18368 15108 18420
rect 15160 18408 15166 18420
rect 15160 18380 15424 18408
rect 15160 18368 15166 18380
rect 11088 18343 11146 18349
rect 11088 18309 11100 18343
rect 11134 18340 11146 18343
rect 11974 18340 11980 18352
rect 11134 18312 11980 18340
rect 11134 18309 11146 18312
rect 11088 18303 11146 18309
rect 11974 18300 11980 18312
rect 12032 18300 12038 18352
rect 15194 18340 15200 18352
rect 13648 18312 15200 18340
rect 9916 18244 9996 18272
rect 9916 18232 9922 18244
rect 10502 18232 10508 18284
rect 10560 18272 10566 18284
rect 12250 18272 12256 18284
rect 10560 18244 12256 18272
rect 10560 18232 10566 18244
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 13170 18232 13176 18284
rect 13228 18232 13234 18284
rect 13648 18281 13676 18312
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18241 13691 18275
rect 13889 18275 13947 18281
rect 13889 18272 13901 18275
rect 13633 18235 13691 18241
rect 13740 18244 13901 18272
rect 9398 18204 9404 18216
rect 9324 18176 9404 18204
rect 9398 18164 9404 18176
rect 9456 18204 9462 18216
rect 9950 18204 9956 18216
rect 9456 18176 9956 18204
rect 9456 18164 9462 18176
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 11333 18207 11391 18213
rect 11333 18173 11345 18207
rect 11379 18204 11391 18207
rect 11422 18204 11428 18216
rect 11379 18176 11428 18204
rect 11379 18173 11391 18176
rect 11333 18167 11391 18173
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 11517 18207 11575 18213
rect 11517 18173 11529 18207
rect 11563 18204 11575 18207
rect 11606 18204 11612 18216
rect 11563 18176 11612 18204
rect 11563 18173 11575 18176
rect 11517 18167 11575 18173
rect 7650 18096 7656 18148
rect 7708 18136 7714 18148
rect 8113 18139 8171 18145
rect 8113 18136 8125 18139
rect 7708 18108 8125 18136
rect 7708 18096 7714 18108
rect 8113 18105 8125 18108
rect 8159 18105 8171 18139
rect 10134 18136 10140 18148
rect 8113 18099 8171 18105
rect 9048 18108 10140 18136
rect 7282 18028 7288 18080
rect 7340 18068 7346 18080
rect 7561 18071 7619 18077
rect 7561 18068 7573 18071
rect 7340 18040 7573 18068
rect 7340 18028 7346 18040
rect 7561 18037 7573 18040
rect 7607 18068 7619 18071
rect 8018 18068 8024 18080
rect 7607 18040 8024 18068
rect 7607 18037 7619 18040
rect 7561 18031 7619 18037
rect 8018 18028 8024 18040
rect 8076 18068 8082 18080
rect 9048 18068 9076 18108
rect 10134 18096 10140 18108
rect 10192 18096 10198 18148
rect 8076 18040 9076 18068
rect 8076 18028 8082 18040
rect 9122 18028 9128 18080
rect 9180 18028 9186 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 11054 18068 11060 18080
rect 9447 18040 11060 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 11054 18028 11060 18040
rect 11112 18068 11118 18080
rect 11532 18068 11560 18167
rect 11606 18164 11612 18176
rect 11664 18164 11670 18216
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 12002 18207 12060 18213
rect 12002 18204 12014 18207
rect 11756 18176 12014 18204
rect 11756 18164 11762 18176
rect 12002 18173 12014 18176
rect 12048 18173 12060 18207
rect 12002 18167 12060 18173
rect 13078 18164 13084 18216
rect 13136 18164 13142 18216
rect 13541 18207 13599 18213
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 13740 18204 13768 18244
rect 13889 18241 13901 18244
rect 13935 18241 13947 18275
rect 13889 18235 13947 18241
rect 15102 18232 15108 18284
rect 15160 18232 15166 18284
rect 15396 18281 15424 18380
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 21358 18408 21364 18420
rect 19208 18380 21364 18408
rect 19208 18368 19214 18380
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 21818 18368 21824 18420
rect 21876 18368 21882 18420
rect 22094 18368 22100 18420
rect 22152 18368 22158 18420
rect 22554 18368 22560 18420
rect 22612 18368 22618 18420
rect 27154 18368 27160 18420
rect 27212 18368 27218 18420
rect 28442 18368 28448 18420
rect 28500 18368 28506 18420
rect 28626 18368 28632 18420
rect 28684 18368 28690 18420
rect 29178 18408 29184 18420
rect 28736 18380 29184 18408
rect 18601 18343 18659 18349
rect 18601 18309 18613 18343
rect 18647 18340 18659 18343
rect 19061 18343 19119 18349
rect 19061 18340 19073 18343
rect 18647 18312 19073 18340
rect 18647 18309 18659 18312
rect 18601 18303 18659 18309
rect 19061 18309 19073 18312
rect 19107 18309 19119 18343
rect 19061 18303 19119 18309
rect 19334 18300 19340 18352
rect 19392 18340 19398 18352
rect 22112 18340 22140 18368
rect 24581 18343 24639 18349
rect 19392 18312 19748 18340
rect 19392 18300 19398 18312
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15304 18204 15332 18235
rect 18874 18232 18880 18284
rect 18932 18232 18938 18284
rect 18966 18232 18972 18284
rect 19024 18232 19030 18284
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18272 19303 18275
rect 19426 18272 19432 18284
rect 19291 18244 19432 18272
rect 19291 18241 19303 18244
rect 19245 18235 19303 18241
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 19610 18232 19616 18284
rect 19668 18232 19674 18284
rect 19720 18281 19748 18312
rect 21468 18312 24348 18340
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 19886 18232 19892 18284
rect 19944 18232 19950 18284
rect 20714 18232 20720 18284
rect 20772 18272 20778 18284
rect 21468 18281 21496 18312
rect 21453 18275 21511 18281
rect 21453 18272 21465 18275
rect 20772 18244 21465 18272
rect 20772 18232 20778 18244
rect 21453 18241 21465 18244
rect 21499 18241 21511 18275
rect 21453 18235 21511 18241
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 13587 18176 13768 18204
rect 15028 18176 15332 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 11112 18040 11560 18068
rect 12161 18071 12219 18077
rect 11112 18028 11118 18040
rect 12161 18037 12173 18071
rect 12207 18068 12219 18071
rect 12894 18068 12900 18080
rect 12207 18040 12900 18068
rect 12207 18037 12219 18040
rect 12161 18031 12219 18037
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 15028 18077 15056 18176
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 17313 18207 17371 18213
rect 17313 18204 17325 18207
rect 16632 18176 17325 18204
rect 16632 18164 16638 18176
rect 17313 18173 17325 18176
rect 17359 18204 17371 18207
rect 17954 18204 17960 18216
rect 17359 18176 17960 18204
rect 17359 18173 17371 18176
rect 17313 18167 17371 18173
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18046 18164 18052 18216
rect 18104 18164 18110 18216
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18204 19579 18207
rect 19797 18207 19855 18213
rect 19797 18204 19809 18207
rect 19567 18176 19809 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 19797 18173 19809 18176
rect 19843 18204 19855 18207
rect 20346 18204 20352 18216
rect 19843 18176 20352 18204
rect 19843 18173 19855 18176
rect 19797 18167 19855 18173
rect 19352 18136 19380 18167
rect 20346 18164 20352 18176
rect 20404 18164 20410 18216
rect 20070 18136 20076 18148
rect 19352 18108 20076 18136
rect 20070 18096 20076 18108
rect 20128 18096 20134 18148
rect 22020 18136 22048 18235
rect 22112 18204 22140 18235
rect 22186 18232 22192 18284
rect 22244 18232 22250 18284
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18272 22431 18275
rect 22554 18272 22560 18284
rect 22419 18244 22560 18272
rect 22419 18241 22431 18244
rect 22373 18235 22431 18241
rect 22554 18232 22560 18244
rect 22612 18232 22618 18284
rect 22646 18232 22652 18284
rect 22704 18272 22710 18284
rect 22704 18244 23428 18272
rect 22704 18232 22710 18244
rect 23400 18216 23428 18244
rect 23474 18232 23480 18284
rect 23532 18232 23538 18284
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 23658 18232 23664 18284
rect 23716 18232 23722 18284
rect 23842 18232 23848 18284
rect 23900 18232 23906 18284
rect 23937 18275 23995 18281
rect 23937 18241 23949 18275
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 22278 18204 22284 18216
rect 22112 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18164 22342 18216
rect 23201 18207 23259 18213
rect 23201 18173 23213 18207
rect 23247 18173 23259 18207
rect 23201 18167 23259 18173
rect 23216 18136 23244 18167
rect 23382 18164 23388 18216
rect 23440 18204 23446 18216
rect 23952 18204 23980 18235
rect 24118 18232 24124 18284
rect 24176 18232 24182 18284
rect 24320 18281 24348 18312
rect 24581 18309 24593 18343
rect 24627 18340 24639 18343
rect 24854 18340 24860 18352
rect 24627 18312 24860 18340
rect 24627 18309 24639 18312
rect 24581 18303 24639 18309
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 25038 18300 25044 18352
rect 25096 18300 25102 18352
rect 27172 18340 27200 18368
rect 28736 18340 28764 18380
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 31202 18368 31208 18420
rect 31260 18368 31266 18420
rect 32677 18411 32735 18417
rect 32677 18377 32689 18411
rect 32723 18408 32735 18411
rect 32723 18380 33088 18408
rect 32723 18377 32735 18380
rect 32677 18371 32735 18377
rect 27172 18312 27476 18340
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18241 24363 18275
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 24305 18235 24363 18241
rect 25976 18244 26985 18272
rect 23440 18176 23980 18204
rect 23440 18164 23446 18176
rect 25314 18164 25320 18216
rect 25372 18204 25378 18216
rect 25976 18204 26004 18244
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 25372 18176 26004 18204
rect 26053 18207 26111 18213
rect 25372 18164 25378 18176
rect 26053 18173 26065 18207
rect 26099 18204 26111 18207
rect 26697 18207 26755 18213
rect 26697 18204 26709 18207
rect 26099 18176 26709 18204
rect 26099 18173 26111 18176
rect 26053 18167 26111 18173
rect 26697 18173 26709 18176
rect 26743 18173 26755 18207
rect 26988 18204 27016 18235
rect 27062 18232 27068 18284
rect 27120 18272 27126 18284
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 27120 18244 27169 18272
rect 27120 18232 27126 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27246 18232 27252 18284
rect 27304 18232 27310 18284
rect 27448 18281 27476 18312
rect 28460 18312 28764 18340
rect 28460 18281 28488 18312
rect 29454 18300 29460 18352
rect 29512 18300 29518 18352
rect 30098 18300 30104 18352
rect 30156 18300 30162 18352
rect 30469 18343 30527 18349
rect 30469 18309 30481 18343
rect 30515 18340 30527 18343
rect 30558 18340 30564 18352
rect 30515 18312 30564 18340
rect 30515 18309 30527 18312
rect 30469 18303 30527 18309
rect 30558 18300 30564 18312
rect 30616 18300 30622 18352
rect 30650 18300 30656 18352
rect 30708 18300 30714 18352
rect 31478 18300 31484 18352
rect 31536 18300 31542 18352
rect 31662 18300 31668 18352
rect 31720 18349 31726 18352
rect 31720 18343 31749 18349
rect 31737 18309 31749 18343
rect 31720 18303 31749 18309
rect 32309 18343 32367 18349
rect 32309 18309 32321 18343
rect 32355 18340 32367 18343
rect 32582 18340 32588 18352
rect 32355 18312 32588 18340
rect 32355 18309 32367 18312
rect 32309 18303 32367 18309
rect 31720 18300 31726 18303
rect 32582 18300 32588 18312
rect 32640 18300 32646 18352
rect 33060 18349 33088 18380
rect 35434 18368 35440 18420
rect 35492 18368 35498 18420
rect 37369 18411 37427 18417
rect 37369 18377 37381 18411
rect 37415 18408 37427 18411
rect 37734 18408 37740 18420
rect 37415 18380 37740 18408
rect 37415 18377 37427 18380
rect 37369 18371 37427 18377
rect 37734 18368 37740 18380
rect 37792 18368 37798 18420
rect 38378 18368 38384 18420
rect 38436 18408 38442 18420
rect 38473 18411 38531 18417
rect 38473 18408 38485 18411
rect 38436 18380 38485 18408
rect 38436 18368 38442 18380
rect 38473 18377 38485 18380
rect 38519 18377 38531 18411
rect 38473 18371 38531 18377
rect 41049 18411 41107 18417
rect 41049 18377 41061 18411
rect 41095 18408 41107 18411
rect 41598 18408 41604 18420
rect 41095 18380 41604 18408
rect 41095 18377 41107 18380
rect 41049 18371 41107 18377
rect 41598 18368 41604 18380
rect 41656 18368 41662 18420
rect 41782 18368 41788 18420
rect 41840 18368 41846 18420
rect 33045 18343 33103 18349
rect 33045 18309 33057 18343
rect 33091 18309 33103 18343
rect 35452 18340 35480 18368
rect 37458 18340 37464 18352
rect 34270 18312 35480 18340
rect 36846 18312 37464 18340
rect 33045 18303 33103 18309
rect 37458 18300 37464 18312
rect 37516 18300 37522 18352
rect 40494 18300 40500 18352
rect 40552 18340 40558 18352
rect 41322 18340 41328 18352
rect 40552 18312 41328 18340
rect 40552 18300 40558 18312
rect 41322 18300 41328 18312
rect 41380 18300 41386 18352
rect 41417 18343 41475 18349
rect 41417 18309 41429 18343
rect 41463 18340 41475 18343
rect 41506 18340 41512 18352
rect 41463 18312 41512 18340
rect 41463 18309 41475 18312
rect 41417 18303 41475 18309
rect 41506 18300 41512 18312
rect 41564 18300 41570 18352
rect 41708 18312 42012 18340
rect 27433 18275 27491 18281
rect 27433 18241 27445 18275
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 28261 18275 28319 18281
rect 28261 18241 28273 18275
rect 28307 18241 28319 18275
rect 28261 18235 28319 18241
rect 28445 18275 28503 18281
rect 28445 18241 28457 18275
rect 28491 18241 28503 18275
rect 28445 18235 28503 18241
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 27341 18207 27399 18213
rect 27341 18204 27353 18207
rect 26988 18176 27353 18204
rect 26697 18167 26755 18173
rect 27341 18173 27353 18176
rect 27387 18173 27399 18207
rect 27341 18167 27399 18173
rect 23293 18139 23351 18145
rect 23293 18136 23305 18139
rect 22020 18108 22094 18136
rect 23216 18108 23305 18136
rect 15013 18071 15071 18077
rect 15013 18068 15025 18071
rect 14608 18040 15025 18068
rect 14608 18028 14614 18040
rect 15013 18037 15025 18040
rect 15059 18037 15071 18071
rect 15013 18031 15071 18037
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15286 18068 15292 18080
rect 15151 18040 15292 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16632 18040 16681 18068
rect 16632 18028 16638 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 18693 18071 18751 18077
rect 18693 18037 18705 18071
rect 18739 18068 18751 18071
rect 18782 18068 18788 18080
rect 18739 18040 18788 18068
rect 18739 18037 18751 18040
rect 18693 18031 18751 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19429 18071 19487 18077
rect 19429 18068 19441 18071
rect 19392 18040 19441 18068
rect 19392 18028 19398 18040
rect 19429 18037 19441 18040
rect 19475 18037 19487 18071
rect 19429 18031 19487 18037
rect 21910 18028 21916 18080
rect 21968 18068 21974 18080
rect 22066 18068 22094 18108
rect 23293 18105 23305 18108
rect 23339 18105 23351 18139
rect 23293 18099 23351 18105
rect 23658 18096 23664 18148
rect 23716 18136 23722 18148
rect 23842 18136 23848 18148
rect 23716 18108 23848 18136
rect 23716 18096 23722 18108
rect 23842 18096 23848 18108
rect 23900 18096 23906 18148
rect 23937 18139 23995 18145
rect 23937 18105 23949 18139
rect 23983 18136 23995 18139
rect 24118 18136 24124 18148
rect 23983 18108 24124 18136
rect 23983 18105 23995 18108
rect 23937 18099 23995 18105
rect 24118 18096 24124 18108
rect 24176 18096 24182 18148
rect 26142 18096 26148 18148
rect 26200 18096 26206 18148
rect 25590 18068 25596 18080
rect 21968 18040 25596 18068
rect 21968 18028 21974 18040
rect 25590 18028 25596 18040
rect 25648 18028 25654 18080
rect 25682 18028 25688 18080
rect 25740 18068 25746 18080
rect 27065 18071 27123 18077
rect 27065 18068 27077 18071
rect 25740 18040 27077 18068
rect 25740 18028 25746 18040
rect 27065 18037 27077 18040
rect 27111 18037 27123 18071
rect 28276 18068 28304 18235
rect 28552 18204 28580 18235
rect 30374 18232 30380 18284
rect 30432 18232 30438 18284
rect 31389 18275 31447 18281
rect 31389 18241 31401 18275
rect 31435 18241 31447 18275
rect 31389 18235 31447 18241
rect 31573 18275 31631 18281
rect 31573 18241 31585 18275
rect 31619 18241 31631 18275
rect 31573 18235 31631 18241
rect 32125 18275 32183 18281
rect 32125 18241 32137 18275
rect 32171 18272 32183 18275
rect 32214 18272 32220 18284
rect 32171 18244 32220 18272
rect 32171 18241 32183 18244
rect 32125 18235 32183 18241
rect 29086 18204 29092 18216
rect 28552 18176 29092 18204
rect 29086 18164 29092 18176
rect 29144 18164 29150 18216
rect 31404 18136 31432 18235
rect 31478 18164 31484 18216
rect 31536 18204 31542 18216
rect 31588 18204 31616 18235
rect 32214 18232 32220 18244
rect 32272 18232 32278 18284
rect 32401 18275 32459 18281
rect 32401 18241 32413 18275
rect 32447 18241 32459 18275
rect 32401 18235 32459 18241
rect 31536 18176 31616 18204
rect 31849 18207 31907 18213
rect 31536 18164 31542 18176
rect 31849 18173 31861 18207
rect 31895 18204 31907 18207
rect 32416 18204 32444 18235
rect 32490 18232 32496 18284
rect 32548 18232 32554 18284
rect 38013 18275 38071 18281
rect 38013 18241 38025 18275
rect 38059 18272 38071 18275
rect 38102 18272 38108 18284
rect 38059 18244 38108 18272
rect 38059 18241 38071 18244
rect 38013 18235 38071 18241
rect 31895 18176 32076 18204
rect 32416 18176 32536 18204
rect 31895 18173 31907 18176
rect 31849 18167 31907 18173
rect 31938 18136 31944 18148
rect 31404 18108 31944 18136
rect 31938 18096 31944 18108
rect 31996 18096 32002 18148
rect 32048 18136 32076 18176
rect 32306 18136 32312 18148
rect 32048 18108 32312 18136
rect 32306 18096 32312 18108
rect 32364 18096 32370 18148
rect 28902 18068 28908 18080
rect 28276 18040 28908 18068
rect 27065 18031 27123 18037
rect 28902 18028 28908 18040
rect 28960 18028 28966 18080
rect 30282 18028 30288 18080
rect 30340 18068 30346 18080
rect 30837 18071 30895 18077
rect 30837 18068 30849 18071
rect 30340 18040 30849 18068
rect 30340 18028 30346 18040
rect 30837 18037 30849 18040
rect 30883 18037 30895 18071
rect 32508 18068 32536 18176
rect 32766 18164 32772 18216
rect 32824 18164 32830 18216
rect 34606 18164 34612 18216
rect 34664 18204 34670 18216
rect 35345 18207 35403 18213
rect 35345 18204 35357 18207
rect 34664 18176 35357 18204
rect 34664 18164 34670 18176
rect 35345 18173 35357 18176
rect 35391 18173 35403 18207
rect 35345 18167 35403 18173
rect 35621 18207 35679 18213
rect 35621 18173 35633 18207
rect 35667 18204 35679 18207
rect 37274 18204 37280 18216
rect 35667 18176 37280 18204
rect 35667 18173 35679 18176
rect 35621 18167 35679 18173
rect 37274 18164 37280 18176
rect 37332 18164 37338 18216
rect 37093 18139 37151 18145
rect 37093 18105 37105 18139
rect 37139 18136 37151 18139
rect 38028 18136 38056 18235
rect 38102 18232 38108 18244
rect 38160 18232 38166 18284
rect 39022 18232 39028 18284
rect 39080 18232 39086 18284
rect 39853 18275 39911 18281
rect 39853 18241 39865 18275
rect 39899 18272 39911 18275
rect 40034 18272 40040 18284
rect 39899 18244 40040 18272
rect 39899 18241 39911 18244
rect 39853 18235 39911 18241
rect 40034 18232 40040 18244
rect 40092 18232 40098 18284
rect 41138 18232 41144 18284
rect 41196 18272 41202 18284
rect 41708 18281 41736 18312
rect 41984 18281 42012 18312
rect 41233 18275 41291 18281
rect 41233 18272 41245 18275
rect 41196 18244 41245 18272
rect 41196 18232 41202 18244
rect 41233 18241 41245 18244
rect 41279 18241 41291 18275
rect 41233 18235 41291 18241
rect 41601 18275 41659 18281
rect 41601 18241 41613 18275
rect 41647 18241 41659 18275
rect 41601 18235 41659 18241
rect 41693 18275 41751 18281
rect 41693 18241 41705 18275
rect 41739 18241 41751 18275
rect 41693 18235 41751 18241
rect 41877 18275 41935 18281
rect 41877 18241 41889 18275
rect 41923 18241 41935 18275
rect 41877 18235 41935 18241
rect 41969 18275 42027 18281
rect 41969 18241 41981 18275
rect 42015 18272 42027 18275
rect 42058 18272 42064 18284
rect 42015 18244 42064 18272
rect 42015 18241 42027 18244
rect 41969 18235 42027 18241
rect 39758 18164 39764 18216
rect 39816 18164 39822 18216
rect 40218 18164 40224 18216
rect 40276 18164 40282 18216
rect 40770 18204 40776 18216
rect 40328 18176 40776 18204
rect 37139 18108 38056 18136
rect 37139 18105 37151 18108
rect 37093 18099 37151 18105
rect 40126 18096 40132 18148
rect 40184 18136 40190 18148
rect 40328 18136 40356 18176
rect 40770 18164 40776 18176
rect 40828 18204 40834 18216
rect 41616 18204 41644 18235
rect 40828 18176 41644 18204
rect 41892 18204 41920 18235
rect 42058 18232 42064 18244
rect 42116 18232 42122 18284
rect 42150 18232 42156 18284
rect 42208 18232 42214 18284
rect 42168 18204 42196 18232
rect 41892 18176 42196 18204
rect 40828 18164 40834 18176
rect 40184 18108 40356 18136
rect 40184 18096 40190 18108
rect 40402 18096 40408 18148
rect 40460 18136 40466 18148
rect 42061 18139 42119 18145
rect 42061 18136 42073 18139
rect 40460 18108 42073 18136
rect 40460 18096 40466 18108
rect 42061 18105 42073 18108
rect 42107 18105 42119 18139
rect 42061 18099 42119 18105
rect 33134 18068 33140 18080
rect 32508 18040 33140 18068
rect 30837 18031 30895 18037
rect 33134 18028 33140 18040
rect 33192 18028 33198 18080
rect 33686 18028 33692 18080
rect 33744 18068 33750 18080
rect 34517 18071 34575 18077
rect 34517 18068 34529 18071
rect 33744 18040 34529 18068
rect 33744 18028 33750 18040
rect 34517 18037 34529 18040
rect 34563 18037 34575 18071
rect 34517 18031 34575 18037
rect 1104 17978 42504 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 42504 17978
rect 1104 17904 42504 17926
rect 3786 17824 3792 17876
rect 3844 17824 3850 17876
rect 5350 17824 5356 17876
rect 5408 17824 5414 17876
rect 5629 17867 5687 17873
rect 5629 17833 5641 17867
rect 5675 17864 5687 17867
rect 5718 17864 5724 17876
rect 5675 17836 5724 17864
rect 5675 17833 5687 17836
rect 5629 17827 5687 17833
rect 5718 17824 5724 17836
rect 5776 17824 5782 17876
rect 7558 17864 7564 17876
rect 6748 17836 7564 17864
rect 5442 17756 5448 17808
rect 5500 17796 5506 17808
rect 5813 17799 5871 17805
rect 5813 17796 5825 17799
rect 5500 17768 5825 17796
rect 5500 17756 5506 17768
rect 5813 17765 5825 17768
rect 5859 17765 5871 17799
rect 5813 17759 5871 17765
rect 1394 17688 1400 17740
rect 1452 17688 1458 17740
rect 4801 17731 4859 17737
rect 4801 17697 4813 17731
rect 4847 17728 4859 17731
rect 5626 17728 5632 17740
rect 4847 17700 5632 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 5718 17688 5724 17740
rect 5776 17688 5782 17740
rect 6748 17737 6776 17836
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 8018 17824 8024 17876
rect 8076 17864 8082 17876
rect 9125 17867 9183 17873
rect 9125 17864 9137 17867
rect 8076 17836 9137 17864
rect 8076 17824 8082 17836
rect 9125 17833 9137 17836
rect 9171 17833 9183 17867
rect 9125 17827 9183 17833
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10042 17864 10048 17876
rect 9732 17836 10048 17864
rect 9732 17824 9738 17836
rect 10042 17824 10048 17836
rect 10100 17864 10106 17876
rect 10413 17867 10471 17873
rect 10413 17864 10425 17867
rect 10100 17836 10425 17864
rect 10100 17824 10106 17836
rect 10413 17833 10425 17836
rect 10459 17864 10471 17867
rect 10502 17864 10508 17876
rect 10459 17836 10508 17864
rect 10459 17833 10471 17836
rect 10413 17827 10471 17833
rect 10502 17824 10508 17836
rect 10560 17824 10566 17876
rect 10594 17824 10600 17876
rect 10652 17824 10658 17876
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13998 17864 14004 17876
rect 13035 17836 14004 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 14182 17824 14188 17876
rect 14240 17824 14246 17876
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17864 17371 17867
rect 18046 17864 18052 17876
rect 17359 17836 18052 17864
rect 17359 17833 17371 17836
rect 17313 17827 17371 17833
rect 18046 17824 18052 17836
rect 18104 17864 18110 17876
rect 19242 17864 19248 17876
rect 18104 17836 19248 17864
rect 18104 17824 18110 17836
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 21545 17867 21603 17873
rect 21545 17864 21557 17867
rect 20864 17836 21557 17864
rect 20864 17824 20870 17836
rect 21545 17833 21557 17836
rect 21591 17833 21603 17867
rect 21545 17827 21603 17833
rect 22186 17824 22192 17876
rect 22244 17864 22250 17876
rect 22281 17867 22339 17873
rect 22281 17864 22293 17867
rect 22244 17836 22293 17864
rect 22244 17824 22250 17836
rect 22281 17833 22293 17836
rect 22327 17833 22339 17867
rect 22281 17827 22339 17833
rect 24854 17824 24860 17876
rect 24912 17824 24918 17876
rect 28350 17824 28356 17876
rect 28408 17864 28414 17876
rect 28721 17867 28779 17873
rect 28721 17864 28733 17867
rect 28408 17836 28733 17864
rect 28408 17824 28414 17836
rect 28721 17833 28733 17836
rect 28767 17833 28779 17867
rect 28721 17827 28779 17833
rect 29546 17824 29552 17876
rect 29604 17824 29610 17876
rect 30929 17867 30987 17873
rect 30929 17833 30941 17867
rect 30975 17864 30987 17867
rect 33229 17867 33287 17873
rect 33229 17864 33241 17867
rect 30975 17836 33241 17864
rect 30975 17833 30987 17836
rect 30929 17827 30987 17833
rect 33229 17833 33241 17836
rect 33275 17833 33287 17867
rect 33229 17827 33287 17833
rect 33505 17867 33563 17873
rect 33505 17833 33517 17867
rect 33551 17864 33563 17867
rect 36170 17864 36176 17876
rect 33551 17836 36176 17864
rect 33551 17833 33563 17836
rect 33505 17827 33563 17833
rect 36170 17824 36176 17836
rect 36228 17824 36234 17876
rect 37274 17824 37280 17876
rect 37332 17824 37338 17876
rect 37550 17824 37556 17876
rect 37608 17864 37614 17876
rect 37921 17867 37979 17873
rect 37921 17864 37933 17867
rect 37608 17836 37933 17864
rect 37608 17824 37614 17836
rect 37921 17833 37933 17836
rect 37967 17833 37979 17867
rect 37921 17827 37979 17833
rect 7190 17756 7196 17808
rect 7248 17756 7254 17808
rect 8754 17756 8760 17808
rect 8812 17796 8818 17808
rect 9490 17796 9496 17808
rect 8812 17768 9496 17796
rect 8812 17756 8818 17768
rect 9490 17756 9496 17768
rect 9548 17796 9554 17808
rect 10226 17796 10232 17808
rect 9548 17768 10232 17796
rect 9548 17756 9554 17768
rect 10226 17756 10232 17768
rect 10284 17756 10290 17808
rect 10321 17799 10379 17805
rect 10321 17765 10333 17799
rect 10367 17796 10379 17799
rect 12158 17796 12164 17808
rect 10367 17768 12164 17796
rect 10367 17765 10379 17768
rect 10321 17759 10379 17765
rect 12158 17756 12164 17768
rect 12216 17756 12222 17808
rect 14645 17799 14703 17805
rect 14645 17796 14657 17799
rect 12820 17768 14657 17796
rect 6733 17731 6791 17737
rect 6733 17697 6745 17731
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17728 6883 17731
rect 7282 17728 7288 17740
rect 6871 17700 7288 17728
rect 6871 17697 6883 17700
rect 6825 17691 6883 17697
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 10060 17728 10180 17736
rect 11514 17728 11520 17740
rect 9324 17708 11520 17728
rect 9324 17700 10088 17708
rect 10152 17700 11520 17708
rect 1762 17620 1768 17672
rect 1820 17620 1826 17672
rect 3191 17663 3249 17669
rect 3191 17629 3203 17663
rect 3237 17660 3249 17663
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 3237 17632 4353 17660
rect 3237 17629 3249 17632
rect 3191 17623 3249 17629
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4614 17620 4620 17672
rect 4672 17660 4678 17672
rect 5166 17660 5172 17672
rect 4672 17632 5172 17660
rect 4672 17620 4678 17632
rect 5166 17620 5172 17632
rect 5224 17660 5230 17672
rect 5445 17663 5503 17669
rect 5445 17660 5457 17663
rect 5224 17632 5457 17660
rect 5224 17620 5230 17632
rect 5445 17629 5457 17632
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17660 5595 17663
rect 5813 17663 5871 17669
rect 5813 17660 5825 17663
rect 5583 17632 5825 17660
rect 5583 17629 5595 17632
rect 5537 17623 5595 17629
rect 5644 17604 5672 17632
rect 5813 17629 5825 17632
rect 5859 17629 5871 17663
rect 5813 17623 5871 17629
rect 5997 17663 6055 17669
rect 5997 17629 6009 17663
rect 6043 17629 6055 17663
rect 5997 17623 6055 17629
rect 2590 17552 2596 17604
rect 2648 17552 2654 17604
rect 4893 17595 4951 17601
rect 4893 17561 4905 17595
rect 4939 17592 4951 17595
rect 5350 17592 5356 17604
rect 4939 17564 5356 17592
rect 4939 17561 4951 17564
rect 4893 17555 4951 17561
rect 5350 17552 5356 17564
rect 5408 17552 5414 17604
rect 5626 17552 5632 17604
rect 5684 17552 5690 17604
rect 6012 17592 6040 17623
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17660 7435 17663
rect 9324 17660 9352 17700
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 12820 17737 12848 17768
rect 14645 17765 14657 17768
rect 14691 17765 14703 17799
rect 14645 17759 14703 17765
rect 20993 17799 21051 17805
rect 20993 17765 21005 17799
rect 21039 17796 21051 17799
rect 21450 17796 21456 17808
rect 21039 17768 21456 17796
rect 21039 17765 21051 17768
rect 20993 17759 21051 17765
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 21637 17799 21695 17805
rect 21637 17765 21649 17799
rect 21683 17796 21695 17799
rect 21683 17768 21956 17796
rect 21683 17765 21695 17768
rect 21637 17759 21695 17765
rect 12805 17731 12863 17737
rect 12805 17697 12817 17731
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 13909 17731 13967 17737
rect 13909 17697 13921 17731
rect 13955 17728 13967 17731
rect 15102 17728 15108 17740
rect 13955 17700 15108 17728
rect 13955 17697 13967 17700
rect 13909 17691 13967 17697
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15473 17731 15531 17737
rect 15473 17728 15485 17731
rect 15252 17700 15485 17728
rect 15252 17688 15258 17700
rect 15473 17697 15485 17700
rect 15519 17697 15531 17731
rect 15473 17691 15531 17697
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 18690 17728 18696 17740
rect 15795 17700 18696 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 18782 17688 18788 17740
rect 18840 17688 18846 17740
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17728 19119 17731
rect 20714 17728 20720 17740
rect 19107 17700 20720 17728
rect 19107 17697 19119 17700
rect 19061 17691 19119 17697
rect 20714 17688 20720 17700
rect 20772 17688 20778 17740
rect 21192 17700 21680 17728
rect 7423 17632 9352 17660
rect 7423 17629 7435 17632
rect 7377 17623 7435 17629
rect 9398 17620 9404 17672
rect 9456 17620 9462 17672
rect 9490 17620 9496 17672
rect 9548 17620 9554 17672
rect 9858 17620 9864 17672
rect 9916 17620 9922 17672
rect 9950 17620 9956 17672
rect 10008 17620 10014 17672
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 7622 17595 7680 17601
rect 7622 17592 7634 17595
rect 5736 17564 6040 17592
rect 7300 17564 7634 17592
rect 5736 17536 5764 17564
rect 4985 17527 5043 17533
rect 4985 17493 4997 17527
rect 5031 17524 5043 17527
rect 5718 17524 5724 17536
rect 5031 17496 5724 17524
rect 5031 17493 5043 17496
rect 4985 17487 5043 17493
rect 5718 17484 5724 17496
rect 5776 17484 5782 17536
rect 6365 17527 6423 17533
rect 6365 17493 6377 17527
rect 6411 17524 6423 17527
rect 6454 17524 6460 17536
rect 6411 17496 6460 17524
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 7300 17533 7328 17564
rect 7622 17561 7634 17564
rect 7668 17561 7680 17595
rect 7622 17555 7680 17561
rect 9033 17595 9091 17601
rect 9033 17561 9045 17595
rect 9079 17592 9091 17595
rect 9582 17592 9588 17604
rect 9079 17564 9588 17592
rect 9079 17561 9091 17564
rect 9033 17555 9091 17561
rect 9582 17552 9588 17564
rect 9640 17592 9646 17604
rect 10060 17592 10088 17623
rect 10134 17620 10140 17672
rect 10192 17620 10198 17672
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10284 17632 10609 17660
rect 10284 17620 10290 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 10686 17620 10692 17672
rect 10744 17620 10750 17672
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 12667 17632 13277 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 13265 17629 13277 17632
rect 13311 17660 13323 17663
rect 13446 17660 13452 17672
rect 13311 17632 13452 17660
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 14090 17620 14096 17672
rect 14148 17620 14154 17672
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14550 17660 14556 17672
rect 14507 17632 14556 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 14829 17663 14887 17669
rect 14829 17629 14841 17663
rect 14875 17660 14887 17663
rect 15286 17660 15292 17672
rect 14875 17632 15292 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 17678 17660 17684 17672
rect 16882 17632 17684 17660
rect 17678 17620 17684 17632
rect 17736 17620 17742 17672
rect 19242 17620 19248 17672
rect 19300 17620 19306 17672
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19886 17660 19892 17672
rect 19475 17632 19892 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20404 17632 20913 17660
rect 20404 17620 20410 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 21192 17669 21220 17700
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 21048 17632 21097 17660
rect 21048 17620 21054 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17629 21235 17663
rect 21177 17623 21235 17629
rect 21266 17620 21272 17672
rect 21324 17660 21330 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 21324 17632 21373 17660
rect 21324 17620 21330 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 21652 17660 21680 17700
rect 21726 17688 21732 17740
rect 21784 17688 21790 17740
rect 21928 17737 21956 17768
rect 22554 17756 22560 17808
rect 22612 17796 22618 17808
rect 22612 17768 24900 17796
rect 22612 17756 22618 17768
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17697 21971 17731
rect 23477 17731 23535 17737
rect 23477 17728 23489 17731
rect 21913 17691 21971 17697
rect 22756 17700 23489 17728
rect 22756 17669 22784 17700
rect 23477 17697 23489 17700
rect 23523 17697 23535 17731
rect 24872 17728 24900 17768
rect 24946 17756 24952 17808
rect 25004 17796 25010 17808
rect 25682 17796 25688 17808
rect 25004 17768 25688 17796
rect 25004 17756 25010 17768
rect 25682 17756 25688 17768
rect 25740 17756 25746 17808
rect 28534 17756 28540 17808
rect 28592 17796 28598 17808
rect 29362 17796 29368 17808
rect 28592 17768 29368 17796
rect 28592 17756 28598 17768
rect 29362 17756 29368 17768
rect 29420 17756 29426 17808
rect 30285 17799 30343 17805
rect 30285 17765 30297 17799
rect 30331 17796 30343 17799
rect 30331 17768 30696 17796
rect 30331 17765 30343 17768
rect 30285 17759 30343 17765
rect 25130 17728 25136 17740
rect 24872 17700 25136 17728
rect 23477 17691 23535 17697
rect 25130 17688 25136 17700
rect 25188 17688 25194 17740
rect 26050 17728 26056 17740
rect 25358 17700 26056 17728
rect 22005 17663 22063 17669
rect 21652 17632 21956 17660
rect 9640 17564 10088 17592
rect 10873 17595 10931 17601
rect 9640 17552 9646 17564
rect 10873 17561 10885 17595
rect 10919 17561 10931 17595
rect 10873 17555 10931 17561
rect 7285 17527 7343 17533
rect 7285 17493 7297 17527
rect 7331 17493 7343 17527
rect 7285 17487 7343 17493
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 9398 17524 9404 17536
rect 7800 17496 9404 17524
rect 7800 17484 7806 17496
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9674 17484 9680 17536
rect 9732 17484 9738 17536
rect 10888 17524 10916 17555
rect 11698 17552 11704 17604
rect 11756 17592 11762 17604
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 11756 17564 13093 17592
rect 11756 17552 11762 17564
rect 13081 17561 13093 17564
rect 13127 17561 13139 17595
rect 13081 17555 13139 17561
rect 20717 17595 20775 17601
rect 20717 17561 20729 17595
rect 20763 17592 20775 17595
rect 21928 17592 21956 17632
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22465 17663 22523 17669
rect 22465 17660 22477 17663
rect 22051 17632 22477 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 22465 17629 22477 17632
rect 22511 17629 22523 17663
rect 22740 17663 22798 17669
rect 22740 17660 22752 17663
rect 22465 17623 22523 17629
rect 22664 17632 22752 17660
rect 22664 17592 22692 17632
rect 22740 17629 22752 17632
rect 22786 17629 22798 17663
rect 22740 17623 22798 17629
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17629 22891 17663
rect 22833 17623 22891 17629
rect 20763 17564 21864 17592
rect 21928 17564 22692 17592
rect 22848 17592 22876 17623
rect 23382 17620 23388 17672
rect 23440 17620 23446 17672
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 24026 17660 24032 17672
rect 23615 17632 24032 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 24946 17660 24952 17672
rect 24811 17632 24952 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 25041 17663 25099 17669
rect 25041 17629 25053 17663
rect 25087 17629 25099 17663
rect 25148 17660 25176 17688
rect 25358 17669 25386 17700
rect 26050 17688 26056 17700
rect 26108 17688 26114 17740
rect 27341 17731 27399 17737
rect 27341 17697 27353 17731
rect 27387 17728 27399 17731
rect 28350 17728 28356 17740
rect 27387 17700 28356 17728
rect 27387 17697 27399 17700
rect 27341 17691 27399 17697
rect 28350 17688 28356 17700
rect 28408 17688 28414 17740
rect 28626 17688 28632 17740
rect 28684 17728 28690 17740
rect 28684 17700 30512 17728
rect 28684 17688 28690 17700
rect 25225 17663 25283 17669
rect 25225 17660 25237 17663
rect 25148 17632 25237 17660
rect 25041 17623 25099 17629
rect 25225 17629 25237 17632
rect 25271 17629 25283 17663
rect 25225 17623 25283 17629
rect 25343 17663 25401 17669
rect 25343 17629 25355 17663
rect 25389 17629 25401 17663
rect 25343 17623 25401 17629
rect 24118 17592 24124 17604
rect 22848 17564 24124 17592
rect 20763 17561 20775 17564
rect 20717 17555 20775 17561
rect 12437 17527 12495 17533
rect 12437 17524 12449 17527
rect 10888 17496 12449 17524
rect 12437 17493 12449 17496
rect 12483 17493 12495 17527
rect 12437 17487 12495 17493
rect 15378 17484 15384 17536
rect 15436 17484 15442 17536
rect 17218 17484 17224 17536
rect 17276 17484 17282 17536
rect 19610 17484 19616 17536
rect 19668 17524 19674 17536
rect 20162 17524 20168 17536
rect 19668 17496 20168 17524
rect 19668 17484 19674 17496
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 21726 17524 21732 17536
rect 21324 17496 21732 17524
rect 21324 17484 21330 17496
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 21836 17524 21864 17564
rect 24118 17552 24124 17564
rect 24176 17552 24182 17604
rect 24673 17595 24731 17601
rect 24673 17561 24685 17595
rect 24719 17592 24731 17595
rect 25056 17592 25084 17623
rect 25498 17620 25504 17672
rect 25556 17620 25562 17672
rect 27433 17663 27491 17669
rect 27433 17629 27445 17663
rect 27479 17629 27491 17663
rect 27433 17623 27491 17629
rect 24719 17564 25084 17592
rect 24719 17561 24731 17564
rect 24673 17555 24731 17561
rect 25130 17552 25136 17604
rect 25188 17552 25194 17604
rect 26510 17552 26516 17604
rect 26568 17552 26574 17604
rect 27062 17552 27068 17604
rect 27120 17552 27126 17604
rect 23474 17524 23480 17536
rect 21836 17496 23480 17524
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 24394 17484 24400 17536
rect 24452 17524 24458 17536
rect 25314 17524 25320 17536
rect 24452 17496 25320 17524
rect 24452 17484 24458 17496
rect 25314 17484 25320 17496
rect 25372 17484 25378 17536
rect 25593 17527 25651 17533
rect 25593 17493 25605 17527
rect 25639 17524 25651 17527
rect 26418 17524 26424 17536
rect 25639 17496 26424 17524
rect 25639 17493 25651 17496
rect 25593 17487 25651 17493
rect 26418 17484 26424 17496
rect 26476 17484 26482 17536
rect 26970 17484 26976 17536
rect 27028 17524 27034 17536
rect 27338 17524 27344 17536
rect 27028 17496 27344 17524
rect 27028 17484 27034 17496
rect 27338 17484 27344 17496
rect 27396 17524 27402 17536
rect 27448 17524 27476 17623
rect 27706 17620 27712 17672
rect 27764 17660 27770 17672
rect 28261 17663 28319 17669
rect 28261 17660 28273 17663
rect 27764 17632 28273 17660
rect 27764 17620 27770 17632
rect 28261 17629 28273 17632
rect 28307 17629 28319 17663
rect 28261 17623 28319 17629
rect 28445 17663 28503 17669
rect 28445 17629 28457 17663
rect 28491 17660 28503 17663
rect 28810 17660 28816 17672
rect 28491 17632 28816 17660
rect 28491 17629 28503 17632
rect 28445 17623 28503 17629
rect 27890 17552 27896 17604
rect 27948 17592 27954 17604
rect 28460 17592 28488 17623
rect 28810 17620 28816 17632
rect 28868 17620 28874 17672
rect 28902 17620 28908 17672
rect 28960 17620 28966 17672
rect 29178 17620 29184 17672
rect 29236 17620 29242 17672
rect 29730 17620 29736 17672
rect 29788 17620 29794 17672
rect 29914 17620 29920 17672
rect 29972 17620 29978 17672
rect 30098 17620 30104 17672
rect 30156 17620 30162 17672
rect 30193 17663 30251 17669
rect 30193 17629 30205 17663
rect 30239 17660 30251 17663
rect 30282 17660 30288 17672
rect 30239 17632 30288 17660
rect 30239 17629 30251 17632
rect 30193 17623 30251 17629
rect 27948 17564 28488 17592
rect 27948 17552 27954 17564
rect 29822 17552 29828 17604
rect 29880 17552 29886 17604
rect 27396 17496 27476 17524
rect 27396 17484 27402 17496
rect 27522 17484 27528 17536
rect 27580 17484 27586 17536
rect 28353 17527 28411 17533
rect 28353 17493 28365 17527
rect 28399 17524 28411 17527
rect 28994 17524 29000 17536
rect 28399 17496 29000 17524
rect 28399 17493 28411 17496
rect 28353 17487 28411 17493
rect 28994 17484 29000 17496
rect 29052 17484 29058 17536
rect 29086 17484 29092 17536
rect 29144 17524 29150 17536
rect 30208 17524 30236 17623
rect 30282 17620 30288 17632
rect 30340 17620 30346 17672
rect 30484 17601 30512 17700
rect 30668 17669 30696 17768
rect 30834 17756 30840 17808
rect 30892 17796 30898 17808
rect 31757 17799 31815 17805
rect 31757 17796 31769 17799
rect 30892 17768 31769 17796
rect 30892 17756 30898 17768
rect 31757 17765 31769 17768
rect 31803 17765 31815 17799
rect 31757 17759 31815 17765
rect 31849 17799 31907 17805
rect 31849 17765 31861 17799
rect 31895 17796 31907 17799
rect 32122 17796 32128 17808
rect 31895 17768 32128 17796
rect 31895 17765 31907 17768
rect 31849 17759 31907 17765
rect 32122 17756 32128 17768
rect 32180 17756 32186 17808
rect 32214 17756 32220 17808
rect 32272 17796 32278 17808
rect 32490 17796 32496 17808
rect 32272 17768 32496 17796
rect 32272 17756 32278 17768
rect 32490 17756 32496 17768
rect 32548 17756 32554 17808
rect 37182 17756 37188 17808
rect 37240 17796 37246 17808
rect 38013 17799 38071 17805
rect 38013 17796 38025 17799
rect 37240 17768 38025 17796
rect 37240 17756 37246 17768
rect 38013 17765 38025 17768
rect 38059 17765 38071 17799
rect 38013 17759 38071 17765
rect 31205 17731 31263 17737
rect 31205 17697 31217 17731
rect 31251 17728 31263 17731
rect 31941 17731 31999 17737
rect 31941 17728 31953 17731
rect 31251 17700 31524 17728
rect 31251 17697 31263 17700
rect 31205 17691 31263 17697
rect 30653 17663 30711 17669
rect 30653 17629 30665 17663
rect 30699 17660 30711 17663
rect 31113 17663 31171 17669
rect 31113 17660 31125 17663
rect 30699 17632 31125 17660
rect 30699 17629 30711 17632
rect 30653 17623 30711 17629
rect 31113 17629 31125 17632
rect 31159 17629 31171 17663
rect 31113 17623 31171 17629
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17629 31355 17663
rect 31297 17623 31355 17629
rect 31389 17663 31447 17669
rect 31389 17629 31401 17663
rect 31435 17629 31447 17663
rect 31389 17623 31447 17629
rect 30469 17595 30527 17601
rect 30469 17561 30481 17595
rect 30515 17592 30527 17595
rect 31312 17592 31340 17623
rect 30515 17564 31340 17592
rect 30515 17561 30527 17564
rect 30469 17555 30527 17561
rect 29144 17496 30236 17524
rect 31404 17524 31432 17623
rect 31496 17592 31524 17700
rect 31588 17700 31953 17728
rect 31588 17669 31616 17700
rect 31941 17697 31953 17700
rect 31987 17728 31999 17731
rect 32582 17728 32588 17740
rect 31987 17700 32588 17728
rect 31987 17697 31999 17700
rect 31941 17691 31999 17697
rect 32582 17688 32588 17700
rect 32640 17688 32646 17740
rect 37918 17688 37924 17740
rect 37976 17728 37982 17740
rect 38381 17731 38439 17737
rect 38381 17728 38393 17731
rect 37976 17700 38393 17728
rect 37976 17688 37982 17700
rect 38381 17697 38393 17700
rect 38427 17697 38439 17731
rect 38381 17691 38439 17697
rect 31573 17663 31631 17669
rect 31573 17629 31585 17663
rect 31619 17629 31631 17663
rect 31573 17623 31631 17629
rect 31662 17620 31668 17672
rect 31720 17660 31726 17672
rect 31720 17620 31734 17660
rect 33410 17620 33416 17672
rect 33468 17660 33474 17672
rect 33505 17663 33563 17669
rect 33505 17660 33517 17663
rect 33468 17632 33517 17660
rect 33468 17620 33474 17632
rect 33505 17629 33517 17632
rect 33551 17629 33563 17663
rect 33505 17623 33563 17629
rect 33686 17620 33692 17672
rect 33744 17620 33750 17672
rect 34701 17663 34759 17669
rect 34701 17629 34713 17663
rect 34747 17629 34759 17663
rect 37093 17663 37151 17669
rect 37093 17660 37105 17663
rect 34701 17623 34759 17629
rect 36464 17632 37105 17660
rect 31706 17592 31734 17620
rect 31496 17564 31734 17592
rect 32033 17595 32091 17601
rect 32033 17561 32045 17595
rect 32079 17592 32091 17595
rect 32214 17592 32220 17604
rect 32079 17564 32220 17592
rect 32079 17561 32091 17564
rect 32033 17555 32091 17561
rect 32214 17552 32220 17564
rect 32272 17552 32278 17604
rect 32766 17552 32772 17604
rect 32824 17592 32830 17604
rect 34606 17592 34612 17604
rect 32824 17564 34612 17592
rect 32824 17552 32830 17564
rect 34606 17552 34612 17564
rect 34664 17592 34670 17604
rect 34716 17592 34744 17623
rect 34664 17564 34744 17592
rect 34664 17552 34670 17564
rect 34974 17552 34980 17604
rect 35032 17552 35038 17604
rect 35434 17552 35440 17604
rect 35492 17552 35498 17604
rect 36464 17536 36492 17632
rect 37093 17629 37105 17632
rect 37139 17629 37151 17663
rect 37093 17623 37151 17629
rect 37461 17663 37519 17669
rect 37461 17629 37473 17663
rect 37507 17629 37519 17663
rect 37461 17623 37519 17629
rect 37476 17536 37504 17623
rect 37642 17620 37648 17672
rect 37700 17620 37706 17672
rect 37829 17663 37887 17669
rect 37829 17629 37841 17663
rect 37875 17660 37887 17663
rect 38102 17660 38108 17672
rect 37875 17632 38108 17660
rect 37875 17629 37887 17632
rect 37829 17623 37887 17629
rect 38102 17620 38108 17632
rect 38160 17660 38166 17672
rect 40586 17660 40592 17672
rect 38160 17632 40592 17660
rect 38160 17620 38166 17632
rect 40586 17620 40592 17632
rect 40644 17620 40650 17672
rect 41141 17663 41199 17669
rect 41141 17629 41153 17663
rect 41187 17660 41199 17663
rect 41782 17660 41788 17672
rect 41187 17632 41788 17660
rect 41187 17629 41199 17632
rect 41141 17623 41199 17629
rect 41782 17620 41788 17632
rect 41840 17620 41846 17672
rect 37553 17595 37611 17601
rect 37553 17561 37565 17595
rect 37599 17592 37611 17595
rect 37734 17592 37740 17604
rect 37599 17564 37740 17592
rect 37599 17561 37611 17564
rect 37553 17555 37611 17561
rect 37734 17552 37740 17564
rect 37792 17552 37798 17604
rect 41325 17595 41383 17601
rect 41325 17561 41337 17595
rect 41371 17592 41383 17595
rect 41874 17592 41880 17604
rect 41371 17564 41880 17592
rect 41371 17561 41383 17564
rect 41325 17555 41383 17561
rect 41874 17552 41880 17564
rect 41932 17552 41938 17604
rect 33042 17524 33048 17536
rect 31404 17496 33048 17524
rect 29144 17484 29150 17496
rect 33042 17484 33048 17496
rect 33100 17484 33106 17536
rect 36446 17484 36452 17536
rect 36504 17484 36510 17536
rect 36538 17484 36544 17536
rect 36596 17484 36602 17536
rect 37458 17484 37464 17536
rect 37516 17524 37522 17536
rect 38010 17524 38016 17536
rect 37516 17496 38016 17524
rect 37516 17484 37522 17496
rect 38010 17484 38016 17496
rect 38068 17484 38074 17536
rect 40770 17484 40776 17536
rect 40828 17524 40834 17536
rect 40957 17527 41015 17533
rect 40957 17524 40969 17527
rect 40828 17496 40969 17524
rect 40828 17484 40834 17496
rect 40957 17493 40969 17496
rect 41003 17493 41015 17527
rect 40957 17487 41015 17493
rect 1104 17434 42504 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 42504 17434
rect 1104 17360 42504 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 1762 17320 1768 17332
rect 1627 17292 1768 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2590 17280 2596 17332
rect 2648 17320 2654 17332
rect 5077 17323 5135 17329
rect 2648 17292 3280 17320
rect 2648 17280 2654 17292
rect 3252 17252 3280 17292
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 5258 17320 5264 17332
rect 5123 17292 5264 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5445 17323 5503 17329
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5534 17320 5540 17332
rect 5491 17292 5540 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 5813 17323 5871 17329
rect 5813 17289 5825 17323
rect 5859 17320 5871 17323
rect 6546 17320 6552 17332
rect 5859 17292 6552 17320
rect 5859 17289 5871 17292
rect 5813 17283 5871 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7248 17292 7849 17320
rect 7248 17280 7254 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 9677 17323 9735 17329
rect 9677 17289 9689 17323
rect 9723 17320 9735 17323
rect 10686 17320 10692 17332
rect 9723 17292 10692 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 13446 17280 13452 17332
rect 13504 17280 13510 17332
rect 15473 17323 15531 17329
rect 15473 17320 15485 17323
rect 14844 17292 15485 17320
rect 3252 17224 3358 17252
rect 4706 17212 4712 17264
rect 4764 17252 4770 17264
rect 4764 17224 5304 17252
rect 4764 17212 4770 17224
rect 5276 17196 5304 17224
rect 6178 17212 6184 17264
rect 6236 17212 6242 17264
rect 6288 17224 6769 17252
rect 842 17144 848 17196
rect 900 17184 906 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 900 17156 1409 17184
rect 900 17144 906 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 2406 17144 2412 17196
rect 2464 17184 2470 17196
rect 2593 17187 2651 17193
rect 2593 17184 2605 17187
rect 2464 17156 2605 17184
rect 2464 17144 2470 17156
rect 2593 17153 2605 17156
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 4387 17187 4445 17193
rect 4387 17153 4399 17187
rect 4433 17184 4445 17187
rect 4525 17187 4583 17193
rect 4525 17184 4537 17187
rect 4433 17156 4537 17184
rect 4433 17153 4445 17156
rect 4387 17147 4445 17153
rect 4525 17153 4537 17156
rect 4571 17184 4583 17187
rect 4571 17156 4752 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 2958 17076 2964 17128
rect 3016 17076 3022 17128
rect 4724 17048 4752 17156
rect 4798 17144 4804 17196
rect 4856 17144 4862 17196
rect 5169 17187 5227 17193
rect 5169 17153 5181 17187
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 5184 17116 5212 17147
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5316 17156 5365 17184
rect 5316 17144 5322 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 5902 17184 5908 17196
rect 5675 17156 5908 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 5442 17116 5448 17128
rect 5184 17088 5448 17116
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 5644 17048 5672 17147
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6288 17184 6316 17224
rect 6043 17156 6316 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 6621 17187 6679 17193
rect 6621 17184 6633 17187
rect 6512 17156 6633 17184
rect 6512 17144 6518 17156
rect 6621 17153 6633 17156
rect 6667 17153 6679 17187
rect 6741 17184 6769 17224
rect 7760 17224 8524 17252
rect 7650 17184 7656 17196
rect 6741 17156 7656 17184
rect 6621 17147 6679 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 6362 17076 6368 17128
rect 6420 17076 6426 17128
rect 7760 17116 7788 17224
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 8496 17193 8524 17224
rect 9122 17212 9128 17264
rect 9180 17252 9186 17264
rect 9217 17255 9275 17261
rect 9217 17252 9229 17255
rect 9180 17224 9229 17252
rect 9180 17212 9186 17224
rect 9217 17221 9229 17224
rect 9263 17221 9275 17255
rect 9217 17215 9275 17221
rect 9769 17255 9827 17261
rect 9769 17221 9781 17255
rect 9815 17252 9827 17255
rect 9858 17252 9864 17264
rect 9815 17224 9864 17252
rect 9815 17221 9827 17224
rect 9769 17215 9827 17221
rect 9858 17212 9864 17224
rect 9916 17212 9922 17264
rect 13464 17252 13492 17280
rect 14090 17252 14096 17264
rect 13464 17224 14096 17252
rect 14090 17212 14096 17224
rect 14148 17252 14154 17264
rect 14584 17255 14642 17261
rect 14148 17224 14504 17252
rect 14148 17212 14154 17224
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7892 17156 8125 17184
rect 7892 17144 7898 17156
rect 8113 17153 8125 17156
rect 8159 17184 8171 17187
rect 8481 17187 8539 17193
rect 8159 17156 8432 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7392 17088 8033 17116
rect 4724 17020 5672 17048
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4764 16952 4905 16980
rect 4764 16940 4770 16952
rect 4893 16949 4905 16952
rect 4939 16980 4951 16983
rect 5626 16980 5632 16992
rect 4939 16952 5632 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 6178 16940 6184 16992
rect 6236 16980 6242 16992
rect 7392 16980 7420 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17085 8263 17119
rect 8205 17079 8263 17085
rect 7650 17008 7656 17060
rect 7708 17048 7714 17060
rect 7745 17051 7803 17057
rect 7745 17048 7757 17051
rect 7708 17020 7757 17048
rect 7708 17008 7714 17020
rect 7745 17017 7757 17020
rect 7791 17048 7803 17051
rect 8220 17048 8248 17079
rect 8294 17076 8300 17128
rect 8352 17076 8358 17128
rect 8404 17116 8432 17156
rect 8481 17153 8493 17187
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 9490 17184 9496 17196
rect 8720 17156 9496 17184
rect 8720 17144 8726 17156
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 13998 17184 14004 17196
rect 13096 17156 14004 17184
rect 8754 17116 8760 17128
rect 8404 17088 8760 17116
rect 8754 17076 8760 17088
rect 8812 17116 8818 17128
rect 9309 17119 9367 17125
rect 9309 17116 9321 17119
rect 8812 17088 9321 17116
rect 8812 17076 8818 17088
rect 9309 17085 9321 17088
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 9916 17119 9974 17125
rect 9916 17116 9928 17119
rect 9732 17088 9928 17116
rect 9732 17076 9738 17088
rect 9916 17085 9928 17088
rect 9962 17085 9974 17119
rect 9916 17079 9974 17085
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10594 17116 10600 17128
rect 10183 17088 10600 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 13096 17116 13124 17156
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 14476 17184 14504 17224
rect 14584 17221 14596 17255
rect 14630 17252 14642 17255
rect 14844 17252 14872 17292
rect 15473 17289 15485 17292
rect 15519 17289 15531 17323
rect 15473 17283 15531 17289
rect 17126 17280 17132 17332
rect 17184 17280 17190 17332
rect 18690 17280 18696 17332
rect 18748 17280 18754 17332
rect 18874 17320 18880 17332
rect 18800 17292 18880 17320
rect 14630 17224 14872 17252
rect 14921 17255 14979 17261
rect 14630 17221 14642 17224
rect 14584 17215 14642 17221
rect 14921 17221 14933 17255
rect 14967 17221 14979 17255
rect 14921 17215 14979 17221
rect 14936 17184 14964 17215
rect 15010 17212 15016 17264
rect 15068 17252 15074 17264
rect 15121 17255 15179 17261
rect 15121 17252 15133 17255
rect 15068 17224 15133 17252
rect 15068 17212 15074 17224
rect 15121 17221 15133 17224
rect 15167 17221 15179 17255
rect 15121 17215 15179 17221
rect 17218 17212 17224 17264
rect 17276 17252 17282 17264
rect 18601 17255 18659 17261
rect 17276 17224 18000 17252
rect 17276 17212 17282 17224
rect 14476 17156 14964 17184
rect 15378 17144 15384 17196
rect 15436 17144 15442 17196
rect 15565 17187 15623 17193
rect 15565 17153 15577 17187
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 12667 17088 13124 17116
rect 14829 17119 14887 17125
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 15194 17116 15200 17128
rect 14875 17088 15200 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 15580 17116 15608 17147
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17972 17193 18000 17224
rect 18601 17221 18613 17255
rect 18647 17252 18659 17255
rect 18800 17252 18828 17292
rect 18874 17280 18880 17292
rect 18932 17320 18938 17332
rect 19150 17320 19156 17332
rect 18932 17292 19156 17320
rect 18932 17280 18938 17292
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 19242 17280 19248 17332
rect 19300 17320 19306 17332
rect 19300 17292 19748 17320
rect 19300 17280 19306 17292
rect 19334 17252 19340 17264
rect 18647 17224 18828 17252
rect 18892 17224 19340 17252
rect 18647 17221 18659 17224
rect 18601 17215 18659 17221
rect 18892 17193 18920 17224
rect 19334 17212 19340 17224
rect 19392 17212 19398 17264
rect 19720 17261 19748 17292
rect 20806 17280 20812 17332
rect 20864 17280 20870 17332
rect 21450 17320 21456 17332
rect 21376 17292 21456 17320
rect 19705 17255 19763 17261
rect 19705 17221 19717 17255
rect 19751 17221 19763 17255
rect 19705 17215 19763 17221
rect 19886 17212 19892 17264
rect 19944 17212 19950 17264
rect 21376 17261 21404 17292
rect 21450 17280 21456 17292
rect 21508 17320 21514 17332
rect 21913 17323 21971 17329
rect 21913 17320 21925 17323
rect 21508 17292 21925 17320
rect 21508 17280 21514 17292
rect 21913 17289 21925 17292
rect 21959 17289 21971 17323
rect 21913 17283 21971 17289
rect 23937 17323 23995 17329
rect 23937 17289 23949 17323
rect 23983 17320 23995 17323
rect 24486 17320 24492 17332
rect 23983 17292 24492 17320
rect 23983 17289 23995 17292
rect 23937 17283 23995 17289
rect 24486 17280 24492 17292
rect 24544 17280 24550 17332
rect 24578 17280 24584 17332
rect 24636 17320 24642 17332
rect 24636 17292 24992 17320
rect 24636 17280 24642 17292
rect 20625 17255 20683 17261
rect 20625 17252 20637 17255
rect 20364 17224 20637 17252
rect 19485 17196 19543 17199
rect 20364 17196 20392 17224
rect 20625 17221 20637 17224
rect 20671 17221 20683 17255
rect 20625 17215 20683 17221
rect 21361 17255 21419 17261
rect 21361 17221 21373 17255
rect 21407 17221 21419 17255
rect 21361 17215 21419 17221
rect 21652 17224 22048 17252
rect 17957 17187 18015 17193
rect 17957 17153 17969 17187
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 18969 17147 19027 17153
rect 15304 17088 15608 17116
rect 17313 17119 17371 17125
rect 8662 17048 8668 17060
rect 7791 17020 8668 17048
rect 7791 17017 7803 17020
rect 7745 17011 7803 17017
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 10045 17051 10103 17057
rect 10045 17017 10057 17051
rect 10091 17048 10103 17051
rect 12345 17051 12403 17057
rect 12345 17048 12357 17051
rect 10091 17020 12357 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 12345 17017 12357 17020
rect 12391 17017 12403 17051
rect 13814 17048 13820 17060
rect 12345 17011 12403 17017
rect 12820 17020 13820 17048
rect 6236 16952 7420 16980
rect 6236 16940 6242 16952
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 8573 16983 8631 16989
rect 8573 16980 8585 16983
rect 7616 16952 8585 16980
rect 7616 16940 7622 16952
rect 8573 16949 8585 16952
rect 8619 16949 8631 16983
rect 8573 16943 8631 16949
rect 9398 16940 9404 16992
rect 9456 16940 9462 16992
rect 10410 16940 10416 16992
rect 10468 16940 10474 16992
rect 12820 16989 12848 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 15304 16992 15332 17088
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17770 17116 17776 17128
rect 17359 17088 17776 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17770 17076 17776 17088
rect 17828 17076 17834 17128
rect 18984 17048 19012 17147
rect 19058 17144 19064 17196
rect 19116 17144 19122 17196
rect 19150 17144 19156 17196
rect 19208 17193 19214 17196
rect 19208 17187 19237 17193
rect 19225 17153 19237 17187
rect 19208 17147 19237 17153
rect 19208 17144 19214 17147
rect 19426 17144 19432 17196
rect 19484 17193 19543 17196
rect 19484 17159 19497 17193
rect 19531 17159 19543 17193
rect 19484 17153 19543 17159
rect 19484 17144 19490 17153
rect 19610 17144 19616 17196
rect 19668 17144 19674 17196
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 20128 17156 20177 17184
rect 20128 17144 20134 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 20346 17144 20352 17196
rect 20404 17144 20410 17196
rect 20441 17187 20499 17193
rect 20441 17153 20453 17187
rect 20487 17184 20499 17187
rect 20990 17184 20996 17196
rect 20487 17156 20996 17184
rect 20487 17153 20499 17156
rect 20441 17147 20499 17153
rect 19334 17076 19340 17128
rect 19392 17076 19398 17128
rect 19981 17051 20039 17057
rect 19981 17048 19993 17051
rect 18984 17020 19472 17048
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16949 12863 16983
rect 12805 16943 12863 16949
rect 13906 16940 13912 16992
rect 13964 16980 13970 16992
rect 14182 16980 14188 16992
rect 13964 16952 14188 16980
rect 13964 16940 13970 16952
rect 14182 16940 14188 16952
rect 14240 16940 14246 16992
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 14608 16952 15117 16980
rect 14608 16940 14614 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 15105 16943 15163 16949
rect 15286 16940 15292 16992
rect 15344 16940 15350 16992
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 15620 16952 16681 16980
rect 15620 16940 15626 16952
rect 16669 16949 16681 16952
rect 16715 16949 16727 16983
rect 19444 16980 19472 17020
rect 19628 17020 19993 17048
rect 19628 16980 19656 17020
rect 19981 17017 19993 17020
rect 20027 17017 20039 17051
rect 19981 17011 20039 17017
rect 20088 17020 20300 17048
rect 19444 16952 19656 16980
rect 19889 16983 19947 16989
rect 16669 16943 16727 16949
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20088 16980 20116 17020
rect 19935 16952 20116 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20162 16940 20168 16992
rect 20220 16940 20226 16992
rect 20272 16980 20300 17020
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 20622 17048 20628 17060
rect 20404 17020 20628 17048
rect 20404 17008 20410 17020
rect 20622 17008 20628 17020
rect 20680 17008 20686 17060
rect 20732 16980 20760 17156
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17184 21511 17187
rect 21542 17184 21548 17196
rect 21499 17156 21548 17184
rect 21499 17153 21511 17156
rect 21453 17147 21511 17153
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 21652 17193 21680 17224
rect 22020 17196 22048 17224
rect 23474 17212 23480 17264
rect 23532 17212 23538 17264
rect 23845 17255 23903 17261
rect 23845 17221 23857 17255
rect 23891 17252 23903 17255
rect 24964 17252 24992 17292
rect 25130 17280 25136 17332
rect 25188 17320 25194 17332
rect 25593 17323 25651 17329
rect 25593 17320 25605 17323
rect 25188 17292 25605 17320
rect 25188 17280 25194 17292
rect 25593 17289 25605 17292
rect 25639 17289 25651 17323
rect 25593 17283 25651 17289
rect 27338 17280 27344 17332
rect 27396 17280 27402 17332
rect 29178 17320 29184 17332
rect 28185 17292 29184 17320
rect 25225 17255 25283 17261
rect 25225 17252 25237 17255
rect 23891 17224 24808 17252
rect 24964 17224 25237 17252
rect 23891 17221 23903 17224
rect 23845 17215 23903 17221
rect 21637 17187 21695 17193
rect 21637 17153 21649 17187
rect 21683 17153 21695 17187
rect 21637 17147 21695 17153
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 21560 17116 21588 17144
rect 21836 17116 21864 17147
rect 22002 17144 22008 17196
rect 22060 17144 22066 17196
rect 21560 17088 21864 17116
rect 23492 17116 23520 17212
rect 24780 17196 24808 17224
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17184 23719 17187
rect 24118 17184 24124 17196
rect 23707 17156 24124 17184
rect 23707 17153 23719 17156
rect 23661 17147 23719 17153
rect 24118 17144 24124 17156
rect 24176 17144 24182 17196
rect 24394 17144 24400 17196
rect 24452 17144 24458 17196
rect 24581 17187 24639 17193
rect 24581 17153 24593 17187
rect 24627 17153 24639 17187
rect 24581 17147 24639 17153
rect 24305 17119 24363 17125
rect 24305 17116 24317 17119
rect 23492 17088 24317 17116
rect 24305 17085 24317 17088
rect 24351 17085 24363 17119
rect 24305 17079 24363 17085
rect 21085 17051 21143 17057
rect 21085 17017 21097 17051
rect 21131 17048 21143 17051
rect 21266 17048 21272 17060
rect 21131 17020 21272 17048
rect 21131 17017 21143 17020
rect 21085 17011 21143 17017
rect 21266 17008 21272 17020
rect 21324 17048 21330 17060
rect 21545 17051 21603 17057
rect 21545 17048 21557 17051
rect 21324 17020 21557 17048
rect 21324 17008 21330 17020
rect 21545 17017 21557 17020
rect 21591 17017 21603 17051
rect 21545 17011 21603 17017
rect 24026 17008 24032 17060
rect 24084 17048 24090 17060
rect 24213 17051 24271 17057
rect 24213 17048 24225 17051
rect 24084 17020 24225 17048
rect 24084 17008 24090 17020
rect 24213 17017 24225 17020
rect 24259 17048 24271 17051
rect 24596 17048 24624 17147
rect 24762 17144 24768 17196
rect 24820 17144 24826 17196
rect 24946 17144 24952 17196
rect 25004 17144 25010 17196
rect 25148 17193 25176 17224
rect 25225 17221 25237 17224
rect 25271 17221 25283 17255
rect 25225 17215 25283 17221
rect 25409 17255 25467 17261
rect 25409 17221 25421 17255
rect 25455 17252 25467 17255
rect 25682 17252 25688 17264
rect 25455 17224 25688 17252
rect 25455 17221 25467 17224
rect 25409 17215 25467 17221
rect 25682 17212 25688 17224
rect 25740 17212 25746 17264
rect 27157 17255 27215 17261
rect 27157 17252 27169 17255
rect 26620 17224 27169 17252
rect 25133 17187 25191 17193
rect 25133 17153 25145 17187
rect 25179 17184 25191 17187
rect 25179 17156 25213 17184
rect 25179 17153 25191 17156
rect 25133 17147 25191 17153
rect 26418 17144 26424 17196
rect 26476 17184 26482 17196
rect 26620 17184 26648 17224
rect 27157 17221 27169 17224
rect 27203 17252 27215 17255
rect 27246 17252 27252 17264
rect 27203 17224 27252 17252
rect 27203 17221 27215 17224
rect 27157 17215 27215 17221
rect 27246 17212 27252 17224
rect 27304 17212 27310 17264
rect 26476 17156 26648 17184
rect 26973 17187 27031 17193
rect 26476 17144 26482 17156
rect 26973 17153 26985 17187
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 24670 17076 24676 17128
rect 24728 17076 24734 17128
rect 24854 17076 24860 17128
rect 24912 17116 24918 17128
rect 26988 17116 27016 17147
rect 27706 17144 27712 17196
rect 27764 17144 27770 17196
rect 27890 17144 27896 17196
rect 27948 17144 27954 17196
rect 28185 17193 28213 17292
rect 29178 17280 29184 17292
rect 29236 17280 29242 17332
rect 31938 17280 31944 17332
rect 31996 17320 32002 17332
rect 32125 17323 32183 17329
rect 32125 17320 32137 17323
rect 31996 17292 32137 17320
rect 31996 17280 32002 17292
rect 32125 17289 32137 17292
rect 32171 17289 32183 17323
rect 32125 17283 32183 17289
rect 32493 17323 32551 17329
rect 32493 17289 32505 17323
rect 32539 17320 32551 17323
rect 32674 17320 32680 17332
rect 32539 17292 32680 17320
rect 32539 17289 32551 17292
rect 32493 17283 32551 17289
rect 32674 17280 32680 17292
rect 32732 17320 32738 17332
rect 32769 17323 32827 17329
rect 32769 17320 32781 17323
rect 32732 17292 32781 17320
rect 32732 17280 32738 17292
rect 32769 17289 32781 17292
rect 32815 17289 32827 17323
rect 32769 17283 32827 17289
rect 34701 17323 34759 17329
rect 34701 17289 34713 17323
rect 34747 17320 34759 17323
rect 34974 17320 34980 17332
rect 34747 17292 34980 17320
rect 34747 17289 34759 17292
rect 34701 17283 34759 17289
rect 34974 17280 34980 17292
rect 35032 17280 35038 17332
rect 35069 17323 35127 17329
rect 35069 17289 35081 17323
rect 35115 17320 35127 17323
rect 36538 17320 36544 17332
rect 35115 17292 36544 17320
rect 35115 17289 35127 17292
rect 35069 17283 35127 17289
rect 36538 17280 36544 17292
rect 36596 17280 36602 17332
rect 36630 17280 36636 17332
rect 36688 17320 36694 17332
rect 38197 17323 38255 17329
rect 38197 17320 38209 17323
rect 36688 17292 38209 17320
rect 36688 17280 36694 17292
rect 38197 17289 38209 17292
rect 38243 17289 38255 17323
rect 40037 17323 40095 17329
rect 40037 17320 40049 17323
rect 38197 17283 38255 17289
rect 39408 17292 40049 17320
rect 28905 17255 28963 17261
rect 28905 17252 28917 17255
rect 28460 17224 28917 17252
rect 28460 17196 28488 17224
rect 28905 17221 28917 17224
rect 28951 17221 28963 17255
rect 28905 17215 28963 17221
rect 32953 17255 33011 17261
rect 32953 17221 32965 17255
rect 32999 17252 33011 17255
rect 33686 17252 33692 17264
rect 32999 17224 33692 17252
rect 32999 17221 33011 17224
rect 32953 17215 33011 17221
rect 33686 17212 33692 17224
rect 33744 17212 33750 17264
rect 34790 17212 34796 17264
rect 34848 17252 34854 17264
rect 35161 17255 35219 17261
rect 35161 17252 35173 17255
rect 34848 17224 35173 17252
rect 34848 17212 34854 17224
rect 35161 17221 35173 17224
rect 35207 17221 35219 17255
rect 35161 17215 35219 17221
rect 38102 17212 38108 17264
rect 38160 17252 38166 17264
rect 39408 17261 39436 17292
rect 40037 17289 40049 17292
rect 40083 17289 40095 17323
rect 40037 17283 40095 17289
rect 40144 17292 40908 17320
rect 39301 17255 39359 17261
rect 39301 17252 39313 17255
rect 38160 17224 39313 17252
rect 38160 17212 38166 17224
rect 39301 17221 39313 17224
rect 39347 17221 39359 17255
rect 39301 17215 39359 17221
rect 39393 17255 39451 17261
rect 39393 17221 39405 17255
rect 39439 17221 39451 17255
rect 39393 17215 39451 17221
rect 39850 17212 39856 17264
rect 39908 17252 39914 17264
rect 40144 17261 40172 17292
rect 40129 17255 40187 17261
rect 40129 17252 40141 17255
rect 39908 17224 40141 17252
rect 39908 17212 39914 17224
rect 40129 17221 40141 17224
rect 40175 17221 40187 17255
rect 40129 17215 40187 17221
rect 40310 17212 40316 17264
rect 40368 17252 40374 17264
rect 40368 17224 40632 17252
rect 40368 17212 40374 17224
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28169 17187 28227 17193
rect 28169 17153 28181 17187
rect 28215 17153 28227 17187
rect 28169 17147 28227 17153
rect 27154 17116 27160 17128
rect 24912 17088 26924 17116
rect 26988 17088 27160 17116
rect 24912 17076 24918 17088
rect 24946 17048 24952 17060
rect 24259 17020 24348 17048
rect 24596 17020 24952 17048
rect 24259 17017 24271 17020
rect 24213 17011 24271 17017
rect 20272 16952 20760 16980
rect 20898 16940 20904 16992
rect 20956 16940 20962 16992
rect 24320 16980 24348 17020
rect 24946 17008 24952 17020
rect 25004 17008 25010 17060
rect 26896 17048 26924 17088
rect 27154 17076 27160 17088
rect 27212 17076 27218 17128
rect 27801 17119 27859 17125
rect 27801 17085 27813 17119
rect 27847 17116 27859 17119
rect 28000 17116 28028 17147
rect 28442 17144 28448 17196
rect 28500 17144 28506 17196
rect 28534 17144 28540 17196
rect 28592 17184 28598 17196
rect 28721 17187 28779 17193
rect 28721 17184 28733 17187
rect 28592 17156 28733 17184
rect 28592 17144 28598 17156
rect 28721 17153 28733 17156
rect 28767 17153 28779 17187
rect 28721 17147 28779 17153
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 29454 17184 29460 17196
rect 29052 17156 29460 17184
rect 29052 17144 29058 17156
rect 29454 17144 29460 17156
rect 29512 17144 29518 17196
rect 30929 17187 30987 17193
rect 30929 17153 30941 17187
rect 30975 17153 30987 17187
rect 30929 17147 30987 17153
rect 29178 17116 29184 17128
rect 27847 17088 29184 17116
rect 27847 17085 27859 17088
rect 27801 17079 27859 17085
rect 29178 17076 29184 17088
rect 29236 17076 29242 17128
rect 30834 17076 30840 17128
rect 30892 17076 30898 17128
rect 30944 17116 30972 17147
rect 32122 17144 32128 17196
rect 32180 17184 32186 17196
rect 32309 17187 32367 17193
rect 32309 17184 32321 17187
rect 32180 17156 32321 17184
rect 32180 17144 32186 17156
rect 32309 17153 32321 17156
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 32585 17187 32643 17193
rect 32585 17153 32597 17187
rect 32631 17184 32643 17187
rect 33042 17184 33048 17196
rect 32631 17156 33048 17184
rect 32631 17153 32643 17156
rect 32585 17147 32643 17153
rect 33042 17144 33048 17156
rect 33100 17144 33106 17196
rect 33137 17187 33195 17193
rect 33137 17153 33149 17187
rect 33183 17184 33195 17187
rect 33410 17184 33416 17196
rect 33183 17156 33416 17184
rect 33183 17153 33195 17156
rect 33137 17147 33195 17153
rect 33410 17144 33416 17156
rect 33468 17144 33474 17196
rect 38470 17184 38476 17196
rect 38028 17156 38476 17184
rect 31389 17119 31447 17125
rect 31389 17116 31401 17119
rect 30944 17088 31401 17116
rect 31389 17085 31401 17088
rect 31435 17085 31447 17119
rect 31389 17079 31447 17085
rect 31662 17076 31668 17128
rect 31720 17116 31726 17128
rect 31849 17119 31907 17125
rect 31849 17116 31861 17119
rect 31720 17088 31861 17116
rect 31720 17076 31726 17088
rect 31849 17085 31861 17088
rect 31895 17116 31907 17119
rect 33226 17116 33232 17128
rect 31895 17088 33232 17116
rect 31895 17085 31907 17088
rect 31849 17079 31907 17085
rect 33226 17076 33232 17088
rect 33284 17076 33290 17128
rect 35345 17119 35403 17125
rect 35345 17085 35357 17119
rect 35391 17116 35403 17119
rect 37090 17116 37096 17128
rect 35391 17088 37096 17116
rect 35391 17085 35403 17088
rect 35345 17079 35403 17085
rect 37090 17076 37096 17088
rect 37148 17076 37154 17128
rect 38028 17125 38056 17156
rect 38470 17144 38476 17156
rect 38528 17144 38534 17196
rect 39163 17187 39221 17193
rect 39163 17184 39175 17187
rect 38764 17156 39175 17184
rect 38764 17128 38792 17156
rect 39163 17153 39175 17156
rect 39209 17153 39221 17187
rect 39163 17147 39221 17153
rect 39485 17187 39543 17193
rect 39485 17153 39497 17187
rect 39531 17153 39543 17187
rect 39485 17147 39543 17153
rect 40037 17187 40095 17193
rect 40037 17153 40049 17187
rect 40083 17184 40095 17187
rect 40218 17184 40224 17196
rect 40083 17156 40224 17184
rect 40083 17153 40095 17156
rect 40037 17147 40095 17153
rect 38013 17119 38071 17125
rect 38013 17085 38025 17119
rect 38059 17085 38071 17119
rect 38013 17079 38071 17085
rect 38105 17119 38163 17125
rect 38105 17085 38117 17119
rect 38151 17116 38163 17119
rect 38746 17116 38752 17128
rect 38151 17088 38752 17116
rect 38151 17085 38163 17088
rect 38105 17079 38163 17085
rect 38746 17076 38752 17088
rect 38804 17076 38810 17128
rect 39025 17119 39083 17125
rect 39025 17085 39037 17119
rect 39071 17085 39083 17119
rect 39500 17116 39528 17147
rect 40218 17144 40224 17156
rect 40276 17184 40282 17196
rect 40604 17193 40632 17224
rect 40770 17212 40776 17264
rect 40828 17212 40834 17264
rect 40589 17187 40647 17193
rect 40276 17156 40540 17184
rect 40276 17144 40282 17156
rect 40405 17119 40463 17125
rect 40405 17116 40417 17119
rect 39500 17088 40417 17116
rect 39025 17079 39083 17085
rect 40405 17085 40417 17088
rect 40451 17085 40463 17119
rect 40512 17116 40540 17156
rect 40589 17153 40601 17187
rect 40635 17153 40647 17187
rect 40589 17147 40647 17153
rect 40788 17116 40816 17212
rect 40880 17193 40908 17292
rect 41800 17224 42196 17252
rect 41800 17196 41828 17224
rect 42168 17196 42196 17224
rect 40865 17187 40923 17193
rect 40865 17153 40877 17187
rect 40911 17153 40923 17187
rect 40865 17147 40923 17153
rect 40512 17088 40816 17116
rect 40880 17116 40908 17147
rect 41782 17144 41788 17196
rect 41840 17144 41846 17196
rect 41874 17144 41880 17196
rect 41932 17184 41938 17196
rect 41969 17187 42027 17193
rect 41969 17184 41981 17187
rect 41932 17156 41981 17184
rect 41932 17144 41938 17156
rect 41969 17153 41981 17156
rect 42015 17153 42027 17187
rect 41969 17147 42027 17153
rect 42150 17144 42156 17196
rect 42208 17144 42214 17196
rect 42061 17119 42119 17125
rect 42061 17116 42073 17119
rect 40880 17088 42073 17116
rect 40405 17079 40463 17085
rect 42061 17085 42073 17088
rect 42107 17085 42119 17119
rect 42061 17079 42119 17085
rect 28261 17051 28319 17057
rect 28261 17048 28273 17051
rect 26896 17020 28273 17048
rect 28261 17017 28273 17020
rect 28307 17017 28319 17051
rect 28261 17011 28319 17017
rect 28353 17051 28411 17057
rect 28353 17017 28365 17051
rect 28399 17048 28411 17051
rect 28994 17048 29000 17060
rect 28399 17020 29000 17048
rect 28399 17017 28411 17020
rect 28353 17011 28411 17017
rect 24670 16980 24676 16992
rect 24320 16952 24676 16980
rect 24670 16940 24676 16952
rect 24728 16940 24734 16992
rect 25777 16983 25835 16989
rect 25777 16949 25789 16983
rect 25823 16980 25835 16983
rect 25958 16980 25964 16992
rect 25823 16952 25964 16980
rect 25823 16949 25835 16952
rect 25777 16943 25835 16949
rect 25958 16940 25964 16952
rect 26016 16940 26022 16992
rect 28276 16980 28304 17011
rect 28994 17008 29000 17020
rect 29052 17008 29058 17060
rect 29086 17008 29092 17060
rect 29144 17048 29150 17060
rect 29365 17051 29423 17057
rect 29365 17048 29377 17051
rect 29144 17020 29377 17048
rect 29144 17008 29150 17020
rect 29365 17017 29377 17020
rect 29411 17017 29423 17051
rect 29365 17011 29423 17017
rect 31297 17051 31355 17057
rect 31297 17017 31309 17051
rect 31343 17048 31355 17051
rect 31478 17048 31484 17060
rect 31343 17020 31484 17048
rect 31343 17017 31355 17020
rect 31297 17011 31355 17017
rect 31478 17008 31484 17020
rect 31536 17008 31542 17060
rect 31573 17051 31631 17057
rect 31573 17017 31585 17051
rect 31619 17048 31631 17051
rect 31754 17048 31760 17060
rect 31619 17020 31760 17048
rect 31619 17017 31631 17020
rect 31573 17011 31631 17017
rect 31754 17008 31760 17020
rect 31812 17008 31818 17060
rect 32306 17008 32312 17060
rect 32364 17048 32370 17060
rect 38838 17048 38844 17060
rect 32364 17020 38844 17048
rect 32364 17008 32370 17020
rect 38838 17008 38844 17020
rect 38896 17048 38902 17060
rect 39040 17048 39068 17079
rect 38896 17020 39068 17048
rect 38896 17008 38902 17020
rect 28534 16980 28540 16992
rect 28276 16952 28540 16980
rect 28534 16940 28540 16952
rect 28592 16940 28598 16992
rect 28626 16940 28632 16992
rect 28684 16940 28690 16992
rect 28902 16940 28908 16992
rect 28960 16980 28966 16992
rect 29273 16983 29331 16989
rect 29273 16980 29285 16983
rect 28960 16952 29285 16980
rect 28960 16940 28966 16952
rect 29273 16949 29285 16952
rect 29319 16949 29331 16983
rect 31772 16980 31800 17008
rect 32582 16980 32588 16992
rect 31772 16952 32588 16980
rect 29273 16943 29331 16949
rect 32582 16940 32588 16952
rect 32640 16940 32646 16992
rect 38378 16940 38384 16992
rect 38436 16980 38442 16992
rect 38565 16983 38623 16989
rect 38565 16980 38577 16983
rect 38436 16952 38577 16980
rect 38436 16940 38442 16952
rect 38565 16949 38577 16952
rect 38611 16949 38623 16983
rect 38565 16943 38623 16949
rect 38654 16940 38660 16992
rect 38712 16980 38718 16992
rect 39669 16983 39727 16989
rect 39669 16980 39681 16983
rect 38712 16952 39681 16980
rect 38712 16940 38718 16952
rect 39669 16949 39681 16952
rect 39715 16949 39727 16983
rect 39669 16943 39727 16949
rect 41230 16940 41236 16992
rect 41288 16940 41294 16992
rect 1104 16890 42504 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 42504 16890
rect 1104 16816 42504 16838
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3016 16748 3801 16776
rect 3016 16736 3022 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 5350 16736 5356 16788
rect 5408 16736 5414 16788
rect 7558 16776 7564 16788
rect 7116 16748 7564 16776
rect 7116 16708 7144 16748
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8754 16736 8760 16788
rect 8812 16736 8818 16788
rect 9398 16736 9404 16788
rect 9456 16776 9462 16788
rect 9493 16779 9551 16785
rect 9493 16776 9505 16779
rect 9456 16748 9505 16776
rect 9456 16736 9462 16748
rect 9493 16745 9505 16748
rect 9539 16745 9551 16779
rect 9493 16739 9551 16745
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12805 16779 12863 16785
rect 12805 16776 12817 16779
rect 12768 16748 12817 16776
rect 12768 16736 12774 16748
rect 12805 16745 12817 16748
rect 12851 16745 12863 16779
rect 12805 16739 12863 16745
rect 7024 16680 7144 16708
rect 12820 16708 12848 16739
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 14093 16779 14151 16785
rect 14093 16776 14105 16779
rect 13872 16748 14105 16776
rect 13872 16736 13878 16748
rect 14093 16745 14105 16748
rect 14139 16745 14151 16779
rect 14093 16739 14151 16745
rect 14550 16736 14556 16788
rect 14608 16736 14614 16788
rect 17034 16736 17040 16788
rect 17092 16776 17098 16788
rect 17129 16779 17187 16785
rect 17129 16776 17141 16779
rect 17092 16748 17141 16776
rect 17092 16736 17098 16748
rect 17129 16745 17141 16748
rect 17175 16745 17187 16779
rect 17129 16739 17187 16745
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 20162 16776 20168 16788
rect 19392 16748 20168 16776
rect 19392 16736 19398 16748
rect 20162 16736 20168 16748
rect 20220 16736 20226 16788
rect 24946 16776 24952 16788
rect 24044 16748 24952 16776
rect 12820 16680 13768 16708
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 7024 16649 7052 16680
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3292 16612 4353 16640
rect 3292 16600 3298 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 9953 16643 10011 16649
rect 9953 16609 9965 16643
rect 9999 16640 10011 16643
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 9999 16612 12449 16640
rect 9999 16609 10011 16612
rect 9953 16603 10011 16609
rect 12437 16609 12449 16612
rect 12483 16640 12495 16643
rect 12802 16640 12808 16652
rect 12483 16612 12808 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13740 16649 13768 16680
rect 17954 16668 17960 16720
rect 18012 16708 18018 16720
rect 24044 16717 24072 16748
rect 24946 16736 24952 16748
rect 25004 16776 25010 16788
rect 25133 16779 25191 16785
rect 25133 16776 25145 16779
rect 25004 16748 25145 16776
rect 25004 16736 25010 16748
rect 25133 16745 25145 16748
rect 25179 16745 25191 16779
rect 25133 16739 25191 16745
rect 26329 16779 26387 16785
rect 26329 16745 26341 16779
rect 26375 16776 26387 16779
rect 27062 16776 27068 16788
rect 26375 16748 27068 16776
rect 26375 16745 26387 16748
rect 26329 16739 26387 16745
rect 27062 16736 27068 16748
rect 27120 16736 27126 16788
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 29086 16776 29092 16788
rect 28960 16748 29092 16776
rect 28960 16736 28966 16748
rect 29086 16736 29092 16748
rect 29144 16736 29150 16788
rect 31754 16736 31760 16788
rect 31812 16776 31818 16788
rect 31849 16779 31907 16785
rect 31849 16776 31861 16779
rect 31812 16748 31861 16776
rect 31812 16736 31818 16748
rect 31849 16745 31861 16748
rect 31895 16745 31907 16779
rect 31849 16739 31907 16745
rect 32122 16736 32128 16788
rect 32180 16776 32186 16788
rect 32306 16776 32312 16788
rect 32180 16748 32312 16776
rect 32180 16736 32186 16748
rect 32306 16736 32312 16748
rect 32364 16736 32370 16788
rect 33226 16736 33232 16788
rect 33284 16736 33290 16788
rect 36630 16736 36636 16788
rect 36688 16776 36694 16788
rect 36909 16779 36967 16785
rect 36909 16776 36921 16779
rect 36688 16748 36921 16776
rect 36688 16736 36694 16748
rect 36909 16745 36921 16748
rect 36955 16745 36967 16779
rect 36909 16739 36967 16745
rect 38746 16736 38752 16788
rect 38804 16736 38810 16788
rect 42150 16736 42156 16788
rect 42208 16736 42214 16788
rect 24029 16711 24087 16717
rect 18012 16680 23704 16708
rect 18012 16668 18018 16680
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 13771 16612 14596 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 4856 16544 5089 16572
rect 4856 16532 4862 16544
rect 5077 16541 5089 16544
rect 5123 16541 5135 16575
rect 5077 16535 5135 16541
rect 6914 16532 6920 16584
rect 6972 16532 6978 16584
rect 7374 16532 7380 16584
rect 7432 16532 7438 16584
rect 9490 16532 9496 16584
rect 9548 16532 9554 16584
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 11330 16572 11336 16584
rect 9907 16544 11336 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 11330 16532 11336 16544
rect 11388 16572 11394 16584
rect 12529 16575 12587 16581
rect 12529 16572 12541 16575
rect 11388 16544 12541 16572
rect 11388 16532 11394 16544
rect 12529 16541 12541 16544
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 13814 16572 13820 16584
rect 12943 16544 13820 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 5169 16507 5227 16513
rect 5169 16504 5181 16507
rect 4672 16476 5181 16504
rect 4672 16464 4678 16476
rect 5169 16473 5181 16476
rect 5215 16473 5227 16507
rect 5169 16467 5227 16473
rect 5350 16464 5356 16516
rect 5408 16504 5414 16516
rect 5718 16504 5724 16516
rect 5408 16476 5724 16504
rect 5408 16464 5414 16476
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 7622 16507 7680 16513
rect 7622 16504 7634 16507
rect 7300 16476 7634 16504
rect 7300 16445 7328 16476
rect 7622 16473 7634 16476
rect 7668 16473 7680 16507
rect 7622 16467 7680 16473
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 12912 16504 12940 16535
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14568 16581 14596 16612
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15289 16643 15347 16649
rect 15289 16640 15301 16643
rect 15252 16612 15301 16640
rect 15252 16600 15258 16612
rect 15289 16609 15301 16612
rect 15335 16609 15347 16643
rect 15289 16603 15347 16609
rect 15562 16600 15568 16652
rect 15620 16600 15626 16652
rect 18524 16649 18552 16680
rect 18509 16643 18567 16649
rect 18509 16609 18521 16643
rect 18555 16609 18567 16643
rect 19426 16640 19432 16652
rect 18509 16603 18567 16609
rect 18800 16612 19432 16640
rect 14237 16575 14295 16581
rect 14237 16572 14249 16575
rect 14148 16544 14249 16572
rect 14148 16532 14154 16544
rect 14237 16541 14249 16544
rect 14283 16541 14295 16575
rect 14237 16535 14295 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 13906 16504 13912 16516
rect 12032 16476 12940 16504
rect 13096 16476 13912 16504
rect 12032 16464 12038 16476
rect 7285 16439 7343 16445
rect 7285 16405 7297 16439
rect 7331 16405 7343 16439
rect 7285 16399 7343 16405
rect 9309 16439 9367 16445
rect 9309 16405 9321 16439
rect 9355 16436 9367 16439
rect 9858 16436 9864 16448
rect 9355 16408 9864 16436
rect 9355 16405 9367 16408
rect 9309 16399 9367 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 13096 16445 13124 16476
rect 13906 16464 13912 16476
rect 13964 16464 13970 16516
rect 14384 16504 14412 16535
rect 14734 16504 14740 16516
rect 14384 16476 14740 16504
rect 13081 16439 13139 16445
rect 13081 16405 13093 16439
rect 13127 16405 13139 16439
rect 13081 16399 13139 16405
rect 13170 16396 13176 16448
rect 13228 16396 13234 16448
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14384 16436 14412 16476
rect 14734 16464 14740 16476
rect 14792 16464 14798 16516
rect 16298 16464 16304 16516
rect 16356 16464 16362 16516
rect 17788 16504 17816 16535
rect 17862 16532 17868 16584
rect 17920 16532 17926 16584
rect 18800 16581 18828 16612
rect 19426 16600 19432 16612
rect 19484 16640 19490 16652
rect 19610 16640 19616 16652
rect 19484 16612 19616 16640
rect 19484 16600 19490 16612
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 20806 16600 20812 16652
rect 20864 16600 20870 16652
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16541 18843 16575
rect 18785 16535 18843 16541
rect 18969 16575 19027 16581
rect 18969 16541 18981 16575
rect 19015 16572 19027 16575
rect 19150 16572 19156 16584
rect 19015 16544 19156 16572
rect 19015 16541 19027 16544
rect 18969 16535 19027 16541
rect 18984 16504 19012 16535
rect 19150 16532 19156 16544
rect 19208 16532 19214 16584
rect 20898 16532 20904 16584
rect 20956 16532 20962 16584
rect 23676 16572 23704 16680
rect 24029 16677 24041 16711
rect 24075 16677 24087 16711
rect 24029 16671 24087 16677
rect 24320 16680 26372 16708
rect 24320 16572 24348 16680
rect 26344 16652 26372 16680
rect 28626 16668 28632 16720
rect 28684 16668 28690 16720
rect 28718 16668 28724 16720
rect 28776 16668 28782 16720
rect 28810 16668 28816 16720
rect 28868 16708 28874 16720
rect 28868 16680 29113 16708
rect 28868 16668 28874 16680
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16640 24731 16643
rect 24762 16640 24768 16652
rect 24719 16612 24768 16640
rect 24719 16609 24731 16612
rect 24673 16603 24731 16609
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 24854 16600 24860 16652
rect 24912 16640 24918 16652
rect 24912 16612 25084 16640
rect 24912 16600 24918 16612
rect 25056 16581 25084 16612
rect 26326 16600 26332 16652
rect 26384 16600 26390 16652
rect 28353 16643 28411 16649
rect 28353 16609 28365 16643
rect 28399 16640 28411 16643
rect 28442 16640 28448 16652
rect 28399 16612 28448 16640
rect 28399 16609 28411 16612
rect 28353 16603 28411 16609
rect 28442 16600 28448 16612
rect 28500 16600 28506 16652
rect 29085 16640 29113 16680
rect 29178 16668 29184 16720
rect 29236 16708 29242 16720
rect 29641 16711 29699 16717
rect 29641 16708 29653 16711
rect 29236 16680 29653 16708
rect 29236 16668 29242 16680
rect 29641 16677 29653 16680
rect 29687 16677 29699 16711
rect 29641 16671 29699 16677
rect 31864 16680 33272 16708
rect 31864 16652 31892 16680
rect 29085 16612 29132 16640
rect 24581 16575 24639 16581
rect 24581 16572 24593 16575
rect 23676 16544 24348 16572
rect 24412 16544 24593 16572
rect 17788 16476 19012 16504
rect 23753 16507 23811 16513
rect 13872 16408 14412 16436
rect 17037 16439 17095 16445
rect 13872 16396 13878 16408
rect 17037 16405 17049 16439
rect 17083 16436 17095 16439
rect 17788 16436 17816 16476
rect 23753 16473 23765 16507
rect 23799 16504 23811 16507
rect 24026 16504 24032 16516
rect 23799 16476 24032 16504
rect 23799 16473 23811 16476
rect 23753 16467 23811 16473
rect 24026 16464 24032 16476
rect 24084 16464 24090 16516
rect 17083 16408 17816 16436
rect 17083 16405 17095 16408
rect 17037 16399 17095 16405
rect 18782 16396 18788 16448
rect 18840 16436 18846 16448
rect 20070 16436 20076 16448
rect 18840 16408 20076 16436
rect 18840 16396 18846 16408
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20438 16396 20444 16448
rect 20496 16436 20502 16448
rect 20533 16439 20591 16445
rect 20533 16436 20545 16439
rect 20496 16408 20545 16436
rect 20496 16396 20502 16408
rect 20533 16405 20545 16408
rect 20579 16405 20591 16439
rect 20533 16399 20591 16405
rect 24213 16439 24271 16445
rect 24213 16405 24225 16439
rect 24259 16436 24271 16439
rect 24412 16436 24440 16544
rect 24581 16541 24593 16544
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 25041 16575 25099 16581
rect 25041 16541 25053 16575
rect 25087 16541 25099 16575
rect 25041 16535 25099 16541
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 25590 16532 25596 16584
rect 25648 16572 25654 16584
rect 25777 16575 25835 16581
rect 25777 16572 25789 16575
rect 25648 16544 25789 16572
rect 25648 16532 25654 16544
rect 25777 16541 25789 16544
rect 25823 16541 25835 16575
rect 25777 16535 25835 16541
rect 25958 16532 25964 16584
rect 26016 16532 26022 16584
rect 26142 16532 26148 16584
rect 26200 16532 26206 16584
rect 28902 16581 28908 16586
rect 28261 16575 28319 16581
rect 28261 16541 28273 16575
rect 28307 16572 28319 16575
rect 28881 16575 28908 16581
rect 28307 16544 28764 16572
rect 28307 16541 28319 16544
rect 28261 16535 28319 16541
rect 26053 16507 26111 16513
rect 26053 16473 26065 16507
rect 26099 16473 26111 16507
rect 26053 16467 26111 16473
rect 24259 16408 24440 16436
rect 24259 16405 24271 16408
rect 24213 16399 24271 16405
rect 24854 16396 24860 16448
rect 24912 16436 24918 16448
rect 24949 16439 25007 16445
rect 24949 16436 24961 16439
rect 24912 16408 24961 16436
rect 24912 16396 24918 16408
rect 24949 16405 24961 16408
rect 24995 16405 25007 16439
rect 24949 16399 25007 16405
rect 25958 16396 25964 16448
rect 26016 16436 26022 16448
rect 26068 16436 26096 16467
rect 26016 16408 26096 16436
rect 28736 16436 28764 16544
rect 28881 16541 28893 16575
rect 28881 16535 28908 16541
rect 28902 16534 28908 16535
rect 28960 16534 28966 16586
rect 29104 16581 29132 16612
rect 29454 16600 29460 16652
rect 29512 16640 29518 16652
rect 30009 16643 30067 16649
rect 30009 16640 30021 16643
rect 29512 16612 30021 16640
rect 29512 16600 29518 16612
rect 30009 16609 30021 16612
rect 30055 16609 30067 16643
rect 30009 16603 30067 16609
rect 31846 16600 31852 16652
rect 31904 16600 31910 16652
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16640 32275 16643
rect 32306 16640 32312 16652
rect 32263 16612 32312 16640
rect 32263 16609 32275 16612
rect 32217 16603 32275 16609
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 33134 16600 33140 16652
rect 33192 16600 33198 16652
rect 29089 16575 29147 16581
rect 29089 16541 29101 16575
rect 29135 16541 29147 16575
rect 29089 16535 29147 16541
rect 29273 16575 29331 16581
rect 29273 16541 29285 16575
rect 29319 16572 29331 16575
rect 29362 16572 29368 16584
rect 29319 16544 29368 16572
rect 29319 16541 29331 16544
rect 29273 16535 29331 16541
rect 29362 16532 29368 16544
rect 29420 16572 29426 16584
rect 29730 16572 29736 16584
rect 29420 16544 29736 16572
rect 29420 16532 29426 16544
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30926 16532 30932 16584
rect 30984 16572 30990 16584
rect 31297 16575 31355 16581
rect 31297 16572 31309 16575
rect 30984 16544 31309 16572
rect 30984 16532 30990 16544
rect 31297 16541 31309 16544
rect 31343 16541 31355 16575
rect 31297 16535 31355 16541
rect 31389 16575 31447 16581
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 31435 16544 31616 16572
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 28997 16507 29055 16513
rect 28997 16473 29009 16507
rect 29043 16504 29055 16507
rect 29178 16504 29184 16516
rect 29043 16476 29184 16504
rect 29043 16473 29055 16476
rect 28997 16467 29055 16473
rect 29178 16464 29184 16476
rect 29236 16464 29242 16516
rect 29454 16464 29460 16516
rect 29512 16504 29518 16516
rect 29822 16504 29828 16516
rect 29512 16476 29828 16504
rect 29512 16464 29518 16476
rect 29822 16464 29828 16476
rect 29880 16464 29886 16516
rect 31478 16464 31484 16516
rect 31536 16464 31542 16516
rect 31588 16504 31616 16544
rect 31662 16532 31668 16584
rect 31720 16532 31726 16584
rect 31757 16575 31815 16581
rect 31757 16541 31769 16575
rect 31803 16572 31815 16575
rect 31864 16572 31892 16600
rect 33244 16581 33272 16680
rect 34330 16668 34336 16720
rect 34388 16708 34394 16720
rect 35342 16708 35348 16720
rect 34388 16680 35348 16708
rect 34388 16668 34394 16680
rect 35342 16668 35348 16680
rect 35400 16668 35406 16720
rect 36446 16708 36452 16720
rect 35452 16680 36452 16708
rect 35452 16649 35480 16680
rect 36446 16668 36452 16680
rect 36504 16668 36510 16720
rect 40034 16708 40040 16720
rect 39316 16680 40040 16708
rect 35437 16643 35495 16649
rect 35437 16609 35449 16643
rect 35483 16609 35495 16643
rect 35437 16603 35495 16609
rect 35713 16643 35771 16649
rect 35713 16609 35725 16643
rect 35759 16640 35771 16643
rect 36078 16640 36084 16652
rect 35759 16612 36084 16640
rect 35759 16609 35771 16612
rect 35713 16603 35771 16609
rect 36078 16600 36084 16612
rect 36136 16600 36142 16652
rect 38378 16600 38384 16652
rect 38436 16600 38442 16652
rect 38657 16643 38715 16649
rect 38657 16609 38669 16643
rect 38703 16640 38715 16643
rect 39206 16640 39212 16652
rect 38703 16612 39212 16640
rect 38703 16609 38715 16612
rect 38657 16603 38715 16609
rect 39206 16600 39212 16612
rect 39264 16600 39270 16652
rect 39316 16649 39344 16680
rect 40034 16668 40040 16680
rect 40092 16668 40098 16720
rect 39301 16643 39359 16649
rect 39301 16609 39313 16643
rect 39347 16609 39359 16643
rect 40405 16643 40463 16649
rect 40405 16640 40417 16643
rect 39301 16603 39359 16609
rect 39776 16612 40417 16640
rect 31803 16544 31892 16572
rect 31941 16575 31999 16581
rect 31803 16541 31815 16544
rect 31757 16535 31815 16541
rect 31941 16541 31953 16575
rect 31987 16541 31999 16575
rect 33229 16575 33287 16581
rect 31941 16535 31999 16541
rect 32876 16544 33180 16572
rect 31956 16504 31984 16535
rect 32674 16504 32680 16516
rect 31588 16476 31892 16504
rect 31956 16476 32680 16504
rect 29549 16439 29607 16445
rect 29549 16436 29561 16439
rect 28736 16408 29561 16436
rect 26016 16396 26022 16408
rect 29549 16405 29561 16408
rect 29595 16405 29607 16439
rect 29549 16399 29607 16405
rect 31110 16396 31116 16448
rect 31168 16396 31174 16448
rect 31864 16436 31892 16476
rect 32674 16464 32680 16476
rect 32732 16504 32738 16516
rect 32876 16504 32904 16544
rect 32732 16476 32904 16504
rect 32732 16464 32738 16476
rect 32950 16464 32956 16516
rect 33008 16464 33014 16516
rect 33152 16504 33180 16544
rect 33229 16541 33241 16575
rect 33275 16541 33287 16575
rect 33229 16535 33287 16541
rect 33413 16575 33471 16581
rect 33413 16541 33425 16575
rect 33459 16541 33471 16575
rect 33413 16535 33471 16541
rect 35345 16575 35403 16581
rect 35345 16541 35357 16575
rect 35391 16572 35403 16575
rect 36354 16572 36360 16584
rect 35391 16544 36360 16572
rect 35391 16541 35403 16544
rect 35345 16535 35403 16541
rect 33428 16504 33456 16535
rect 36354 16532 36360 16544
rect 36412 16532 36418 16584
rect 33152 16476 33456 16504
rect 37826 16464 37832 16516
rect 37884 16464 37890 16516
rect 38286 16464 38292 16516
rect 38344 16504 38350 16516
rect 39776 16504 39804 16612
rect 40405 16609 40417 16612
rect 40451 16609 40463 16643
rect 40405 16603 40463 16609
rect 39850 16532 39856 16584
rect 39908 16532 39914 16584
rect 40218 16532 40224 16584
rect 40276 16532 40282 16584
rect 40310 16532 40316 16584
rect 40368 16532 40374 16584
rect 38344 16476 39804 16504
rect 38344 16464 38350 16476
rect 40678 16464 40684 16516
rect 40736 16464 40742 16516
rect 42058 16504 42064 16516
rect 41906 16476 42064 16504
rect 42058 16464 42064 16476
rect 42116 16464 42122 16516
rect 32769 16439 32827 16445
rect 32769 16436 32781 16439
rect 31864 16408 32781 16436
rect 32769 16405 32781 16408
rect 32815 16436 32827 16439
rect 33226 16436 33232 16448
rect 32815 16408 33232 16436
rect 32815 16405 32827 16408
rect 32769 16399 32827 16405
rect 33226 16396 33232 16408
rect 33284 16396 33290 16448
rect 33318 16396 33324 16448
rect 33376 16436 33382 16448
rect 37734 16436 37740 16448
rect 33376 16408 37740 16436
rect 33376 16396 33382 16408
rect 37734 16396 37740 16408
rect 37792 16436 37798 16448
rect 38102 16436 38108 16448
rect 37792 16408 38108 16436
rect 37792 16396 37798 16408
rect 38102 16396 38108 16408
rect 38160 16396 38166 16448
rect 40129 16439 40187 16445
rect 40129 16405 40141 16439
rect 40175 16436 40187 16439
rect 40586 16436 40592 16448
rect 40175 16408 40592 16436
rect 40175 16405 40187 16408
rect 40129 16399 40187 16405
rect 40586 16396 40592 16408
rect 40644 16396 40650 16448
rect 1104 16346 42504 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 42504 16346
rect 1104 16272 42504 16294
rect 2590 16192 2596 16244
rect 2648 16232 2654 16244
rect 4387 16235 4445 16241
rect 2648 16204 3280 16232
rect 2648 16192 2654 16204
rect 3252 16164 3280 16204
rect 4387 16201 4399 16235
rect 4433 16232 4445 16235
rect 4798 16232 4804 16244
rect 4433 16204 4804 16232
rect 4433 16201 4445 16204
rect 4387 16195 4445 16201
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 6972 16204 7941 16232
rect 6972 16192 6978 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16201 11391 16235
rect 11333 16195 11391 16201
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17310 16232 17316 16244
rect 17083 16204 17316 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 3252 16136 3358 16164
rect 10870 16124 10876 16176
rect 10928 16164 10934 16176
rect 10965 16167 11023 16173
rect 10965 16164 10977 16167
rect 10928 16136 10977 16164
rect 10928 16124 10934 16136
rect 10965 16133 10977 16136
rect 11011 16133 11023 16167
rect 11165 16167 11223 16173
rect 11165 16164 11177 16167
rect 10965 16127 11023 16133
rect 11164 16133 11177 16164
rect 11211 16133 11223 16167
rect 11348 16164 11376 16195
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 19518 16192 19524 16244
rect 19576 16192 19582 16244
rect 24026 16192 24032 16244
rect 24084 16232 24090 16244
rect 24213 16235 24271 16241
rect 24213 16232 24225 16235
rect 24084 16204 24225 16232
rect 24084 16192 24090 16204
rect 24213 16201 24225 16204
rect 24259 16201 24271 16235
rect 25222 16232 25228 16244
rect 24213 16195 24271 16201
rect 24320 16204 25228 16232
rect 11762 16167 11820 16173
rect 11762 16164 11774 16167
rect 11348 16136 11774 16164
rect 11164 16127 11223 16133
rect 11762 16133 11774 16136
rect 11808 16133 11820 16167
rect 11762 16127 11820 16133
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 900 16068 1409 16096
rect 900 16056 906 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 1670 16056 1676 16108
rect 1728 16056 1734 16108
rect 2406 16056 2412 16108
rect 2464 16096 2470 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 2464 16068 2605 16096
rect 2464 16056 2470 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 4706 16056 4712 16108
rect 4764 16056 4770 16108
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 8754 16096 8760 16108
rect 8619 16068 8760 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 8754 16056 8760 16068
rect 8812 16056 8818 16108
rect 11164 16096 11192 16127
rect 12158 16124 12164 16176
rect 12216 16164 12222 16176
rect 13081 16167 13139 16173
rect 12216 16136 13032 16164
rect 12216 16124 12222 16136
rect 12894 16096 12900 16108
rect 11164 16068 12900 16096
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 13004 16105 13032 16136
rect 13081 16133 13093 16167
rect 13127 16164 13139 16167
rect 14400 16167 14458 16173
rect 13127 16136 13952 16164
rect 13127 16133 13139 16136
rect 13081 16127 13139 16133
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 3786 16028 3792 16040
rect 3007 16000 3792 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 3936 16000 4537 16028
rect 3936 15988 3942 16000
rect 4525 15997 4537 16000
rect 4571 16028 4583 16031
rect 5350 16028 5356 16040
rect 4571 16000 5356 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 11514 15988 11520 16040
rect 11572 15988 11578 16040
rect 13004 16028 13032 16059
rect 13170 16056 13176 16108
rect 13228 16056 13234 16108
rect 13924 16096 13952 16136
rect 14400 16133 14412 16167
rect 14446 16164 14458 16167
rect 14829 16167 14887 16173
rect 14829 16164 14841 16167
rect 14446 16136 14841 16164
rect 14446 16133 14458 16136
rect 14400 16127 14458 16133
rect 14829 16133 14841 16136
rect 14875 16133 14887 16167
rect 18719 16167 18777 16173
rect 18719 16164 18731 16167
rect 14829 16127 14887 16133
rect 18156 16136 18731 16164
rect 14737 16099 14795 16105
rect 14737 16096 14749 16099
rect 13924 16068 14749 16096
rect 14737 16065 14749 16068
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 14918 16056 14924 16108
rect 14976 16056 14982 16108
rect 18156 16105 18184 16136
rect 18719 16133 18731 16136
rect 18765 16164 18777 16167
rect 19536 16164 19564 16192
rect 19978 16164 19984 16176
rect 18765 16136 19472 16164
rect 19536 16136 19984 16164
rect 18765 16133 18777 16136
rect 18719 16127 18777 16133
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17175 16068 18153 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 18141 16065 18153 16068
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 18509 16099 18567 16105
rect 18509 16065 18521 16099
rect 18555 16065 18567 16099
rect 18509 16059 18567 16065
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16096 18659 16099
rect 19058 16096 19064 16108
rect 18647 16068 19064 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 14645 16031 14703 16037
rect 13004 16000 13676 16028
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 11388 15932 11560 15960
rect 11388 15920 11394 15932
rect 1581 15895 1639 15901
rect 1581 15861 1593 15895
rect 1627 15892 1639 15895
rect 1762 15892 1768 15904
rect 1627 15864 1768 15892
rect 1627 15861 1639 15864
rect 1581 15855 1639 15861
rect 1762 15852 1768 15864
rect 1820 15852 1826 15904
rect 1854 15852 1860 15904
rect 1912 15852 1918 15904
rect 4893 15895 4951 15901
rect 4893 15861 4905 15895
rect 4939 15892 4951 15895
rect 5258 15892 5264 15904
rect 4939 15864 5264 15892
rect 4939 15861 4951 15864
rect 4893 15855 4951 15861
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11422 15892 11428 15904
rect 11195 15864 11428 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 11422 15852 11428 15864
rect 11480 15852 11486 15904
rect 11532 15892 11560 15932
rect 12710 15920 12716 15972
rect 12768 15960 12774 15972
rect 13262 15960 13268 15972
rect 12768 15932 13268 15960
rect 12768 15920 12774 15932
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 12250 15892 12256 15904
rect 11532 15864 12256 15892
rect 12250 15852 12256 15864
rect 12308 15892 12314 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12308 15864 12909 15892
rect 12308 15852 12314 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 13648 15892 13676 16000
rect 14645 15997 14657 16031
rect 14691 16028 14703 16031
rect 15194 16028 15200 16040
rect 14691 16000 15200 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 17034 15988 17040 16040
rect 17092 16028 17098 16040
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 17092 16000 17233 16028
rect 17092 15988 17098 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 17497 16031 17555 16037
rect 17497 16028 17509 16031
rect 17368 16000 17509 16028
rect 17368 15988 17374 16000
rect 17497 15997 17509 16000
rect 17543 15997 17555 16031
rect 18524 16028 18552 16059
rect 19058 16056 19064 16068
rect 19116 16096 19122 16108
rect 19444 16105 19472 16136
rect 19429 16099 19487 16105
rect 19116 16068 19334 16096
rect 19116 16056 19122 16068
rect 18782 16028 18788 16040
rect 18524 16000 18788 16028
rect 17497 15991 17555 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 18877 16031 18935 16037
rect 18877 15997 18889 16031
rect 18923 15997 18935 16031
rect 19306 16028 19334 16068
rect 19429 16065 19441 16099
rect 19475 16065 19487 16099
rect 19429 16059 19487 16065
rect 19518 16056 19524 16108
rect 19576 16056 19582 16108
rect 19610 16056 19616 16108
rect 19668 16056 19674 16108
rect 19812 16105 19840 16136
rect 19978 16124 19984 16136
rect 20036 16124 20042 16176
rect 20162 16124 20168 16176
rect 20220 16164 20226 16176
rect 20220 16136 20392 16164
rect 20220 16124 20226 16136
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 19886 16056 19892 16108
rect 19944 16056 19950 16108
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16065 20315 16099
rect 20364 16096 20392 16136
rect 20438 16124 20444 16176
rect 20496 16124 20502 16176
rect 20530 16124 20536 16176
rect 20588 16164 20594 16176
rect 20901 16167 20959 16173
rect 20901 16164 20913 16167
rect 20588 16136 20913 16164
rect 20588 16124 20594 16136
rect 20901 16133 20913 16136
rect 20947 16133 20959 16167
rect 20901 16127 20959 16133
rect 23934 16124 23940 16176
rect 23992 16164 23998 16176
rect 24320 16164 24348 16204
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 26234 16192 26240 16244
rect 26292 16232 26298 16244
rect 27338 16232 27344 16244
rect 26292 16204 27344 16232
rect 26292 16192 26298 16204
rect 27338 16192 27344 16204
rect 27396 16192 27402 16244
rect 27433 16235 27491 16241
rect 27433 16201 27445 16235
rect 27479 16232 27491 16235
rect 28902 16232 28908 16244
rect 27479 16204 28908 16232
rect 27479 16201 27491 16204
rect 27433 16195 27491 16201
rect 28902 16192 28908 16204
rect 28960 16192 28966 16244
rect 29914 16232 29920 16244
rect 29012 16204 29920 16232
rect 23992 16136 24348 16164
rect 23992 16124 23998 16136
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 20364 16068 20637 16096
rect 20257 16059 20315 16065
rect 20625 16065 20637 16068
rect 20671 16096 20683 16099
rect 21910 16096 21916 16108
rect 20671 16068 21916 16096
rect 20671 16065 20683 16068
rect 20625 16059 20683 16065
rect 20272 16028 20300 16059
rect 21910 16056 21916 16068
rect 21968 16056 21974 16108
rect 24320 16105 24348 16136
rect 24670 16124 24676 16176
rect 24728 16124 24734 16176
rect 24765 16167 24823 16173
rect 24765 16133 24777 16167
rect 24811 16164 24823 16167
rect 24854 16164 24860 16176
rect 24811 16136 24860 16164
rect 24811 16133 24823 16136
rect 24765 16127 24823 16133
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 29012 16164 29040 16204
rect 29914 16192 29920 16204
rect 29972 16232 29978 16244
rect 31386 16232 31392 16244
rect 29972 16204 31392 16232
rect 29972 16192 29978 16204
rect 31386 16192 31392 16204
rect 31444 16232 31450 16244
rect 31662 16232 31668 16244
rect 31444 16204 31668 16232
rect 31444 16192 31450 16204
rect 31662 16192 31668 16204
rect 31720 16192 31726 16244
rect 33962 16192 33968 16244
rect 34020 16232 34026 16244
rect 34517 16235 34575 16241
rect 34517 16232 34529 16235
rect 34020 16204 34529 16232
rect 34020 16192 34026 16204
rect 34517 16201 34529 16204
rect 34563 16201 34575 16235
rect 34517 16195 34575 16201
rect 36354 16192 36360 16244
rect 36412 16192 36418 16244
rect 37826 16192 37832 16244
rect 37884 16232 37890 16244
rect 37884 16204 38792 16232
rect 37884 16192 37890 16204
rect 24964 16136 29040 16164
rect 24964 16105 24992 16136
rect 29638 16124 29644 16176
rect 29696 16124 29702 16176
rect 30469 16167 30527 16173
rect 30469 16133 30481 16167
rect 30515 16164 30527 16167
rect 32582 16164 32588 16176
rect 30515 16136 32588 16164
rect 30515 16133 30527 16136
rect 30469 16127 30527 16133
rect 32582 16124 32588 16136
rect 32640 16124 32646 16176
rect 33318 16124 33324 16176
rect 33376 16164 33382 16176
rect 35342 16164 35348 16176
rect 33376 16136 33534 16164
rect 34532 16136 35348 16164
rect 33376 16124 33382 16136
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16065 24179 16099
rect 24121 16059 24179 16065
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 24949 16099 25007 16105
rect 24627 16068 24900 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 20438 16028 20444 16040
rect 19306 16000 20444 16028
rect 18877 15991 18935 15997
rect 18892 15960 18920 15991
rect 20438 15988 20444 16000
rect 20496 15988 20502 16040
rect 21450 15988 21456 16040
rect 21508 15988 21514 16040
rect 24136 16028 24164 16059
rect 24762 16028 24768 16040
rect 24136 16000 24768 16028
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 24872 16028 24900 16068
rect 24949 16065 24961 16099
rect 24995 16065 25007 16099
rect 25498 16096 25504 16108
rect 24949 16059 25007 16065
rect 25056 16068 25504 16096
rect 25056 16028 25084 16068
rect 25498 16056 25504 16068
rect 25556 16096 25562 16108
rect 25556 16068 28028 16096
rect 25556 16056 25562 16068
rect 24872 16000 25084 16028
rect 25682 15988 25688 16040
rect 25740 16028 25746 16040
rect 27525 16031 27583 16037
rect 27525 16028 27537 16031
rect 25740 16000 27537 16028
rect 25740 15988 25746 16000
rect 27525 15997 27537 16000
rect 27571 16028 27583 16031
rect 27893 16031 27951 16037
rect 27893 16028 27905 16031
rect 27571 16000 27905 16028
rect 27571 15997 27583 16000
rect 27525 15991 27583 15997
rect 27893 15997 27905 16000
rect 27939 15997 27951 16031
rect 28000 16028 28028 16068
rect 28074 16056 28080 16108
rect 28132 16096 28138 16108
rect 28169 16099 28227 16105
rect 28169 16096 28181 16099
rect 28132 16068 28181 16096
rect 28132 16056 28138 16068
rect 28169 16065 28181 16068
rect 28215 16065 28227 16099
rect 28169 16059 28227 16065
rect 28350 16056 28356 16108
rect 28408 16056 28414 16108
rect 30282 16096 30288 16108
rect 29840 16068 30288 16096
rect 29086 16028 29092 16040
rect 28000 16000 29092 16028
rect 27893 15991 27951 15997
rect 29086 15988 29092 16000
rect 29144 16028 29150 16040
rect 29362 16028 29368 16040
rect 29144 16000 29368 16028
rect 29144 15988 29150 16000
rect 29362 15988 29368 16000
rect 29420 15988 29426 16040
rect 19334 15960 19340 15972
rect 18892 15932 19340 15960
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 19978 15920 19984 15972
rect 20036 15960 20042 15972
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 20036 15932 20085 15960
rect 20036 15920 20042 15932
rect 20073 15929 20085 15932
rect 20119 15960 20131 15963
rect 23658 15960 23664 15972
rect 20119 15932 23664 15960
rect 20119 15929 20131 15932
rect 20073 15923 20131 15929
rect 23658 15920 23664 15932
rect 23716 15920 23722 15972
rect 24397 15963 24455 15969
rect 24397 15929 24409 15963
rect 24443 15960 24455 15963
rect 26418 15960 26424 15972
rect 24443 15932 26424 15960
rect 24443 15929 24455 15932
rect 24397 15923 24455 15929
rect 26418 15920 26424 15932
rect 26476 15920 26482 15972
rect 15194 15892 15200 15904
rect 13648 15864 15200 15892
rect 12897 15855 12955 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 15804 15864 16681 15892
rect 15804 15852 15810 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 18233 15895 18291 15901
rect 18233 15861 18245 15895
rect 18279 15892 18291 15895
rect 18782 15892 18788 15904
rect 18279 15864 18788 15892
rect 18279 15861 18291 15864
rect 18233 15855 18291 15861
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 19245 15895 19303 15901
rect 19245 15861 19257 15895
rect 19291 15892 19303 15895
rect 19518 15892 19524 15904
rect 19291 15864 19524 15892
rect 19291 15861 19303 15864
rect 19245 15855 19303 15861
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 20806 15852 20812 15904
rect 20864 15852 20870 15904
rect 26050 15852 26056 15904
rect 26108 15892 26114 15904
rect 26973 15895 27031 15901
rect 26973 15892 26985 15895
rect 26108 15864 26985 15892
rect 26108 15852 26114 15864
rect 26973 15861 26985 15864
rect 27019 15861 27031 15895
rect 26973 15855 27031 15861
rect 28616 15895 28674 15901
rect 28616 15861 28628 15895
rect 28662 15892 28674 15895
rect 28718 15892 28724 15904
rect 28662 15864 28724 15892
rect 28662 15861 28674 15864
rect 28616 15855 28674 15861
rect 28718 15852 28724 15864
rect 28776 15852 28782 15904
rect 29178 15852 29184 15904
rect 29236 15892 29242 15904
rect 29840 15892 29868 16068
rect 30282 16056 30288 16068
rect 30340 16056 30346 16108
rect 30558 16056 30564 16108
rect 30616 16056 30622 16108
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 29236 15864 29868 15892
rect 30101 15895 30159 15901
rect 29236 15852 29242 15864
rect 30101 15861 30113 15895
rect 30147 15892 30159 15895
rect 30466 15892 30472 15904
rect 30147 15864 30472 15892
rect 30147 15861 30159 15864
rect 30101 15855 30159 15861
rect 30466 15852 30472 15864
rect 30524 15852 30530 15904
rect 30668 15892 30696 16059
rect 32214 16056 32220 16108
rect 32272 16056 32278 16108
rect 31113 16031 31171 16037
rect 31113 15997 31125 16031
rect 31159 15997 31171 16031
rect 31113 15991 31171 15997
rect 30837 15963 30895 15969
rect 30837 15929 30849 15963
rect 30883 15960 30895 15963
rect 31128 15960 31156 15991
rect 31202 15988 31208 16040
rect 31260 16028 31266 16040
rect 32766 16028 32772 16040
rect 31260 16000 32772 16028
rect 31260 15988 31266 16000
rect 32766 15988 32772 16000
rect 32824 15988 32830 16040
rect 33045 16031 33103 16037
rect 33045 15997 33057 16031
rect 33091 16028 33103 16031
rect 33594 16028 33600 16040
rect 33091 16000 33600 16028
rect 33091 15997 33103 16000
rect 33045 15991 33103 15997
rect 33594 15988 33600 16000
rect 33652 15988 33658 16040
rect 32306 15960 32312 15972
rect 30883 15932 31156 15960
rect 31220 15932 32312 15960
rect 30883 15929 30895 15932
rect 30837 15923 30895 15929
rect 31220 15892 31248 15932
rect 32306 15920 32312 15932
rect 32364 15920 32370 15972
rect 30668 15864 31248 15892
rect 31478 15852 31484 15904
rect 31536 15892 31542 15904
rect 31757 15895 31815 15901
rect 31757 15892 31769 15895
rect 31536 15864 31769 15892
rect 31536 15852 31542 15864
rect 31757 15861 31769 15864
rect 31803 15861 31815 15895
rect 31757 15855 31815 15861
rect 33410 15852 33416 15904
rect 33468 15892 33474 15904
rect 34532 15892 34560 16136
rect 35342 16124 35348 16136
rect 35400 16124 35406 16176
rect 34606 16056 34612 16108
rect 34664 16056 34670 16108
rect 36372 16096 36400 16192
rect 37553 16167 37611 16173
rect 37553 16164 37565 16167
rect 37108 16136 37565 16164
rect 37001 16099 37059 16105
rect 37001 16096 37013 16099
rect 36372 16068 37013 16096
rect 37001 16065 37013 16068
rect 37047 16065 37059 16099
rect 37001 16059 37059 16065
rect 34885 16031 34943 16037
rect 34885 15997 34897 16031
rect 34931 16028 34943 16031
rect 35434 16028 35440 16040
rect 34931 16000 35440 16028
rect 34931 15997 34943 16000
rect 34885 15991 34943 15997
rect 35434 15988 35440 16000
rect 35492 15988 35498 16040
rect 35526 15988 35532 16040
rect 35584 16028 35590 16040
rect 37108 16028 37136 16136
rect 37553 16133 37565 16136
rect 37599 16133 37611 16167
rect 37553 16127 37611 16133
rect 38565 16167 38623 16173
rect 38565 16133 38577 16167
rect 38611 16164 38623 16167
rect 38654 16164 38660 16176
rect 38611 16136 38660 16164
rect 38611 16133 38623 16136
rect 38565 16127 38623 16133
rect 38654 16124 38660 16136
rect 38712 16124 38718 16176
rect 38764 16164 38792 16204
rect 40034 16192 40040 16244
rect 40092 16192 40098 16244
rect 40678 16192 40684 16244
rect 40736 16232 40742 16244
rect 40773 16235 40831 16241
rect 40773 16232 40785 16235
rect 40736 16204 40785 16232
rect 40736 16192 40742 16204
rect 40773 16201 40785 16204
rect 40819 16201 40831 16235
rect 40773 16195 40831 16201
rect 40313 16167 40371 16173
rect 38764 16136 39054 16164
rect 40313 16133 40325 16167
rect 40359 16164 40371 16167
rect 41230 16164 41236 16176
rect 40359 16136 41236 16164
rect 40359 16133 40371 16136
rect 40313 16127 40371 16133
rect 41230 16124 41236 16136
rect 41288 16124 41294 16176
rect 37458 16056 37464 16108
rect 37516 16056 37522 16108
rect 37642 16056 37648 16108
rect 37700 16056 37706 16108
rect 37734 16056 37740 16108
rect 37792 16096 37798 16108
rect 37829 16099 37887 16105
rect 37829 16096 37841 16099
rect 37792 16068 37841 16096
rect 37792 16056 37798 16068
rect 37829 16065 37841 16068
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 40126 16056 40132 16108
rect 40184 16056 40190 16108
rect 40402 16056 40408 16108
rect 40460 16056 40466 16108
rect 40497 16099 40555 16105
rect 40497 16065 40509 16099
rect 40543 16065 40555 16099
rect 40497 16059 40555 16065
rect 38286 16028 38292 16040
rect 35584 16000 37136 16028
rect 37476 16000 38292 16028
rect 35584 15988 35590 16000
rect 37476 15972 37504 16000
rect 38286 15988 38292 16000
rect 38344 15988 38350 16040
rect 40034 15988 40040 16040
rect 40092 16028 40098 16040
rect 40512 16028 40540 16059
rect 40586 16056 40592 16108
rect 40644 16096 40650 16108
rect 41509 16099 41567 16105
rect 41509 16096 41521 16099
rect 40644 16068 41521 16096
rect 40644 16056 40650 16068
rect 41509 16065 41521 16068
rect 41555 16065 41567 16099
rect 41509 16059 41567 16065
rect 40092 16000 40540 16028
rect 41325 16031 41383 16037
rect 40092 15988 40098 16000
rect 41325 15997 41337 16031
rect 41371 15997 41383 16031
rect 41325 15991 41383 15997
rect 37458 15920 37464 15972
rect 37516 15920 37522 15972
rect 40681 15963 40739 15969
rect 40681 15929 40693 15963
rect 40727 15960 40739 15963
rect 41340 15960 41368 15991
rect 41598 15988 41604 16040
rect 41656 15988 41662 16040
rect 40727 15932 41368 15960
rect 40727 15929 40739 15932
rect 40681 15923 40739 15929
rect 33468 15864 34560 15892
rect 33468 15852 33474 15864
rect 35342 15852 35348 15904
rect 35400 15892 35406 15904
rect 36449 15895 36507 15901
rect 36449 15892 36461 15895
rect 35400 15864 36461 15892
rect 35400 15852 35406 15864
rect 36449 15861 36461 15864
rect 36495 15861 36507 15895
rect 36449 15855 36507 15861
rect 37182 15852 37188 15904
rect 37240 15892 37246 15904
rect 37277 15895 37335 15901
rect 37277 15892 37289 15895
rect 37240 15864 37289 15892
rect 37240 15852 37246 15864
rect 37277 15861 37289 15864
rect 37323 15861 37335 15895
rect 37277 15855 37335 15861
rect 38102 15852 38108 15904
rect 38160 15892 38166 15904
rect 39758 15892 39764 15904
rect 38160 15864 39764 15892
rect 38160 15852 38166 15864
rect 39758 15852 39764 15864
rect 39816 15852 39822 15904
rect 40218 15852 40224 15904
rect 40276 15892 40282 15904
rect 41509 15895 41567 15901
rect 41509 15892 41521 15895
rect 40276 15864 41521 15892
rect 40276 15852 40282 15864
rect 41509 15861 41521 15864
rect 41555 15861 41567 15895
rect 41509 15855 41567 15861
rect 41690 15852 41696 15904
rect 41748 15892 41754 15904
rect 41877 15895 41935 15901
rect 41877 15892 41889 15895
rect 41748 15864 41889 15892
rect 41748 15852 41754 15864
rect 41877 15861 41889 15864
rect 41923 15861 41935 15895
rect 41877 15855 41935 15861
rect 1104 15802 42504 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 42504 15802
rect 1104 15728 42504 15750
rect 3786 15648 3792 15700
rect 3844 15648 3850 15700
rect 11330 15648 11336 15700
rect 11388 15648 11394 15700
rect 11422 15648 11428 15700
rect 11480 15688 11486 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11480 15660 11621 15688
rect 11480 15648 11486 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 11756 15660 12848 15688
rect 11756 15648 11762 15660
rect 12253 15623 12311 15629
rect 12253 15620 12265 15623
rect 11072 15592 12265 15620
rect 1394 15512 1400 15564
rect 1452 15552 1458 15564
rect 2314 15552 2320 15564
rect 1452 15524 2320 15552
rect 1452 15512 1458 15524
rect 2314 15512 2320 15524
rect 2372 15512 2378 15564
rect 5718 15512 5724 15564
rect 5776 15512 5782 15564
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 6454 15552 6460 15564
rect 6227 15524 6460 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 10870 15552 10876 15564
rect 10827 15524 10876 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 1762 15444 1768 15496
rect 1820 15444 1826 15496
rect 3191 15487 3249 15493
rect 3191 15453 3203 15487
rect 3237 15484 3249 15487
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 3237 15456 4353 15484
rect 3237 15453 3249 15456
rect 3191 15447 3249 15453
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 5810 15444 5816 15496
rect 5868 15444 5874 15496
rect 6641 15487 6699 15493
rect 6641 15453 6653 15487
rect 6687 15484 6699 15487
rect 6730 15484 6736 15496
rect 6687 15456 6736 15484
rect 6687 15453 6699 15456
rect 6641 15447 6699 15453
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15484 6883 15487
rect 8478 15484 8484 15496
rect 6871 15456 8484 15484
rect 6871 15453 6883 15456
rect 6825 15447 6883 15453
rect 8478 15444 8484 15456
rect 8536 15484 8542 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 8536 15456 8953 15484
rect 8536 15444 8542 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15484 9183 15487
rect 9214 15484 9220 15496
rect 9171 15456 9220 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9585 15487 9643 15493
rect 9355 15456 9536 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 2590 15376 2596 15428
rect 2648 15376 2654 15428
rect 6638 15308 6644 15360
rect 6696 15348 6702 15360
rect 9508 15357 9536 15456
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 10042 15484 10048 15496
rect 9631 15456 10048 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 11072 15493 11100 15592
rect 12253 15589 12265 15592
rect 12299 15589 12311 15623
rect 12253 15583 12311 15589
rect 11793 15555 11851 15561
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12158 15552 12164 15564
rect 11839 15524 12164 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 12820 15552 12848 15660
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 13081 15691 13139 15697
rect 13081 15688 13093 15691
rect 12952 15660 13093 15688
rect 12952 15648 12958 15660
rect 13081 15657 13093 15660
rect 13127 15657 13139 15691
rect 13081 15651 13139 15657
rect 17218 15648 17224 15700
rect 17276 15648 17282 15700
rect 17310 15648 17316 15700
rect 17368 15648 17374 15700
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 18472 15660 19257 15688
rect 18472 15648 18478 15660
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 19245 15651 19303 15657
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 19668 15660 19809 15688
rect 19668 15648 19674 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 19797 15651 19855 15657
rect 23658 15648 23664 15700
rect 23716 15688 23722 15700
rect 25590 15688 25596 15700
rect 23716 15660 25596 15688
rect 23716 15648 23722 15660
rect 25590 15648 25596 15660
rect 25648 15688 25654 15700
rect 25648 15660 27292 15688
rect 25648 15648 25654 15660
rect 14918 15620 14924 15632
rect 13372 15592 14924 15620
rect 13372 15561 13400 15592
rect 14918 15580 14924 15592
rect 14976 15620 14982 15632
rect 15197 15623 15255 15629
rect 15197 15620 15209 15623
rect 14976 15592 15209 15620
rect 14976 15580 14982 15592
rect 15197 15589 15209 15592
rect 15243 15589 15255 15623
rect 25682 15620 25688 15632
rect 15197 15583 15255 15589
rect 23860 15592 25688 15620
rect 13357 15555 13415 15561
rect 13357 15552 13369 15555
rect 12820 15524 13369 15552
rect 13357 15521 13369 15524
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 13817 15555 13875 15561
rect 13817 15521 13829 15555
rect 13863 15552 13875 15555
rect 13906 15552 13912 15564
rect 13863 15524 13912 15552
rect 13863 15521 13875 15524
rect 13817 15515 13875 15521
rect 13906 15512 13912 15524
rect 13964 15512 13970 15564
rect 19061 15555 19119 15561
rect 19061 15552 19073 15555
rect 15488 15524 19073 15552
rect 15488 15496 15516 15524
rect 19061 15521 19073 15524
rect 19107 15521 19119 15555
rect 19061 15515 19119 15521
rect 20622 15512 20628 15564
rect 20680 15512 20686 15564
rect 21450 15512 21456 15564
rect 21508 15552 21514 15564
rect 22373 15555 22431 15561
rect 22373 15552 22385 15555
rect 21508 15524 22385 15552
rect 21508 15512 21514 15524
rect 22373 15521 22385 15524
rect 22419 15521 22431 15555
rect 22373 15515 22431 15521
rect 23198 15512 23204 15564
rect 23256 15552 23262 15564
rect 23860 15561 23888 15592
rect 25682 15580 25688 15592
rect 25740 15580 25746 15632
rect 23845 15555 23903 15561
rect 23845 15552 23857 15555
rect 23256 15524 23857 15552
rect 23256 15512 23262 15524
rect 23845 15521 23857 15524
rect 23891 15521 23903 15555
rect 23845 15515 23903 15521
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 25777 15555 25835 15561
rect 25777 15552 25789 15555
rect 24912 15524 25789 15552
rect 24912 15512 24918 15524
rect 25777 15521 25789 15524
rect 25823 15552 25835 15555
rect 26142 15552 26148 15564
rect 25823 15524 26148 15552
rect 25823 15521 25835 15524
rect 25777 15515 25835 15521
rect 26142 15512 26148 15524
rect 26200 15512 26206 15564
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 11698 15484 11704 15496
rect 11057 15447 11115 15453
rect 11440 15456 11704 15484
rect 10980 15416 11008 15447
rect 11317 15419 11375 15425
rect 10980 15388 11192 15416
rect 11164 15360 11192 15388
rect 11317 15385 11329 15419
rect 11363 15416 11375 15419
rect 11440 15416 11468 15456
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 11363 15388 11468 15416
rect 11517 15419 11575 15425
rect 11363 15385 11375 15388
rect 11317 15379 11375 15385
rect 11517 15385 11529 15419
rect 11563 15385 11575 15419
rect 11900 15416 11928 15447
rect 11974 15444 11980 15496
rect 12032 15444 12038 15496
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 12250 15484 12256 15496
rect 12115 15456 12256 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12894 15444 12900 15496
rect 12952 15444 12958 15496
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15484 13507 15487
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13495 15456 14105 15484
rect 13495 15453 13507 15456
rect 13449 15447 13507 15453
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 12710 15416 12716 15428
rect 11900 15388 12716 15416
rect 11517 15379 11575 15385
rect 6733 15351 6791 15357
rect 6733 15348 6745 15351
rect 6696 15320 6745 15348
rect 6696 15308 6702 15320
rect 6733 15317 6745 15320
rect 6779 15317 6791 15351
rect 6733 15311 6791 15317
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9858 15348 9864 15360
rect 9539 15320 9864 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 10781 15351 10839 15357
rect 10781 15317 10793 15351
rect 10827 15348 10839 15351
rect 11054 15348 11060 15360
rect 10827 15320 11060 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11146 15308 11152 15360
rect 11204 15308 11210 15360
rect 11532 15348 11560 15379
rect 12710 15376 12716 15388
rect 12768 15376 12774 15428
rect 11974 15348 11980 15360
rect 11532 15320 11980 15348
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 13004 15348 13032 15447
rect 14734 15444 14740 15496
rect 14792 15444 14798 15496
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15484 15071 15487
rect 15194 15484 15200 15496
rect 15059 15456 15200 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 14844 15416 14872 15447
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 15470 15444 15476 15496
rect 15528 15444 15534 15496
rect 17678 15444 17684 15496
rect 17736 15444 17742 15496
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19208 15456 19625 15484
rect 19208 15444 19214 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 24302 15484 24308 15496
rect 23707 15456 24308 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 13320 15388 14872 15416
rect 13320 15376 13326 15388
rect 15746 15376 15752 15428
rect 15804 15376 15810 15428
rect 16298 15376 16304 15428
rect 16356 15376 16362 15428
rect 18782 15376 18788 15428
rect 18840 15376 18846 15428
rect 19426 15376 19432 15428
rect 19484 15416 19490 15428
rect 20364 15416 20392 15447
rect 24302 15444 24308 15456
rect 24360 15444 24366 15496
rect 24946 15444 24952 15496
rect 25004 15484 25010 15496
rect 25409 15487 25467 15493
rect 25409 15484 25421 15487
rect 25004 15456 25421 15484
rect 25004 15444 25010 15456
rect 25409 15453 25421 15456
rect 25455 15453 25467 15487
rect 27264 15484 27292 15660
rect 27338 15648 27344 15700
rect 27396 15688 27402 15700
rect 27525 15691 27583 15697
rect 27525 15688 27537 15691
rect 27396 15660 27537 15688
rect 27396 15648 27402 15660
rect 27525 15657 27537 15660
rect 27571 15657 27583 15691
rect 27525 15651 27583 15657
rect 28537 15691 28595 15697
rect 28537 15657 28549 15691
rect 28583 15688 28595 15691
rect 28994 15688 29000 15700
rect 28583 15660 29000 15688
rect 28583 15657 28595 15660
rect 28537 15651 28595 15657
rect 28994 15648 29000 15660
rect 29052 15648 29058 15700
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 30190 15688 30196 15700
rect 29144 15660 30196 15688
rect 29144 15648 29150 15660
rect 30190 15648 30196 15660
rect 30248 15688 30254 15700
rect 30248 15660 30880 15688
rect 30248 15648 30254 15660
rect 28261 15623 28319 15629
rect 28261 15589 28273 15623
rect 28307 15620 28319 15623
rect 30650 15620 30656 15632
rect 28307 15592 30656 15620
rect 28307 15589 28319 15592
rect 28261 15583 28319 15589
rect 30650 15580 30656 15592
rect 30708 15580 30714 15632
rect 27706 15512 27712 15564
rect 27764 15512 27770 15564
rect 28350 15512 28356 15564
rect 28408 15552 28414 15564
rect 28408 15524 30788 15552
rect 28408 15512 28414 15524
rect 29086 15484 29092 15496
rect 27264 15456 29092 15484
rect 25409 15447 25467 15453
rect 29086 15444 29092 15456
rect 29144 15444 29150 15496
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15484 29239 15487
rect 29914 15484 29920 15496
rect 29227 15456 29920 15484
rect 29227 15453 29239 15456
rect 29181 15447 29239 15453
rect 29914 15444 29920 15456
rect 29972 15444 29978 15496
rect 30193 15487 30251 15493
rect 30193 15453 30205 15487
rect 30239 15453 30251 15487
rect 30193 15447 30251 15453
rect 19484 15388 20392 15416
rect 19484 15376 19490 15388
rect 20806 15376 20812 15428
rect 20864 15416 20870 15428
rect 20901 15419 20959 15425
rect 20901 15416 20913 15419
rect 20864 15388 20913 15416
rect 20864 15376 20870 15388
rect 20901 15385 20913 15388
rect 20947 15385 20959 15419
rect 20901 15379 20959 15385
rect 20990 15376 20996 15428
rect 21048 15416 21054 15428
rect 23753 15419 23811 15425
rect 21048 15388 21390 15416
rect 22572 15388 23704 15416
rect 21048 15376 21054 15388
rect 12124 15320 13032 15348
rect 12124 15308 12130 15320
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 22572 15348 22600 15388
rect 19944 15320 22600 15348
rect 19944 15308 19950 15320
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 23293 15351 23351 15357
rect 23293 15348 23305 15351
rect 22704 15320 23305 15348
rect 22704 15308 22710 15320
rect 23293 15317 23305 15320
rect 23339 15317 23351 15351
rect 23676 15348 23704 15388
rect 23753 15385 23765 15419
rect 23799 15416 23811 15419
rect 24670 15416 24676 15428
rect 23799 15388 24676 15416
rect 23799 15385 23811 15388
rect 23753 15379 23811 15385
rect 24670 15376 24676 15388
rect 24728 15416 24734 15428
rect 24857 15419 24915 15425
rect 24857 15416 24869 15419
rect 24728 15388 24869 15416
rect 24728 15376 24734 15388
rect 24857 15385 24869 15388
rect 24903 15385 24915 15419
rect 24857 15379 24915 15385
rect 26050 15376 26056 15428
rect 26108 15376 26114 15428
rect 27522 15416 27528 15428
rect 27278 15388 27528 15416
rect 27522 15376 27528 15388
rect 27580 15376 27586 15428
rect 29454 15376 29460 15428
rect 29512 15416 29518 15428
rect 30208 15416 30236 15447
rect 30466 15444 30472 15496
rect 30524 15444 30530 15496
rect 30650 15444 30656 15496
rect 30708 15444 30714 15496
rect 30561 15419 30619 15425
rect 29512 15388 30052 15416
rect 30208 15388 30328 15416
rect 29512 15376 29518 15388
rect 28442 15348 28448 15360
rect 23676 15320 28448 15348
rect 23293 15311 23351 15317
rect 28442 15308 28448 15320
rect 28500 15348 28506 15360
rect 29178 15348 29184 15360
rect 28500 15320 29184 15348
rect 28500 15308 28506 15320
rect 29178 15308 29184 15320
rect 29236 15308 29242 15360
rect 29546 15308 29552 15360
rect 29604 15308 29610 15360
rect 30024 15348 30052 15388
rect 30190 15348 30196 15360
rect 30024 15320 30196 15348
rect 30190 15308 30196 15320
rect 30248 15308 30254 15360
rect 30300 15357 30328 15388
rect 30561 15385 30573 15419
rect 30607 15385 30619 15419
rect 30760 15416 30788 15524
rect 30852 15493 30880 15660
rect 32582 15648 32588 15700
rect 32640 15688 32646 15700
rect 32769 15691 32827 15697
rect 32769 15688 32781 15691
rect 32640 15660 32781 15688
rect 32640 15648 32646 15660
rect 32769 15657 32781 15660
rect 32815 15657 32827 15691
rect 32769 15651 32827 15657
rect 33594 15648 33600 15700
rect 33652 15648 33658 15700
rect 35434 15648 35440 15700
rect 35492 15648 35498 15700
rect 35544 15660 37412 15688
rect 32674 15580 32680 15632
rect 32732 15620 32738 15632
rect 32732 15592 33364 15620
rect 32732 15580 32738 15592
rect 31202 15552 31208 15564
rect 30944 15524 31208 15552
rect 30944 15493 30972 15524
rect 31202 15512 31208 15524
rect 31260 15512 31266 15564
rect 33336 15561 33364 15592
rect 34238 15580 34244 15632
rect 34296 15620 34302 15632
rect 35544 15620 35572 15660
rect 34296 15592 35572 15620
rect 34296 15580 34302 15592
rect 33321 15555 33379 15561
rect 33321 15521 33333 15555
rect 33367 15521 33379 15555
rect 33321 15515 33379 15521
rect 33410 15512 33416 15564
rect 33468 15552 33474 15564
rect 34149 15555 34207 15561
rect 34149 15552 34161 15555
rect 33468 15524 34161 15552
rect 33468 15512 33474 15524
rect 34149 15521 34161 15524
rect 34195 15552 34207 15555
rect 34195 15524 35848 15552
rect 34195 15521 34207 15524
rect 34149 15515 34207 15521
rect 30837 15487 30895 15493
rect 30837 15453 30849 15487
rect 30883 15453 30895 15487
rect 30837 15447 30895 15453
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15453 30987 15487
rect 30929 15447 30987 15453
rect 30944 15416 30972 15447
rect 33962 15444 33968 15496
rect 34020 15444 34026 15496
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 34793 15487 34851 15493
rect 34793 15484 34805 15487
rect 34756 15456 34805 15484
rect 34756 15444 34762 15456
rect 34793 15453 34805 15456
rect 34839 15453 34851 15487
rect 34793 15447 34851 15453
rect 34882 15444 34888 15496
rect 34940 15484 34946 15496
rect 35526 15484 35532 15496
rect 34940 15456 35532 15484
rect 34940 15444 34946 15456
rect 35526 15444 35532 15456
rect 35584 15444 35590 15496
rect 30760 15388 30972 15416
rect 31205 15419 31263 15425
rect 30561 15379 30619 15385
rect 31205 15385 31217 15419
rect 31251 15416 31263 15419
rect 31478 15416 31484 15428
rect 31251 15388 31484 15416
rect 31251 15385 31263 15388
rect 31205 15379 31263 15385
rect 30285 15351 30343 15357
rect 30285 15317 30297 15351
rect 30331 15317 30343 15351
rect 30285 15311 30343 15317
rect 30374 15308 30380 15360
rect 30432 15348 30438 15360
rect 30576 15348 30604 15379
rect 31478 15376 31484 15388
rect 31536 15376 31542 15428
rect 32490 15416 32496 15428
rect 32430 15388 32496 15416
rect 32490 15376 32496 15388
rect 32548 15416 32554 15428
rect 33318 15416 33324 15428
rect 32548 15388 33324 15416
rect 32548 15376 32554 15388
rect 33318 15376 33324 15388
rect 33376 15376 33382 15428
rect 34057 15419 34115 15425
rect 34057 15385 34069 15419
rect 34103 15416 34115 15419
rect 34900 15416 34928 15444
rect 34103 15388 34928 15416
rect 34103 15385 34115 15388
rect 34057 15379 34115 15385
rect 30432 15320 30604 15348
rect 30432 15308 30438 15320
rect 31846 15308 31852 15360
rect 31904 15348 31910 15360
rect 32950 15348 32956 15360
rect 31904 15320 32956 15348
rect 31904 15308 31910 15320
rect 32950 15308 32956 15320
rect 33008 15308 33014 15360
rect 35434 15308 35440 15360
rect 35492 15348 35498 15360
rect 35713 15351 35771 15357
rect 35713 15348 35725 15351
rect 35492 15320 35725 15348
rect 35492 15308 35498 15320
rect 35713 15317 35725 15320
rect 35759 15317 35771 15351
rect 35820 15348 35848 15524
rect 37182 15512 37188 15564
rect 37240 15512 37246 15564
rect 37384 15552 37412 15660
rect 40218 15648 40224 15700
rect 40276 15648 40282 15700
rect 41966 15620 41972 15632
rect 40604 15592 41972 15620
rect 40604 15561 40632 15592
rect 41966 15580 41972 15592
rect 42024 15620 42030 15632
rect 42024 15592 42104 15620
rect 42024 15580 42030 15592
rect 42076 15561 42104 15592
rect 40589 15555 40647 15561
rect 37384 15524 40540 15552
rect 37458 15444 37464 15496
rect 37516 15484 37522 15496
rect 38562 15484 38568 15496
rect 37516 15456 38568 15484
rect 37516 15444 37522 15456
rect 38562 15444 38568 15456
rect 38620 15484 38626 15496
rect 39025 15487 39083 15493
rect 39025 15484 39037 15487
rect 38620 15456 39037 15484
rect 38620 15444 38626 15456
rect 39025 15453 39037 15456
rect 39071 15453 39083 15487
rect 39025 15447 39083 15453
rect 40402 15444 40408 15496
rect 40460 15444 40466 15496
rect 40512 15484 40540 15524
rect 40589 15521 40601 15555
rect 40635 15521 40647 15555
rect 41509 15555 41567 15561
rect 41509 15552 41521 15555
rect 40589 15515 40647 15521
rect 40972 15524 41521 15552
rect 40972 15493 41000 15524
rect 41509 15521 41521 15524
rect 41555 15521 41567 15555
rect 41509 15515 41567 15521
rect 42061 15555 42119 15561
rect 42061 15521 42073 15555
rect 42107 15521 42119 15555
rect 42061 15515 42119 15521
rect 40773 15487 40831 15493
rect 40773 15484 40785 15487
rect 40512 15456 40785 15484
rect 40773 15453 40785 15456
rect 40819 15453 40831 15487
rect 40773 15447 40831 15453
rect 40957 15487 41015 15493
rect 40957 15453 40969 15487
rect 41003 15453 41015 15487
rect 40957 15447 41015 15453
rect 41141 15487 41199 15493
rect 41141 15453 41153 15487
rect 41187 15453 41199 15487
rect 41141 15447 41199 15453
rect 37826 15416 37832 15428
rect 36754 15388 37832 15416
rect 37826 15376 37832 15388
rect 37884 15376 37890 15428
rect 38286 15376 38292 15428
rect 38344 15376 38350 15428
rect 40494 15376 40500 15428
rect 40552 15416 40558 15428
rect 40862 15416 40868 15428
rect 40552 15388 40868 15416
rect 40552 15376 40558 15388
rect 40862 15376 40868 15388
rect 40920 15416 40926 15428
rect 41049 15419 41107 15425
rect 41049 15416 41061 15419
rect 40920 15388 41061 15416
rect 40920 15376 40926 15388
rect 41049 15385 41061 15388
rect 41095 15385 41107 15419
rect 41156 15416 41184 15447
rect 41506 15416 41512 15428
rect 41156 15388 41512 15416
rect 41049 15379 41107 15385
rect 41506 15376 41512 15388
rect 41564 15376 41570 15428
rect 38470 15348 38476 15360
rect 35820 15320 38476 15348
rect 35713 15311 35771 15317
rect 38470 15308 38476 15320
rect 38528 15308 38534 15360
rect 41325 15351 41383 15357
rect 41325 15317 41337 15351
rect 41371 15348 41383 15351
rect 41414 15348 41420 15360
rect 41371 15320 41420 15348
rect 41371 15317 41383 15320
rect 41325 15311 41383 15317
rect 41414 15308 41420 15320
rect 41472 15308 41478 15360
rect 1104 15258 42504 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 42504 15258
rect 1104 15184 42504 15206
rect 3234 15153 3240 15156
rect 3191 15147 3240 15153
rect 3191 15113 3203 15147
rect 3237 15113 3240 15147
rect 3191 15107 3240 15113
rect 3234 15104 3240 15107
rect 3292 15104 3298 15156
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 6089 15147 6147 15153
rect 6089 15144 6101 15147
rect 5868 15116 6101 15144
rect 5868 15104 5874 15116
rect 6089 15113 6101 15116
rect 6135 15113 6147 15147
rect 6089 15107 6147 15113
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 6822 15144 6828 15156
rect 6236 15116 6828 15144
rect 6236 15104 6242 15116
rect 6822 15104 6828 15116
rect 6880 15144 6886 15156
rect 10226 15144 10232 15156
rect 6880 15116 7972 15144
rect 6880 15104 6886 15116
rect 2590 15036 2596 15088
rect 2648 15036 2654 15088
rect 7024 15076 7052 15116
rect 7944 15076 7972 15116
rect 8404 15116 10232 15144
rect 8404 15076 8432 15116
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 12066 15144 12072 15156
rect 11204 15116 12072 15144
rect 11204 15104 11210 15116
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14792 15116 15025 15144
rect 14792 15104 14798 15116
rect 15013 15113 15025 15116
rect 15059 15113 15071 15147
rect 15013 15107 15071 15113
rect 18049 15147 18107 15153
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 19426 15144 19432 15156
rect 18095 15116 19432 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 20625 15147 20683 15153
rect 20625 15113 20637 15147
rect 20671 15144 20683 15147
rect 20714 15144 20720 15156
rect 20671 15116 20720 15144
rect 20671 15113 20683 15116
rect 20625 15107 20683 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 21358 15144 21364 15156
rect 20864 15116 21364 15144
rect 20864 15104 20870 15116
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 23290 15104 23296 15156
rect 23348 15144 23354 15156
rect 23348 15116 32168 15144
rect 23348 15104 23354 15116
rect 11241 15079 11299 15085
rect 7024 15048 7130 15076
rect 7944 15048 8510 15076
rect 11241 15045 11253 15079
rect 11287 15076 11299 15079
rect 11762 15079 11820 15085
rect 11762 15076 11774 15079
rect 11287 15048 11774 15076
rect 11287 15045 11299 15048
rect 11241 15039 11299 15045
rect 11762 15045 11774 15048
rect 11808 15045 11820 15079
rect 11762 15039 11820 15045
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 17736 15048 18354 15076
rect 17736 15036 17742 15048
rect 19518 15036 19524 15088
rect 19576 15036 19582 15088
rect 20257 15079 20315 15085
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 20303 15048 21833 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 21821 15039 21879 15045
rect 23106 15036 23112 15088
rect 23164 15076 23170 15088
rect 23164 15062 23414 15076
rect 23164 15048 23428 15062
rect 23164 15036 23170 15048
rect 1394 14968 1400 15020
rect 1452 14968 1458 15020
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 1854 15008 1860 15020
rect 1811 14980 1860 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 11112 14980 11161 15008
rect 11112 14968 11118 14980
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 11330 14968 11336 15020
rect 11388 14968 11394 15020
rect 11514 14968 11520 15020
rect 11572 14968 11578 15020
rect 13906 15017 13912 15020
rect 13900 15008 13912 15017
rect 13867 14980 13912 15008
rect 13900 14971 13912 14980
rect 13906 14968 13912 14971
rect 13964 14968 13970 15020
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 20036 14980 20085 15008
rect 20036 14968 20042 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20162 14968 20168 15020
rect 20220 15008 20226 15020
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20220 14980 20361 15008
rect 20220 14968 20226 14980
rect 20349 14977 20361 14980
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 15008 20499 15011
rect 21450 15008 21456 15020
rect 20487 14980 21456 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14940 5595 14943
rect 5810 14940 5816 14952
rect 5583 14912 5816 14940
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 6362 14900 6368 14952
rect 6420 14900 6426 14952
rect 6638 14900 6644 14952
rect 6696 14900 6702 14952
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9953 14943 10011 14949
rect 9723 14912 9904 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 9876 14872 9904 14912
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 11532 14940 11560 14968
rect 9999 14912 11560 14940
rect 13633 14943 13691 14949
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 13633 14909 13645 14943
rect 13679 14909 13691 14943
rect 19797 14943 19855 14949
rect 19797 14940 19809 14943
rect 13633 14903 13691 14909
rect 19720 14912 19809 14940
rect 10318 14872 10324 14884
rect 9876 14844 10324 14872
rect 10318 14832 10324 14844
rect 10376 14832 10382 14884
rect 8110 14764 8116 14816
rect 8168 14764 8174 14816
rect 8205 14807 8263 14813
rect 8205 14773 8217 14807
rect 8251 14804 8263 14807
rect 9674 14804 9680 14816
rect 8251 14776 9680 14804
rect 8251 14773 8263 14776
rect 8205 14767 8263 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 12894 14764 12900 14816
rect 12952 14764 12958 14816
rect 13648 14804 13676 14903
rect 15470 14872 15476 14884
rect 14936 14844 15476 14872
rect 13906 14804 13912 14816
rect 13648 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14804 13970 14816
rect 14936 14804 14964 14844
rect 15470 14832 15476 14844
rect 15528 14832 15534 14884
rect 13964 14776 14964 14804
rect 13964 14764 13970 14776
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19720 14804 19748 14912
rect 19797 14909 19809 14912
rect 19843 14909 19855 14943
rect 20364 14940 20392 14971
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 22060 14980 22385 15008
rect 22060 14968 22066 14980
rect 22373 14977 22385 14980
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 20364 14912 20668 14940
rect 19797 14903 19855 14909
rect 20640 14872 20668 14912
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 21269 14943 21327 14949
rect 21269 14940 21281 14943
rect 20772 14912 21281 14940
rect 20772 14900 20778 14912
rect 21269 14909 21281 14912
rect 21315 14909 21327 14943
rect 23400 14940 23428 15048
rect 24486 15036 24492 15088
rect 24544 15076 24550 15088
rect 24544 15048 25254 15076
rect 24544 15036 24550 15048
rect 26142 15036 26148 15088
rect 26200 15076 26206 15088
rect 28813 15079 28871 15085
rect 26200 15048 26740 15076
rect 26200 15036 26206 15048
rect 26712 15017 26740 15048
rect 28813 15045 28825 15079
rect 28859 15076 28871 15079
rect 29546 15076 29552 15088
rect 28859 15048 29552 15076
rect 28859 15045 28871 15048
rect 28813 15039 28871 15045
rect 29546 15036 29552 15048
rect 29604 15036 29610 15088
rect 29638 15036 29644 15088
rect 29696 15076 29702 15088
rect 29696 15048 29946 15076
rect 29696 15036 29702 15048
rect 31202 15036 31208 15088
rect 31260 15076 31266 15088
rect 32140 15085 32168 15116
rect 32214 15104 32220 15156
rect 32272 15144 32278 15156
rect 36538 15144 36544 15156
rect 32272 15116 36544 15144
rect 32272 15104 32278 15116
rect 33888 15085 33916 15116
rect 36538 15104 36544 15116
rect 36596 15144 36602 15156
rect 38286 15144 38292 15156
rect 36596 15116 38292 15144
rect 36596 15104 36602 15116
rect 38286 15104 38292 15116
rect 38344 15104 38350 15156
rect 38562 15104 38568 15156
rect 38620 15144 38626 15156
rect 38620 15116 39528 15144
rect 38620 15104 38626 15116
rect 32125 15079 32183 15085
rect 31260 15048 31432 15076
rect 31260 15036 31266 15048
rect 26697 15011 26755 15017
rect 26697 14977 26709 15011
rect 26743 14977 26755 15011
rect 26697 14971 26755 14977
rect 27522 14968 27528 15020
rect 27580 15008 27586 15020
rect 27580 14994 27738 15008
rect 27580 14980 27752 14994
rect 27580 14968 27586 14980
rect 24486 14940 24492 14952
rect 23400 14912 24492 14940
rect 21269 14903 21327 14909
rect 24486 14900 24492 14912
rect 24544 14900 24550 14952
rect 24578 14900 24584 14952
rect 24636 14900 24642 14952
rect 24854 14900 24860 14952
rect 24912 14900 24918 14952
rect 24946 14900 24952 14952
rect 25004 14900 25010 14952
rect 26418 14900 26424 14952
rect 26476 14900 26482 14952
rect 27341 14943 27399 14949
rect 27341 14909 27353 14943
rect 27387 14940 27399 14943
rect 27614 14940 27620 14952
rect 27387 14912 27620 14940
rect 27387 14909 27399 14912
rect 27341 14903 27399 14909
rect 27614 14900 27620 14912
rect 27672 14900 27678 14952
rect 27724 14940 27752 14980
rect 29178 14968 29184 15020
rect 29236 14968 29242 15020
rect 27724 14912 29040 14940
rect 23566 14872 23572 14884
rect 20640 14844 23572 14872
rect 23566 14832 23572 14844
rect 23624 14832 23630 14884
rect 29012 14872 29040 14912
rect 29086 14900 29092 14952
rect 29144 14900 29150 14952
rect 29546 14940 29552 14952
rect 29196 14912 29552 14940
rect 29196 14872 29224 14912
rect 29546 14900 29552 14912
rect 29604 14940 29610 14952
rect 29656 14940 29684 15036
rect 31404 15017 31432 15048
rect 32125 15045 32137 15079
rect 32171 15045 32183 15079
rect 32125 15039 32183 15045
rect 33873 15079 33931 15085
rect 33873 15045 33885 15079
rect 33919 15045 33931 15079
rect 33873 15039 33931 15045
rect 34425 15079 34483 15085
rect 34425 15045 34437 15079
rect 34471 15076 34483 15079
rect 35342 15076 35348 15088
rect 34471 15048 35348 15076
rect 34471 15045 34483 15048
rect 34425 15039 34483 15045
rect 35342 15036 35348 15048
rect 35400 15036 35406 15088
rect 37826 15036 37832 15088
rect 37884 15076 37890 15088
rect 37884 15048 38042 15076
rect 37884 15036 37890 15048
rect 31389 15011 31447 15017
rect 31389 14977 31401 15011
rect 31435 14977 31447 15011
rect 31389 14971 31447 14977
rect 31570 14968 31576 15020
rect 31628 14968 31634 15020
rect 34238 14968 34244 15020
rect 34296 14968 34302 15020
rect 34517 15011 34575 15017
rect 34517 14977 34529 15011
rect 34563 14977 34575 15011
rect 34517 14971 34575 14977
rect 34609 15011 34667 15017
rect 34609 14977 34621 15011
rect 34655 15008 34667 15011
rect 35434 15008 35440 15020
rect 34655 14980 35440 15008
rect 34655 14977 34667 14980
rect 34609 14971 34667 14977
rect 29604 14912 29684 14940
rect 31113 14943 31171 14949
rect 29604 14900 29610 14912
rect 31113 14909 31125 14943
rect 31159 14940 31171 14943
rect 32766 14940 32772 14952
rect 31159 14912 32772 14940
rect 31159 14909 31171 14912
rect 31113 14903 31171 14909
rect 32766 14900 32772 14912
rect 32824 14900 32830 14952
rect 33134 14900 33140 14952
rect 33192 14940 33198 14952
rect 34532 14940 34560 14971
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 35989 15011 36047 15017
rect 35989 14977 36001 15011
rect 36035 15008 36047 15011
rect 36078 15008 36084 15020
rect 36035 14980 36084 15008
rect 36035 14977 36047 14980
rect 35989 14971 36047 14977
rect 36078 14968 36084 14980
rect 36136 14968 36142 15020
rect 39500 15017 39528 15116
rect 40034 15104 40040 15156
rect 40092 15144 40098 15156
rect 40402 15144 40408 15156
rect 40092 15116 40408 15144
rect 40092 15104 40098 15116
rect 40402 15104 40408 15116
rect 40460 15144 40466 15156
rect 40460 15116 41828 15144
rect 40460 15104 40466 15116
rect 39485 15011 39543 15017
rect 39485 14977 39497 15011
rect 39531 14977 39543 15011
rect 39485 14971 39543 14977
rect 40218 14968 40224 15020
rect 40276 15008 40282 15020
rect 40497 15011 40555 15017
rect 40497 15008 40509 15011
rect 40276 14980 40509 15008
rect 40276 14968 40282 14980
rect 40497 14977 40509 14980
rect 40543 14977 40555 15011
rect 40497 14971 40555 14977
rect 40586 14968 40592 15020
rect 40644 15008 40650 15020
rect 40773 15011 40831 15017
rect 40773 15008 40785 15011
rect 40644 14980 40785 15008
rect 40644 14968 40650 14980
rect 40773 14977 40785 14980
rect 40819 14977 40831 15011
rect 40773 14971 40831 14977
rect 40957 15011 41015 15017
rect 40957 14977 40969 15011
rect 41003 14977 41015 15011
rect 40957 14971 41015 14977
rect 33192 14912 34560 14940
rect 33192 14900 33198 14912
rect 34882 14900 34888 14952
rect 34940 14900 34946 14952
rect 35897 14943 35955 14949
rect 35897 14909 35909 14943
rect 35943 14909 35955 14943
rect 35897 14903 35955 14909
rect 29641 14875 29699 14881
rect 29012 14844 29224 14872
rect 29288 14844 29592 14872
rect 19484 14776 19748 14804
rect 19484 14764 19490 14776
rect 20714 14764 20720 14816
rect 20772 14764 20778 14816
rect 23109 14807 23167 14813
rect 23109 14773 23121 14807
rect 23155 14804 23167 14807
rect 24762 14804 24768 14816
rect 23155 14776 24768 14804
rect 23155 14773 23167 14776
rect 23109 14767 23167 14773
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 28074 14764 28080 14816
rect 28132 14804 28138 14816
rect 29288 14804 29316 14844
rect 28132 14776 29316 14804
rect 29365 14807 29423 14813
rect 28132 14764 28138 14776
rect 29365 14773 29377 14807
rect 29411 14804 29423 14807
rect 29454 14804 29460 14816
rect 29411 14776 29460 14804
rect 29411 14773 29423 14776
rect 29365 14767 29423 14773
rect 29454 14764 29460 14776
rect 29512 14764 29518 14816
rect 29564 14804 29592 14844
rect 29641 14841 29653 14875
rect 29687 14872 29699 14875
rect 29914 14872 29920 14884
rect 29687 14844 29920 14872
rect 29687 14841 29699 14844
rect 29641 14835 29699 14841
rect 29914 14832 29920 14844
rect 29972 14832 29978 14884
rect 31849 14875 31907 14881
rect 31849 14872 31861 14875
rect 31726 14844 31861 14872
rect 31726 14804 31754 14844
rect 31849 14841 31861 14844
rect 31895 14872 31907 14875
rect 33410 14872 33416 14884
rect 31895 14844 33416 14872
rect 31895 14841 31907 14844
rect 31849 14835 31907 14841
rect 33410 14832 33416 14844
rect 33468 14832 33474 14884
rect 34698 14832 34704 14884
rect 34756 14872 34762 14884
rect 34793 14875 34851 14881
rect 34793 14872 34805 14875
rect 34756 14844 34805 14872
rect 34756 14832 34762 14844
rect 34793 14841 34805 14844
rect 34839 14841 34851 14875
rect 35912 14872 35940 14903
rect 36446 14900 36452 14952
rect 36504 14900 36510 14952
rect 37093 14943 37151 14949
rect 37093 14909 37105 14943
rect 37139 14940 37151 14943
rect 37274 14940 37280 14952
rect 37139 14912 37280 14940
rect 37139 14909 37151 14912
rect 37093 14903 37151 14909
rect 37274 14900 37280 14912
rect 37332 14900 37338 14952
rect 37737 14943 37795 14949
rect 37737 14909 37749 14943
rect 37783 14940 37795 14943
rect 37826 14940 37832 14952
rect 37783 14912 37832 14940
rect 37783 14909 37795 14912
rect 37737 14903 37795 14909
rect 37826 14900 37832 14912
rect 37884 14900 37890 14952
rect 39209 14943 39267 14949
rect 39209 14909 39221 14943
rect 39255 14940 39267 14943
rect 39577 14943 39635 14949
rect 39577 14940 39589 14943
rect 39255 14912 39589 14940
rect 39255 14909 39267 14912
rect 39209 14903 39267 14909
rect 39577 14909 39589 14912
rect 39623 14909 39635 14943
rect 39577 14903 39635 14909
rect 40126 14900 40132 14952
rect 40184 14900 40190 14952
rect 35912 14844 37872 14872
rect 34793 14835 34851 14841
rect 29564 14776 31754 14804
rect 36265 14807 36323 14813
rect 36265 14773 36277 14807
rect 36311 14804 36323 14807
rect 37642 14804 37648 14816
rect 36311 14776 37648 14804
rect 36311 14773 36323 14776
rect 36265 14767 36323 14773
rect 37642 14764 37648 14776
rect 37700 14764 37706 14816
rect 37844 14804 37872 14844
rect 39850 14832 39856 14884
rect 39908 14872 39914 14884
rect 40972 14872 41000 14971
rect 41414 14968 41420 15020
rect 41472 15008 41478 15020
rect 41800 15017 41828 15116
rect 41601 15011 41659 15017
rect 41601 15008 41613 15011
rect 41472 14980 41613 15008
rect 41472 14968 41478 14980
rect 41601 14977 41613 14980
rect 41647 14977 41659 15011
rect 41601 14971 41659 14977
rect 41785 15011 41843 15017
rect 41785 14977 41797 15011
rect 41831 14977 41843 15011
rect 41785 14971 41843 14977
rect 41966 14968 41972 15020
rect 42024 14968 42030 15020
rect 41598 14872 41604 14884
rect 39908 14844 41604 14872
rect 39908 14832 39914 14844
rect 41598 14832 41604 14844
rect 41656 14872 41662 14884
rect 41785 14875 41843 14881
rect 41785 14872 41797 14875
rect 41656 14844 41797 14872
rect 41656 14832 41662 14844
rect 41785 14841 41797 14844
rect 41831 14841 41843 14875
rect 41785 14835 41843 14841
rect 40313 14807 40371 14813
rect 40313 14804 40325 14807
rect 37844 14776 40325 14804
rect 40313 14773 40325 14776
rect 40359 14773 40371 14807
rect 40313 14767 40371 14773
rect 40678 14764 40684 14816
rect 40736 14804 40742 14816
rect 41049 14807 41107 14813
rect 41049 14804 41061 14807
rect 40736 14776 41061 14804
rect 40736 14764 40742 14776
rect 41049 14773 41061 14776
rect 41095 14773 41107 14807
rect 41049 14767 41107 14773
rect 1104 14714 42504 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 42504 14714
rect 1104 14640 42504 14662
rect 4985 14603 5043 14609
rect 4985 14569 4997 14603
rect 5031 14600 5043 14603
rect 5810 14600 5816 14612
rect 5031 14572 5816 14600
rect 5031 14569 5043 14572
rect 4985 14563 5043 14569
rect 5810 14560 5816 14572
rect 5868 14600 5874 14612
rect 6638 14600 6644 14612
rect 5868 14572 6644 14600
rect 5868 14560 5874 14572
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 9858 14560 9864 14612
rect 9916 14560 9922 14612
rect 10318 14560 10324 14612
rect 10376 14560 10382 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 11388 14572 11529 14600
rect 11388 14560 11394 14572
rect 11517 14569 11529 14572
rect 11563 14600 11575 14603
rect 11974 14600 11980 14612
rect 11563 14572 11980 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 14921 14603 14979 14609
rect 14921 14600 14933 14603
rect 14700 14572 14933 14600
rect 14700 14560 14706 14572
rect 14921 14569 14933 14572
rect 14967 14600 14979 14603
rect 14967 14572 17264 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 10410 14532 10416 14544
rect 7760 14504 10416 14532
rect 2225 14467 2283 14473
rect 2225 14433 2237 14467
rect 2271 14464 2283 14467
rect 7760 14464 7788 14504
rect 10410 14492 10416 14504
rect 10468 14492 10474 14544
rect 2271 14436 7788 14464
rect 2271 14433 2283 14436
rect 2225 14427 2283 14433
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 8389 14467 8447 14473
rect 8389 14464 8401 14467
rect 8168 14436 8401 14464
rect 8168 14424 8174 14436
rect 8389 14433 8401 14436
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 11885 14467 11943 14473
rect 8711 14436 10180 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2498 14396 2504 14408
rect 2179 14368 2504 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2498 14356 2504 14368
rect 2556 14396 2562 14408
rect 3970 14396 3976 14408
rect 2556 14368 3976 14396
rect 2556 14356 2562 14368
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 7374 14396 7380 14408
rect 6779 14368 7380 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 4672 14300 5290 14328
rect 4672 14288 4678 14300
rect 6454 14288 6460 14340
rect 6512 14288 6518 14340
rect 6546 14288 6552 14340
rect 6604 14328 6610 14340
rect 6748 14328 6776 14359
rect 7374 14356 7380 14368
rect 7432 14396 7438 14408
rect 7561 14399 7619 14405
rect 7561 14396 7573 14399
rect 7432 14368 7573 14396
rect 7432 14356 7438 14368
rect 7561 14365 7573 14368
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 8573 14399 8631 14405
rect 8573 14396 8585 14399
rect 8536 14368 8585 14396
rect 8536 14356 8542 14368
rect 8573 14365 8585 14368
rect 8619 14365 8631 14399
rect 8573 14359 8631 14365
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14396 8815 14399
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8803 14368 8953 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 9490 14356 9496 14408
rect 9548 14356 9554 14408
rect 9646 14396 9904 14398
rect 9600 14370 9904 14396
rect 9600 14368 9674 14370
rect 6604 14300 6776 14328
rect 6825 14331 6883 14337
rect 6604 14288 6610 14300
rect 6825 14297 6837 14331
rect 6871 14297 6883 14331
rect 9600 14328 9628 14368
rect 6825 14291 6883 14297
rect 7668 14300 9628 14328
rect 2501 14263 2559 14269
rect 2501 14229 2513 14263
rect 2547 14260 2559 14263
rect 2682 14260 2688 14272
rect 2547 14232 2688 14260
rect 2547 14229 2559 14232
rect 2501 14223 2559 14229
rect 2682 14220 2688 14232
rect 2740 14220 2746 14272
rect 5442 14220 5448 14272
rect 5500 14260 5506 14272
rect 6840 14260 6868 14291
rect 7668 14260 7696 14300
rect 9699 14288 9705 14340
rect 9757 14328 9763 14340
rect 9876 14328 9904 14370
rect 9950 14356 9956 14408
rect 10008 14356 10014 14408
rect 10152 14405 10180 14436
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12894 14464 12900 14476
rect 11931 14436 12900 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 17236 14473 17264 14572
rect 22002 14560 22008 14612
rect 22060 14600 22066 14612
rect 24121 14603 24179 14609
rect 22060 14560 22094 14600
rect 24121 14569 24133 14603
rect 24167 14600 24179 14603
rect 24302 14600 24308 14612
rect 24167 14572 24308 14600
rect 24167 14569 24179 14572
rect 24121 14563 24179 14569
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 24578 14560 24584 14612
rect 24636 14600 24642 14612
rect 25041 14603 25099 14609
rect 25041 14600 25053 14603
rect 24636 14572 25053 14600
rect 24636 14560 24642 14572
rect 25041 14569 25053 14572
rect 25087 14569 25099 14603
rect 25041 14563 25099 14569
rect 25682 14560 25688 14612
rect 25740 14600 25746 14612
rect 26878 14600 26884 14612
rect 25740 14572 26884 14600
rect 25740 14560 25746 14572
rect 26878 14560 26884 14572
rect 26936 14600 26942 14612
rect 27706 14600 27712 14612
rect 26936 14572 27712 14600
rect 26936 14560 26942 14572
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 28258 14560 28264 14612
rect 28316 14600 28322 14612
rect 32214 14600 32220 14612
rect 28316 14572 32220 14600
rect 28316 14560 28322 14572
rect 32214 14560 32220 14572
rect 32272 14560 32278 14612
rect 32306 14560 32312 14612
rect 32364 14600 32370 14612
rect 32677 14603 32735 14609
rect 32677 14600 32689 14603
rect 32364 14572 32689 14600
rect 32364 14560 32370 14572
rect 32677 14569 32689 14572
rect 32723 14569 32735 14603
rect 32677 14563 32735 14569
rect 32766 14560 32772 14612
rect 32824 14560 32830 14612
rect 36262 14600 36268 14612
rect 36188 14572 36268 14600
rect 22066 14532 22094 14560
rect 22189 14535 22247 14541
rect 22189 14532 22201 14535
rect 22066 14504 22201 14532
rect 22189 14501 22201 14504
rect 22235 14501 22247 14535
rect 22189 14495 22247 14501
rect 24486 14492 24492 14544
rect 24544 14532 24550 14544
rect 26237 14535 26295 14541
rect 26237 14532 26249 14535
rect 24544 14504 26249 14532
rect 24544 14492 24550 14504
rect 26237 14501 26249 14504
rect 26283 14532 26295 14535
rect 26510 14532 26516 14544
rect 26283 14504 26516 14532
rect 26283 14501 26295 14504
rect 26237 14495 26295 14501
rect 26510 14492 26516 14504
rect 26568 14492 26574 14544
rect 26697 14535 26755 14541
rect 26697 14501 26709 14535
rect 26743 14532 26755 14535
rect 27246 14532 27252 14544
rect 26743 14504 27252 14532
rect 26743 14501 26755 14504
rect 26697 14495 26755 14501
rect 27246 14492 27252 14504
rect 27304 14492 27310 14544
rect 29362 14492 29368 14544
rect 29420 14532 29426 14544
rect 29549 14535 29607 14541
rect 29549 14532 29561 14535
rect 29420 14504 29561 14532
rect 29420 14492 29426 14504
rect 29549 14501 29561 14504
rect 29595 14501 29607 14535
rect 29549 14495 29607 14501
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14433 17279 14467
rect 17221 14427 17279 14433
rect 17402 14424 17408 14476
rect 17460 14424 17466 14476
rect 20714 14424 20720 14476
rect 20772 14424 20778 14476
rect 22373 14467 22431 14473
rect 22373 14433 22385 14467
rect 22419 14464 22431 14467
rect 24854 14464 24860 14476
rect 22419 14436 24860 14464
rect 22419 14433 22431 14436
rect 22373 14427 22431 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 25130 14424 25136 14476
rect 25188 14464 25194 14476
rect 25188 14436 26004 14464
rect 25188 14424 25194 14436
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10318 14356 10324 14408
rect 10376 14356 10382 14408
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14396 11759 14399
rect 12066 14396 12072 14408
rect 11747 14368 12072 14396
rect 11747 14365 11759 14368
rect 11701 14359 11759 14365
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 18509 14399 18567 14405
rect 18509 14365 18521 14399
rect 18555 14396 18567 14399
rect 18598 14396 18604 14408
rect 18555 14368 18604 14396
rect 18555 14365 18567 14368
rect 18509 14359 18567 14365
rect 18598 14356 18604 14368
rect 18656 14396 18662 14408
rect 19886 14396 19892 14408
rect 18656 14368 19892 14396
rect 18656 14356 18662 14368
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 9968 14328 9996 14356
rect 11422 14328 11428 14340
rect 9757 14300 9802 14328
rect 9876 14300 11428 14328
rect 9757 14288 9763 14300
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 16393 14331 16451 14337
rect 15962 14300 16344 14328
rect 16316 14272 16344 14300
rect 16393 14297 16405 14331
rect 16439 14297 16451 14331
rect 16393 14291 16451 14297
rect 5500 14232 7696 14260
rect 5500 14220 5506 14232
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 7837 14263 7895 14269
rect 7837 14260 7849 14263
rect 7800 14232 7849 14260
rect 7800 14220 7806 14232
rect 7837 14229 7849 14232
rect 7883 14229 7895 14263
rect 7837 14223 7895 14229
rect 9214 14220 9220 14272
rect 9272 14260 9278 14272
rect 9877 14263 9935 14269
rect 9877 14260 9889 14263
rect 9272 14232 9889 14260
rect 9272 14220 9278 14232
rect 9877 14229 9889 14232
rect 9923 14229 9935 14263
rect 9877 14223 9935 14229
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10318 14260 10324 14272
rect 10100 14232 10324 14260
rect 10100 14220 10106 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 13722 14260 13728 14272
rect 13679 14232 13728 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 16298 14220 16304 14272
rect 16356 14220 16362 14272
rect 16408 14260 16436 14291
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 18141 14331 18199 14337
rect 18141 14328 18153 14331
rect 18012 14300 18153 14328
rect 18012 14288 18018 14300
rect 18141 14297 18153 14300
rect 18187 14297 18199 14331
rect 18141 14291 18199 14297
rect 18877 14331 18935 14337
rect 18877 14297 18889 14331
rect 18923 14297 18935 14331
rect 20456 14328 20484 14359
rect 24394 14356 24400 14408
rect 24452 14356 24458 14408
rect 24762 14356 24768 14408
rect 24820 14396 24826 14408
rect 25976 14405 26004 14436
rect 26142 14424 26148 14476
rect 26200 14464 26206 14476
rect 30929 14467 30987 14473
rect 26200 14436 27200 14464
rect 26200 14424 26206 14436
rect 25685 14399 25743 14405
rect 25685 14396 25697 14399
rect 24820 14368 25697 14396
rect 24820 14356 24826 14368
rect 25685 14365 25697 14368
rect 25731 14365 25743 14399
rect 25685 14359 25743 14365
rect 25961 14399 26019 14405
rect 25961 14365 25973 14399
rect 26007 14365 26019 14399
rect 25961 14359 26019 14365
rect 26326 14356 26332 14408
rect 26384 14396 26390 14408
rect 26421 14399 26479 14405
rect 26421 14396 26433 14399
rect 26384 14368 26433 14396
rect 26384 14356 26390 14368
rect 26421 14365 26433 14368
rect 26467 14365 26479 14399
rect 26421 14359 26479 14365
rect 26697 14399 26755 14405
rect 26697 14365 26709 14399
rect 26743 14396 26755 14399
rect 27062 14396 27068 14408
rect 26743 14368 27068 14396
rect 26743 14365 26755 14368
rect 26697 14359 26755 14365
rect 27062 14356 27068 14368
rect 27120 14356 27126 14408
rect 27172 14405 27200 14436
rect 30929 14433 30941 14467
rect 30975 14464 30987 14467
rect 31202 14464 31208 14476
rect 30975 14436 31208 14464
rect 30975 14433 30987 14436
rect 30929 14427 30987 14433
rect 31202 14424 31208 14436
rect 31260 14424 31266 14476
rect 33226 14424 33232 14476
rect 33284 14424 33290 14476
rect 33410 14424 33416 14476
rect 33468 14424 33474 14476
rect 34517 14467 34575 14473
rect 34517 14433 34529 14467
rect 34563 14464 34575 14467
rect 34698 14464 34704 14476
rect 34563 14436 34704 14464
rect 34563 14433 34575 14436
rect 34517 14427 34575 14433
rect 34698 14424 34704 14436
rect 34756 14424 34762 14476
rect 36188 14473 36216 14572
rect 36262 14560 36268 14572
rect 36320 14560 36326 14612
rect 38197 14603 38255 14609
rect 38197 14569 38209 14603
rect 38243 14600 38255 14603
rect 40126 14600 40132 14612
rect 38243 14572 40132 14600
rect 38243 14569 38255 14572
rect 38197 14563 38255 14569
rect 40126 14560 40132 14572
rect 40184 14560 40190 14612
rect 40494 14560 40500 14612
rect 40552 14560 40558 14612
rect 41966 14560 41972 14612
rect 42024 14600 42030 14612
rect 42153 14603 42211 14609
rect 42153 14600 42165 14603
rect 42024 14572 42165 14600
rect 42024 14560 42030 14572
rect 42153 14569 42165 14572
rect 42199 14569 42211 14603
rect 42153 14563 42211 14569
rect 39945 14535 40003 14541
rect 39945 14501 39957 14535
rect 39991 14532 40003 14535
rect 40218 14532 40224 14544
rect 39991 14504 40224 14532
rect 39991 14501 40003 14504
rect 39945 14495 40003 14501
rect 40218 14492 40224 14504
rect 40276 14492 40282 14544
rect 36173 14467 36231 14473
rect 36173 14433 36185 14467
rect 36219 14433 36231 14467
rect 36173 14427 36231 14433
rect 36354 14424 36360 14476
rect 36412 14464 36418 14476
rect 37093 14467 37151 14473
rect 37093 14464 37105 14467
rect 36412 14436 37105 14464
rect 36412 14424 36418 14436
rect 37093 14433 37105 14436
rect 37139 14433 37151 14467
rect 37093 14427 37151 14433
rect 37182 14424 37188 14476
rect 37240 14464 37246 14476
rect 37553 14467 37611 14473
rect 37553 14464 37565 14467
rect 37240 14436 37565 14464
rect 37240 14424 37246 14436
rect 37553 14433 37565 14436
rect 37599 14433 37611 14467
rect 37553 14427 37611 14433
rect 37737 14467 37795 14473
rect 37737 14433 37749 14467
rect 37783 14464 37795 14467
rect 38194 14464 38200 14476
rect 37783 14436 38200 14464
rect 37783 14433 37795 14436
rect 37737 14427 37795 14433
rect 38194 14424 38200 14436
rect 38252 14424 38258 14476
rect 40129 14467 40187 14473
rect 40129 14433 40141 14467
rect 40175 14464 40187 14467
rect 40512 14464 40540 14560
rect 40175 14436 40540 14464
rect 40175 14433 40187 14436
rect 40129 14427 40187 14433
rect 40678 14424 40684 14476
rect 40736 14424 40742 14476
rect 27157 14399 27215 14405
rect 27157 14365 27169 14399
rect 27203 14365 27215 14399
rect 27157 14359 27215 14365
rect 28258 14356 28264 14408
rect 28316 14356 28322 14408
rect 28350 14356 28356 14408
rect 28408 14396 28414 14408
rect 29454 14396 29460 14408
rect 28408 14368 29460 14396
rect 28408 14356 28414 14368
rect 29454 14356 29460 14368
rect 29512 14356 29518 14408
rect 32490 14396 32496 14408
rect 32338 14368 32496 14396
rect 32490 14356 32496 14368
rect 32548 14396 32554 14408
rect 33962 14396 33968 14408
rect 32548 14368 33968 14396
rect 32548 14356 32554 14368
rect 33962 14356 33968 14368
rect 34020 14356 34026 14408
rect 34330 14356 34336 14408
rect 34388 14396 34394 14408
rect 35253 14399 35311 14405
rect 35253 14396 35265 14399
rect 34388 14368 35265 14396
rect 34388 14356 34394 14368
rect 35253 14365 35265 14368
rect 35299 14365 35311 14399
rect 35253 14359 35311 14365
rect 36081 14399 36139 14405
rect 36081 14365 36093 14399
rect 36127 14396 36139 14399
rect 36446 14396 36452 14408
rect 36127 14368 36452 14396
rect 36127 14365 36139 14368
rect 36081 14359 36139 14365
rect 36446 14356 36452 14368
rect 36504 14356 36510 14408
rect 36722 14356 36728 14408
rect 36780 14396 36786 14408
rect 37001 14399 37059 14405
rect 37001 14396 37013 14399
rect 36780 14368 37013 14396
rect 36780 14356 36786 14368
rect 37001 14365 37013 14368
rect 37047 14365 37059 14399
rect 37001 14359 37059 14365
rect 37458 14356 37464 14408
rect 37516 14396 37522 14408
rect 38378 14396 38384 14408
rect 37516 14368 38384 14396
rect 37516 14356 37522 14368
rect 38378 14356 38384 14368
rect 38436 14356 38442 14408
rect 39850 14356 39856 14408
rect 39908 14356 39914 14408
rect 40405 14399 40463 14405
rect 40405 14365 40417 14399
rect 40451 14365 40463 14399
rect 40405 14359 40463 14365
rect 20622 14328 20628 14340
rect 20456 14300 20628 14328
rect 18877 14291 18935 14297
rect 16761 14263 16819 14269
rect 16761 14260 16773 14263
rect 16408 14232 16773 14260
rect 16761 14229 16773 14232
rect 16807 14229 16819 14263
rect 16761 14223 16819 14229
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17129 14263 17187 14269
rect 17129 14260 17141 14263
rect 17092 14232 17141 14260
rect 17092 14220 17098 14232
rect 17129 14229 17141 14232
rect 17175 14229 17187 14263
rect 17129 14223 17187 14229
rect 18782 14220 18788 14272
rect 18840 14220 18846 14272
rect 18892 14260 18920 14291
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 21174 14328 21180 14340
rect 21048 14300 21180 14328
rect 21048 14288 21054 14300
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 22646 14288 22652 14340
rect 22704 14288 22710 14340
rect 23106 14288 23112 14340
rect 23164 14288 23170 14340
rect 28994 14288 29000 14340
rect 29052 14288 29058 14340
rect 29730 14288 29736 14340
rect 29788 14328 29794 14340
rect 30926 14328 30932 14340
rect 29788 14300 30932 14328
rect 29788 14288 29794 14300
rect 30926 14288 30932 14300
rect 30984 14288 30990 14340
rect 31110 14288 31116 14340
rect 31168 14328 31174 14340
rect 31205 14331 31263 14337
rect 31205 14328 31217 14331
rect 31168 14300 31217 14328
rect 31168 14288 31174 14300
rect 31205 14297 31217 14300
rect 31251 14297 31263 14331
rect 33137 14331 33195 14337
rect 33137 14328 33149 14331
rect 31205 14291 31263 14297
rect 32508 14300 33149 14328
rect 20530 14260 20536 14272
rect 18892 14232 20536 14260
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 25130 14220 25136 14272
rect 25188 14220 25194 14272
rect 26510 14220 26516 14272
rect 26568 14220 26574 14272
rect 29914 14220 29920 14272
rect 29972 14260 29978 14272
rect 32508 14260 32536 14300
rect 33137 14297 33149 14300
rect 33183 14297 33195 14331
rect 33137 14291 33195 14297
rect 33410 14288 33416 14340
rect 33468 14328 33474 14340
rect 34701 14331 34759 14337
rect 34701 14328 34713 14331
rect 33468 14300 34713 14328
rect 33468 14288 33474 14300
rect 34701 14297 34713 14300
rect 34747 14297 34759 14331
rect 38396 14328 38424 14356
rect 40420 14328 40448 14359
rect 41966 14328 41972 14340
rect 38396 14300 40448 14328
rect 41906 14300 41972 14328
rect 34701 14291 34759 14297
rect 41966 14288 41972 14300
rect 42024 14288 42030 14340
rect 29972 14232 32536 14260
rect 33873 14263 33931 14269
rect 29972 14220 29978 14232
rect 33873 14229 33885 14263
rect 33919 14260 33931 14263
rect 34238 14260 34244 14272
rect 33919 14232 34244 14260
rect 33919 14229 33931 14232
rect 33873 14223 33931 14229
rect 34238 14220 34244 14232
rect 34296 14220 34302 14272
rect 35434 14220 35440 14272
rect 35492 14260 35498 14272
rect 35713 14263 35771 14269
rect 35713 14260 35725 14263
rect 35492 14232 35725 14260
rect 35492 14220 35498 14232
rect 35713 14229 35725 14232
rect 35759 14229 35771 14263
rect 35713 14223 35771 14229
rect 36262 14220 36268 14272
rect 36320 14260 36326 14272
rect 36541 14263 36599 14269
rect 36541 14260 36553 14263
rect 36320 14232 36553 14260
rect 36320 14220 36326 14232
rect 36541 14229 36553 14232
rect 36587 14229 36599 14263
rect 36541 14223 36599 14229
rect 36906 14220 36912 14272
rect 36964 14220 36970 14272
rect 37826 14220 37832 14272
rect 37884 14260 37890 14272
rect 39942 14260 39948 14272
rect 37884 14232 39948 14260
rect 37884 14220 37890 14232
rect 39942 14220 39948 14232
rect 40000 14220 40006 14272
rect 40034 14220 40040 14272
rect 40092 14260 40098 14272
rect 40129 14263 40187 14269
rect 40129 14260 40141 14263
rect 40092 14232 40141 14260
rect 40092 14220 40098 14232
rect 40129 14229 40141 14232
rect 40175 14229 40187 14263
rect 40129 14223 40187 14229
rect 1104 14170 42504 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 42504 14170
rect 1104 14096 42504 14118
rect 5718 14056 5724 14068
rect 5368 14028 5724 14056
rect 2682 13948 2688 14000
rect 2740 13948 2746 14000
rect 3970 13948 3976 14000
rect 4028 13988 4034 14000
rect 4433 13991 4491 13997
rect 4433 13988 4445 13991
rect 4028 13960 4445 13988
rect 4028 13948 4034 13960
rect 4433 13957 4445 13960
rect 4479 13957 4491 13991
rect 4433 13951 4491 13957
rect 5368 13929 5396 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6730 14065 6736 14068
rect 6726 14056 6736 14065
rect 6691 14028 6736 14056
rect 6726 14019 6736 14028
rect 6730 14016 6736 14019
rect 6788 14016 6794 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7156 14028 7849 14056
rect 7156 14016 7162 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 12614 14059 12672 14065
rect 12614 14025 12626 14059
rect 12660 14056 12672 14059
rect 12986 14056 12992 14068
rect 12660 14028 12992 14056
rect 12660 14025 12672 14028
rect 12614 14019 12672 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 16574 14056 16580 14068
rect 15488 14028 16580 14056
rect 6825 13991 6883 13997
rect 5552 13960 6776 13988
rect 5552 13929 5580 13960
rect 5353 13923 5411 13929
rect 2406 13812 2412 13864
rect 2464 13812 2470 13864
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3804 13852 3832 13906
rect 5353 13889 5365 13923
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6178 13920 6184 13932
rect 6043 13892 6184 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 5368 13852 5396 13883
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6362 13852 6368 13864
rect 2740 13824 4384 13852
rect 5368 13824 6368 13852
rect 2740 13812 2746 13824
rect 4356 13784 4384 13824
rect 6362 13812 6368 13824
rect 6420 13852 6426 13864
rect 6564 13852 6592 13883
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6748 13920 6776 13960
rect 6825 13957 6837 13991
rect 6871 13988 6883 13991
rect 7742 13988 7748 14000
rect 6871 13960 7748 13988
rect 6871 13957 6883 13960
rect 6825 13951 6883 13957
rect 7742 13948 7748 13960
rect 7800 13948 7806 14000
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 10321 13991 10379 13997
rect 10321 13988 10333 13991
rect 10284 13960 10333 13988
rect 10284 13948 10290 13960
rect 10321 13957 10333 13960
rect 10367 13957 10379 13991
rect 10321 13951 10379 13957
rect 7561 13923 7619 13929
rect 6748 13892 7052 13920
rect 6420 13824 6592 13852
rect 6917 13855 6975 13861
rect 6420 13812 6426 13824
rect 6917 13821 6929 13855
rect 6963 13821 6975 13855
rect 7024 13852 7052 13892
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7653 13923 7711 13929
rect 7653 13920 7665 13923
rect 7607 13892 7665 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 7653 13889 7665 13892
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 11882 13920 11888 13932
rect 10551 13892 11888 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 7024 13824 7696 13852
rect 6917 13815 6975 13821
rect 4614 13784 4620 13796
rect 4356 13756 4620 13784
rect 4614 13744 4620 13756
rect 4672 13784 4678 13796
rect 5721 13787 5779 13793
rect 5721 13784 5733 13787
rect 4672 13756 5733 13784
rect 4672 13744 4678 13756
rect 5721 13753 5733 13756
rect 5767 13753 5779 13787
rect 6932 13784 6960 13815
rect 7374 13784 7380 13796
rect 6932 13756 7380 13784
rect 5721 13747 5779 13753
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 7668 13793 7696 13824
rect 7653 13787 7711 13793
rect 7653 13753 7665 13787
rect 7699 13753 7711 13787
rect 7653 13747 7711 13753
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 4764 13688 5365 13716
rect 4764 13676 4770 13688
rect 5353 13685 5365 13688
rect 5399 13685 5411 13719
rect 5353 13679 5411 13685
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7944 13716 7972 13883
rect 11882 13880 11888 13892
rect 11940 13880 11946 13932
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 12032 13892 12449 13920
rect 12032 13880 12038 13892
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 12526 13880 12532 13932
rect 12584 13880 12590 13932
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 12805 13923 12863 13929
rect 12805 13920 12817 13923
rect 12759 13892 12817 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 12805 13889 12817 13892
rect 12851 13889 12863 13923
rect 12805 13883 12863 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13044 13892 13553 13920
rect 13044 13880 13050 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15488 13920 15516 14028
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 18598 14016 18604 14068
rect 18656 14016 18662 14068
rect 18969 14059 19027 14065
rect 18969 14025 18981 14059
rect 19015 14056 19027 14059
rect 19794 14056 19800 14068
rect 19015 14028 19800 14056
rect 19015 14025 19027 14028
rect 18969 14019 19027 14025
rect 19794 14016 19800 14028
rect 19852 14016 19858 14068
rect 20993 14059 21051 14065
rect 20993 14025 21005 14059
rect 21039 14056 21051 14059
rect 22281 14059 22339 14065
rect 21039 14028 22094 14056
rect 21039 14025 21051 14028
rect 20993 14019 21051 14025
rect 17034 13988 17040 14000
rect 15764 13960 17040 13988
rect 15764 13929 15792 13960
rect 17034 13948 17040 13960
rect 17092 13948 17098 14000
rect 17678 13948 17684 14000
rect 17736 13948 17742 14000
rect 19886 13988 19892 14000
rect 18800 13960 19892 13988
rect 18800 13929 18828 13960
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20346 13948 20352 14000
rect 20404 13988 20410 14000
rect 20533 13991 20591 13997
rect 20533 13988 20545 13991
rect 20404 13960 20545 13988
rect 20404 13948 20410 13960
rect 20533 13957 20545 13960
rect 20579 13957 20591 13991
rect 21266 13988 21272 14000
rect 20533 13951 20591 13957
rect 21008 13960 21272 13988
rect 21008 13932 21036 13960
rect 21266 13948 21272 13960
rect 21324 13948 21330 14000
rect 22066 13988 22094 14028
rect 22281 14025 22293 14059
rect 22327 14056 22339 14059
rect 22462 14056 22468 14068
rect 22327 14028 22468 14056
rect 22327 14025 22339 14028
rect 22281 14019 22339 14025
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 24394 14016 24400 14068
rect 24452 14016 24458 14068
rect 24946 14056 24952 14068
rect 24596 14028 24952 14056
rect 22066 13960 24532 13988
rect 15335 13892 15516 13920
rect 15565 13923 15623 13929
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 15749 13923 15807 13929
rect 15611 13892 15700 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13852 10287 13855
rect 10686 13852 10692 13864
rect 10275 13824 10692 13852
rect 10275 13821 10287 13824
rect 10229 13815 10287 13821
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 15105 13855 15163 13861
rect 15105 13821 15117 13855
rect 15151 13852 15163 13855
rect 15378 13852 15384 13864
rect 15151 13824 15384 13852
rect 15151 13821 15163 13824
rect 15105 13815 15163 13821
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 13372 13784 13400 13815
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15672 13852 15700 13892
rect 15749 13889 15761 13923
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13920 19395 13923
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19383 13892 19809 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 20806 13880 20812 13932
rect 20864 13880 20870 13932
rect 20990 13880 20996 13932
rect 21048 13880 21054 13932
rect 21634 13880 21640 13932
rect 21692 13880 21698 13932
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13920 22247 13923
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 22235 13892 22661 13920
rect 22235 13889 22247 13892
rect 22189 13883 22247 13889
rect 22649 13889 22661 13892
rect 22695 13889 22707 13923
rect 22649 13883 22707 13889
rect 15841 13855 15899 13861
rect 15841 13852 15853 13855
rect 15672 13824 15853 13852
rect 15841 13821 15853 13824
rect 15887 13852 15899 13855
rect 16485 13855 16543 13861
rect 15887 13824 16436 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 12768 13756 13400 13784
rect 16408 13784 16436 13824
rect 16485 13821 16497 13855
rect 16531 13852 16543 13855
rect 16574 13852 16580 13864
rect 16531 13824 16580 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 16666 13812 16672 13864
rect 16724 13812 16730 13864
rect 16942 13812 16948 13864
rect 17000 13812 17006 13864
rect 17678 13812 17684 13864
rect 17736 13852 17742 13864
rect 18966 13852 18972 13864
rect 17736 13824 18972 13852
rect 17736 13812 17742 13824
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19429 13815 19487 13821
rect 19444 13784 19472 13815
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19576 13824 19625 13852
rect 19576 13812 19582 13824
rect 19613 13821 19625 13824
rect 19659 13852 19671 13855
rect 20162 13852 20168 13864
rect 19659 13824 20168 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20349 13855 20407 13861
rect 20349 13852 20361 13855
rect 20312 13824 20361 13852
rect 20312 13812 20318 13824
rect 20349 13821 20361 13824
rect 20395 13821 20407 13855
rect 20349 13815 20407 13821
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 20898 13852 20904 13864
rect 20763 13824 20904 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 22465 13855 22523 13861
rect 22465 13821 22477 13855
rect 22511 13821 22523 13855
rect 22465 13815 22523 13821
rect 19702 13784 19708 13796
rect 16408 13756 16804 13784
rect 19444 13756 19708 13784
rect 12768 13744 12774 13756
rect 16776 13728 16804 13756
rect 19702 13744 19708 13756
rect 19760 13784 19766 13796
rect 19760 13756 20668 13784
rect 19760 13744 19766 13756
rect 6972 13688 7972 13716
rect 6972 13676 6978 13688
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 9585 13719 9643 13725
rect 9585 13716 9597 13719
rect 8444 13688 9597 13716
rect 8444 13676 8450 13688
rect 9585 13685 9597 13688
rect 9631 13685 9643 13719
rect 9585 13679 9643 13685
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 13725 13719 13783 13725
rect 13725 13716 13737 13719
rect 13688 13688 13737 13716
rect 13688 13676 13694 13688
rect 13725 13685 13737 13688
rect 13771 13685 13783 13719
rect 13725 13679 13783 13685
rect 16758 13676 16764 13728
rect 16816 13676 16822 13728
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 20640 13725 20668 13756
rect 21266 13744 21272 13796
rect 21324 13784 21330 13796
rect 22480 13784 22508 13815
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 24504 13852 24532 13960
rect 24596 13929 24624 14028
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 26142 14016 26148 14068
rect 26200 14016 26206 14068
rect 28721 14059 28779 14065
rect 26988 14028 28580 14056
rect 24765 13991 24823 13997
rect 24765 13957 24777 13991
rect 24811 13988 24823 13991
rect 25130 13988 25136 14000
rect 24811 13960 25136 13988
rect 24811 13957 24823 13960
rect 24765 13951 24823 13957
rect 25130 13948 25136 13960
rect 25188 13948 25194 14000
rect 25593 13991 25651 13997
rect 25593 13957 25605 13991
rect 25639 13988 25651 13991
rect 25884 13988 25912 14016
rect 25639 13960 25912 13988
rect 26160 13988 26188 14016
rect 26988 13988 27016 14028
rect 26160 13960 27016 13988
rect 25639 13957 25651 13960
rect 25593 13951 25651 13957
rect 24581 13923 24639 13929
rect 24581 13889 24593 13923
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 24670 13880 24676 13932
rect 24728 13880 24734 13932
rect 24949 13923 25007 13929
rect 24949 13889 24961 13923
rect 24995 13920 25007 13923
rect 25498 13920 25504 13932
rect 24995 13892 25504 13920
rect 24995 13889 25007 13892
rect 24949 13883 25007 13889
rect 25498 13880 25504 13892
rect 25556 13880 25562 13932
rect 25608 13892 25820 13920
rect 25608 13852 25636 13892
rect 24504 13824 25636 13852
rect 25682 13812 25688 13864
rect 25740 13812 25746 13864
rect 25792 13852 25820 13892
rect 25866 13880 25872 13932
rect 25924 13880 25930 13932
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13920 26203 13923
rect 26191 13892 26280 13920
rect 26191 13889 26203 13892
rect 26145 13883 26203 13889
rect 26252 13852 26280 13892
rect 26326 13880 26332 13932
rect 26384 13880 26390 13932
rect 26418 13880 26424 13932
rect 26476 13880 26482 13932
rect 26988 13929 27016 13960
rect 27246 13948 27252 14000
rect 27304 13948 27310 14000
rect 26513 13923 26571 13929
rect 26513 13889 26525 13923
rect 26559 13920 26571 13923
rect 26973 13923 27031 13929
rect 26559 13892 26924 13920
rect 26559 13889 26571 13892
rect 26513 13883 26571 13889
rect 26786 13852 26792 13864
rect 25792 13824 26188 13852
rect 26252 13824 26792 13852
rect 25866 13784 25872 13796
rect 21324 13756 25872 13784
rect 21324 13744 21330 13756
rect 25866 13744 25872 13756
rect 25924 13744 25930 13796
rect 18417 13719 18475 13725
rect 18417 13716 18429 13719
rect 18104 13688 18429 13716
rect 18104 13676 18110 13688
rect 18417 13685 18429 13688
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 20625 13719 20683 13725
rect 20625 13685 20637 13719
rect 20671 13685 20683 13719
rect 20625 13679 20683 13685
rect 21542 13676 21548 13728
rect 21600 13716 21606 13728
rect 21821 13719 21879 13725
rect 21821 13716 21833 13719
rect 21600 13688 21833 13716
rect 21600 13676 21606 13688
rect 21821 13685 21833 13688
rect 21867 13685 21879 13719
rect 21821 13679 21879 13685
rect 25682 13676 25688 13728
rect 25740 13676 25746 13728
rect 26050 13676 26056 13728
rect 26108 13676 26114 13728
rect 26160 13716 26188 13824
rect 26786 13812 26792 13824
rect 26844 13812 26850 13864
rect 26896 13852 26924 13892
rect 26973 13889 26985 13923
rect 27019 13889 27031 13923
rect 28552 13920 28580 14028
rect 28721 14025 28733 14059
rect 28767 14056 28779 14059
rect 29454 14056 29460 14068
rect 28767 14028 29460 14056
rect 28767 14025 28779 14028
rect 28721 14019 28779 14025
rect 29454 14016 29460 14028
rect 29512 14016 29518 14068
rect 30561 14059 30619 14065
rect 30561 14025 30573 14059
rect 30607 14056 30619 14059
rect 31570 14056 31576 14068
rect 30607 14028 31576 14056
rect 30607 14025 30619 14028
rect 30561 14019 30619 14025
rect 31570 14016 31576 14028
rect 31628 14016 31634 14068
rect 33410 14016 33416 14068
rect 33468 14016 33474 14068
rect 33502 14016 33508 14068
rect 33560 14016 33566 14068
rect 34238 14016 34244 14068
rect 34296 14016 34302 14068
rect 34333 14059 34391 14065
rect 34333 14025 34345 14059
rect 34379 14056 34391 14059
rect 34422 14056 34428 14068
rect 34379 14028 34428 14056
rect 34379 14025 34391 14028
rect 34333 14019 34391 14025
rect 34422 14016 34428 14028
rect 34480 14016 34486 14068
rect 35434 14016 35440 14068
rect 35492 14016 35498 14068
rect 37001 14059 37059 14065
rect 37001 14025 37013 14059
rect 37047 14056 37059 14059
rect 37274 14056 37280 14068
rect 37047 14028 37280 14056
rect 37047 14025 37059 14028
rect 37001 14019 37059 14025
rect 37274 14016 37280 14028
rect 37332 14056 37338 14068
rect 37550 14056 37556 14068
rect 37332 14028 37556 14056
rect 37332 14016 37338 14028
rect 37550 14016 37556 14028
rect 37608 14016 37614 14068
rect 38212 14028 39160 14056
rect 28994 13988 29000 14000
rect 28828 13960 29000 13988
rect 28828 13929 28856 13960
rect 28994 13948 29000 13960
rect 29052 13948 29058 14000
rect 29546 13948 29552 14000
rect 29604 13948 29610 14000
rect 31018 13948 31024 14000
rect 31076 13988 31082 14000
rect 31113 13991 31171 13997
rect 31113 13988 31125 13991
rect 31076 13960 31125 13988
rect 31076 13948 31082 13960
rect 31113 13957 31125 13960
rect 31159 13957 31171 13991
rect 31113 13951 31171 13957
rect 31478 13948 31484 14000
rect 31536 13948 31542 14000
rect 34514 13948 34520 14000
rect 34572 13988 34578 14000
rect 35452 13988 35480 14016
rect 35529 13991 35587 13997
rect 35529 13988 35541 13991
rect 34572 13960 35020 13988
rect 35452 13960 35541 13988
rect 34572 13948 34578 13960
rect 28813 13923 28871 13929
rect 28813 13920 28825 13923
rect 26973 13883 27031 13889
rect 27982 13852 27988 13864
rect 26896 13824 27988 13852
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 28368 13852 28396 13906
rect 28552 13892 28825 13920
rect 28813 13889 28825 13892
rect 28859 13889 28871 13923
rect 28813 13883 28871 13889
rect 30745 13923 30803 13929
rect 30745 13889 30757 13923
rect 30791 13920 30803 13923
rect 31849 13923 31907 13929
rect 30791 13892 31754 13920
rect 30791 13889 30803 13892
rect 30745 13883 30803 13889
rect 29546 13852 29552 13864
rect 28368 13824 29552 13852
rect 29546 13812 29552 13824
rect 29604 13812 29610 13864
rect 31726 13852 31754 13892
rect 31849 13889 31861 13923
rect 31895 13920 31907 13923
rect 31938 13920 31944 13932
rect 31895 13892 31944 13920
rect 31895 13889 31907 13892
rect 31849 13883 31907 13889
rect 31938 13880 31944 13892
rect 31996 13880 32002 13932
rect 34054 13880 34060 13932
rect 34112 13920 34118 13932
rect 34992 13929 35020 13960
rect 35529 13957 35541 13960
rect 35575 13957 35587 13991
rect 35529 13951 35587 13957
rect 37918 13948 37924 14000
rect 37976 13988 37982 14000
rect 38212 13988 38240 14028
rect 39132 13988 39160 14028
rect 39298 14016 39304 14068
rect 39356 14016 39362 14068
rect 41417 14059 41475 14065
rect 40328 14028 41276 14056
rect 40328 13988 40356 14028
rect 41248 13988 41276 14028
rect 41417 14025 41429 14059
rect 41463 14056 41475 14059
rect 41506 14056 41512 14068
rect 41463 14028 41512 14056
rect 41463 14025 41475 14028
rect 41417 14019 41475 14025
rect 41506 14016 41512 14028
rect 41564 14056 41570 14068
rect 41564 14028 42104 14056
rect 41564 14016 41570 14028
rect 41966 13988 41972 14000
rect 37976 13960 38318 13988
rect 39132 13960 40434 13988
rect 41248 13960 41972 13988
rect 37976 13948 37982 13960
rect 41966 13948 41972 13960
rect 42024 13948 42030 14000
rect 34701 13923 34759 13929
rect 34701 13920 34713 13923
rect 34112 13892 34713 13920
rect 34112 13880 34118 13892
rect 34701 13889 34713 13892
rect 34747 13889 34759 13923
rect 34701 13883 34759 13889
rect 34977 13923 35035 13929
rect 34977 13889 34989 13923
rect 35023 13889 35035 13923
rect 34977 13883 35035 13889
rect 36630 13880 36636 13932
rect 36688 13880 36694 13932
rect 42076 13929 42104 14028
rect 42061 13923 42119 13929
rect 42061 13889 42073 13923
rect 42107 13889 42119 13923
rect 42061 13883 42119 13889
rect 32306 13852 32312 13864
rect 31726 13824 32312 13852
rect 32306 13812 32312 13824
rect 32364 13812 32370 13864
rect 32398 13812 32404 13864
rect 32456 13812 32462 13864
rect 33689 13855 33747 13861
rect 33689 13821 33701 13855
rect 33735 13821 33747 13855
rect 33689 13815 33747 13821
rect 34517 13855 34575 13861
rect 34517 13821 34529 13855
rect 34563 13821 34575 13855
rect 34517 13815 34575 13821
rect 32858 13744 32864 13796
rect 32916 13784 32922 13796
rect 33045 13787 33103 13793
rect 33045 13784 33057 13787
rect 32916 13756 33057 13784
rect 32916 13744 32922 13756
rect 33045 13753 33057 13756
rect 33091 13753 33103 13787
rect 33045 13747 33103 13753
rect 33134 13744 33140 13796
rect 33192 13784 33198 13796
rect 33704 13784 33732 13815
rect 34422 13784 34428 13796
rect 33192 13756 34428 13784
rect 33192 13744 33198 13756
rect 34422 13744 34428 13756
rect 34480 13784 34486 13796
rect 34532 13784 34560 13815
rect 34606 13812 34612 13864
rect 34664 13852 34670 13864
rect 34793 13855 34851 13861
rect 34793 13852 34805 13855
rect 34664 13824 34805 13852
rect 34664 13812 34670 13824
rect 34793 13821 34805 13824
rect 34839 13821 34851 13855
rect 34793 13815 34851 13821
rect 35250 13812 35256 13864
rect 35308 13852 35314 13864
rect 37458 13852 37464 13864
rect 35308 13824 37464 13852
rect 35308 13812 35314 13824
rect 37458 13812 37464 13824
rect 37516 13852 37522 13864
rect 37553 13855 37611 13861
rect 37553 13852 37565 13855
rect 37516 13824 37565 13852
rect 37516 13812 37522 13824
rect 37553 13821 37565 13824
rect 37599 13821 37611 13855
rect 37553 13815 37611 13821
rect 37826 13812 37832 13864
rect 37884 13812 37890 13864
rect 38378 13812 38384 13864
rect 38436 13852 38442 13864
rect 39669 13855 39727 13861
rect 39669 13852 39681 13855
rect 38436 13824 39681 13852
rect 38436 13812 38442 13824
rect 39669 13821 39681 13824
rect 39715 13821 39727 13855
rect 39669 13815 39727 13821
rect 39942 13812 39948 13864
rect 40000 13812 40006 13864
rect 40402 13812 40408 13864
rect 40460 13852 40466 13864
rect 41509 13855 41567 13861
rect 41509 13852 41521 13855
rect 40460 13824 41521 13852
rect 40460 13812 40466 13824
rect 41509 13821 41521 13824
rect 41555 13821 41567 13855
rect 41509 13815 41567 13821
rect 34480 13756 34560 13784
rect 34480 13744 34486 13756
rect 26234 13716 26240 13728
rect 26160 13688 26240 13716
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 26697 13719 26755 13725
rect 26697 13685 26709 13719
rect 26743 13716 26755 13719
rect 28810 13716 28816 13728
rect 26743 13688 28816 13716
rect 26743 13685 26755 13688
rect 26697 13679 26755 13685
rect 28810 13676 28816 13688
rect 28868 13676 28874 13728
rect 28902 13676 28908 13728
rect 28960 13716 28966 13728
rect 29070 13719 29128 13725
rect 29070 13716 29082 13719
rect 28960 13688 29082 13716
rect 28960 13676 28966 13688
rect 29070 13685 29082 13688
rect 29116 13685 29128 13719
rect 29070 13679 29128 13685
rect 32950 13676 32956 13728
rect 33008 13676 33014 13728
rect 33410 13676 33416 13728
rect 33468 13716 33474 13728
rect 33873 13719 33931 13725
rect 33873 13716 33885 13719
rect 33468 13688 33885 13716
rect 33468 13676 33474 13688
rect 33873 13685 33885 13688
rect 33919 13685 33931 13719
rect 33873 13679 33931 13685
rect 34882 13676 34888 13728
rect 34940 13676 34946 13728
rect 35161 13719 35219 13725
rect 35161 13685 35173 13719
rect 35207 13716 35219 13719
rect 35526 13716 35532 13728
rect 35207 13688 35532 13716
rect 35207 13685 35219 13688
rect 35161 13679 35219 13685
rect 35526 13676 35532 13688
rect 35584 13676 35590 13728
rect 1104 13626 42504 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 42504 13626
rect 1104 13552 42504 13574
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 5537 13515 5595 13521
rect 5537 13512 5549 13515
rect 4120 13484 5549 13512
rect 4120 13472 4126 13484
rect 5537 13481 5549 13484
rect 5583 13512 5595 13515
rect 5626 13512 5632 13524
rect 5583 13484 5632 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 5994 13512 6000 13524
rect 5767 13484 6000 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 7098 13472 7104 13524
rect 7156 13472 7162 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7208 13484 7849 13512
rect 6546 13444 6552 13456
rect 3252 13416 3832 13444
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 3252 13385 3280 13416
rect 3804 13385 3832 13416
rect 6104 13416 6552 13444
rect 3237 13379 3295 13385
rect 3237 13376 3249 13379
rect 2464 13348 3249 13376
rect 2464 13336 2470 13348
rect 3237 13345 3249 13348
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13376 3571 13379
rect 3789 13379 3847 13385
rect 3559 13348 3740 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 3605 13311 3663 13317
rect 3605 13277 3617 13311
rect 3651 13277 3663 13311
rect 3605 13271 3663 13277
rect 2682 13240 2688 13252
rect 2530 13212 2688 13240
rect 2682 13200 2688 13212
rect 2740 13200 2746 13252
rect 2958 13200 2964 13252
rect 3016 13200 3022 13252
rect 1489 13175 1547 13181
rect 1489 13141 1501 13175
rect 1535 13172 1547 13175
rect 2222 13172 2228 13184
rect 1535 13144 2228 13172
rect 1535 13141 1547 13144
rect 1489 13135 1547 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 3620 13172 3648 13271
rect 3712 13240 3740 13348
rect 3789 13345 3801 13379
rect 3835 13376 3847 13379
rect 6104 13376 6132 13416
rect 6546 13404 6552 13416
rect 6604 13444 6610 13456
rect 6604 13416 6868 13444
rect 6604 13404 6610 13416
rect 3835 13348 6132 13376
rect 6181 13379 6239 13385
rect 3835 13345 3847 13348
rect 3789 13339 3847 13345
rect 6181 13345 6193 13379
rect 6227 13376 6239 13379
rect 6730 13376 6736 13388
rect 6227 13348 6736 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 6840 13376 6868 13416
rect 7208 13385 7236 13484
rect 7837 13481 7849 13484
rect 7883 13512 7895 13515
rect 8110 13512 8116 13524
rect 7883 13484 8116 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9198 13515 9256 13521
rect 9198 13512 9210 13515
rect 8803 13484 9210 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9198 13481 9210 13484
rect 9244 13481 9256 13515
rect 9198 13475 9256 13481
rect 10686 13472 10692 13524
rect 10744 13472 10750 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17083 13515 17141 13521
rect 17083 13512 17095 13515
rect 16632 13484 17095 13512
rect 16632 13472 16638 13484
rect 17083 13481 17095 13484
rect 17129 13481 17141 13515
rect 19518 13512 19524 13524
rect 17083 13475 17141 13481
rect 18892 13484 19524 13512
rect 17678 13404 17684 13456
rect 17736 13444 17742 13456
rect 18892 13444 18920 13484
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 21634 13512 21640 13524
rect 19760 13484 21640 13512
rect 19760 13472 19766 13484
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 23017 13515 23075 13521
rect 23017 13481 23029 13515
rect 23063 13512 23075 13515
rect 23198 13512 23204 13524
rect 23063 13484 23204 13512
rect 23063 13481 23075 13484
rect 23017 13475 23075 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 26326 13472 26332 13524
rect 26384 13472 26390 13524
rect 26510 13472 26516 13524
rect 26568 13472 26574 13524
rect 28629 13515 28687 13521
rect 28629 13481 28641 13515
rect 28675 13512 28687 13515
rect 28902 13512 28908 13524
rect 28675 13484 28908 13512
rect 28675 13481 28687 13484
rect 28629 13475 28687 13481
rect 28902 13472 28908 13484
rect 28960 13472 28966 13524
rect 34701 13515 34759 13521
rect 34701 13512 34713 13515
rect 29012 13484 34713 13512
rect 17736 13416 18920 13444
rect 17736 13404 17742 13416
rect 7193 13379 7251 13385
rect 6840 13348 6960 13376
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 6822 13308 6828 13320
rect 6135 13280 6828 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 6822 13268 6828 13280
rect 6880 13268 6886 13320
rect 6932 13317 6960 13348
rect 7193 13345 7205 13379
rect 7239 13345 7251 13379
rect 7193 13339 7251 13345
rect 8481 13379 8539 13385
rect 8481 13345 8493 13379
rect 8527 13345 8539 13379
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 8481 13339 8539 13345
rect 8956 13348 11069 13376
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7282 13308 7288 13320
rect 6963 13280 7288 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7432 13280 8064 13308
rect 7432 13268 7438 13280
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 3712 13212 4077 13240
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4614 13200 4620 13252
rect 4672 13200 4678 13252
rect 6638 13200 6644 13252
rect 6696 13240 6702 13252
rect 8036 13249 8064 13280
rect 8386 13268 8392 13320
rect 8444 13268 8450 13320
rect 7101 13243 7159 13249
rect 7101 13240 7113 13243
rect 6696 13212 7113 13240
rect 6696 13200 6702 13212
rect 7101 13209 7113 13212
rect 7147 13240 7159 13243
rect 7805 13243 7863 13249
rect 7805 13240 7817 13243
rect 7147 13212 7817 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 7805 13209 7817 13212
rect 7851 13209 7863 13243
rect 7805 13203 7863 13209
rect 8021 13243 8079 13249
rect 8021 13209 8033 13243
rect 8067 13209 8079 13243
rect 8021 13203 8079 13209
rect 4338 13172 4344 13184
rect 3620 13144 4344 13172
rect 4338 13132 4344 13144
rect 4396 13132 4402 13184
rect 7558 13132 7564 13184
rect 7616 13132 7622 13184
rect 7650 13132 7656 13184
rect 7708 13132 7714 13184
rect 8496 13172 8524 13339
rect 8662 13268 8668 13320
rect 8720 13308 8726 13320
rect 8956 13317 8984 13348
rect 11057 13345 11069 13348
rect 11103 13345 11115 13379
rect 11057 13339 11115 13345
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 13964 13348 15301 13376
rect 13964 13336 13970 13348
rect 15289 13345 15301 13348
rect 15335 13376 15347 13379
rect 16666 13376 16672 13388
rect 15335 13348 16672 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 16666 13336 16672 13348
rect 16724 13376 16730 13388
rect 17862 13376 17868 13388
rect 16724 13348 17868 13376
rect 16724 13336 16730 13348
rect 17862 13336 17868 13348
rect 17920 13376 17926 13388
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 17920 13348 17969 13376
rect 17920 13336 17926 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8720 13280 8953 13308
rect 8720 13268 8726 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 13630 13268 13636 13320
rect 13688 13317 13694 13320
rect 13688 13308 13700 13317
rect 14093 13311 14151 13317
rect 13688 13280 13733 13308
rect 13688 13271 13700 13280
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 13688 13268 13694 13271
rect 10226 13200 10232 13252
rect 10284 13200 10290 13252
rect 11324 13243 11382 13249
rect 11324 13209 11336 13243
rect 11370 13240 11382 13243
rect 11514 13240 11520 13252
rect 11370 13212 11520 13240
rect 11370 13209 11382 13212
rect 11324 13203 11382 13209
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 13170 13200 13176 13252
rect 13228 13240 13234 13252
rect 14108 13240 14136 13271
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 15378 13268 15384 13320
rect 15436 13308 15442 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 15436 13280 15669 13308
rect 15436 13268 15442 13280
rect 15657 13277 15669 13280
rect 15703 13277 15715 13311
rect 15657 13271 15715 13277
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 17972 13308 18000 13339
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 18892 13385 18920 13416
rect 26234 13404 26240 13456
rect 26292 13404 26298 13456
rect 29012 13444 29040 13484
rect 34701 13481 34713 13484
rect 34747 13481 34759 13515
rect 34701 13475 34759 13481
rect 34974 13472 34980 13524
rect 35032 13472 35038 13524
rect 36170 13512 36176 13524
rect 35084 13484 36176 13512
rect 26344 13416 29040 13444
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 18564 13348 18705 13376
rect 18564 13336 18570 13348
rect 18693 13345 18705 13348
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 18877 13379 18935 13385
rect 18877 13345 18889 13379
rect 18923 13345 18935 13379
rect 18877 13339 18935 13345
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 21269 13379 21327 13385
rect 21269 13376 21281 13379
rect 20772 13348 21281 13376
rect 20772 13336 20778 13348
rect 21269 13345 21281 13348
rect 21315 13345 21327 13379
rect 21269 13339 21327 13345
rect 21542 13336 21548 13388
rect 21600 13336 21606 13388
rect 26050 13336 26056 13388
rect 26108 13336 26114 13388
rect 19426 13308 19432 13320
rect 16540 13280 17356 13308
rect 17972 13280 19432 13308
rect 16540 13268 16546 13280
rect 13228 13212 14136 13240
rect 16684 13226 16712 13280
rect 13228 13200 13234 13212
rect 17218 13200 17224 13252
rect 17276 13200 17282 13252
rect 17328 13240 17356 13280
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 21174 13268 21180 13320
rect 21232 13268 21238 13320
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 26344 13317 26372 13416
rect 29546 13404 29552 13456
rect 29604 13444 29610 13456
rect 30193 13447 30251 13453
rect 30193 13444 30205 13447
rect 29604 13416 30205 13444
rect 29604 13404 29610 13416
rect 30193 13413 30205 13416
rect 30239 13413 30251 13447
rect 30193 13407 30251 13413
rect 34330 13404 34336 13456
rect 34388 13404 34394 13456
rect 28350 13376 28356 13388
rect 26436 13348 28356 13376
rect 26436 13320 26464 13348
rect 28350 13336 28356 13348
rect 28408 13336 28414 13388
rect 28994 13336 29000 13388
rect 29052 13376 29058 13388
rect 30745 13379 30803 13385
rect 30745 13376 30757 13379
rect 29052 13348 30757 13376
rect 29052 13336 29058 13348
rect 30745 13345 30757 13348
rect 30791 13345 30803 13379
rect 30745 13339 30803 13345
rect 32398 13336 32404 13388
rect 32456 13376 32462 13388
rect 32493 13379 32551 13385
rect 32493 13376 32505 13379
rect 32456 13348 32505 13376
rect 32456 13336 32462 13348
rect 32493 13345 32505 13348
rect 32539 13345 32551 13379
rect 32493 13339 32551 13345
rect 32858 13336 32864 13388
rect 32916 13336 32922 13388
rect 35084 13385 35112 13484
rect 36170 13472 36176 13484
rect 36228 13472 36234 13524
rect 36906 13472 36912 13524
rect 36964 13512 36970 13524
rect 37185 13515 37243 13521
rect 37185 13512 37197 13515
rect 36964 13484 37197 13512
rect 36964 13472 36970 13484
rect 37185 13481 37197 13484
rect 37231 13481 37243 13515
rect 37185 13475 37243 13481
rect 37826 13472 37832 13524
rect 37884 13512 37890 13524
rect 38289 13515 38347 13521
rect 38289 13512 38301 13515
rect 37884 13484 38301 13512
rect 37884 13472 37890 13484
rect 38289 13481 38301 13484
rect 38335 13481 38347 13515
rect 38289 13475 38347 13481
rect 39853 13515 39911 13521
rect 39853 13481 39865 13515
rect 39899 13512 39911 13515
rect 39942 13512 39948 13524
rect 39899 13484 39948 13512
rect 39899 13481 39911 13484
rect 39853 13475 39911 13481
rect 39942 13472 39948 13484
rect 40000 13472 40006 13524
rect 38654 13404 38660 13456
rect 38712 13404 38718 13456
rect 40402 13444 40408 13456
rect 39408 13416 40408 13444
rect 35069 13379 35127 13385
rect 35069 13345 35081 13379
rect 35115 13345 35127 13379
rect 35069 13339 35127 13345
rect 35342 13336 35348 13388
rect 35400 13336 35406 13388
rect 35621 13379 35679 13385
rect 35621 13345 35633 13379
rect 35667 13376 35679 13379
rect 36262 13376 36268 13388
rect 35667 13348 36268 13376
rect 35667 13345 35679 13348
rect 35621 13339 35679 13345
rect 36262 13336 36268 13348
rect 36320 13336 36326 13388
rect 36630 13336 36636 13388
rect 36688 13376 36694 13388
rect 37918 13376 37924 13388
rect 36688 13348 37924 13376
rect 36688 13336 36694 13348
rect 25041 13311 25099 13317
rect 25041 13308 25053 13311
rect 24820 13280 25053 13308
rect 24820 13268 24826 13280
rect 25041 13277 25053 13280
rect 25087 13277 25099 13311
rect 25041 13271 25099 13277
rect 26329 13311 26387 13317
rect 26329 13277 26341 13311
rect 26375 13277 26387 13311
rect 26329 13271 26387 13277
rect 26418 13268 26424 13320
rect 26476 13268 26482 13320
rect 28166 13268 28172 13320
rect 28224 13268 28230 13320
rect 28810 13268 28816 13320
rect 28868 13268 28874 13320
rect 29089 13311 29147 13317
rect 29089 13277 29101 13311
rect 29135 13277 29147 13311
rect 29089 13271 29147 13277
rect 19610 13240 19616 13252
rect 17328 13212 19616 13240
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 19705 13243 19763 13249
rect 19705 13209 19717 13243
rect 19751 13240 19763 13243
rect 19978 13240 19984 13252
rect 19751 13212 19984 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 21192 13240 21220 13268
rect 23106 13240 23112 13252
rect 20088 13212 20194 13240
rect 21100 13212 21220 13240
rect 22770 13212 23112 13240
rect 10042 13172 10048 13184
rect 8496 13144 10048 13172
rect 10042 13132 10048 13144
rect 10100 13172 10106 13184
rect 11146 13172 11152 13184
rect 10100 13144 11152 13172
rect 10100 13132 10106 13144
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12434 13132 12440 13184
rect 12492 13132 12498 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12710 13172 12716 13184
rect 12575 13144 12716 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 14366 13132 14372 13184
rect 14424 13172 14430 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14424 13144 14473 13172
rect 14424 13132 14430 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 18230 13132 18236 13184
rect 18288 13132 18294 13184
rect 18598 13132 18604 13184
rect 18656 13132 18662 13184
rect 18966 13132 18972 13184
rect 19024 13172 19030 13184
rect 20088 13172 20116 13212
rect 21100 13172 21128 13212
rect 23106 13200 23112 13212
rect 23164 13200 23170 13252
rect 29104 13240 29132 13271
rect 29454 13268 29460 13320
rect 29512 13308 29518 13320
rect 29641 13311 29699 13317
rect 29641 13308 29653 13311
rect 29512 13280 29653 13308
rect 29512 13268 29518 13280
rect 29641 13277 29653 13280
rect 29687 13277 29699 13311
rect 29641 13271 29699 13277
rect 29822 13268 29828 13320
rect 29880 13308 29886 13320
rect 30009 13311 30067 13317
rect 30009 13308 30021 13311
rect 29880 13280 30021 13308
rect 29880 13268 29886 13280
rect 30009 13277 30021 13280
rect 30055 13277 30067 13311
rect 30009 13271 30067 13277
rect 32122 13268 32128 13320
rect 32180 13268 32186 13320
rect 32585 13311 32643 13317
rect 32585 13277 32597 13311
rect 32631 13277 32643 13311
rect 32585 13271 32643 13277
rect 30469 13243 30527 13249
rect 29104 13212 29776 13240
rect 19024 13144 21128 13172
rect 21177 13175 21235 13181
rect 19024 13132 19030 13144
rect 21177 13141 21189 13175
rect 21223 13172 21235 13175
rect 22462 13172 22468 13184
rect 21223 13144 22468 13172
rect 21223 13141 21235 13144
rect 21177 13135 21235 13141
rect 22462 13132 22468 13144
rect 22520 13132 22526 13184
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 24489 13175 24547 13181
rect 24489 13172 24501 13175
rect 24084 13144 24501 13172
rect 24084 13132 24090 13144
rect 24489 13141 24501 13144
rect 24535 13141 24547 13175
rect 24489 13135 24547 13141
rect 24670 13132 24676 13184
rect 24728 13172 24734 13184
rect 25958 13172 25964 13184
rect 24728 13144 25964 13172
rect 24728 13132 24734 13144
rect 25958 13132 25964 13144
rect 26016 13172 26022 13184
rect 26418 13172 26424 13184
rect 26016 13144 26424 13172
rect 26016 13132 26022 13144
rect 26418 13132 26424 13144
rect 26476 13132 26482 13184
rect 27430 13132 27436 13184
rect 27488 13172 27494 13184
rect 27617 13175 27675 13181
rect 27617 13172 27629 13175
rect 27488 13144 27629 13172
rect 27488 13132 27494 13144
rect 27617 13141 27629 13144
rect 27663 13141 27675 13175
rect 27617 13135 27675 13141
rect 28997 13175 29055 13181
rect 28997 13141 29009 13175
rect 29043 13172 29055 13175
rect 29638 13172 29644 13184
rect 29043 13144 29644 13172
rect 29043 13141 29055 13144
rect 28997 13135 29055 13141
rect 29638 13132 29644 13144
rect 29696 13132 29702 13184
rect 29748 13172 29776 13212
rect 30469 13209 30481 13243
rect 30515 13240 30527 13243
rect 30926 13240 30932 13252
rect 30515 13212 30932 13240
rect 30515 13209 30527 13212
rect 30469 13203 30527 13209
rect 30926 13200 30932 13212
rect 30984 13200 30990 13252
rect 31018 13200 31024 13252
rect 31076 13200 31082 13252
rect 32600 13240 32628 13271
rect 34146 13268 34152 13320
rect 34204 13308 34210 13320
rect 34885 13311 34943 13317
rect 34885 13308 34897 13311
rect 34204 13280 34897 13308
rect 34204 13268 34210 13280
rect 34885 13277 34897 13280
rect 34931 13277 34943 13311
rect 36740 13294 36768 13348
rect 37918 13336 37924 13348
rect 37976 13336 37982 13388
rect 38672 13376 38700 13404
rect 38841 13379 38899 13385
rect 38841 13376 38853 13379
rect 38672 13348 38853 13376
rect 38841 13345 38853 13348
rect 38887 13345 38899 13379
rect 38841 13339 38899 13345
rect 37737 13311 37795 13317
rect 37737 13308 37749 13311
rect 34885 13271 34943 13277
rect 37108 13280 37749 13308
rect 32858 13240 32864 13252
rect 32600 13212 32864 13240
rect 32858 13200 32864 13212
rect 32916 13200 32922 13252
rect 34422 13240 34428 13252
rect 34086 13212 34428 13240
rect 34422 13200 34428 13212
rect 34480 13200 34486 13252
rect 35161 13243 35219 13249
rect 35161 13209 35173 13243
rect 35207 13240 35219 13243
rect 35526 13240 35532 13252
rect 35207 13212 35532 13240
rect 35207 13209 35219 13212
rect 35161 13203 35219 13209
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 30558 13172 30564 13184
rect 29748 13144 30564 13172
rect 30558 13132 30564 13144
rect 30616 13172 30622 13184
rect 36262 13172 36268 13184
rect 30616 13144 36268 13172
rect 30616 13132 30622 13144
rect 36262 13132 36268 13144
rect 36320 13132 36326 13184
rect 36998 13132 37004 13184
rect 37056 13172 37062 13184
rect 37108 13181 37136 13280
rect 37737 13277 37749 13280
rect 37783 13277 37795 13311
rect 37737 13271 37795 13277
rect 38657 13311 38715 13317
rect 38657 13277 38669 13311
rect 38703 13308 38715 13311
rect 39298 13308 39304 13320
rect 38703 13280 39304 13308
rect 38703 13277 38715 13280
rect 38657 13271 38715 13277
rect 39298 13268 39304 13280
rect 39356 13268 39362 13320
rect 38749 13243 38807 13249
rect 38749 13209 38761 13243
rect 38795 13240 38807 13243
rect 39408 13240 39436 13416
rect 39482 13336 39488 13388
rect 39540 13376 39546 13388
rect 39758 13376 39764 13388
rect 39540 13348 39764 13376
rect 39540 13336 39546 13348
rect 39758 13336 39764 13348
rect 39816 13376 39822 13388
rect 39816 13348 40264 13376
rect 39816 13336 39822 13348
rect 40034 13268 40040 13320
rect 40092 13268 40098 13320
rect 40236 13317 40264 13348
rect 40328 13317 40356 13416
rect 40402 13404 40408 13416
rect 40460 13404 40466 13456
rect 41966 13404 41972 13456
rect 42024 13404 42030 13456
rect 40221 13311 40279 13317
rect 40221 13277 40233 13311
rect 40267 13277 40279 13311
rect 40328 13311 40397 13317
rect 40328 13280 40351 13311
rect 40221 13271 40279 13277
rect 40339 13277 40351 13280
rect 40385 13277 40397 13311
rect 40339 13271 40397 13277
rect 40494 13268 40500 13320
rect 40552 13268 40558 13320
rect 41782 13268 41788 13320
rect 41840 13268 41846 13320
rect 38795 13212 39436 13240
rect 40129 13243 40187 13249
rect 38795 13209 38807 13212
rect 38749 13203 38807 13209
rect 40129 13209 40141 13243
rect 40175 13209 40187 13243
rect 40129 13203 40187 13209
rect 37093 13175 37151 13181
rect 37093 13172 37105 13175
rect 37056 13144 37105 13172
rect 37056 13132 37062 13144
rect 37093 13141 37105 13144
rect 37139 13141 37151 13175
rect 40144 13172 40172 13203
rect 41690 13172 41696 13184
rect 40144 13144 41696 13172
rect 37093 13135 37151 13141
rect 41690 13132 41696 13144
rect 41748 13132 41754 13184
rect 1104 13082 42504 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 42504 13082
rect 1104 13008 42504 13030
rect 2498 12928 2504 12980
rect 2556 12928 2562 12980
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 2958 12968 2964 12980
rect 2823 12940 2964 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 3782 12971 3840 12977
rect 3782 12968 3794 12971
rect 3476 12940 3794 12968
rect 3476 12928 3482 12940
rect 3782 12937 3794 12940
rect 3828 12937 3840 12971
rect 3782 12931 3840 12937
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 6181 12971 6239 12977
rect 4672 12940 4844 12968
rect 4672 12928 4678 12940
rect 2222 12860 2228 12912
rect 2280 12900 2286 12912
rect 2317 12903 2375 12909
rect 2317 12900 2329 12903
rect 2280 12872 2329 12900
rect 2280 12860 2286 12872
rect 2317 12869 2329 12872
rect 2363 12869 2375 12903
rect 2317 12863 2375 12869
rect 3881 12903 3939 12909
rect 3881 12869 3893 12903
rect 3927 12900 3939 12903
rect 4062 12900 4068 12912
rect 3927 12872 4068 12900
rect 3927 12869 3939 12872
rect 3881 12863 3939 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 4706 12860 4712 12912
rect 4764 12860 4770 12912
rect 4816 12900 4844 12940
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6227 12940 6776 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6748 12909 6776 12940
rect 6822 12928 6828 12980
rect 6880 12928 6886 12980
rect 11146 12977 11152 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11133 12971 11152 12977
rect 11133 12937 11145 12971
rect 11133 12931 11152 12937
rect 6533 12903 6591 12909
rect 4816 12872 5198 12900
rect 6533 12869 6545 12903
rect 6579 12900 6591 12903
rect 6733 12903 6791 12909
rect 6579 12869 6592 12900
rect 6533 12863 6592 12869
rect 6733 12869 6745 12903
rect 6779 12900 6791 12903
rect 7374 12900 7380 12912
rect 6779 12872 7380 12900
rect 6779 12869 6791 12872
rect 6733 12863 6791 12869
rect 1670 12792 1676 12844
rect 1728 12792 1734 12844
rect 2590 12792 2596 12844
rect 2648 12792 2654 12844
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2685 12795 2743 12801
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3510 12832 3516 12844
rect 2915 12804 3516 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 2700 12764 2728 12795
rect 3510 12792 3516 12804
rect 3568 12832 3574 12844
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3568 12804 3617 12832
rect 3568 12792 3574 12804
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 3970 12832 3976 12844
rect 3743 12804 3976 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 6564 12832 6592 12863
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 8662 12900 8668 12912
rect 8128 12872 8668 12900
rect 6914 12832 6920 12844
rect 6564 12804 6920 12832
rect 2332 12736 2728 12764
rect 4433 12767 4491 12773
rect 2332 12705 2360 12736
rect 4433 12733 4445 12767
rect 4479 12733 4491 12767
rect 4433 12727 4491 12733
rect 2317 12699 2375 12705
rect 2317 12665 2329 12699
rect 2363 12665 2375 12699
rect 2317 12659 2375 12665
rect 1486 12588 1492 12640
rect 1544 12588 1550 12640
rect 4448 12628 4476 12727
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 6564 12764 6592 12804
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 8128 12841 8156 12872
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 9858 12900 9864 12912
rect 9614 12872 9864 12900
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 10594 12900 10600 12912
rect 9968 12872 10600 12900
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 7340 12804 8125 12832
rect 7340 12792 7346 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 9968 12841 9996 12872
rect 10594 12860 10600 12872
rect 10652 12900 10658 12912
rect 10980 12900 11008 12931
rect 11146 12928 11152 12931
rect 11204 12928 11210 12980
rect 13170 12928 13176 12980
rect 13228 12928 13234 12980
rect 13998 12928 14004 12980
rect 14056 12928 14062 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17037 12971 17095 12977
rect 17037 12968 17049 12971
rect 17000 12940 17049 12968
rect 17000 12928 17006 12940
rect 17037 12937 17049 12940
rect 17083 12937 17095 12971
rect 17037 12931 17095 12937
rect 17402 12928 17408 12980
rect 17460 12928 17466 12980
rect 17678 12928 17684 12980
rect 17736 12968 17742 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17736 12940 17785 12968
rect 17736 12928 17742 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 19242 12968 19248 12980
rect 18012 12940 19248 12968
rect 18012 12928 18018 12940
rect 19242 12928 19248 12940
rect 19300 12928 19306 12980
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20625 12971 20683 12977
rect 20625 12968 20637 12971
rect 20036 12940 20637 12968
rect 20036 12928 20042 12940
rect 20625 12937 20637 12940
rect 20671 12937 20683 12971
rect 20625 12931 20683 12937
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 22741 12971 22799 12977
rect 22741 12968 22753 12971
rect 21232 12940 22753 12968
rect 21232 12928 21238 12940
rect 22741 12937 22753 12940
rect 22787 12937 22799 12971
rect 22741 12931 22799 12937
rect 24026 12928 24032 12980
rect 24084 12928 24090 12980
rect 24118 12928 24124 12980
rect 24176 12928 24182 12980
rect 25038 12928 25044 12980
rect 25096 12928 25102 12980
rect 25148 12940 30696 12968
rect 10652 12872 11008 12900
rect 11333 12903 11391 12909
rect 10652 12860 10658 12872
rect 11333 12869 11345 12903
rect 11379 12869 11391 12903
rect 13906 12900 13912 12912
rect 11333 12863 11391 12869
rect 13832 12872 13912 12900
rect 9953 12835 10011 12841
rect 9953 12832 9965 12835
rect 9824 12804 9965 12832
rect 9824 12792 9830 12804
rect 9953 12801 9965 12804
rect 9999 12801 10011 12835
rect 9953 12795 10011 12801
rect 10134 12792 10140 12844
rect 10192 12792 10198 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11348 12832 11376 12863
rect 10744 12804 11376 12832
rect 11885 12835 11943 12841
rect 10744 12792 10750 12804
rect 11885 12801 11897 12835
rect 11931 12832 11943 12835
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 11931 12804 12265 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12986 12792 12992 12844
rect 13044 12792 13050 12844
rect 13832 12841 13860 12872
rect 13906 12860 13912 12872
rect 13964 12900 13970 12912
rect 14461 12903 14519 12909
rect 14461 12900 14473 12903
rect 13964 12872 14473 12900
rect 13964 12860 13970 12872
rect 14461 12869 14473 12872
rect 14507 12869 14519 12903
rect 18138 12900 18144 12912
rect 14461 12863 14519 12869
rect 17420 12872 18144 12900
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12832 13231 12835
rect 13265 12835 13323 12841
rect 13265 12832 13277 12835
rect 13219 12804 13277 12832
rect 13219 12801 13231 12804
rect 13173 12795 13231 12801
rect 13265 12801 13277 12804
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12801 13875 12835
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13817 12795 13875 12801
rect 13924 12804 14197 12832
rect 4764 12736 6592 12764
rect 4764 12724 4770 12736
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 7156 12736 7389 12764
rect 7156 12724 7162 12736
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 8435 12736 10057 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 10045 12733 10057 12736
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 6362 12656 6368 12708
rect 6420 12656 6426 12708
rect 10796 12696 10824 12727
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 11974 12724 11980 12776
rect 12032 12724 12038 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 9876 12668 10824 12696
rect 4706 12628 4712 12640
rect 4448 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 7098 12628 7104 12640
rect 6595 12600 7104 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 9876 12637 9904 12668
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9732 12600 9873 12628
rect 9732 12588 9738 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 10226 12588 10232 12640
rect 10284 12588 10290 12640
rect 10796 12628 10824 12668
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 10796 12600 11161 12628
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 12636 12628 12664 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 13924 12696 13952 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 17420 12841 17448 12872
rect 18138 12860 18144 12872
rect 18196 12900 18202 12912
rect 18782 12900 18788 12912
rect 18196 12872 18788 12900
rect 18196 12860 18202 12872
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 18966 12860 18972 12912
rect 19024 12860 19030 12912
rect 20162 12900 20168 12912
rect 20088 12872 20168 12900
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16816 12804 16865 12832
rect 16816 12792 16822 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17589 12835 17647 12841
rect 17589 12801 17601 12835
rect 17635 12832 17647 12835
rect 17954 12832 17960 12844
rect 17635 12804 17960 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 20088 12841 20116 12872
rect 20162 12860 20168 12872
rect 20220 12900 20226 12912
rect 21266 12900 21272 12912
rect 20220 12872 21272 12900
rect 20220 12860 20226 12872
rect 21266 12860 21272 12872
rect 21324 12860 21330 12912
rect 21634 12860 21640 12912
rect 21692 12900 21698 12912
rect 22649 12903 22707 12909
rect 22649 12900 22661 12903
rect 21692 12872 22661 12900
rect 21692 12860 21698 12872
rect 22649 12869 22661 12872
rect 22695 12869 22707 12903
rect 25148 12900 25176 12940
rect 26418 12900 26424 12912
rect 22649 12863 22707 12869
rect 23584 12872 25176 12900
rect 25700 12872 26424 12900
rect 23584 12844 23612 12872
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12801 20315 12835
rect 20257 12795 20315 12801
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 21039 12804 21833 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 14090 12724 14096 12776
rect 14148 12764 14154 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 14148 12736 14289 12764
rect 14148 12724 14154 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 14550 12724 14556 12776
rect 14608 12724 14614 12776
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12764 16727 12767
rect 17770 12764 17776 12776
rect 16715 12736 17776 12764
rect 16715 12733 16727 12736
rect 16669 12727 16727 12733
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 17920 12736 18245 12764
rect 17920 12724 17926 12736
rect 18233 12733 18245 12736
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 19242 12764 19248 12776
rect 18555 12736 19248 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 19242 12724 19248 12736
rect 19300 12724 19306 12776
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 20162 12764 20168 12776
rect 20027 12736 20168 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 20162 12724 20168 12736
rect 20220 12724 20226 12776
rect 12768 12668 13952 12696
rect 12768 12656 12774 12668
rect 20272 12640 20300 12795
rect 23566 12792 23572 12844
rect 23624 12792 23630 12844
rect 24949 12835 25007 12841
rect 24949 12801 24961 12835
rect 24995 12832 25007 12835
rect 25593 12835 25651 12841
rect 25593 12832 25605 12835
rect 24995 12804 25605 12832
rect 24995 12801 25007 12804
rect 24949 12795 25007 12801
rect 25593 12801 25605 12804
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 21266 12724 21272 12776
rect 21324 12724 21330 12776
rect 22462 12724 22468 12776
rect 22520 12764 22526 12776
rect 22738 12764 22744 12776
rect 22520 12736 22744 12764
rect 22520 12724 22526 12736
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 24305 12767 24363 12773
rect 24305 12764 24317 12767
rect 23400 12736 24317 12764
rect 23400 12705 23428 12736
rect 24305 12733 24317 12736
rect 24351 12764 24363 12767
rect 25225 12767 25283 12773
rect 25225 12764 25237 12767
rect 24351 12736 25237 12764
rect 24351 12733 24363 12736
rect 24305 12727 24363 12733
rect 25225 12733 25237 12736
rect 25271 12764 25283 12767
rect 25700 12764 25728 12872
rect 26418 12860 26424 12872
rect 26476 12900 26482 12912
rect 26786 12900 26792 12912
rect 26476 12872 26792 12900
rect 26476 12860 26482 12872
rect 26786 12860 26792 12872
rect 26844 12860 26850 12912
rect 27430 12860 27436 12912
rect 27488 12860 27494 12912
rect 28902 12900 28908 12912
rect 28658 12872 28908 12900
rect 28902 12860 28908 12872
rect 28960 12860 28966 12912
rect 30668 12900 30696 12940
rect 31018 12928 31024 12980
rect 31076 12968 31082 12980
rect 32125 12971 32183 12977
rect 32125 12968 32137 12971
rect 31076 12940 32137 12968
rect 31076 12928 31082 12940
rect 32125 12937 32137 12940
rect 32171 12937 32183 12971
rect 32125 12931 32183 12937
rect 32493 12971 32551 12977
rect 32493 12937 32505 12971
rect 32539 12968 32551 12971
rect 32950 12968 32956 12980
rect 32539 12940 32956 12968
rect 32539 12937 32551 12940
rect 32493 12931 32551 12937
rect 32950 12928 32956 12940
rect 33008 12928 33014 12980
rect 33060 12940 34652 12968
rect 31938 12900 31944 12912
rect 30668 12872 31944 12900
rect 31938 12860 31944 12872
rect 31996 12900 32002 12912
rect 33060 12900 33088 12940
rect 31996 12872 33088 12900
rect 33321 12903 33379 12909
rect 31996 12860 32002 12872
rect 33321 12869 33333 12903
rect 33367 12900 33379 12903
rect 33410 12900 33416 12912
rect 33367 12872 33416 12900
rect 33367 12869 33379 12872
rect 33321 12863 33379 12869
rect 33410 12860 33416 12872
rect 33468 12860 33474 12912
rect 25774 12792 25780 12844
rect 25832 12832 25838 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 25832 12804 27169 12832
rect 25832 12792 25838 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 29457 12835 29515 12841
rect 29457 12801 29469 12835
rect 29503 12832 29515 12835
rect 29822 12832 29828 12844
rect 29503 12804 29828 12832
rect 29503 12801 29515 12804
rect 29457 12795 29515 12801
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 30558 12792 30564 12844
rect 30616 12841 30622 12844
rect 30616 12832 30625 12841
rect 30745 12835 30803 12841
rect 30616 12804 30661 12832
rect 30616 12795 30625 12804
rect 30745 12801 30757 12835
rect 30791 12832 30803 12835
rect 31018 12832 31024 12844
rect 30791 12804 31024 12832
rect 30791 12801 30803 12804
rect 30745 12795 30803 12801
rect 30616 12792 30622 12795
rect 25271 12736 25728 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 26234 12724 26240 12776
rect 26292 12724 26298 12776
rect 29641 12767 29699 12773
rect 29641 12764 29653 12767
rect 26344 12736 29653 12764
rect 23385 12699 23443 12705
rect 23385 12665 23397 12699
rect 23431 12665 23443 12699
rect 26344 12696 26372 12736
rect 29641 12733 29653 12736
rect 29687 12733 29699 12767
rect 29641 12727 29699 12733
rect 29917 12767 29975 12773
rect 29917 12733 29929 12767
rect 29963 12764 29975 12767
rect 30760 12764 30788 12795
rect 31018 12792 31024 12804
rect 31076 12792 31082 12844
rect 32490 12792 32496 12844
rect 32548 12832 32554 12844
rect 32585 12835 32643 12841
rect 32585 12832 32597 12835
rect 32548 12804 32597 12832
rect 32548 12792 32554 12804
rect 32585 12801 32597 12804
rect 32631 12801 32643 12835
rect 32950 12832 32956 12844
rect 32585 12795 32643 12801
rect 32692 12804 32956 12832
rect 29963 12736 30788 12764
rect 29963 12733 29975 12736
rect 29917 12727 29975 12733
rect 30834 12724 30840 12776
rect 30892 12724 30898 12776
rect 31478 12724 31484 12776
rect 31536 12764 31542 12776
rect 32692 12773 32720 12804
rect 32950 12792 32956 12804
rect 33008 12792 33014 12844
rect 34422 12792 34428 12844
rect 34480 12792 34486 12844
rect 34624 12832 34652 12940
rect 35158 12928 35164 12980
rect 35216 12928 35222 12980
rect 35345 12971 35403 12977
rect 35345 12937 35357 12971
rect 35391 12968 35403 12971
rect 37182 12968 37188 12980
rect 35391 12940 37188 12968
rect 35391 12937 35403 12940
rect 35345 12931 35403 12937
rect 37182 12928 37188 12940
rect 37240 12928 37246 12980
rect 35713 12903 35771 12909
rect 35713 12869 35725 12903
rect 35759 12900 35771 12903
rect 36078 12900 36084 12912
rect 35759 12872 36084 12900
rect 35759 12869 35771 12872
rect 35713 12863 35771 12869
rect 36078 12860 36084 12872
rect 36136 12860 36142 12912
rect 36538 12860 36544 12912
rect 36596 12860 36602 12912
rect 36998 12860 37004 12912
rect 37056 12900 37062 12912
rect 37056 12872 37872 12900
rect 37056 12860 37062 12872
rect 34977 12835 35035 12841
rect 34977 12832 34989 12835
rect 34624 12804 34989 12832
rect 34977 12801 34989 12804
rect 35023 12801 35035 12835
rect 34977 12795 35035 12801
rect 35526 12792 35532 12844
rect 35584 12792 35590 12844
rect 35805 12835 35863 12841
rect 35805 12801 35817 12835
rect 35851 12832 35863 12835
rect 35894 12832 35900 12844
rect 35851 12804 35900 12832
rect 35851 12801 35863 12804
rect 35805 12795 35863 12801
rect 35894 12792 35900 12804
rect 35952 12832 35958 12844
rect 36556 12832 36584 12860
rect 35952 12804 36584 12832
rect 37461 12835 37519 12841
rect 35952 12792 35958 12804
rect 37461 12801 37473 12835
rect 37507 12801 37519 12835
rect 37461 12795 37519 12801
rect 32677 12767 32735 12773
rect 32677 12764 32689 12767
rect 31536 12736 32689 12764
rect 31536 12724 31542 12736
rect 32677 12733 32689 12736
rect 32723 12733 32735 12767
rect 32677 12727 32735 12733
rect 32858 12724 32864 12776
rect 32916 12764 32922 12776
rect 33045 12767 33103 12773
rect 33045 12764 33057 12767
rect 32916 12736 33057 12764
rect 32916 12724 32922 12736
rect 33045 12733 33057 12736
rect 33091 12733 33103 12767
rect 33045 12727 33103 12733
rect 33962 12724 33968 12776
rect 34020 12764 34026 12776
rect 34440 12764 34468 12792
rect 34020 12736 34919 12764
rect 34020 12724 34026 12736
rect 23385 12659 23443 12665
rect 23492 12668 26372 12696
rect 14185 12631 14243 12637
rect 14185 12628 14197 12631
rect 12636 12600 14197 12628
rect 11149 12591 11207 12597
rect 14185 12597 14197 12600
rect 14231 12597 14243 12631
rect 14185 12591 14243 12597
rect 15194 12588 15200 12640
rect 15252 12588 15258 12640
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 19702 12628 19708 12640
rect 18104 12600 19708 12628
rect 18104 12588 18110 12600
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 19886 12588 19892 12640
rect 19944 12628 19950 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 19944 12600 20085 12628
rect 19944 12588 19950 12600
rect 20073 12597 20085 12600
rect 20119 12597 20131 12631
rect 20073 12591 20131 12597
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 20530 12588 20536 12640
rect 20588 12628 20594 12640
rect 23492 12628 23520 12668
rect 34698 12656 34704 12708
rect 34756 12696 34762 12708
rect 34793 12699 34851 12705
rect 34793 12696 34805 12699
rect 34756 12668 34805 12696
rect 34756 12656 34762 12668
rect 34793 12665 34805 12668
rect 34839 12665 34851 12699
rect 34891 12696 34919 12736
rect 36538 12724 36544 12776
rect 36596 12724 36602 12776
rect 37366 12724 37372 12776
rect 37424 12724 37430 12776
rect 37476 12764 37504 12795
rect 37550 12792 37556 12844
rect 37608 12792 37614 12844
rect 37844 12841 37872 12872
rect 37918 12860 37924 12912
rect 37976 12860 37982 12912
rect 38289 12903 38347 12909
rect 38289 12869 38301 12903
rect 38335 12900 38347 12903
rect 38654 12900 38660 12912
rect 38335 12872 38660 12900
rect 38335 12869 38347 12872
rect 38289 12863 38347 12869
rect 38654 12860 38660 12872
rect 38712 12900 38718 12912
rect 41782 12900 41788 12912
rect 38712 12872 41788 12900
rect 38712 12860 38718 12872
rect 41782 12860 41788 12872
rect 41840 12860 41846 12912
rect 37829 12835 37887 12841
rect 37829 12801 37841 12835
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 38473 12835 38531 12841
rect 38473 12801 38485 12835
rect 38519 12832 38531 12835
rect 38838 12832 38844 12844
rect 38519 12804 38844 12832
rect 38519 12801 38531 12804
rect 38473 12795 38531 12801
rect 38838 12792 38844 12804
rect 38896 12792 38902 12844
rect 37642 12764 37648 12776
rect 37476 12736 37648 12764
rect 37642 12724 37648 12736
rect 37700 12724 37706 12776
rect 36630 12696 36636 12708
rect 34891 12668 36636 12696
rect 34793 12659 34851 12665
rect 36630 12656 36636 12668
rect 36688 12656 36694 12708
rect 37384 12696 37412 12724
rect 37918 12696 37924 12708
rect 37384 12668 37924 12696
rect 37918 12656 37924 12668
rect 37976 12696 37982 12708
rect 38657 12699 38715 12705
rect 38657 12696 38669 12699
rect 37976 12668 38669 12696
rect 37976 12656 37982 12668
rect 38657 12665 38669 12668
rect 38703 12696 38715 12699
rect 40494 12696 40500 12708
rect 38703 12668 40500 12696
rect 38703 12665 38715 12668
rect 38657 12659 38715 12665
rect 40494 12656 40500 12668
rect 40552 12656 40558 12708
rect 20588 12600 23520 12628
rect 20588 12588 20594 12600
rect 23566 12588 23572 12640
rect 23624 12628 23630 12640
rect 23661 12631 23719 12637
rect 23661 12628 23673 12631
rect 23624 12600 23673 12628
rect 23624 12588 23630 12600
rect 23661 12597 23673 12600
rect 23707 12597 23719 12631
rect 23661 12591 23719 12597
rect 24581 12631 24639 12637
rect 24581 12597 24593 12631
rect 24627 12628 24639 12631
rect 24670 12628 24676 12640
rect 24627 12600 24676 12628
rect 24627 12597 24639 12600
rect 24581 12591 24639 12597
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 28810 12588 28816 12640
rect 28868 12628 28874 12640
rect 28905 12631 28963 12637
rect 28905 12628 28917 12631
rect 28868 12600 28917 12628
rect 28868 12588 28874 12600
rect 28905 12597 28917 12600
rect 28951 12597 28963 12631
rect 28905 12591 28963 12597
rect 29178 12588 29184 12640
rect 29236 12628 29242 12640
rect 29365 12631 29423 12637
rect 29365 12628 29377 12631
rect 29236 12600 29377 12628
rect 29236 12588 29242 12600
rect 29365 12597 29377 12600
rect 29411 12628 29423 12631
rect 29638 12628 29644 12640
rect 29411 12600 29644 12628
rect 29411 12597 29423 12600
rect 29365 12591 29423 12597
rect 29638 12588 29644 12600
rect 29696 12588 29702 12640
rect 30558 12588 30564 12640
rect 30616 12588 30622 12640
rect 31481 12631 31539 12637
rect 31481 12597 31493 12631
rect 31527 12628 31539 12631
rect 31754 12628 31760 12640
rect 31527 12600 31760 12628
rect 31527 12597 31539 12600
rect 31481 12591 31539 12597
rect 31754 12588 31760 12600
rect 31812 12588 31818 12640
rect 37277 12631 37335 12637
rect 37277 12597 37289 12631
rect 37323 12628 37335 12631
rect 37366 12628 37372 12640
rect 37323 12600 37372 12628
rect 37323 12597 37335 12600
rect 37277 12591 37335 12597
rect 37366 12588 37372 12600
rect 37424 12588 37430 12640
rect 37737 12631 37795 12637
rect 37737 12597 37749 12631
rect 37783 12628 37795 12631
rect 37826 12628 37832 12640
rect 37783 12600 37832 12628
rect 37783 12597 37795 12600
rect 37737 12591 37795 12597
rect 37826 12588 37832 12600
rect 37884 12588 37890 12640
rect 1104 12538 42504 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 42504 12538
rect 1104 12464 42504 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1765 12427 1823 12433
rect 1765 12424 1777 12427
rect 1728 12396 1777 12424
rect 1728 12384 1734 12396
rect 1765 12393 1777 12396
rect 1811 12393 1823 12427
rect 1765 12387 1823 12393
rect 1946 12384 1952 12436
rect 2004 12384 2010 12436
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 4614 12424 4620 12436
rect 4571 12396 4620 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 4709 12427 4767 12433
rect 4709 12393 4721 12427
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 4724 12356 4752 12387
rect 7098 12384 7104 12436
rect 7156 12424 7162 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7156 12396 7481 12424
rect 7156 12384 7162 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 7469 12387 7527 12393
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10192 12396 10241 12424
rect 10192 12384 10198 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 11701 12427 11759 12433
rect 11701 12424 11713 12427
rect 11572 12396 11713 12424
rect 11572 12384 11578 12396
rect 11701 12393 11713 12396
rect 11747 12424 11759 12427
rect 17218 12424 17224 12436
rect 11747 12396 17224 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 17218 12384 17224 12396
rect 17276 12424 17282 12436
rect 20714 12424 20720 12436
rect 17276 12396 20720 12424
rect 17276 12384 17282 12396
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 24670 12433 24676 12436
rect 24660 12427 24676 12433
rect 21284 12396 21588 12424
rect 14090 12356 14096 12368
rect 2832 12328 4752 12356
rect 13924 12328 14096 12356
rect 2832 12316 2838 12328
rect 2222 12288 2228 12300
rect 1964 12260 2228 12288
rect 1964 12229 1992 12260
rect 2222 12248 2228 12260
rect 2280 12288 2286 12300
rect 3786 12288 3792 12300
rect 2280 12260 3792 12288
rect 2280 12248 2286 12260
rect 3786 12248 3792 12260
rect 3844 12288 3850 12300
rect 4338 12288 4344 12300
rect 3844 12260 4344 12288
rect 3844 12248 3850 12260
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 4672 12260 5733 12288
rect 4672 12248 4678 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 5994 12248 6000 12300
rect 6052 12248 6058 12300
rect 10042 12288 10048 12300
rect 9968 12260 10048 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2133 12223 2191 12229
rect 2133 12220 2145 12223
rect 2096 12192 2145 12220
rect 2096 12180 2102 12192
rect 2133 12189 2145 12192
rect 2179 12220 2191 12223
rect 5534 12220 5540 12232
rect 2179 12192 5540 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 9766 12220 9772 12232
rect 9539 12192 9772 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 9968 12229 9996 12260
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10594 12248 10600 12300
rect 10652 12248 10658 12300
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 11882 12288 11888 12300
rect 10919 12260 11888 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 13924 12297 13952 12328
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 21284 12356 21312 12396
rect 18524 12328 21312 12356
rect 21560 12356 21588 12396
rect 24660 12393 24672 12427
rect 24660 12387 24676 12393
rect 24670 12384 24676 12387
rect 24728 12384 24734 12436
rect 26145 12427 26203 12433
rect 26145 12393 26157 12427
rect 26191 12424 26203 12427
rect 26234 12424 26240 12436
rect 26191 12396 26240 12424
rect 26191 12393 26203 12396
rect 26145 12387 26203 12393
rect 26234 12384 26240 12396
rect 26292 12384 26298 12436
rect 27709 12427 27767 12433
rect 27709 12393 27721 12427
rect 27755 12424 27767 12427
rect 28166 12424 28172 12436
rect 27755 12396 28172 12424
rect 27755 12393 27767 12396
rect 27709 12387 27767 12393
rect 28166 12384 28172 12396
rect 28224 12384 28230 12436
rect 31297 12427 31355 12433
rect 31297 12393 31309 12427
rect 31343 12424 31355 12427
rect 31846 12424 31852 12436
rect 31343 12396 31852 12424
rect 31343 12393 31355 12396
rect 31297 12387 31355 12393
rect 31846 12384 31852 12396
rect 31904 12384 31910 12436
rect 35434 12384 35440 12436
rect 35492 12424 35498 12436
rect 35894 12424 35900 12436
rect 35492 12396 35900 12424
rect 35492 12384 35498 12396
rect 35894 12384 35900 12396
rect 35952 12384 35958 12436
rect 23290 12356 23296 12368
rect 21560 12328 23296 12356
rect 13909 12291 13967 12297
rect 13909 12257 13921 12291
rect 13955 12257 13967 12291
rect 18524 12288 18552 12328
rect 23290 12316 23296 12328
rect 23348 12316 23354 12368
rect 26418 12316 26424 12368
rect 26476 12356 26482 12368
rect 26476 12328 26832 12356
rect 26476 12316 26482 12328
rect 13909 12251 13967 12257
rect 15396 12260 18552 12288
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12220 13047 12223
rect 15396 12220 15424 12260
rect 19242 12248 19248 12300
rect 19300 12248 19306 12300
rect 19794 12248 19800 12300
rect 19852 12248 19858 12300
rect 20530 12248 20536 12300
rect 20588 12248 20594 12300
rect 22738 12288 22744 12300
rect 20640 12260 21404 12288
rect 13035 12192 15424 12220
rect 15473 12223 15531 12229
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 16850 12220 16856 12232
rect 15519 12192 16856 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 16850 12180 16856 12192
rect 16908 12220 16914 12232
rect 17221 12223 17279 12229
rect 17221 12220 17233 12223
rect 16908 12192 17233 12220
rect 16908 12180 16914 12192
rect 17221 12189 17233 12192
rect 17267 12189 17279 12223
rect 17221 12183 17279 12189
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20640 12229 20668 12260
rect 21376 12232 21404 12260
rect 21928 12260 22744 12288
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20496 12192 20637 12220
rect 20496 12180 20502 12192
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21358 12180 21364 12232
rect 21416 12180 21422 12232
rect 21928 12229 21956 12260
rect 22738 12248 22744 12260
rect 22796 12248 22802 12300
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12288 23443 12291
rect 24762 12288 24768 12300
rect 23431 12260 24768 12288
rect 23431 12257 23443 12260
rect 23385 12251 23443 12257
rect 24762 12248 24768 12260
rect 24820 12248 24826 12300
rect 25866 12248 25872 12300
rect 25924 12248 25930 12300
rect 26694 12248 26700 12300
rect 26752 12248 26758 12300
rect 26804 12297 26832 12328
rect 26878 12316 26884 12368
rect 26936 12356 26942 12368
rect 29178 12356 29184 12368
rect 26936 12328 29184 12356
rect 26936 12316 26942 12328
rect 29178 12316 29184 12328
rect 29236 12316 29242 12368
rect 38838 12316 38844 12368
rect 38896 12356 38902 12368
rect 39117 12359 39175 12365
rect 39117 12356 39129 12359
rect 38896 12328 39129 12356
rect 38896 12316 38902 12328
rect 39117 12325 39129 12328
rect 39163 12325 39175 12359
rect 39117 12319 39175 12325
rect 26789 12291 26847 12297
rect 26789 12257 26801 12291
rect 26835 12257 26847 12291
rect 28261 12291 28319 12297
rect 28261 12288 28273 12291
rect 26789 12251 26847 12257
rect 26896 12260 28273 12288
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12189 21511 12223
rect 21453 12183 21511 12189
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 2409 12155 2467 12161
rect 2409 12121 2421 12155
rect 2455 12152 2467 12155
rect 2498 12152 2504 12164
rect 2455 12124 2504 12152
rect 2455 12121 2467 12124
rect 2409 12115 2467 12121
rect 2498 12112 2504 12124
rect 2556 12112 2562 12164
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 4893 12155 4951 12161
rect 4893 12152 4905 12155
rect 4856 12124 4905 12152
rect 4856 12112 4862 12124
rect 4893 12121 4905 12124
rect 4939 12152 4951 12155
rect 5258 12152 5264 12164
rect 4939 12124 5264 12152
rect 4939 12121 4951 12124
rect 4893 12115 4951 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 7282 12152 7288 12164
rect 7222 12124 7288 12152
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 9861 12155 9919 12161
rect 9861 12121 9873 12155
rect 9907 12121 9919 12155
rect 9861 12115 9919 12121
rect 4154 12044 4160 12096
rect 4212 12084 4218 12096
rect 4693 12087 4751 12093
rect 4693 12084 4705 12087
rect 4212 12056 4705 12084
rect 4212 12044 4218 12056
rect 4693 12053 4705 12056
rect 4739 12084 4751 12087
rect 5350 12084 5356 12096
rect 4739 12056 5356 12084
rect 4739 12053 4751 12056
rect 4693 12047 4751 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5718 12044 5724 12096
rect 5776 12084 5782 12096
rect 9214 12084 9220 12096
rect 5776 12056 9220 12084
rect 5776 12044 5782 12056
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9306 12044 9312 12096
rect 9364 12044 9370 12096
rect 9582 12044 9588 12096
rect 9640 12044 9646 12096
rect 9674 12044 9680 12096
rect 9732 12044 9738 12096
rect 9876 12084 9904 12115
rect 15194 12112 15200 12164
rect 15252 12161 15258 12164
rect 15252 12115 15264 12161
rect 17497 12155 17555 12161
rect 17497 12121 17509 12155
rect 17543 12121 17555 12155
rect 17497 12115 17555 12121
rect 15252 12112 15258 12115
rect 9950 12084 9956 12096
rect 9876 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12084 10014 12096
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 10008 12056 10057 12084
rect 10008 12044 10014 12056
rect 10045 12053 10057 12056
rect 10091 12084 10103 12087
rect 10686 12084 10692 12096
rect 10091 12056 10692 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 13265 12087 13323 12093
rect 13265 12053 13277 12087
rect 13311 12084 13323 12087
rect 13538 12084 13544 12096
rect 13311 12056 13544 12084
rect 13311 12053 13323 12056
rect 13265 12047 13323 12053
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 17512 12084 17540 12115
rect 17954 12112 17960 12164
rect 18012 12112 18018 12164
rect 19981 12155 20039 12161
rect 19981 12121 19993 12155
rect 20027 12121 20039 12155
rect 19981 12115 20039 12121
rect 20165 12155 20223 12161
rect 20165 12121 20177 12155
rect 20211 12152 20223 12155
rect 20530 12152 20536 12164
rect 20211 12124 20536 12152
rect 20211 12121 20223 12124
rect 20165 12115 20223 12121
rect 18230 12084 18236 12096
rect 17512 12056 18236 12084
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 18969 12087 19027 12093
rect 18969 12053 18981 12087
rect 19015 12084 19027 12087
rect 19518 12084 19524 12096
rect 19015 12056 19524 12084
rect 19015 12053 19027 12056
rect 18969 12047 19027 12053
rect 19518 12044 19524 12056
rect 19576 12084 19582 12096
rect 19996 12084 20024 12115
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 21266 12112 21272 12164
rect 21324 12112 21330 12164
rect 21468 12152 21496 12183
rect 22094 12180 22100 12232
rect 22152 12180 22158 12232
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12220 22247 12223
rect 22278 12220 22284 12232
rect 22235 12192 22284 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 23109 12223 23167 12229
rect 23109 12220 23121 12223
rect 22520 12192 23121 12220
rect 22520 12180 22526 12192
rect 23109 12189 23121 12192
rect 23155 12189 23167 12223
rect 23109 12183 23167 12189
rect 23293 12223 23351 12229
rect 23293 12189 23305 12223
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23014 12152 23020 12164
rect 21468 12124 23020 12152
rect 23014 12112 23020 12124
rect 23072 12112 23078 12164
rect 19576 12056 20024 12084
rect 19576 12044 19582 12056
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 20349 12087 20407 12093
rect 20349 12084 20361 12087
rect 20128 12056 20361 12084
rect 20128 12044 20134 12056
rect 20349 12053 20361 12056
rect 20395 12053 20407 12087
rect 20349 12047 20407 12053
rect 21634 12044 21640 12096
rect 21692 12044 21698 12096
rect 21729 12087 21787 12093
rect 21729 12053 21741 12087
rect 21775 12084 21787 12087
rect 21818 12084 21824 12096
rect 21775 12056 21824 12084
rect 21775 12053 21787 12056
rect 21729 12047 21787 12053
rect 21818 12044 21824 12056
rect 21876 12044 21882 12096
rect 23308 12084 23336 12183
rect 23474 12180 23480 12232
rect 23532 12180 23538 12232
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12189 24455 12223
rect 25884 12220 25912 12248
rect 26896 12220 26924 12260
rect 28261 12257 28273 12260
rect 28307 12257 28319 12291
rect 28261 12251 28319 12257
rect 28994 12248 29000 12300
rect 29052 12288 29058 12300
rect 29549 12291 29607 12297
rect 29549 12288 29561 12291
rect 29052 12260 29561 12288
rect 29052 12248 29058 12260
rect 29549 12257 29561 12260
rect 29595 12257 29607 12291
rect 29549 12251 29607 12257
rect 29825 12291 29883 12297
rect 29825 12257 29837 12291
rect 29871 12288 29883 12291
rect 30558 12288 30564 12300
rect 29871 12260 30564 12288
rect 29871 12257 29883 12260
rect 29825 12251 29883 12257
rect 30558 12248 30564 12260
rect 30616 12248 30622 12300
rect 31478 12248 31484 12300
rect 31536 12288 31542 12300
rect 31941 12291 31999 12297
rect 31941 12288 31953 12291
rect 31536 12260 31953 12288
rect 31536 12248 31542 12260
rect 31941 12257 31953 12260
rect 31987 12257 31999 12291
rect 31941 12251 31999 12257
rect 37090 12248 37096 12300
rect 37148 12288 37154 12300
rect 37148 12260 39712 12288
rect 37148 12248 37154 12260
rect 25884 12192 26924 12220
rect 24397 12183 24455 12189
rect 23382 12112 23388 12164
rect 23440 12152 23446 12164
rect 23676 12152 23704 12183
rect 23440 12124 23704 12152
rect 23440 12112 23446 12124
rect 23658 12084 23664 12096
rect 23308 12056 23664 12084
rect 23658 12044 23664 12056
rect 23716 12044 23722 12096
rect 23845 12087 23903 12093
rect 23845 12053 23857 12087
rect 23891 12084 23903 12087
rect 24302 12084 24308 12096
rect 23891 12056 24308 12084
rect 23891 12053 23903 12056
rect 23845 12047 23903 12053
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 24412 12084 24440 12183
rect 27706 12180 27712 12232
rect 27764 12220 27770 12232
rect 28169 12223 28227 12229
rect 28169 12220 28181 12223
rect 27764 12192 28181 12220
rect 27764 12180 27770 12192
rect 28169 12189 28181 12192
rect 28215 12189 28227 12223
rect 28169 12183 28227 12189
rect 28810 12180 28816 12232
rect 28868 12220 28874 12232
rect 29089 12223 29147 12229
rect 29089 12220 29101 12223
rect 28868 12192 29101 12220
rect 28868 12180 28874 12192
rect 29089 12189 29101 12192
rect 29135 12189 29147 12223
rect 29089 12183 29147 12189
rect 31754 12180 31760 12232
rect 31812 12180 31818 12232
rect 31849 12223 31907 12229
rect 31849 12189 31861 12223
rect 31895 12220 31907 12223
rect 32030 12220 32036 12232
rect 31895 12192 32036 12220
rect 31895 12189 31907 12192
rect 31849 12183 31907 12189
rect 32030 12180 32036 12192
rect 32088 12180 32094 12232
rect 34698 12180 34704 12232
rect 34756 12220 34762 12232
rect 35437 12223 35495 12229
rect 35437 12220 35449 12223
rect 34756 12192 35449 12220
rect 34756 12180 34762 12192
rect 35437 12189 35449 12192
rect 35483 12189 35495 12223
rect 35437 12183 35495 12189
rect 35989 12223 36047 12229
rect 35989 12189 36001 12223
rect 36035 12220 36047 12223
rect 36538 12220 36544 12232
rect 36035 12192 36544 12220
rect 36035 12189 36047 12192
rect 35989 12183 36047 12189
rect 24578 12112 24584 12164
rect 24636 12152 24642 12164
rect 28077 12155 28135 12161
rect 24636 12124 25162 12152
rect 24636 12112 24642 12124
rect 28077 12121 28089 12155
rect 28123 12152 28135 12155
rect 28537 12155 28595 12161
rect 28537 12152 28549 12155
rect 28123 12124 28549 12152
rect 28123 12121 28135 12124
rect 28077 12115 28135 12121
rect 28537 12121 28549 12124
rect 28583 12121 28595 12155
rect 28537 12115 28595 12121
rect 29914 12112 29920 12164
rect 29972 12152 29978 12164
rect 29972 12124 30314 12152
rect 29972 12112 29978 12124
rect 34514 12112 34520 12164
rect 34572 12152 34578 12164
rect 35342 12152 35348 12164
rect 34572 12124 35348 12152
rect 34572 12112 34578 12124
rect 35342 12112 35348 12124
rect 35400 12152 35406 12164
rect 36004 12152 36032 12183
rect 36538 12180 36544 12192
rect 36596 12220 36602 12232
rect 37274 12220 37280 12232
rect 36596 12192 37280 12220
rect 36596 12180 36602 12192
rect 37274 12180 37280 12192
rect 37332 12180 37338 12232
rect 39482 12180 39488 12232
rect 39540 12180 39546 12232
rect 39684 12229 39712 12260
rect 39669 12223 39727 12229
rect 39669 12189 39681 12223
rect 39715 12189 39727 12223
rect 39669 12183 39727 12189
rect 35400 12124 36032 12152
rect 35400 12112 35406 12124
rect 37550 12112 37556 12164
rect 37608 12112 37614 12164
rect 38838 12152 38844 12164
rect 38778 12124 38844 12152
rect 38838 12112 38844 12124
rect 38896 12112 38902 12164
rect 39301 12155 39359 12161
rect 39301 12121 39313 12155
rect 39347 12152 39359 12155
rect 39577 12155 39635 12161
rect 39577 12152 39589 12155
rect 39347 12124 39589 12152
rect 39347 12121 39359 12124
rect 39301 12115 39359 12121
rect 39577 12121 39589 12124
rect 39623 12121 39635 12155
rect 39577 12115 39635 12121
rect 24854 12084 24860 12096
rect 24412 12056 24860 12084
rect 24854 12044 24860 12056
rect 24912 12044 24918 12096
rect 26234 12044 26240 12096
rect 26292 12044 26298 12096
rect 26605 12087 26663 12093
rect 26605 12053 26617 12087
rect 26651 12084 26663 12087
rect 27154 12084 27160 12096
rect 26651 12056 27160 12084
rect 26651 12053 26663 12056
rect 26605 12047 26663 12053
rect 27154 12044 27160 12056
rect 27212 12044 27218 12096
rect 31386 12044 31392 12096
rect 31444 12044 31450 12096
rect 34790 12044 34796 12096
rect 34848 12084 34854 12096
rect 34885 12087 34943 12093
rect 34885 12084 34897 12087
rect 34848 12056 34897 12084
rect 34848 12044 34854 12056
rect 34885 12053 34897 12056
rect 34931 12053 34943 12087
rect 34885 12047 34943 12053
rect 35526 12044 35532 12096
rect 35584 12084 35590 12096
rect 36170 12084 36176 12096
rect 35584 12056 36176 12084
rect 35584 12044 35590 12056
rect 36170 12044 36176 12056
rect 36228 12044 36234 12096
rect 39025 12087 39083 12093
rect 39025 12053 39037 12087
rect 39071 12084 39083 12087
rect 39482 12084 39488 12096
rect 39071 12056 39488 12084
rect 39071 12053 39083 12056
rect 39025 12047 39083 12053
rect 39482 12044 39488 12056
rect 39540 12044 39546 12096
rect 1104 11994 42504 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 42504 11994
rect 1104 11920 42504 11942
rect 1765 11883 1823 11889
rect 1765 11849 1777 11883
rect 1811 11849 1823 11883
rect 1765 11843 1823 11849
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1780 11744 1808 11843
rect 3510 11840 3516 11892
rect 3568 11840 3574 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3620 11852 3985 11880
rect 1719 11716 1808 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1946 11704 1952 11756
rect 2004 11704 2010 11756
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2317 11747 2375 11753
rect 2317 11744 2329 11747
rect 2280 11716 2329 11744
rect 2280 11704 2286 11716
rect 2317 11713 2329 11716
rect 2363 11713 2375 11747
rect 2317 11707 2375 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2498 11744 2504 11756
rect 2455 11716 2504 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 2832 11716 3157 11744
rect 2832 11704 2838 11716
rect 3145 11713 3157 11716
rect 3191 11713 3203 11747
rect 3145 11707 3203 11713
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3620 11744 3648 11852
rect 3973 11849 3985 11852
rect 4019 11880 4031 11883
rect 4154 11880 4160 11892
rect 4019 11852 4160 11880
rect 4019 11849 4031 11852
rect 3973 11843 4031 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 5077 11883 5135 11889
rect 4632 11852 4936 11880
rect 3375 11716 3648 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 2130 11568 2136 11620
rect 2188 11608 2194 11620
rect 2516 11608 2544 11704
rect 3160 11676 3188 11707
rect 3786 11704 3792 11756
rect 3844 11704 3850 11756
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 4632 11753 4660 11852
rect 4908 11812 4936 11852
rect 5077 11849 5089 11883
rect 5123 11880 5135 11883
rect 5123 11852 6684 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 6656 11821 6684 11852
rect 10502 11840 10508 11892
rect 10560 11840 10566 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12913 11883 12971 11889
rect 12913 11880 12925 11883
rect 12032 11852 12925 11880
rect 12032 11840 12038 11852
rect 12913 11849 12925 11852
rect 12959 11849 12971 11883
rect 12913 11843 12971 11849
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 13906 11880 13912 11892
rect 13311 11852 13912 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18877 11883 18935 11889
rect 18877 11880 18889 11883
rect 18656 11852 18889 11880
rect 18656 11840 18662 11852
rect 18877 11849 18889 11852
rect 18923 11849 18935 11883
rect 18877 11843 18935 11849
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 22278 11880 22284 11892
rect 20947 11852 22284 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 22462 11840 22468 11892
rect 22520 11840 22526 11892
rect 23382 11880 23388 11892
rect 23124 11852 23388 11880
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 4908 11784 5181 11812
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 5169 11775 5227 11781
rect 6641 11815 6699 11821
rect 6641 11781 6653 11815
rect 6687 11812 6699 11815
rect 7006 11812 7012 11824
rect 6687 11784 7012 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 7006 11772 7012 11784
rect 7064 11812 7070 11824
rect 9585 11815 9643 11821
rect 7064 11784 7236 11812
rect 7064 11772 7070 11784
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4212 11716 4445 11744
rect 4212 11704 4218 11716
rect 4433 11713 4445 11716
rect 4479 11744 4491 11747
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4479 11716 4629 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 4893 11747 4951 11753
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 4939 11716 5457 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 3418 11676 3424 11688
rect 3160 11648 3424 11676
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11645 3663 11679
rect 3605 11639 3663 11645
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4908 11676 4936 11707
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7208 11753 7236 11784
rect 9585 11781 9597 11815
rect 9631 11812 9643 11815
rect 9766 11812 9772 11824
rect 9631 11784 9772 11812
rect 9631 11781 9643 11784
rect 9585 11775 9643 11781
rect 9766 11772 9772 11784
rect 9824 11772 9830 11824
rect 11514 11772 11520 11824
rect 11572 11772 11578 11824
rect 12710 11772 12716 11824
rect 12768 11772 12774 11824
rect 14366 11772 14372 11824
rect 14424 11821 14430 11824
rect 14424 11812 14436 11821
rect 14424 11784 14469 11812
rect 14424 11775 14436 11784
rect 14424 11772 14430 11775
rect 18506 11772 18512 11824
rect 18564 11812 18570 11824
rect 19751 11815 19809 11821
rect 19751 11812 19763 11815
rect 18564 11784 19763 11812
rect 18564 11772 18570 11784
rect 19751 11781 19763 11784
rect 19797 11781 19809 11815
rect 19751 11775 19809 11781
rect 19981 11815 20039 11821
rect 19981 11781 19993 11815
rect 20027 11812 20039 11815
rect 20162 11812 20168 11824
rect 20027 11784 20168 11812
rect 20027 11781 20039 11784
rect 19981 11775 20039 11781
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 20530 11772 20536 11824
rect 20588 11772 20594 11824
rect 20749 11815 20807 11821
rect 20749 11781 20761 11815
rect 20795 11812 20807 11815
rect 21358 11812 21364 11824
rect 20795 11784 21364 11812
rect 20795 11781 20807 11784
rect 20749 11775 20807 11781
rect 21358 11772 21364 11784
rect 21416 11772 21422 11824
rect 22189 11815 22247 11821
rect 22189 11781 22201 11815
rect 22235 11812 22247 11815
rect 23124 11812 23152 11852
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 24302 11840 24308 11892
rect 24360 11880 24366 11892
rect 26326 11880 26332 11892
rect 24360 11852 24900 11880
rect 24360 11840 24366 11852
rect 22235 11784 23152 11812
rect 23293 11815 23351 11821
rect 22235 11781 22247 11784
rect 22189 11775 22247 11781
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 23566 11812 23572 11824
rect 23339 11784 23572 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 23566 11772 23572 11784
rect 23624 11772 23630 11824
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 7558 11744 7564 11756
rect 7423 11716 7564 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 9861 11747 9919 11753
rect 9861 11713 9873 11747
rect 9907 11744 9919 11747
rect 9950 11744 9956 11756
rect 9907 11716 9956 11744
rect 9907 11713 9919 11716
rect 9861 11707 9919 11713
rect 9950 11704 9956 11716
rect 10008 11704 10014 11756
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 19576 11716 19625 11744
rect 19576 11704 19582 11716
rect 19613 11713 19625 11716
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 4111 11648 4936 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 3620 11608 3648 11639
rect 2188 11580 3648 11608
rect 2188 11568 2194 11580
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 1489 11543 1547 11549
rect 1489 11540 1501 11543
rect 900 11512 1501 11540
rect 900 11500 906 11512
rect 1489 11509 1501 11512
rect 1535 11509 1547 11543
rect 1489 11503 1547 11509
rect 2038 11500 2044 11552
rect 2096 11500 2102 11552
rect 3620 11540 3648 11580
rect 4080 11540 4108 11639
rect 5350 11636 5356 11688
rect 5408 11636 5414 11688
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 9582 11636 9588 11688
rect 9640 11676 9646 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9640 11648 9689 11676
rect 9640 11636 9646 11648
rect 9677 11645 9689 11648
rect 9723 11676 9735 11679
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 9723 11648 11069 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 14645 11679 14703 11685
rect 14645 11645 14657 11679
rect 14691 11676 14703 11679
rect 16850 11676 16856 11688
rect 14691 11648 16856 11676
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 19904 11676 19932 11707
rect 20070 11704 20076 11756
rect 20128 11704 20134 11756
rect 21818 11704 21824 11756
rect 21876 11704 21882 11756
rect 21914 11747 21972 11753
rect 21914 11713 21926 11747
rect 21960 11713 21972 11747
rect 21914 11707 21972 11713
rect 19536 11648 19932 11676
rect 19536 11620 19564 11648
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4338 11608 4344 11620
rect 4203 11580 4344 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4338 11568 4344 11580
rect 4396 11608 4402 11620
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 4396 11580 4813 11608
rect 4396 11568 4402 11580
rect 4801 11577 4813 11580
rect 4847 11608 4859 11611
rect 7742 11608 7748 11620
rect 4847 11580 5212 11608
rect 4847 11577 4859 11580
rect 4801 11571 4859 11577
rect 3620 11512 4108 11540
rect 4246 11500 4252 11552
rect 4304 11500 4310 11552
rect 4430 11500 4436 11552
rect 4488 11500 4494 11552
rect 5184 11549 5212 11580
rect 6932 11580 7748 11608
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11509 5227 11543
rect 5169 11503 5227 11509
rect 5626 11500 5632 11552
rect 5684 11500 5690 11552
rect 6932 11549 6960 11580
rect 7742 11568 7748 11580
rect 7800 11568 7806 11620
rect 19518 11568 19524 11620
rect 19576 11568 19582 11620
rect 6917 11543 6975 11549
rect 6917 11509 6929 11543
rect 6963 11509 6975 11543
rect 6917 11503 6975 11509
rect 7098 11500 7104 11552
rect 7156 11500 7162 11552
rect 7190 11500 7196 11552
rect 7248 11500 7254 11552
rect 9674 11500 9680 11552
rect 9732 11500 9738 11552
rect 10045 11543 10103 11549
rect 10045 11509 10057 11543
rect 10091 11540 10103 11543
rect 10410 11540 10416 11552
rect 10091 11512 10416 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12492 11512 12909 11540
rect 12492 11500 12498 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 19904 11540 19932 11648
rect 21450 11636 21456 11688
rect 21508 11676 21514 11688
rect 21545 11679 21603 11685
rect 21545 11676 21557 11679
rect 21508 11648 21557 11676
rect 21508 11636 21514 11648
rect 21545 11645 21557 11648
rect 21591 11645 21603 11679
rect 21545 11639 21603 11645
rect 20257 11611 20315 11617
rect 20257 11577 20269 11611
rect 20303 11608 20315 11611
rect 21928 11608 21956 11707
rect 22094 11704 22100 11756
rect 22152 11704 22158 11756
rect 22327 11747 22385 11753
rect 22327 11713 22339 11747
rect 22373 11744 22385 11747
rect 22830 11744 22836 11756
rect 22373 11716 22836 11744
rect 22373 11713 22385 11716
rect 22327 11707 22385 11713
rect 22830 11704 22836 11716
rect 22888 11704 22894 11756
rect 24394 11704 24400 11756
rect 24452 11704 24458 11756
rect 24872 11753 24900 11852
rect 25792 11852 26332 11880
rect 25792 11821 25820 11852
rect 26326 11840 26332 11852
rect 26384 11840 26390 11892
rect 26789 11883 26847 11889
rect 26789 11849 26801 11883
rect 26835 11880 26847 11883
rect 27985 11883 28043 11889
rect 27985 11880 27997 11883
rect 26835 11852 27997 11880
rect 26835 11849 26847 11852
rect 26789 11843 26847 11849
rect 27985 11849 27997 11852
rect 28031 11849 28043 11883
rect 27985 11843 28043 11849
rect 28537 11883 28595 11889
rect 28537 11849 28549 11883
rect 28583 11849 28595 11883
rect 30374 11880 30380 11892
rect 28537 11843 28595 11849
rect 28920 11852 30380 11880
rect 25225 11815 25283 11821
rect 25225 11781 25237 11815
rect 25271 11812 25283 11815
rect 25777 11815 25835 11821
rect 25777 11812 25789 11815
rect 25271 11784 25789 11812
rect 25271 11781 25283 11784
rect 25225 11775 25283 11781
rect 25777 11781 25789 11784
rect 25823 11781 25835 11815
rect 25777 11775 25835 11781
rect 25961 11815 26019 11821
rect 25961 11781 25973 11815
rect 26007 11812 26019 11815
rect 26421 11815 26479 11821
rect 26421 11812 26433 11815
rect 26007 11784 26433 11812
rect 26007 11781 26019 11784
rect 25961 11775 26019 11781
rect 26421 11781 26433 11784
rect 26467 11781 26479 11815
rect 26421 11775 26479 11781
rect 27154 11772 27160 11824
rect 27212 11772 27218 11824
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11713 24915 11747
rect 24857 11707 24915 11713
rect 24950 11747 25008 11753
rect 24950 11713 24962 11747
rect 24996 11713 25008 11747
rect 24950 11707 25008 11713
rect 25133 11747 25191 11753
rect 25133 11713 25145 11747
rect 25179 11713 25191 11747
rect 25133 11707 25191 11713
rect 25363 11747 25421 11753
rect 25363 11713 25375 11747
rect 25409 11744 25421 11747
rect 25498 11744 25504 11756
rect 25409 11716 25504 11744
rect 25409 11713 25421 11716
rect 25363 11707 25421 11713
rect 23017 11679 23075 11685
rect 23017 11645 23029 11679
rect 23063 11676 23075 11679
rect 23063 11648 23152 11676
rect 23063 11645 23075 11648
rect 23017 11639 23075 11645
rect 20303 11580 21956 11608
rect 20303 11577 20315 11580
rect 20257 11571 20315 11577
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 19904 11512 20729 11540
rect 12897 11503 12955 11509
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 20717 11503 20775 11509
rect 20993 11543 21051 11549
rect 20993 11509 21005 11543
rect 21039 11540 21051 11543
rect 21082 11540 21088 11552
rect 21039 11512 21088 11540
rect 21039 11509 21051 11512
rect 20993 11503 21051 11509
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 23124 11540 23152 11648
rect 24762 11636 24768 11688
rect 24820 11676 24826 11688
rect 24965 11676 24993 11707
rect 24820 11648 24993 11676
rect 24820 11636 24826 11648
rect 23382 11540 23388 11552
rect 23124 11512 23388 11540
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 23658 11500 23664 11552
rect 23716 11540 23722 11552
rect 25148 11540 25176 11707
rect 25498 11704 25504 11716
rect 25556 11744 25562 11756
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25556 11716 25605 11744
rect 25556 11704 25562 11716
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11713 26295 11747
rect 26237 11707 26295 11713
rect 26513 11747 26571 11753
rect 26513 11713 26525 11747
rect 26559 11713 26571 11747
rect 26513 11707 26571 11713
rect 26605 11747 26663 11753
rect 26605 11713 26617 11747
rect 26651 11744 26663 11747
rect 27430 11744 27436 11756
rect 26651 11716 27436 11744
rect 26651 11713 26663 11716
rect 26605 11707 26663 11713
rect 26252 11676 26280 11707
rect 25516 11648 26280 11676
rect 26528 11676 26556 11707
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 27890 11704 27896 11756
rect 27948 11704 27954 11756
rect 28169 11747 28227 11753
rect 28169 11713 28181 11747
rect 28215 11744 28227 11747
rect 28552 11744 28580 11843
rect 28920 11821 28948 11852
rect 30374 11840 30380 11852
rect 30432 11840 30438 11892
rect 34606 11880 34612 11892
rect 34532 11852 34612 11880
rect 28905 11815 28963 11821
rect 28905 11781 28917 11815
rect 28951 11781 28963 11815
rect 28905 11775 28963 11781
rect 28994 11772 29000 11824
rect 29052 11812 29058 11824
rect 29914 11812 29920 11824
rect 29052 11784 29920 11812
rect 29052 11772 29058 11784
rect 29914 11772 29920 11784
rect 29972 11812 29978 11824
rect 31297 11815 31355 11821
rect 29972 11784 30130 11812
rect 29972 11772 29978 11784
rect 31297 11781 31309 11815
rect 31343 11812 31355 11815
rect 31386 11812 31392 11824
rect 31343 11784 31392 11812
rect 31343 11781 31355 11784
rect 31297 11775 31355 11781
rect 31386 11772 31392 11784
rect 31444 11772 31450 11824
rect 32398 11772 32404 11824
rect 32456 11772 32462 11824
rect 34330 11812 34336 11824
rect 32692 11784 34336 11812
rect 28215 11716 28580 11744
rect 28215 11713 28227 11716
rect 28169 11707 28227 11713
rect 28718 11704 28724 11756
rect 28776 11704 28782 11756
rect 28810 11704 28816 11756
rect 28868 11704 28874 11756
rect 29089 11747 29147 11753
rect 29089 11713 29101 11747
rect 29135 11744 29147 11747
rect 29135 11716 29868 11744
rect 29135 11713 29147 11716
rect 29089 11707 29147 11713
rect 27522 11676 27528 11688
rect 26528 11648 27528 11676
rect 25516 11617 25544 11648
rect 27522 11636 27528 11648
rect 27580 11676 27586 11688
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 27580 11648 27721 11676
rect 27580 11636 27586 11648
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 27982 11636 27988 11688
rect 28040 11676 28046 11688
rect 28828 11676 28856 11704
rect 28040 11648 28856 11676
rect 28040 11636 28046 11648
rect 25501 11611 25559 11617
rect 25501 11577 25513 11611
rect 25547 11577 25559 11611
rect 25501 11571 25559 11577
rect 23716 11512 25176 11540
rect 23716 11500 23722 11512
rect 28350 11500 28356 11552
rect 28408 11500 28414 11552
rect 29840 11549 29868 11716
rect 31846 11704 31852 11756
rect 31904 11744 31910 11756
rect 32309 11747 32367 11753
rect 32309 11744 32321 11747
rect 31904 11716 32321 11744
rect 31904 11704 31910 11716
rect 32309 11713 32321 11716
rect 32355 11713 32367 11747
rect 32309 11707 32367 11713
rect 32490 11704 32496 11756
rect 32548 11704 32554 11756
rect 32692 11753 32720 11784
rect 34330 11772 34336 11784
rect 34388 11772 34394 11824
rect 32677 11747 32735 11753
rect 32677 11713 32689 11747
rect 32723 11713 32735 11747
rect 32677 11707 32735 11713
rect 33962 11704 33968 11756
rect 34020 11704 34026 11756
rect 34057 11747 34115 11753
rect 34057 11713 34069 11747
rect 34103 11713 34115 11747
rect 34057 11707 34115 11713
rect 34241 11747 34299 11753
rect 34241 11713 34253 11747
rect 34287 11744 34299 11747
rect 34532 11744 34560 11852
rect 34606 11840 34612 11852
rect 34664 11840 34670 11892
rect 36170 11840 36176 11892
rect 36228 11880 36234 11892
rect 36265 11883 36323 11889
rect 36265 11880 36277 11883
rect 36228 11852 36277 11880
rect 36228 11840 36234 11852
rect 36265 11849 36277 11852
rect 36311 11849 36323 11883
rect 36265 11843 36323 11849
rect 34790 11772 34796 11824
rect 34848 11772 34854 11824
rect 34287 11716 34560 11744
rect 36280 11744 36308 11843
rect 37274 11840 37280 11892
rect 37332 11880 37338 11892
rect 37332 11852 40172 11880
rect 37332 11840 37338 11852
rect 38838 11772 38844 11824
rect 38896 11772 38902 11824
rect 36909 11747 36967 11753
rect 36909 11744 36921 11747
rect 34287 11713 34299 11716
rect 34241 11707 34299 11713
rect 31570 11636 31576 11688
rect 31628 11636 31634 11688
rect 32582 11636 32588 11688
rect 32640 11676 32646 11688
rect 34072 11676 34100 11707
rect 32640 11648 34100 11676
rect 32640 11636 32646 11648
rect 34514 11636 34520 11688
rect 34572 11636 34578 11688
rect 35250 11636 35256 11688
rect 35308 11676 35314 11688
rect 35526 11676 35532 11688
rect 35308 11648 35532 11676
rect 35308 11636 35314 11648
rect 35526 11636 35532 11648
rect 35584 11636 35590 11688
rect 35912 11676 35940 11730
rect 36280 11716 36921 11744
rect 36909 11713 36921 11716
rect 36955 11713 36967 11747
rect 36909 11707 36967 11713
rect 37826 11704 37832 11756
rect 37884 11704 37890 11756
rect 37918 11704 37924 11756
rect 37976 11744 37982 11756
rect 40144 11753 40172 11852
rect 40129 11747 40187 11753
rect 37976 11716 38240 11744
rect 37976 11704 37982 11716
rect 38212 11688 38240 11716
rect 40129 11713 40141 11747
rect 40175 11713 40187 11747
rect 40129 11707 40187 11713
rect 36446 11676 36452 11688
rect 35912 11648 36452 11676
rect 36446 11636 36452 11648
rect 36504 11636 36510 11688
rect 37734 11636 37740 11688
rect 37792 11636 37798 11688
rect 38105 11679 38163 11685
rect 38105 11645 38117 11679
rect 38151 11645 38163 11679
rect 38105 11639 38163 11645
rect 32858 11568 32864 11620
rect 32916 11608 32922 11620
rect 34532 11608 34560 11636
rect 32916 11580 34560 11608
rect 32916 11568 32922 11580
rect 37550 11568 37556 11620
rect 37608 11568 37614 11620
rect 38120 11608 38148 11639
rect 38194 11636 38200 11688
rect 38252 11636 38258 11688
rect 39853 11679 39911 11685
rect 39853 11645 39865 11679
rect 39899 11676 39911 11679
rect 40221 11679 40279 11685
rect 40221 11676 40233 11679
rect 39899 11648 40233 11676
rect 39899 11645 39911 11648
rect 39853 11639 39911 11645
rect 40221 11645 40233 11648
rect 40267 11645 40279 11679
rect 40221 11639 40279 11645
rect 40770 11636 40776 11688
rect 40828 11636 40834 11688
rect 38838 11608 38844 11620
rect 38120 11580 38844 11608
rect 38838 11568 38844 11580
rect 38896 11568 38902 11620
rect 29825 11543 29883 11549
rect 29825 11509 29837 11543
rect 29871 11540 29883 11543
rect 30834 11540 30840 11552
rect 29871 11512 30840 11540
rect 29871 11509 29883 11512
rect 29825 11503 29883 11509
rect 30834 11500 30840 11512
rect 30892 11540 30898 11552
rect 31294 11540 31300 11552
rect 30892 11512 31300 11540
rect 30892 11500 30898 11512
rect 31294 11500 31300 11512
rect 31352 11500 31358 11552
rect 32125 11543 32183 11549
rect 32125 11509 32137 11543
rect 32171 11540 32183 11543
rect 32214 11540 32220 11552
rect 32171 11512 32220 11540
rect 32171 11509 32183 11512
rect 32125 11503 32183 11509
rect 32214 11500 32220 11512
rect 32272 11500 32278 11552
rect 34422 11500 34428 11552
rect 34480 11500 34486 11552
rect 36354 11500 36360 11552
rect 36412 11500 36418 11552
rect 38378 11500 38384 11552
rect 38436 11500 38442 11552
rect 1104 11450 42504 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 42504 11450
rect 1104 11376 42504 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2317 11339 2375 11345
rect 2317 11336 2329 11339
rect 2004 11308 2329 11336
rect 2004 11296 2010 11308
rect 2317 11305 2329 11308
rect 2363 11336 2375 11339
rect 5353 11339 5411 11345
rect 2363 11308 3188 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11237 1823 11271
rect 1765 11231 1823 11237
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 1780 11132 1808 11231
rect 2498 11228 2504 11280
rect 2556 11228 2562 11280
rect 2961 11271 3019 11277
rect 2961 11268 2973 11271
rect 2746 11240 2973 11268
rect 2038 11160 2044 11212
rect 2096 11160 2102 11212
rect 2746 11200 2774 11240
rect 2961 11237 2973 11240
rect 3007 11237 3019 11271
rect 2961 11231 3019 11237
rect 3160 11268 3188 11308
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 5399 11308 6377 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 6365 11305 6377 11308
rect 6411 11336 6423 11339
rect 6638 11336 6644 11348
rect 6411 11308 6644 11336
rect 6411 11305 6423 11308
rect 6365 11299 6423 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 9950 11336 9956 11348
rect 9508 11308 9956 11336
rect 4062 11268 4068 11280
rect 3160 11240 4068 11268
rect 3160 11212 3188 11240
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 5537 11271 5595 11277
rect 5537 11237 5549 11271
rect 5583 11268 5595 11271
rect 5718 11268 5724 11280
rect 5583 11240 5724 11268
rect 5583 11237 5595 11240
rect 5537 11231 5595 11237
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 7377 11271 7435 11277
rect 6656 11240 7328 11268
rect 2516 11172 2774 11200
rect 1719 11104 1808 11132
rect 1949 11135 2007 11141
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 1949 11101 1961 11135
rect 1995 11132 2007 11135
rect 2130 11132 2136 11144
rect 1995 11104 2136 11132
rect 1995 11101 2007 11104
rect 1949 11095 2007 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2516 11141 2544 11172
rect 3142 11160 3148 11212
rect 3200 11160 3206 11212
rect 3510 11160 3516 11212
rect 3568 11160 3574 11212
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 6656 11209 6684 11240
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 5684 11172 6653 11200
rect 5684 11160 5690 11172
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 6825 11203 6883 11209
rect 6825 11169 6837 11203
rect 6871 11200 6883 11203
rect 7190 11200 7196 11212
rect 6871 11172 7196 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7300 11200 7328 11240
rect 7377 11237 7389 11271
rect 7423 11268 7435 11271
rect 7558 11268 7564 11280
rect 7423 11240 7564 11268
rect 7423 11237 7435 11240
rect 7377 11231 7435 11237
rect 7558 11228 7564 11240
rect 7616 11228 7622 11280
rect 9508 11277 9536 11308
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10137 11339 10195 11345
rect 10137 11305 10149 11339
rect 10183 11336 10195 11339
rect 10502 11336 10508 11348
rect 10183 11308 10508 11336
rect 10183 11305 10195 11308
rect 10137 11299 10195 11305
rect 9493 11271 9551 11277
rect 9493 11237 9505 11271
rect 9539 11237 9551 11271
rect 9493 11231 9551 11237
rect 9582 11228 9588 11280
rect 9640 11228 9646 11280
rect 10152 11268 10180 11299
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 13173 11339 13231 11345
rect 13173 11305 13185 11339
rect 13219 11336 13231 11339
rect 14274 11336 14280 11348
rect 13219 11308 14280 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 18506 11296 18512 11348
rect 18564 11296 18570 11348
rect 21358 11296 21364 11348
rect 21416 11296 21422 11348
rect 21450 11296 21456 11348
rect 21508 11296 21514 11348
rect 27522 11296 27528 11348
rect 27580 11296 27586 11348
rect 27890 11296 27896 11348
rect 27948 11336 27954 11348
rect 28261 11339 28319 11345
rect 28261 11336 28273 11339
rect 27948 11308 28273 11336
rect 27948 11296 27954 11308
rect 28261 11305 28273 11308
rect 28307 11305 28319 11339
rect 28261 11299 28319 11305
rect 32401 11339 32459 11345
rect 32401 11305 32413 11339
rect 32447 11336 32459 11339
rect 32582 11336 32588 11348
rect 32447 11308 32588 11336
rect 32447 11305 32459 11308
rect 32401 11299 32459 11305
rect 32582 11296 32588 11308
rect 32640 11296 32646 11348
rect 33962 11296 33968 11348
rect 34020 11336 34026 11348
rect 34425 11339 34483 11345
rect 34425 11336 34437 11339
rect 34020 11308 34437 11336
rect 34020 11296 34026 11308
rect 34425 11305 34437 11308
rect 34471 11305 34483 11339
rect 34425 11299 34483 11305
rect 34698 11296 34704 11348
rect 34756 11336 34762 11348
rect 34977 11339 35035 11345
rect 34977 11336 34989 11339
rect 34756 11308 34989 11336
rect 34756 11296 34762 11308
rect 34977 11305 34989 11308
rect 35023 11305 35035 11339
rect 35986 11336 35992 11348
rect 34977 11299 35035 11305
rect 35452 11308 35992 11336
rect 9692 11240 10180 11268
rect 13909 11271 13967 11277
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 7300 11172 7481 11200
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7576 11200 7604 11228
rect 7576 11172 8064 11200
rect 7469 11163 7527 11169
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2280 11104 2421 11132
rect 2280 11092 2286 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11132 3295 11135
rect 3528 11132 3556 11160
rect 3283 11104 3556 11132
rect 3283 11101 3295 11104
rect 3237 11095 3295 11101
rect 2792 11064 2820 11095
rect 3252 11064 3280 11095
rect 3878 11092 3884 11144
rect 3936 11092 3942 11144
rect 6086 11132 6092 11144
rect 4724 11104 6092 11132
rect 2792 11036 3280 11064
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 3513 11067 3571 11073
rect 3513 11064 3525 11067
rect 3476 11036 3525 11064
rect 3476 11024 3482 11036
rect 3513 11033 3525 11036
rect 3559 11033 3571 11067
rect 3513 11027 3571 11033
rect 3605 11067 3663 11073
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 4724 11064 4752 11104
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6549 11135 6607 11141
rect 6549 11101 6561 11135
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 6914 11132 6920 11144
rect 6779 11104 6920 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 3651 11036 4752 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 5169 11067 5227 11073
rect 5169 11064 5181 11067
rect 4856 11036 5181 11064
rect 4856 11024 4862 11036
rect 5169 11033 5181 11036
rect 5215 11033 5227 11067
rect 6564 11064 6592 11095
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7285 11135 7343 11141
rect 7285 11132 7297 11135
rect 7156 11104 7297 11132
rect 7156 11092 7162 11104
rect 7285 11101 7297 11104
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 7374 11064 7380 11076
rect 6564 11036 7380 11064
rect 5169 11027 5227 11033
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 7484 11064 7512 11163
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7742 11132 7748 11144
rect 7607 11104 7748 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 8036 11141 8064 11172
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9398 11132 9404 11144
rect 9355 11104 9404 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 7852 11064 7880 11095
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9490 11102 9496 11154
rect 9548 11102 9554 11154
rect 9585 11135 9643 11141
rect 9493 11101 9505 11102
rect 9539 11101 9551 11102
rect 9493 11095 9551 11101
rect 9585 11101 9597 11135
rect 9631 11101 9643 11135
rect 9585 11095 9643 11101
rect 7484 11036 7880 11064
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 9600 11064 9628 11095
rect 9692 11064 9720 11240
rect 13909 11237 13921 11271
rect 13955 11268 13967 11271
rect 14550 11268 14556 11280
rect 13955 11240 14556 11268
rect 13955 11237 13967 11240
rect 13909 11231 13967 11237
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 9784 11172 10517 11200
rect 9784 11144 9812 11172
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 8168 11036 9720 11064
rect 9876 11064 9904 11092
rect 10336 11073 10364 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11480 11172 12265 11200
rect 11480 11160 11486 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 13170 11160 13176 11212
rect 13228 11200 13234 11212
rect 13449 11203 13507 11209
rect 13449 11200 13461 11203
rect 13228 11172 13461 11200
rect 13228 11160 13234 11172
rect 13449 11169 13461 11172
rect 13495 11169 13507 11203
rect 13449 11163 13507 11169
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 13078 11132 13084 11144
rect 12851 11104 13084 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 18782 11092 18788 11144
rect 18840 11092 18846 11144
rect 18892 11132 18920 11163
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19484 11172 19625 11200
rect 19484 11160 19490 11172
rect 19613 11169 19625 11172
rect 19659 11200 19671 11203
rect 20438 11200 20444 11212
rect 19659 11172 20444 11200
rect 19659 11169 19671 11172
rect 19613 11163 19671 11169
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 21634 11160 21640 11212
rect 21692 11200 21698 11212
rect 22925 11203 22983 11209
rect 22925 11200 22937 11203
rect 21692 11172 22937 11200
rect 21692 11160 21698 11172
rect 22925 11169 22937 11172
rect 22971 11169 22983 11203
rect 22925 11163 22983 11169
rect 26053 11203 26111 11209
rect 26053 11169 26065 11203
rect 26099 11200 26111 11203
rect 26142 11200 26148 11212
rect 26099 11172 26148 11200
rect 26099 11169 26111 11172
rect 26053 11163 26111 11169
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 19518 11132 19524 11144
rect 18892 11104 19524 11132
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 23201 11135 23259 11141
rect 23201 11101 23213 11135
rect 23247 11132 23259 11135
rect 23382 11132 23388 11144
rect 23247 11104 23388 11132
rect 23247 11101 23259 11104
rect 23201 11095 23259 11101
rect 23382 11092 23388 11104
rect 23440 11132 23446 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 23440 11104 24777 11132
rect 23440 11092 23446 11104
rect 24765 11101 24777 11104
rect 24811 11132 24823 11135
rect 24854 11132 24860 11144
rect 24811 11104 24860 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 24854 11092 24860 11104
rect 24912 11132 24918 11144
rect 25774 11132 25780 11144
rect 24912 11104 25780 11132
rect 24912 11092 24918 11104
rect 25774 11092 25780 11104
rect 25832 11092 25838 11144
rect 27540 11132 27568 11296
rect 33413 11271 33471 11277
rect 33413 11237 33425 11271
rect 33459 11268 33471 11271
rect 33594 11268 33600 11280
rect 33459 11240 33600 11268
rect 33459 11237 33471 11240
rect 33413 11231 33471 11237
rect 33594 11228 33600 11240
rect 33652 11228 33658 11280
rect 27801 11203 27859 11209
rect 27801 11169 27813 11203
rect 27847 11169 27859 11203
rect 27801 11163 27859 11169
rect 27709 11135 27767 11141
rect 27709 11132 27721 11135
rect 27540 11104 27721 11132
rect 27709 11101 27721 11104
rect 27755 11101 27767 11135
rect 27709 11095 27767 11101
rect 10105 11067 10163 11073
rect 10105 11064 10117 11067
rect 9876 11036 10117 11064
rect 8168 11024 8174 11036
rect 10105 11033 10117 11036
rect 10151 11033 10163 11067
rect 10105 11027 10163 11033
rect 10321 11067 10379 11073
rect 10321 11033 10333 11067
rect 10367 11033 10379 11067
rect 10321 11027 10379 11033
rect 10428 11036 10810 11064
rect 1486 10956 1492 11008
rect 1544 10956 1550 11008
rect 2685 10999 2743 11005
rect 2685 10965 2697 10999
rect 2731 10996 2743 10999
rect 3142 10996 3148 11008
rect 2731 10968 3148 10996
rect 2731 10965 2743 10968
rect 2685 10959 2743 10965
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 5258 10956 5264 11008
rect 5316 10996 5322 11008
rect 5379 10999 5437 11005
rect 5379 10996 5391 10999
rect 5316 10968 5391 10996
rect 5316 10956 5322 10968
rect 5379 10965 5391 10968
rect 5425 10996 5437 10999
rect 5810 10996 5816 11008
rect 5425 10968 5816 10996
rect 5425 10965 5437 10968
rect 5379 10959 5437 10965
rect 5810 10956 5816 10968
rect 5868 10956 5874 11008
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7616 10968 7757 10996
rect 7616 10956 7622 10968
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 7745 10959 7803 10965
rect 7926 10956 7932 11008
rect 7984 10956 7990 11008
rect 9628 10956 9634 11008
rect 9686 10996 9692 11008
rect 9766 10996 9772 11008
rect 9686 10968 9772 10996
rect 9686 10956 9692 10968
rect 9766 10956 9772 10968
rect 9824 10996 9830 11008
rect 9953 10999 10011 11005
rect 9953 10996 9965 10999
rect 9824 10968 9965 10996
rect 9824 10956 9830 10968
rect 9953 10965 9965 10968
rect 9999 10965 10011 10999
rect 9953 10959 10011 10965
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 10428 10996 10456 11036
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 11977 11067 12035 11073
rect 11977 11064 11989 11067
rect 11940 11036 11989 11064
rect 11940 11024 11946 11036
rect 11977 11033 11989 11036
rect 12023 11033 12035 11067
rect 11977 11027 12035 11033
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 13906 11064 13912 11076
rect 13035 11036 13912 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 19610 11064 19616 11076
rect 19392 11036 19616 11064
rect 19392 11024 19398 11036
rect 19610 11024 19616 11036
rect 19668 11024 19674 11076
rect 19889 11067 19947 11073
rect 19889 11033 19901 11067
rect 19935 11064 19947 11067
rect 20162 11064 20168 11076
rect 19935 11036 20168 11064
rect 19935 11033 19947 11036
rect 19889 11027 19947 11033
rect 20162 11024 20168 11036
rect 20220 11024 20226 11076
rect 24394 11064 24400 11076
rect 20272 11036 20378 11064
rect 22494 11036 24400 11064
rect 10284 10968 10456 10996
rect 10284 10956 10290 10968
rect 18874 10956 18880 11008
rect 18932 10996 18938 11008
rect 20272 10996 20300 11036
rect 24394 11024 24400 11036
rect 24452 11024 24458 11076
rect 27278 11036 27384 11064
rect 20806 10996 20812 11008
rect 18932 10968 20812 10996
rect 18932 10956 18938 10968
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 27356 10996 27384 11036
rect 27430 11024 27436 11076
rect 27488 11064 27494 11076
rect 27816 11064 27844 11163
rect 30374 11160 30380 11212
rect 30432 11200 30438 11212
rect 31389 11203 31447 11209
rect 31389 11200 31401 11203
rect 30432 11172 31401 11200
rect 30432 11160 30438 11172
rect 31389 11169 31401 11172
rect 31435 11169 31447 11203
rect 32398 11200 32404 11212
rect 31389 11163 31447 11169
rect 31588 11172 32404 11200
rect 27982 11092 27988 11144
rect 28040 11092 28046 11144
rect 28074 11092 28080 11144
rect 28132 11132 28138 11144
rect 28718 11132 28724 11144
rect 28132 11104 28724 11132
rect 28132 11092 28138 11104
rect 28718 11092 28724 11104
rect 28776 11092 28782 11144
rect 31294 11092 31300 11144
rect 31352 11092 31358 11144
rect 31588 11141 31616 11172
rect 32398 11160 32404 11172
rect 32456 11160 32462 11212
rect 32490 11160 32496 11212
rect 32548 11200 32554 11212
rect 33965 11203 34023 11209
rect 33965 11200 33977 11203
rect 32548 11172 33977 11200
rect 32548 11160 32554 11172
rect 33965 11169 33977 11172
rect 34011 11169 34023 11203
rect 34330 11200 34336 11212
rect 33965 11163 34023 11169
rect 34072 11172 34336 11200
rect 31573 11135 31631 11141
rect 31573 11101 31585 11135
rect 31619 11101 31631 11135
rect 31573 11095 31631 11101
rect 31665 11135 31723 11141
rect 31665 11101 31677 11135
rect 31711 11132 31723 11135
rect 31754 11132 31760 11144
rect 31711 11104 31760 11132
rect 31711 11101 31723 11104
rect 31665 11095 31723 11101
rect 31754 11092 31760 11104
rect 31812 11092 31818 11144
rect 31849 11135 31907 11141
rect 31849 11101 31861 11135
rect 31895 11132 31907 11135
rect 31941 11135 31999 11141
rect 31941 11132 31953 11135
rect 31895 11104 31953 11132
rect 31895 11101 31907 11104
rect 31849 11095 31907 11101
rect 31941 11101 31953 11104
rect 31987 11101 31999 11135
rect 31941 11095 31999 11101
rect 32214 11092 32220 11144
rect 32272 11092 32278 11144
rect 33229 11135 33287 11141
rect 33229 11101 33241 11135
rect 33275 11101 33287 11135
rect 33229 11095 33287 11101
rect 33873 11135 33931 11141
rect 33873 11101 33885 11135
rect 33919 11132 33931 11135
rect 34072 11132 34100 11172
rect 34330 11160 34336 11172
rect 34388 11160 34394 11212
rect 35452 11209 35480 11308
rect 35986 11296 35992 11308
rect 36044 11296 36050 11348
rect 36262 11296 36268 11348
rect 36320 11296 36326 11348
rect 37366 11336 37372 11348
rect 36464 11308 37372 11336
rect 35437 11203 35495 11209
rect 35437 11169 35449 11203
rect 35483 11169 35495 11203
rect 35437 11163 35495 11169
rect 35526 11160 35532 11212
rect 35584 11160 35590 11212
rect 36354 11200 36360 11212
rect 35820 11172 36360 11200
rect 33919 11104 34100 11132
rect 34149 11135 34207 11141
rect 33919 11101 33931 11104
rect 33873 11095 33931 11101
rect 34149 11101 34161 11135
rect 34195 11101 34207 11135
rect 34149 11095 34207 11101
rect 27488 11036 27844 11064
rect 27488 11024 27494 11036
rect 27890 11024 27896 11076
rect 27948 11024 27954 11076
rect 28350 11024 28356 11076
rect 28408 11064 28414 11076
rect 32033 11067 32091 11073
rect 32033 11064 32045 11067
rect 28408 11036 32045 11064
rect 28408 11024 28414 11036
rect 32033 11033 32045 11036
rect 32079 11033 32091 11067
rect 32033 11027 32091 11033
rect 27908 10996 27936 11024
rect 27356 10968 27936 10996
rect 29270 10956 29276 11008
rect 29328 10996 29334 11008
rect 33244 10996 33272 11095
rect 34164 11064 34192 11095
rect 34238 11092 34244 11144
rect 34296 11092 34302 11144
rect 34514 11132 34520 11144
rect 34348 11104 34520 11132
rect 34348 11064 34376 11104
rect 34514 11092 34520 11104
rect 34572 11132 34578 11144
rect 34790 11132 34796 11144
rect 34572 11104 34796 11132
rect 34572 11092 34578 11104
rect 34790 11092 34796 11104
rect 34848 11092 34854 11144
rect 35345 11135 35403 11141
rect 35345 11101 35357 11135
rect 35391 11132 35403 11135
rect 35820 11132 35848 11172
rect 36354 11160 36360 11172
rect 36412 11160 36418 11212
rect 35391 11104 35848 11132
rect 36265 11135 36323 11141
rect 35391 11101 35403 11104
rect 35345 11095 35403 11101
rect 36265 11101 36277 11135
rect 36311 11132 36323 11135
rect 36464 11132 36492 11308
rect 37366 11296 37372 11308
rect 37424 11296 37430 11348
rect 37826 11296 37832 11348
rect 37884 11296 37890 11348
rect 38838 11296 38844 11348
rect 38896 11336 38902 11348
rect 38933 11339 38991 11345
rect 38933 11336 38945 11339
rect 38896 11308 38945 11336
rect 38896 11296 38902 11308
rect 38933 11305 38945 11308
rect 38979 11305 38991 11339
rect 38933 11299 38991 11305
rect 37737 11271 37795 11277
rect 37737 11268 37749 11271
rect 36556 11240 37749 11268
rect 36556 11141 36584 11240
rect 37737 11237 37749 11240
rect 37783 11237 37795 11271
rect 37737 11231 37795 11237
rect 36998 11200 37004 11212
rect 36832 11172 37004 11200
rect 36832 11141 36860 11172
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 37844 11200 37872 11296
rect 37108 11172 37872 11200
rect 37108 11141 37136 11172
rect 38102 11160 38108 11212
rect 38160 11160 38166 11212
rect 39482 11160 39488 11212
rect 39540 11160 39546 11212
rect 36311 11104 36492 11132
rect 36541 11135 36599 11141
rect 36311 11101 36323 11104
rect 36265 11095 36323 11101
rect 36541 11101 36553 11135
rect 36587 11101 36599 11135
rect 36541 11095 36599 11101
rect 36817 11135 36875 11141
rect 36817 11101 36829 11135
rect 36863 11101 36875 11135
rect 36817 11095 36875 11101
rect 37093 11135 37151 11141
rect 37093 11101 37105 11135
rect 37139 11101 37151 11135
rect 37093 11095 37151 11101
rect 37182 11092 37188 11144
rect 37240 11092 37246 11144
rect 37458 11092 37464 11144
rect 37516 11092 37522 11144
rect 37553 11135 37611 11141
rect 37553 11101 37565 11135
rect 37599 11132 37611 11135
rect 37642 11132 37648 11144
rect 37599 11104 37648 11132
rect 37599 11101 37611 11104
rect 37553 11095 37611 11101
rect 37642 11092 37648 11104
rect 37700 11092 37706 11144
rect 38197 11135 38255 11141
rect 38197 11101 38209 11135
rect 38243 11132 38255 11135
rect 38378 11132 38384 11144
rect 38243 11104 38384 11132
rect 38243 11101 38255 11104
rect 38197 11095 38255 11101
rect 38378 11092 38384 11104
rect 38436 11092 38442 11144
rect 34164 11036 34376 11064
rect 34422 11024 34428 11076
rect 34480 11064 34486 11076
rect 37369 11067 37427 11073
rect 37369 11064 37381 11067
rect 34480 11036 37381 11064
rect 34480 11024 34486 11036
rect 37369 11033 37381 11036
rect 37415 11033 37427 11067
rect 37369 11027 37427 11033
rect 29328 10968 33272 10996
rect 29328 10956 29334 10968
rect 34238 10956 34244 11008
rect 34296 10996 34302 11008
rect 35986 10996 35992 11008
rect 34296 10968 35992 10996
rect 34296 10956 34302 10968
rect 35986 10956 35992 10968
rect 36044 10956 36050 11008
rect 37458 10956 37464 11008
rect 37516 10996 37522 11008
rect 37734 10996 37740 11008
rect 37516 10968 37740 10996
rect 37516 10956 37522 10968
rect 37734 10956 37740 10968
rect 37792 10956 37798 11008
rect 37918 10956 37924 11008
rect 37976 10996 37982 11008
rect 38562 10996 38568 11008
rect 37976 10968 38568 10996
rect 37976 10956 37982 10968
rect 38562 10956 38568 10968
rect 38620 10996 38626 11008
rect 40862 10996 40868 11008
rect 38620 10968 40868 10996
rect 38620 10956 38626 10968
rect 40862 10956 40868 10968
rect 40920 10956 40926 11008
rect 1104 10906 42504 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 42504 10906
rect 1104 10832 42504 10854
rect 2498 10792 2504 10804
rect 1688 10764 2504 10792
rect 1688 10733 1716 10764
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3878 10792 3884 10804
rect 3191 10764 3884 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 5810 10752 5816 10804
rect 5868 10752 5874 10804
rect 6086 10752 6092 10804
rect 6144 10752 6150 10804
rect 7650 10792 7656 10804
rect 6656 10764 7656 10792
rect 1673 10727 1731 10733
rect 1673 10693 1685 10727
rect 1719 10693 1731 10727
rect 2958 10724 2964 10736
rect 2898 10696 2964 10724
rect 1673 10687 1731 10693
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 5353 10727 5411 10733
rect 5353 10693 5365 10727
rect 5399 10724 5411 10727
rect 6656 10724 6684 10764
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8110 10792 8116 10804
rect 7800 10764 8116 10792
rect 7800 10752 7806 10764
rect 8110 10752 8116 10764
rect 8168 10792 8174 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 8168 10764 8493 10792
rect 8168 10752 8174 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 10042 10792 10048 10804
rect 8481 10755 8539 10761
rect 9876 10764 10048 10792
rect 5399 10696 6684 10724
rect 5399 10693 5411 10696
rect 5353 10687 5411 10693
rect 6730 10684 6736 10736
rect 6788 10684 6794 10736
rect 6917 10727 6975 10733
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 7006 10724 7012 10736
rect 6963 10696 7012 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 7006 10684 7012 10696
rect 7064 10684 7070 10736
rect 9876 10724 9904 10764
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 17954 10752 17960 10804
rect 18012 10792 18018 10804
rect 18693 10795 18751 10801
rect 18012 10764 18644 10792
rect 18012 10752 18018 10764
rect 9522 10696 9904 10724
rect 9950 10684 9956 10736
rect 10008 10684 10014 10736
rect 10489 10727 10547 10733
rect 10489 10693 10501 10727
rect 10535 10724 10547 10727
rect 10535 10696 10640 10724
rect 10535 10693 10547 10696
rect 10489 10687 10547 10693
rect 10612 10668 10640 10696
rect 10686 10684 10692 10736
rect 10744 10684 10750 10736
rect 17862 10684 17868 10736
rect 17920 10684 17926 10736
rect 18616 10724 18644 10764
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 18782 10792 18788 10804
rect 18739 10764 18788 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 18782 10752 18788 10764
rect 18840 10792 18846 10804
rect 20530 10792 20536 10804
rect 18840 10764 20536 10792
rect 18840 10752 18846 10764
rect 20530 10752 20536 10764
rect 20588 10792 20594 10804
rect 20625 10795 20683 10801
rect 20625 10792 20637 10795
rect 20588 10764 20637 10792
rect 20588 10752 20594 10764
rect 20625 10761 20637 10764
rect 20671 10761 20683 10795
rect 20625 10755 20683 10761
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 22557 10795 22615 10801
rect 22557 10792 22569 10795
rect 22152 10764 22569 10792
rect 22152 10752 22158 10764
rect 22557 10761 22569 10764
rect 22603 10761 22615 10795
rect 22557 10755 22615 10761
rect 23014 10752 23020 10804
rect 23072 10792 23078 10804
rect 23109 10795 23167 10801
rect 23109 10792 23121 10795
rect 23072 10764 23121 10792
rect 23072 10752 23078 10764
rect 23109 10761 23121 10764
rect 23155 10761 23167 10795
rect 25498 10792 25504 10804
rect 23109 10755 23167 10761
rect 24228 10764 25504 10792
rect 18874 10724 18880 10736
rect 18616 10696 18880 10724
rect 18874 10684 18880 10696
rect 18932 10724 18938 10736
rect 18932 10696 18998 10724
rect 18932 10684 18938 10696
rect 20254 10684 20260 10736
rect 20312 10724 20318 10736
rect 20809 10727 20867 10733
rect 20312 10696 20668 10724
rect 20312 10684 20318 10696
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10656 4215 10659
rect 4614 10656 4620 10668
rect 4203 10628 4620 10656
rect 4203 10625 4215 10628
rect 4157 10619 4215 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10652 10628 12434 10656
rect 10652 10616 10658 10628
rect 1394 10548 1400 10600
rect 1452 10548 1458 10600
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 6822 10588 6828 10600
rect 5951 10560 6828 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7466 10548 7472 10600
rect 7524 10548 7530 10600
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10588 7987 10591
rect 9858 10588 9864 10600
rect 7975 10560 9864 10588
rect 7975 10557 7987 10560
rect 7929 10551 7987 10557
rect 5350 10480 5356 10532
rect 5408 10480 5414 10532
rect 7374 10520 7380 10532
rect 6564 10492 7380 10520
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6564 10461 6592 10492
rect 7374 10480 7380 10492
rect 7432 10520 7438 10532
rect 7852 10520 7880 10551
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10588 10287 10591
rect 11422 10588 11428 10600
rect 10275 10560 11428 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 12406 10588 12434 10628
rect 20438 10616 20444 10668
rect 20496 10616 20502 10668
rect 20533 10659 20591 10665
rect 20533 10625 20545 10659
rect 20579 10625 20591 10659
rect 20533 10619 20591 10625
rect 12894 10588 12900 10600
rect 12406 10560 12900 10588
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 16850 10548 16856 10600
rect 16908 10548 16914 10600
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 18322 10588 18328 10600
rect 17175 10560 18328 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 20162 10548 20168 10600
rect 20220 10548 20226 10600
rect 7432 10492 7880 10520
rect 7432 10480 7438 10492
rect 11698 10480 11704 10532
rect 11756 10520 11762 10532
rect 12989 10523 13047 10529
rect 12989 10520 13001 10523
rect 11756 10492 13001 10520
rect 11756 10480 11762 10492
rect 12989 10489 13001 10492
rect 13035 10489 13047 10523
rect 12989 10483 13047 10489
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 6328 10424 6561 10452
rect 6328 10412 6334 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6549 10415 6607 10421
rect 7285 10455 7343 10461
rect 7285 10421 7297 10455
rect 7331 10452 7343 10455
rect 7834 10452 7840 10464
rect 7331 10424 7840 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9640 10424 10333 10452
rect 9640 10412 9646 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 10502 10412 10508 10464
rect 10560 10412 10566 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 11204 10424 12265 10452
rect 11204 10412 11210 10424
rect 12253 10421 12265 10424
rect 12299 10421 12311 10455
rect 12253 10415 12311 10421
rect 18601 10455 18659 10461
rect 18601 10421 18613 10455
rect 18647 10452 18659 10455
rect 19150 10452 19156 10464
rect 18647 10424 19156 10452
rect 18647 10421 18659 10424
rect 18601 10415 18659 10421
rect 19150 10412 19156 10424
rect 19208 10412 19214 10464
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 20548 10452 20576 10619
rect 20640 10588 20668 10696
rect 20809 10693 20821 10727
rect 20855 10724 20867 10727
rect 21358 10724 21364 10736
rect 20855 10696 21364 10724
rect 20855 10693 20867 10696
rect 20809 10687 20867 10693
rect 21358 10684 21364 10696
rect 21416 10724 21422 10736
rect 21416 10696 22094 10724
rect 21416 10684 21422 10696
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 21177 10659 21235 10665
rect 21177 10625 21189 10659
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10656 21511 10659
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21499 10628 21833 10656
rect 21499 10625 21511 10628
rect 21453 10619 21511 10625
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 22066 10656 22094 10696
rect 24228 10668 24256 10764
rect 25498 10752 25504 10764
rect 25556 10752 25562 10804
rect 28074 10752 28080 10804
rect 28132 10752 28138 10804
rect 28166 10752 28172 10804
rect 28224 10792 28230 10804
rect 29086 10792 29092 10804
rect 28224 10764 29092 10792
rect 28224 10752 28230 10764
rect 29086 10752 29092 10764
rect 29144 10752 29150 10804
rect 29457 10795 29515 10801
rect 29457 10761 29469 10795
rect 29503 10792 29515 10795
rect 29546 10792 29552 10804
rect 29503 10764 29552 10792
rect 29503 10761 29515 10764
rect 29457 10755 29515 10761
rect 29546 10752 29552 10764
rect 29604 10752 29610 10804
rect 32122 10752 32128 10804
rect 32180 10792 32186 10804
rect 32180 10764 33732 10792
rect 32180 10752 32186 10764
rect 24854 10684 24860 10736
rect 24912 10684 24918 10736
rect 25590 10684 25596 10736
rect 25648 10684 25654 10736
rect 33704 10724 33732 10764
rect 34514 10752 34520 10804
rect 34572 10792 34578 10804
rect 34572 10764 35848 10792
rect 34572 10752 34578 10764
rect 34146 10724 34152 10736
rect 28460 10696 30420 10724
rect 33626 10696 34152 10724
rect 22373 10659 22431 10665
rect 22373 10656 22385 10659
rect 22066 10628 22385 10656
rect 21821 10619 21879 10625
rect 22373 10625 22385 10628
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 21192 10588 21220 10619
rect 20640 10560 21220 10588
rect 21174 10480 21180 10532
rect 21232 10520 21238 10532
rect 21284 10520 21312 10619
rect 22738 10616 22744 10668
rect 22796 10616 22802 10668
rect 22925 10659 22983 10665
rect 22925 10625 22937 10659
rect 22971 10656 22983 10659
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22971 10628 23029 10656
rect 22971 10625 22983 10628
rect 22925 10619 22983 10625
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23201 10659 23259 10665
rect 23201 10656 23213 10659
rect 23017 10619 23075 10625
rect 23124 10628 23213 10656
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22940 10588 22968 10619
rect 22244 10560 22968 10588
rect 22244 10548 22250 10560
rect 22922 10520 22928 10532
rect 21232 10492 21312 10520
rect 22756 10492 22928 10520
rect 21232 10480 21238 10492
rect 19576 10424 20576 10452
rect 20809 10455 20867 10461
rect 19576 10412 19582 10424
rect 20809 10421 20821 10455
rect 20855 10452 20867 10455
rect 22186 10452 22192 10464
rect 20855 10424 22192 10452
rect 20855 10421 20867 10424
rect 20809 10415 20867 10421
rect 22186 10412 22192 10424
rect 22244 10412 22250 10464
rect 22278 10412 22284 10464
rect 22336 10452 22342 10464
rect 22756 10461 22784 10492
rect 22922 10480 22928 10492
rect 22980 10520 22986 10532
rect 23124 10520 23152 10628
rect 23201 10625 23213 10628
rect 23247 10625 23259 10659
rect 23201 10619 23259 10625
rect 24210 10616 24216 10668
rect 24268 10616 24274 10668
rect 24489 10659 24547 10665
rect 24489 10625 24501 10659
rect 24535 10656 24547 10659
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 24535 10628 26341 10656
rect 24535 10625 24547 10628
rect 24489 10619 24547 10625
rect 26329 10625 26341 10628
rect 26375 10656 26387 10659
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 26375 10628 27169 10656
rect 26375 10625 26387 10628
rect 26329 10619 26387 10625
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10625 27307 10659
rect 27249 10619 27307 10625
rect 23842 10548 23848 10600
rect 23900 10588 23906 10600
rect 24121 10591 24179 10597
rect 24121 10588 24133 10591
rect 23900 10560 24133 10588
rect 23900 10548 23906 10560
rect 24121 10557 24133 10560
rect 24167 10557 24179 10591
rect 24121 10551 24179 10557
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10588 24639 10591
rect 24670 10588 24676 10600
rect 24627 10560 24676 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 25682 10548 25688 10600
rect 25740 10548 25746 10600
rect 26510 10548 26516 10600
rect 26568 10588 26574 10600
rect 27264 10588 27292 10619
rect 27338 10616 27344 10668
rect 27396 10616 27402 10668
rect 27522 10616 27528 10668
rect 27580 10616 27586 10668
rect 28460 10665 28488 10696
rect 28445 10659 28503 10665
rect 28445 10625 28457 10659
rect 28491 10625 28503 10659
rect 28445 10619 28503 10625
rect 28810 10616 28816 10668
rect 28868 10656 28874 10668
rect 28905 10659 28963 10665
rect 28905 10656 28917 10659
rect 28868 10628 28917 10656
rect 28868 10616 28874 10628
rect 28905 10625 28917 10628
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 28997 10659 29055 10665
rect 28997 10625 29009 10659
rect 29043 10625 29055 10659
rect 28997 10619 29055 10625
rect 26568 10560 27292 10588
rect 26568 10548 26574 10560
rect 22980 10492 23152 10520
rect 27264 10520 27292 10560
rect 27614 10548 27620 10600
rect 27672 10588 27678 10600
rect 28353 10591 28411 10597
rect 28353 10588 28365 10591
rect 27672 10560 28365 10588
rect 27672 10548 27678 10560
rect 28353 10557 28365 10560
rect 28399 10588 28411 10591
rect 28718 10588 28724 10600
rect 28399 10560 28724 10588
rect 28399 10557 28411 10560
rect 28353 10551 28411 10557
rect 28718 10548 28724 10560
rect 28776 10548 28782 10600
rect 29012 10520 29040 10619
rect 29086 10616 29092 10668
rect 29144 10616 29150 10668
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10625 29331 10659
rect 29273 10619 29331 10625
rect 29641 10659 29699 10665
rect 29641 10625 29653 10659
rect 29687 10656 29699 10659
rect 29730 10656 29736 10668
rect 29687 10628 29736 10656
rect 29687 10625 29699 10628
rect 29641 10619 29699 10625
rect 29288 10588 29316 10619
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 30392 10665 30420 10696
rect 34146 10684 34152 10696
rect 34204 10684 34210 10736
rect 34974 10684 34980 10736
rect 35032 10684 35038 10736
rect 35342 10684 35348 10736
rect 35400 10724 35406 10736
rect 35400 10696 35756 10724
rect 35400 10684 35406 10696
rect 30377 10659 30435 10665
rect 30377 10625 30389 10659
rect 30423 10656 30435 10659
rect 30650 10656 30656 10668
rect 30423 10628 30656 10656
rect 30423 10625 30435 10628
rect 30377 10619 30435 10625
rect 30650 10616 30656 10628
rect 30708 10616 30714 10668
rect 35728 10665 35756 10696
rect 35820 10665 35848 10764
rect 36170 10752 36176 10804
rect 36228 10752 36234 10804
rect 37461 10795 37519 10801
rect 37461 10761 37473 10795
rect 37507 10792 37519 10795
rect 38102 10792 38108 10804
rect 37507 10764 38108 10792
rect 37507 10761 37519 10764
rect 37461 10755 37519 10761
rect 38102 10752 38108 10764
rect 38160 10752 38166 10804
rect 38841 10795 38899 10801
rect 38841 10761 38853 10795
rect 38887 10792 38899 10795
rect 40770 10792 40776 10804
rect 38887 10764 40776 10792
rect 38887 10761 38899 10764
rect 38841 10755 38899 10761
rect 40770 10752 40776 10764
rect 40828 10752 40834 10804
rect 35986 10684 35992 10736
rect 36044 10684 36050 10736
rect 36081 10727 36139 10733
rect 36081 10693 36093 10727
rect 36127 10724 36139 10727
rect 36188 10724 36216 10752
rect 40678 10724 40684 10736
rect 36127 10696 36216 10724
rect 37476 10696 40684 10724
rect 36127 10693 36139 10696
rect 36081 10687 36139 10693
rect 35713 10659 35771 10665
rect 35713 10625 35725 10659
rect 35759 10625 35771 10659
rect 35713 10619 35771 10625
rect 35805 10659 35863 10665
rect 35805 10625 35817 10659
rect 35851 10625 35863 10659
rect 35805 10619 35863 10625
rect 36170 10616 36176 10668
rect 36228 10616 36234 10668
rect 36906 10616 36912 10668
rect 36964 10656 36970 10668
rect 37277 10659 37335 10665
rect 37277 10656 37289 10659
rect 36964 10628 37289 10656
rect 36964 10616 36970 10628
rect 37277 10625 37289 10628
rect 37323 10625 37335 10659
rect 37277 10619 37335 10625
rect 37366 10616 37372 10668
rect 37424 10656 37430 10668
rect 37476 10665 37504 10696
rect 40678 10684 40684 10696
rect 40736 10684 40742 10736
rect 37461 10659 37519 10665
rect 37461 10656 37473 10659
rect 37424 10628 37473 10656
rect 37424 10616 37430 10628
rect 37461 10625 37473 10628
rect 37507 10625 37519 10659
rect 37461 10619 37519 10625
rect 37645 10659 37703 10665
rect 37645 10625 37657 10659
rect 37691 10656 37703 10659
rect 37734 10656 37740 10668
rect 37691 10628 37740 10656
rect 37691 10625 37703 10628
rect 37645 10619 37703 10625
rect 37734 10616 37740 10628
rect 37792 10616 37798 10668
rect 37829 10659 37887 10665
rect 37829 10625 37841 10659
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 29825 10591 29883 10597
rect 29825 10588 29837 10591
rect 29288 10560 29837 10588
rect 29825 10557 29837 10560
rect 29871 10557 29883 10591
rect 29825 10551 29883 10557
rect 32125 10591 32183 10597
rect 32125 10557 32137 10591
rect 32171 10557 32183 10591
rect 32125 10551 32183 10557
rect 29086 10520 29092 10532
rect 27264 10492 29092 10520
rect 22980 10480 22986 10492
rect 29086 10480 29092 10492
rect 29144 10480 29150 10532
rect 22741 10455 22799 10461
rect 22741 10452 22753 10455
rect 22336 10424 22753 10452
rect 22336 10412 22342 10424
rect 22741 10421 22753 10424
rect 22787 10421 22799 10455
rect 22741 10415 22799 10421
rect 23934 10412 23940 10464
rect 23992 10412 23998 10464
rect 26970 10412 26976 10464
rect 27028 10412 27034 10464
rect 27338 10412 27344 10464
rect 27396 10452 27402 10464
rect 28166 10452 28172 10464
rect 27396 10424 28172 10452
rect 27396 10412 27402 10424
rect 28166 10412 28172 10424
rect 28224 10412 28230 10464
rect 28721 10455 28779 10461
rect 28721 10421 28733 10455
rect 28767 10452 28779 10455
rect 28902 10452 28908 10464
rect 28767 10424 28908 10452
rect 28767 10421 28779 10424
rect 28721 10415 28779 10421
rect 28902 10412 28908 10424
rect 28960 10412 28966 10464
rect 32140 10452 32168 10551
rect 32398 10548 32404 10600
rect 32456 10548 32462 10600
rect 34790 10548 34796 10600
rect 34848 10588 34854 10600
rect 35437 10591 35495 10597
rect 35437 10588 35449 10591
rect 34848 10560 35449 10588
rect 34848 10548 34854 10560
rect 35437 10557 35449 10560
rect 35483 10557 35495 10591
rect 37844 10588 37872 10619
rect 37918 10616 37924 10668
rect 37976 10616 37982 10668
rect 38010 10616 38016 10668
rect 38068 10616 38074 10668
rect 38289 10659 38347 10665
rect 38289 10625 38301 10659
rect 38335 10656 38347 10659
rect 38378 10656 38384 10668
rect 38335 10628 38384 10656
rect 38335 10625 38347 10628
rect 38289 10619 38347 10625
rect 38378 10616 38384 10628
rect 38436 10616 38442 10668
rect 38470 10616 38476 10668
rect 38528 10616 38534 10668
rect 38562 10616 38568 10668
rect 38620 10616 38626 10668
rect 38657 10659 38715 10665
rect 38657 10625 38669 10659
rect 38703 10656 38715 10659
rect 38838 10656 38844 10668
rect 38703 10628 38844 10656
rect 38703 10625 38715 10628
rect 38657 10619 38715 10625
rect 38838 10616 38844 10628
rect 38896 10616 38902 10668
rect 39577 10659 39635 10665
rect 39577 10625 39589 10659
rect 39623 10656 39635 10659
rect 41874 10656 41880 10668
rect 39623 10628 41880 10656
rect 39623 10625 39635 10628
rect 39577 10619 39635 10625
rect 37844 10560 37964 10588
rect 35437 10551 35495 10557
rect 32582 10452 32588 10464
rect 32140 10424 32588 10452
rect 32582 10412 32588 10424
rect 32640 10412 32646 10464
rect 33870 10412 33876 10464
rect 33928 10412 33934 10464
rect 33965 10455 34023 10461
rect 33965 10421 33977 10455
rect 34011 10452 34023 10455
rect 34146 10452 34152 10464
rect 34011 10424 34152 10452
rect 34011 10421 34023 10424
rect 33965 10415 34023 10421
rect 34146 10412 34152 10424
rect 34204 10412 34210 10464
rect 34698 10412 34704 10464
rect 34756 10452 34762 10464
rect 36357 10455 36415 10461
rect 36357 10452 36369 10455
rect 34756 10424 36369 10452
rect 34756 10412 34762 10424
rect 36357 10421 36369 10424
rect 36403 10421 36415 10455
rect 37936 10452 37964 10560
rect 38102 10548 38108 10600
rect 38160 10588 38166 10600
rect 39592 10588 39620 10619
rect 41874 10616 41880 10628
rect 41932 10616 41938 10668
rect 38160 10560 39620 10588
rect 38160 10548 38166 10560
rect 38197 10523 38255 10529
rect 38197 10489 38209 10523
rect 38243 10520 38255 10523
rect 39390 10520 39396 10532
rect 38243 10492 39396 10520
rect 38243 10489 38255 10492
rect 38197 10483 38255 10489
rect 39390 10480 39396 10492
rect 39448 10480 39454 10532
rect 38470 10452 38476 10464
rect 37936 10424 38476 10452
rect 36357 10415 36415 10421
rect 38470 10412 38476 10424
rect 38528 10412 38534 10464
rect 38930 10412 38936 10464
rect 38988 10452 38994 10464
rect 39485 10455 39543 10461
rect 39485 10452 39497 10455
rect 38988 10424 39497 10452
rect 38988 10412 38994 10424
rect 39485 10421 39497 10424
rect 39531 10421 39543 10455
rect 39485 10415 39543 10421
rect 1104 10362 42504 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 42504 10362
rect 1104 10288 42504 10310
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 3418 10248 3424 10260
rect 3375 10220 3424 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5592 10220 6009 10248
rect 5592 10208 5598 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 5997 10211 6055 10217
rect 6178 10208 6184 10260
rect 6236 10208 6242 10260
rect 7006 10248 7012 10260
rect 6288 10220 7012 10248
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 6288 10112 6316 10220
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7156 10220 7665 10248
rect 7156 10208 7162 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 7653 10211 7711 10217
rect 9858 10208 9864 10260
rect 9916 10208 9922 10260
rect 10413 10251 10471 10257
rect 10413 10217 10425 10251
rect 10459 10248 10471 10251
rect 10594 10248 10600 10260
rect 10459 10220 10600 10248
rect 10459 10217 10471 10220
rect 10413 10211 10471 10217
rect 10594 10208 10600 10220
rect 10652 10208 10658 10260
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 10735 10220 10824 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 6638 10140 6644 10192
rect 6696 10180 6702 10192
rect 6696 10152 7420 10180
rect 6696 10140 6702 10152
rect 2740 10084 3188 10112
rect 2740 10072 2746 10084
rect 3160 9976 3188 10084
rect 4632 10084 6316 10112
rect 6917 10115 6975 10121
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4632 10044 4660 10084
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7190 10112 7196 10124
rect 6963 10084 7196 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 7392 10112 7420 10152
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 9953 10183 10011 10189
rect 9953 10180 9965 10183
rect 7524 10152 9965 10180
rect 7524 10140 7530 10152
rect 7392 10084 7604 10112
rect 3283 10016 4660 10044
rect 4709 10047 4767 10053
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 5442 10044 5448 10056
rect 4755 10016 5448 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 6270 10044 6276 10056
rect 6227 10016 6276 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6365 10047 6423 10053
rect 6365 10013 6377 10047
rect 6411 10044 6423 10047
rect 7009 10047 7067 10053
rect 6411 10016 6960 10044
rect 6411 10013 6423 10016
rect 6365 10007 6423 10013
rect 6932 9988 6960 10016
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 7466 10044 7472 10056
rect 7055 10016 7472 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 3973 9979 4031 9985
rect 3973 9976 3985 9979
rect 3160 9948 3985 9976
rect 3973 9945 3985 9948
rect 4019 9976 4031 9979
rect 4614 9976 4620 9988
rect 4019 9948 4620 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 6638 9936 6644 9988
rect 6696 9936 6702 9988
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 7576 9976 7604 10084
rect 7944 10053 7972 10152
rect 9953 10149 9965 10152
rect 9999 10149 10011 10183
rect 9953 10143 10011 10149
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 9217 10115 9275 10121
rect 9217 10112 9229 10115
rect 8076 10084 9229 10112
rect 8076 10072 8082 10084
rect 9217 10081 9229 10084
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 9493 10115 9551 10121
rect 9493 10112 9505 10115
rect 9364 10084 9505 10112
rect 9364 10072 9370 10084
rect 9493 10081 9505 10084
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9702 10115 9760 10121
rect 9702 10081 9714 10115
rect 9748 10112 9760 10115
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 9748 10084 10333 10112
rect 9748 10081 9760 10084
rect 9702 10075 9760 10081
rect 10321 10081 10333 10084
rect 10367 10112 10379 10115
rect 10796 10112 10824 10220
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 12952 10220 13369 10248
rect 12952 10208 12958 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 13357 10211 13415 10217
rect 18322 10208 18328 10260
rect 18380 10208 18386 10260
rect 19702 10248 19708 10260
rect 18524 10220 19708 10248
rect 10873 10183 10931 10189
rect 10873 10149 10885 10183
rect 10919 10149 10931 10183
rect 10873 10143 10931 10149
rect 10367 10084 10824 10112
rect 10888 10112 10916 10143
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10888 10084 11253 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 7632 9979 7690 9985
rect 7632 9976 7644 9979
rect 7024 9948 7512 9976
rect 7576 9948 7644 9976
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9908 5043 9911
rect 5258 9908 5264 9920
rect 5031 9880 5264 9908
rect 5031 9877 5043 9880
rect 4985 9871 5043 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 6546 9868 6552 9920
rect 6604 9908 6610 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6604 9880 6745 9908
rect 6604 9868 6610 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 7024 9908 7052 9948
rect 6880 9880 7052 9908
rect 6880 9868 6886 9880
rect 7374 9868 7380 9920
rect 7432 9868 7438 9920
rect 7484 9917 7512 9948
rect 7632 9945 7644 9948
rect 7678 9945 7690 9979
rect 7632 9939 7690 9945
rect 7834 9936 7840 9988
rect 7892 9936 7898 9988
rect 10152 9976 10180 10007
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10502 9976 10508 9988
rect 10152 9948 10508 9976
rect 10502 9936 10508 9948
rect 10560 9936 10566 9988
rect 7469 9911 7527 9917
rect 7469 9877 7481 9911
rect 7515 9877 7527 9911
rect 7469 9871 7527 9877
rect 8018 9868 8024 9920
rect 8076 9868 8082 9920
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 10705 9911 10763 9917
rect 10705 9908 10717 9911
rect 9824 9880 10717 9908
rect 9824 9868 9830 9880
rect 10705 9877 10717 9880
rect 10751 9877 10763 9911
rect 10796 9908 10824 10084
rect 11241 10081 11253 10084
rect 11287 10112 11299 10115
rect 11330 10112 11336 10124
rect 11287 10084 11336 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11563 10084 11897 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12032 10084 18092 10112
rect 12032 10072 12038 10084
rect 11146 10004 11152 10056
rect 11204 10004 11210 10056
rect 11422 10004 11428 10056
rect 11480 10044 11486 10056
rect 11609 10047 11667 10053
rect 11609 10044 11621 10047
rect 11480 10016 11621 10044
rect 11480 10004 11486 10016
rect 11609 10013 11621 10016
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 17954 9976 17960 9988
rect 13110 9948 17960 9976
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 18064 9976 18092 10084
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18524 10121 18552 10220
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 19981 10251 20039 10257
rect 19981 10217 19993 10251
rect 20027 10248 20039 10251
rect 20162 10248 20168 10260
rect 20027 10220 20168 10248
rect 20027 10217 20039 10220
rect 19981 10211 20039 10217
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 22002 10248 22008 10260
rect 20266 10220 22008 10248
rect 20266 10180 20294 10220
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 23106 10208 23112 10260
rect 23164 10248 23170 10260
rect 23293 10251 23351 10257
rect 23293 10248 23305 10251
rect 23164 10220 23305 10248
rect 23164 10208 23170 10220
rect 23293 10217 23305 10220
rect 23339 10217 23351 10251
rect 23293 10211 23351 10217
rect 24210 10208 24216 10260
rect 24268 10208 24274 10260
rect 24857 10251 24915 10257
rect 24857 10217 24869 10251
rect 24903 10248 24915 10251
rect 25866 10248 25872 10260
rect 24903 10220 25872 10248
rect 24903 10217 24915 10220
rect 24857 10211 24915 10217
rect 23124 10180 23152 10208
rect 24872 10180 24900 10211
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 26347 10251 26405 10257
rect 26347 10217 26359 10251
rect 26393 10248 26405 10251
rect 26970 10248 26976 10260
rect 26393 10220 26976 10248
rect 26393 10217 26405 10220
rect 26347 10211 26405 10217
rect 26970 10208 26976 10220
rect 27028 10208 27034 10260
rect 27890 10208 27896 10260
rect 27948 10248 27954 10260
rect 28994 10248 29000 10260
rect 27948 10220 29000 10248
rect 27948 10208 27954 10220
rect 28994 10208 29000 10220
rect 29052 10248 29058 10260
rect 29362 10248 29368 10260
rect 29052 10220 29368 10248
rect 29052 10208 29058 10220
rect 29362 10208 29368 10220
rect 29420 10208 29426 10260
rect 30650 10208 30656 10260
rect 30708 10248 30714 10260
rect 31018 10248 31024 10260
rect 30708 10220 31024 10248
rect 30708 10208 30714 10220
rect 31018 10208 31024 10220
rect 31076 10208 31082 10260
rect 32125 10251 32183 10257
rect 32125 10217 32137 10251
rect 32171 10248 32183 10251
rect 32398 10248 32404 10260
rect 32171 10220 32404 10248
rect 32171 10217 32183 10220
rect 32125 10211 32183 10217
rect 32398 10208 32404 10220
rect 32456 10208 32462 10260
rect 32508 10220 37688 10248
rect 19168 10152 20294 10180
rect 22204 10152 23152 10180
rect 23860 10152 24900 10180
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18196 10084 18521 10112
rect 18196 10072 18202 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 19168 10112 19196 10152
rect 18509 10075 18567 10081
rect 18800 10084 19196 10112
rect 18598 10004 18604 10056
rect 18656 10004 18662 10056
rect 18800 9976 18828 10084
rect 19242 10072 19248 10124
rect 19300 10112 19306 10124
rect 19337 10115 19395 10121
rect 19337 10112 19349 10115
rect 19300 10084 19349 10112
rect 19300 10072 19306 10084
rect 19337 10081 19349 10084
rect 19383 10081 19395 10115
rect 19337 10075 19395 10081
rect 18877 10047 18935 10053
rect 18877 10013 18889 10047
rect 18923 10044 18935 10047
rect 19889 10047 19947 10053
rect 19889 10044 19901 10047
rect 18923 10016 19901 10044
rect 18923 10013 18935 10016
rect 18877 10007 18935 10013
rect 19889 10013 19901 10016
rect 19935 10044 19947 10047
rect 20165 10047 20223 10053
rect 20165 10044 20177 10047
rect 19935 10016 20177 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20165 10013 20177 10016
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 20254 10004 20260 10056
rect 20312 10004 20318 10056
rect 20530 10004 20536 10056
rect 20588 10004 20594 10056
rect 22204 10053 22232 10152
rect 23109 10115 23167 10121
rect 23109 10081 23121 10115
rect 23155 10112 23167 10115
rect 23750 10112 23756 10124
rect 23155 10084 23756 10112
rect 23155 10081 23167 10084
rect 23109 10075 23167 10081
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22738 10004 22744 10056
rect 22796 10004 22802 10056
rect 22922 10004 22928 10056
rect 22980 10004 22986 10056
rect 23860 10053 23888 10152
rect 28810 10140 28816 10192
rect 28868 10180 28874 10192
rect 29549 10183 29607 10189
rect 29549 10180 29561 10183
rect 28868 10152 29561 10180
rect 28868 10140 28874 10152
rect 29549 10149 29561 10152
rect 29595 10149 29607 10183
rect 29549 10143 29607 10149
rect 31205 10183 31263 10189
rect 31205 10149 31217 10183
rect 31251 10180 31263 10183
rect 31478 10180 31484 10192
rect 31251 10152 31484 10180
rect 31251 10149 31263 10152
rect 31205 10143 31263 10149
rect 31478 10140 31484 10152
rect 31536 10140 31542 10192
rect 32508 10180 32536 10220
rect 31588 10152 32536 10180
rect 34333 10183 34391 10189
rect 23937 10115 23995 10121
rect 23937 10081 23949 10115
rect 23983 10112 23995 10115
rect 24118 10112 24124 10124
rect 23983 10084 24124 10112
rect 23983 10081 23995 10084
rect 23937 10075 23995 10081
rect 24118 10072 24124 10084
rect 24176 10072 24182 10124
rect 24210 10072 24216 10124
rect 24268 10112 24274 10124
rect 24394 10112 24400 10124
rect 24268 10084 24400 10112
rect 24268 10072 24274 10084
rect 24394 10072 24400 10084
rect 24452 10112 24458 10124
rect 24452 10084 25268 10112
rect 24452 10072 24458 10084
rect 23477 10047 23535 10053
rect 23477 10013 23489 10047
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10013 23903 10047
rect 25240 10030 25268 10084
rect 25774 10072 25780 10124
rect 25832 10112 25838 10124
rect 26605 10115 26663 10121
rect 26605 10112 26617 10115
rect 25832 10084 26617 10112
rect 25832 10072 25838 10084
rect 26605 10081 26617 10084
rect 26651 10112 26663 10115
rect 27157 10115 27215 10121
rect 27157 10112 27169 10115
rect 26651 10084 27169 10112
rect 26651 10081 26663 10084
rect 26605 10075 26663 10081
rect 27157 10081 27169 10084
rect 27203 10081 27215 10115
rect 27157 10075 27215 10081
rect 28905 10115 28963 10121
rect 28905 10081 28917 10115
rect 28951 10112 28963 10115
rect 30101 10115 30159 10121
rect 30101 10112 30113 10115
rect 28951 10084 30113 10112
rect 28951 10081 28963 10084
rect 28905 10075 28963 10081
rect 30101 10081 30113 10084
rect 30147 10081 30159 10115
rect 31588 10112 31616 10152
rect 34333 10149 34345 10183
rect 34379 10180 34391 10183
rect 34698 10180 34704 10192
rect 34379 10152 34704 10180
rect 34379 10149 34391 10152
rect 34333 10143 34391 10149
rect 34698 10140 34704 10152
rect 34756 10140 34762 10192
rect 37185 10183 37243 10189
rect 36832 10152 37136 10180
rect 30101 10075 30159 10081
rect 30208 10084 31616 10112
rect 32309 10115 32367 10121
rect 23845 10007 23903 10013
rect 18064 9948 18828 9976
rect 18969 9979 19027 9985
rect 18969 9945 18981 9979
rect 19015 9945 19027 9979
rect 18969 9939 19027 9945
rect 13538 9908 13544 9920
rect 10796 9880 13544 9908
rect 10705 9871 10763 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 17972 9908 18000 9936
rect 18230 9908 18236 9920
rect 17972 9880 18236 9908
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18984 9908 19012 9939
rect 19610 9936 19616 9988
rect 19668 9976 19674 9988
rect 20349 9979 20407 9985
rect 20349 9976 20361 9979
rect 19668 9948 20361 9976
rect 19668 9936 19674 9948
rect 20349 9945 20361 9948
rect 20395 9976 20407 9979
rect 21174 9976 21180 9988
rect 20395 9948 21180 9976
rect 20395 9945 20407 9948
rect 20349 9939 20407 9945
rect 21174 9936 21180 9948
rect 21232 9936 21238 9988
rect 19794 9908 19800 9920
rect 18984 9880 19800 9908
rect 19794 9868 19800 9880
rect 19852 9908 19858 9920
rect 21266 9908 21272 9920
rect 19852 9880 21272 9908
rect 19852 9868 19858 9880
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 23492 9908 23520 10007
rect 28718 10004 28724 10056
rect 28776 10044 28782 10056
rect 29178 10044 29184 10056
rect 28776 10016 29184 10044
rect 28776 10004 28782 10016
rect 29178 10004 29184 10016
rect 29236 10004 29242 10056
rect 29270 10004 29276 10056
rect 29328 10004 29334 10056
rect 26418 9936 26424 9988
rect 26476 9976 26482 9988
rect 27338 9976 27344 9988
rect 26476 9948 27344 9976
rect 26476 9936 26482 9948
rect 27338 9936 27344 9948
rect 27396 9936 27402 9988
rect 27433 9979 27491 9985
rect 27433 9945 27445 9979
rect 27479 9976 27491 9979
rect 27706 9976 27712 9988
rect 27479 9948 27712 9976
rect 27479 9945 27491 9948
rect 27433 9939 27491 9945
rect 27706 9936 27712 9948
rect 27764 9936 27770 9988
rect 27890 9936 27896 9988
rect 27948 9936 27954 9988
rect 30208 9976 30236 10084
rect 32309 10081 32321 10115
rect 32355 10112 32367 10115
rect 33778 10112 33784 10124
rect 32355 10084 33784 10112
rect 32355 10081 32367 10084
rect 32309 10075 32367 10081
rect 30929 10047 30987 10053
rect 30929 10044 30941 10047
rect 30684 10016 30941 10044
rect 28966 9948 30236 9976
rect 28966 9908 28994 9948
rect 30466 9936 30472 9988
rect 30524 9936 30530 9988
rect 23492 9880 28994 9908
rect 29086 9868 29092 9920
rect 29144 9868 29150 9920
rect 29178 9868 29184 9920
rect 29236 9908 29242 9920
rect 30684 9917 30712 10016
rect 30929 10013 30941 10016
rect 30975 10013 30987 10047
rect 30929 10007 30987 10013
rect 31018 10004 31024 10056
rect 31076 10004 31082 10056
rect 31573 10047 31631 10053
rect 31573 10044 31585 10047
rect 31128 10016 31585 10044
rect 31128 9976 31156 10016
rect 31573 10013 31585 10016
rect 31619 10044 31631 10047
rect 31662 10044 31668 10056
rect 31619 10016 31668 10044
rect 31619 10013 31631 10016
rect 31573 10007 31631 10013
rect 31662 10004 31668 10016
rect 31720 10004 31726 10056
rect 31754 10004 31760 10056
rect 31812 10004 31818 10056
rect 30852 9948 31156 9976
rect 30852 9917 30880 9948
rect 31202 9936 31208 9988
rect 31260 9936 31266 9988
rect 32324 9976 32352 10075
rect 33778 10072 33784 10084
rect 33836 10072 33842 10124
rect 33870 10072 33876 10124
rect 33928 10072 33934 10124
rect 36832 10112 36860 10152
rect 34256 10084 36860 10112
rect 32401 10047 32459 10053
rect 32401 10013 32413 10047
rect 32447 10044 32459 10047
rect 32490 10044 32496 10056
rect 32447 10016 32496 10044
rect 32447 10013 32459 10016
rect 32401 10007 32459 10013
rect 32490 10004 32496 10016
rect 32548 10004 32554 10056
rect 32677 10047 32735 10053
rect 32677 10013 32689 10047
rect 32723 10044 32735 10047
rect 33318 10044 33324 10056
rect 32723 10016 33324 10044
rect 32723 10013 32735 10016
rect 32677 10007 32735 10013
rect 33318 10004 33324 10016
rect 33376 10004 33382 10056
rect 34057 10047 34115 10053
rect 34057 10044 34069 10047
rect 33888 10016 34069 10044
rect 33888 9988 33916 10016
rect 34057 10013 34069 10016
rect 34103 10013 34115 10047
rect 34057 10007 34115 10013
rect 31312 9948 32352 9976
rect 30669 9911 30727 9917
rect 30669 9908 30681 9911
rect 29236 9880 30681 9908
rect 29236 9868 29242 9880
rect 30669 9877 30681 9880
rect 30715 9877 30727 9911
rect 30669 9871 30727 9877
rect 30837 9911 30895 9917
rect 30837 9877 30849 9911
rect 30883 9877 30895 9911
rect 30837 9871 30895 9877
rect 31110 9868 31116 9920
rect 31168 9908 31174 9920
rect 31312 9908 31340 9948
rect 32766 9936 32772 9988
rect 32824 9936 32830 9988
rect 33870 9936 33876 9988
rect 33928 9936 33934 9988
rect 34256 9976 34284 10084
rect 36906 10072 36912 10124
rect 36964 10072 36970 10124
rect 37108 10112 37136 10152
rect 37185 10149 37197 10183
rect 37231 10180 37243 10183
rect 37550 10180 37556 10192
rect 37231 10152 37556 10180
rect 37231 10149 37243 10152
rect 37185 10143 37243 10149
rect 37550 10140 37556 10152
rect 37608 10140 37614 10192
rect 37660 10180 37688 10220
rect 37734 10208 37740 10260
rect 37792 10248 37798 10260
rect 39853 10251 39911 10257
rect 39853 10248 39865 10251
rect 37792 10220 39865 10248
rect 37792 10208 37798 10220
rect 39853 10217 39865 10220
rect 39899 10217 39911 10251
rect 41782 10248 41788 10260
rect 39853 10211 39911 10217
rect 40788 10220 41788 10248
rect 38102 10180 38108 10192
rect 37660 10152 38108 10180
rect 38102 10140 38108 10152
rect 38160 10140 38166 10192
rect 38562 10140 38568 10192
rect 38620 10180 38626 10192
rect 40310 10180 40316 10192
rect 38620 10152 40316 10180
rect 38620 10140 38626 10152
rect 40310 10140 40316 10152
rect 40368 10140 40374 10192
rect 37829 10115 37887 10121
rect 37108 10084 37780 10112
rect 36817 10047 36875 10053
rect 36817 10013 36829 10047
rect 36863 10044 36875 10047
rect 37366 10044 37372 10056
rect 36863 10016 37372 10044
rect 36863 10013 36875 10016
rect 36817 10007 36875 10013
rect 37366 10004 37372 10016
rect 37424 10004 37430 10056
rect 37458 10004 37464 10056
rect 37516 10004 37522 10056
rect 37553 10047 37611 10053
rect 37553 10013 37565 10047
rect 37599 10044 37611 10047
rect 37642 10044 37648 10056
rect 37599 10016 37648 10044
rect 37599 10013 37611 10016
rect 37553 10007 37611 10013
rect 37642 10004 37648 10016
rect 37700 10004 37706 10056
rect 37752 10044 37780 10084
rect 37829 10081 37841 10115
rect 37875 10112 37887 10115
rect 38010 10112 38016 10124
rect 37875 10084 38016 10112
rect 37875 10081 37887 10084
rect 37829 10075 37887 10081
rect 38010 10072 38016 10084
rect 38068 10112 38074 10124
rect 38473 10115 38531 10121
rect 38473 10112 38485 10115
rect 38068 10084 38485 10112
rect 38068 10072 38074 10084
rect 38473 10081 38485 10084
rect 38519 10081 38531 10115
rect 40497 10115 40555 10121
rect 38473 10075 38531 10081
rect 38948 10084 39160 10112
rect 38948 10056 38976 10084
rect 38930 10044 38936 10056
rect 37752 10016 38936 10044
rect 38930 10004 38936 10016
rect 38988 10004 38994 10056
rect 39022 10004 39028 10056
rect 39080 10004 39086 10056
rect 39132 10044 39160 10084
rect 40497 10081 40509 10115
rect 40543 10112 40555 10115
rect 40678 10112 40684 10124
rect 40543 10084 40684 10112
rect 40543 10081 40555 10084
rect 40497 10075 40555 10081
rect 40678 10072 40684 10084
rect 40736 10072 40742 10124
rect 40586 10044 40592 10056
rect 39132 10016 40592 10044
rect 40586 10004 40592 10016
rect 40644 10004 40650 10056
rect 34072 9948 34284 9976
rect 31168 9880 31340 9908
rect 31665 9911 31723 9917
rect 31168 9868 31174 9880
rect 31665 9877 31677 9911
rect 31711 9908 31723 9911
rect 31938 9908 31944 9920
rect 31711 9880 31944 9908
rect 31711 9877 31723 9880
rect 31665 9871 31723 9877
rect 31938 9868 31944 9880
rect 31996 9868 32002 9920
rect 32306 9868 32312 9920
rect 32364 9908 32370 9920
rect 34072 9908 34100 9948
rect 34330 9936 34336 9988
rect 34388 9936 34394 9988
rect 37921 9979 37979 9985
rect 37921 9945 37933 9979
rect 37967 9976 37979 9979
rect 38194 9976 38200 9988
rect 37967 9948 38200 9976
rect 37967 9945 37979 9948
rect 37921 9939 37979 9945
rect 32364 9880 34100 9908
rect 32364 9868 32370 9880
rect 34146 9868 34152 9920
rect 34204 9868 34210 9920
rect 37277 9911 37335 9917
rect 37277 9877 37289 9911
rect 37323 9908 37335 9911
rect 37550 9908 37556 9920
rect 37323 9880 37556 9908
rect 37323 9877 37335 9880
rect 37277 9871 37335 9877
rect 37550 9868 37556 9880
rect 37608 9868 37614 9920
rect 37642 9868 37648 9920
rect 37700 9908 37706 9920
rect 37936 9908 37964 9939
rect 38194 9936 38200 9948
rect 38252 9936 38258 9988
rect 39298 9936 39304 9988
rect 39356 9976 39362 9988
rect 40788 9976 40816 10220
rect 41782 10208 41788 10220
rect 41840 10208 41846 10260
rect 39356 9948 40816 9976
rect 39356 9936 39362 9948
rect 37700 9880 37964 9908
rect 37700 9868 37706 9880
rect 38930 9868 38936 9920
rect 38988 9908 38994 9920
rect 39393 9911 39451 9917
rect 39393 9908 39405 9911
rect 38988 9880 39405 9908
rect 38988 9868 38994 9880
rect 39393 9877 39405 9880
rect 39439 9908 39451 9911
rect 39850 9908 39856 9920
rect 39439 9880 39856 9908
rect 39439 9877 39451 9880
rect 39393 9871 39451 9877
rect 39850 9868 39856 9880
rect 39908 9868 39914 9920
rect 40788 9917 40816 9948
rect 40773 9911 40831 9917
rect 40773 9877 40785 9911
rect 40819 9877 40831 9911
rect 40773 9871 40831 9877
rect 1104 9818 42504 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 42504 9818
rect 1104 9744 42504 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 4893 9707 4951 9713
rect 3476 9676 4476 9704
rect 3476 9664 3482 9676
rect 3234 9596 3240 9648
rect 3292 9636 3298 9648
rect 3292 9608 3634 9636
rect 3292 9596 3298 9608
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 2682 9568 2688 9580
rect 1452 9540 2688 9568
rect 1452 9528 1458 9540
rect 2682 9528 2688 9540
rect 2740 9568 2746 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2740 9540 2881 9568
rect 2740 9528 2746 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 4448 9568 4476 9676
rect 4893 9673 4905 9707
rect 4939 9673 4951 9707
rect 4893 9667 4951 9673
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6638 9704 6644 9716
rect 5859 9676 6644 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 4908 9636 4936 9667
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 7098 9664 7104 9716
rect 7156 9664 7162 9716
rect 7834 9704 7840 9716
rect 7208 9676 7840 9704
rect 5442 9636 5448 9648
rect 4908 9608 5448 9636
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 7208 9636 7236 9676
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 13265 9707 13323 9713
rect 13265 9673 13277 9707
rect 13311 9704 13323 9707
rect 13538 9704 13544 9716
rect 13311 9676 13544 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 25133 9707 25191 9713
rect 25133 9673 25145 9707
rect 25179 9704 25191 9707
rect 25682 9704 25688 9716
rect 25179 9676 25688 9704
rect 25179 9673 25191 9676
rect 25133 9667 25191 9673
rect 25682 9664 25688 9676
rect 25740 9664 25746 9716
rect 25866 9664 25872 9716
rect 25924 9704 25930 9716
rect 27157 9707 27215 9713
rect 27157 9704 27169 9707
rect 25924 9676 27169 9704
rect 25924 9664 25930 9676
rect 6052 9608 7236 9636
rect 6052 9596 6058 9608
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 8018 9636 8024 9648
rect 7616 9608 8024 9636
rect 7616 9596 7622 9608
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 10689 9639 10747 9645
rect 10689 9636 10701 9639
rect 10060 9608 10701 9636
rect 4834 9571 4892 9577
rect 4834 9568 4846 9571
rect 4448 9540 4846 9568
rect 2869 9531 2927 9537
rect 4834 9537 4846 9540
rect 4880 9568 4892 9571
rect 4880 9540 5212 9568
rect 4880 9537 4892 9540
rect 4834 9531 4892 9537
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3191 9472 4752 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 4724 9441 4752 9472
rect 4709 9435 4767 9441
rect 4709 9401 4721 9435
rect 4755 9401 4767 9435
rect 5184 9432 5212 9540
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 5626 9528 5632 9580
rect 5684 9528 5690 9580
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9537 5779 9571
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 5721 9531 5779 9537
rect 5920 9540 6745 9568
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5399 9472 5457 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5736 9500 5764 9531
rect 5445 9463 5503 9469
rect 5552 9472 5764 9500
rect 5552 9432 5580 9472
rect 5184 9404 5580 9432
rect 4709 9395 4767 9401
rect 5626 9392 5632 9444
rect 5684 9432 5690 9444
rect 5920 9432 5948 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7926 9568 7932 9580
rect 7791 9540 7932 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 6546 9460 6552 9512
rect 6604 9460 6610 9512
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 7484 9500 7512 9531
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 10060 9577 10088 9608
rect 10689 9605 10701 9608
rect 10735 9605 10747 9639
rect 11698 9636 11704 9648
rect 10689 9599 10747 9605
rect 10980 9608 11704 9636
rect 10045 9571 10103 9577
rect 10045 9537 10057 9571
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10980 9568 11008 9608
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 12434 9596 12440 9648
rect 12492 9596 12498 9648
rect 23661 9639 23719 9645
rect 23661 9605 23673 9639
rect 23707 9636 23719 9639
rect 23934 9636 23940 9648
rect 23707 9608 23940 9636
rect 23707 9605 23719 9608
rect 23661 9599 23719 9605
rect 23934 9596 23940 9608
rect 23992 9596 23998 9648
rect 24210 9596 24216 9648
rect 24268 9596 24274 9648
rect 26344 9636 26372 9676
rect 27157 9673 27169 9676
rect 27203 9704 27215 9707
rect 27522 9704 27528 9716
rect 27203 9676 27528 9704
rect 27203 9673 27215 9676
rect 27157 9667 27215 9673
rect 27522 9664 27528 9676
rect 27580 9664 27586 9716
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 27893 9707 27951 9713
rect 27893 9704 27905 9707
rect 27764 9676 27905 9704
rect 27764 9664 27770 9676
rect 27893 9673 27905 9676
rect 27939 9673 27951 9707
rect 27893 9667 27951 9673
rect 28258 9664 28264 9716
rect 28316 9704 28322 9716
rect 30377 9707 30435 9713
rect 28316 9676 30236 9704
rect 28316 9664 28322 9676
rect 26160 9608 26372 9636
rect 26973 9639 27031 9645
rect 10643 9540 11008 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 6696 9472 7512 9500
rect 6696 9460 6702 9472
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 9953 9503 10011 9509
rect 9953 9500 9965 9503
rect 9824 9472 9965 9500
rect 9824 9460 9830 9472
rect 9953 9469 9965 9472
rect 9999 9500 10011 9503
rect 10336 9500 10364 9531
rect 9999 9472 10364 9500
rect 10428 9500 10456 9531
rect 20898 9528 20904 9580
rect 20956 9568 20962 9580
rect 22738 9568 22744 9580
rect 20956 9540 22744 9568
rect 20956 9528 20962 9540
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 10502 9500 10508 9512
rect 10428 9472 10508 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10502 9460 10508 9472
rect 10560 9500 10566 9512
rect 10962 9500 10968 9512
rect 10560 9472 10968 9500
rect 10560 9460 10566 9472
rect 10962 9460 10968 9472
rect 11020 9500 11026 9512
rect 11241 9503 11299 9509
rect 11241 9500 11253 9503
rect 11020 9472 11253 9500
rect 11020 9460 11026 9472
rect 11241 9469 11253 9472
rect 11287 9469 11299 9503
rect 11241 9463 11299 9469
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11480 9472 11529 9500
rect 11480 9460 11486 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 5684 9404 5948 9432
rect 10597 9435 10655 9441
rect 5684 9392 5690 9404
rect 10597 9401 10609 9435
rect 10643 9432 10655 9435
rect 11146 9432 11152 9444
rect 10643 9404 11152 9432
rect 10643 9401 10655 9404
rect 10597 9395 10655 9401
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 5534 9364 5540 9376
rect 4663 9336 5540 9364
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 7653 9367 7711 9373
rect 7653 9333 7665 9367
rect 7699 9364 7711 9367
rect 8294 9364 8300 9376
rect 7699 9336 8300 9364
rect 7699 9333 7711 9336
rect 7653 9327 7711 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9674 9324 9680 9376
rect 9732 9324 9738 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 11532 9364 11560 9463
rect 11790 9460 11796 9512
rect 11848 9460 11854 9512
rect 21818 9460 21824 9512
rect 21876 9460 21882 9512
rect 22833 9503 22891 9509
rect 22833 9469 22845 9503
rect 22879 9500 22891 9503
rect 22922 9500 22928 9512
rect 22879 9472 22928 9500
rect 22879 9469 22891 9472
rect 22833 9463 22891 9469
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23382 9460 23388 9512
rect 23440 9460 23446 9512
rect 26160 9432 26188 9608
rect 26973 9605 26985 9639
rect 27019 9605 27031 9639
rect 26973 9599 27031 9605
rect 26512 9571 26570 9577
rect 26512 9537 26524 9571
rect 26558 9548 26570 9571
rect 26602 9548 26608 9580
rect 26558 9537 26608 9548
rect 26512 9531 26608 9537
rect 26528 9528 26608 9531
rect 26660 9528 26666 9580
rect 26988 9569 27016 9599
rect 27338 9596 27344 9648
rect 27396 9596 27402 9648
rect 28074 9596 28080 9648
rect 28132 9636 28138 9648
rect 28445 9639 28503 9645
rect 28132 9608 28212 9636
rect 28132 9596 28138 9608
rect 26988 9541 27108 9569
rect 26528 9520 26648 9528
rect 27080 9512 27108 9541
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 28184 9577 28212 9608
rect 28445 9605 28457 9639
rect 28491 9636 28503 9639
rect 28810 9636 28816 9648
rect 28491 9608 28816 9636
rect 28491 9605 28503 9608
rect 28445 9599 28503 9605
rect 28810 9596 28816 9608
rect 28868 9596 28874 9648
rect 28902 9596 28908 9648
rect 28960 9596 28966 9648
rect 29362 9596 29368 9648
rect 29420 9596 29426 9648
rect 30208 9636 30236 9676
rect 30377 9673 30389 9707
rect 30423 9704 30435 9707
rect 30558 9704 30564 9716
rect 30423 9676 30564 9704
rect 30423 9673 30435 9676
rect 30377 9667 30435 9673
rect 30558 9664 30564 9676
rect 30616 9664 30622 9716
rect 33870 9704 33876 9716
rect 32876 9676 33876 9704
rect 30653 9639 30711 9645
rect 30208 9608 30512 9636
rect 27249 9571 27307 9577
rect 27249 9568 27261 9571
rect 27212 9540 27261 9568
rect 27212 9528 27218 9540
rect 27249 9537 27261 9540
rect 27295 9537 27307 9571
rect 27249 9531 27307 9537
rect 28169 9571 28227 9577
rect 28169 9537 28181 9571
rect 28215 9537 28227 9571
rect 30484 9568 30512 9608
rect 30653 9605 30665 9639
rect 30699 9636 30711 9639
rect 30742 9636 30748 9648
rect 30699 9608 30748 9636
rect 30699 9605 30711 9608
rect 30653 9599 30711 9605
rect 30742 9596 30748 9608
rect 30800 9636 30806 9648
rect 31570 9636 31576 9648
rect 30800 9608 31576 9636
rect 30800 9596 30806 9608
rect 31570 9596 31576 9608
rect 31628 9596 31634 9648
rect 31662 9596 31668 9648
rect 31720 9596 31726 9648
rect 31938 9596 31944 9648
rect 31996 9636 32002 9648
rect 32125 9639 32183 9645
rect 32125 9636 32137 9639
rect 31996 9608 32137 9636
rect 31996 9596 32002 9608
rect 32125 9605 32137 9608
rect 32171 9605 32183 9639
rect 32125 9599 32183 9605
rect 32309 9639 32367 9645
rect 32309 9605 32321 9639
rect 32355 9636 32367 9639
rect 32876 9636 32904 9676
rect 33870 9664 33876 9676
rect 33928 9704 33934 9716
rect 34441 9707 34499 9713
rect 34441 9704 34453 9707
rect 33928 9676 34453 9704
rect 33928 9664 33934 9676
rect 34441 9673 34453 9676
rect 34487 9673 34499 9707
rect 34441 9667 34499 9673
rect 35897 9707 35955 9713
rect 35897 9673 35909 9707
rect 35943 9704 35955 9707
rect 36078 9704 36084 9716
rect 35943 9676 36084 9704
rect 35943 9673 35955 9676
rect 35897 9667 35955 9673
rect 36078 9664 36084 9676
rect 36136 9664 36142 9716
rect 36449 9707 36507 9713
rect 36449 9673 36461 9707
rect 36495 9704 36507 9707
rect 36906 9704 36912 9716
rect 36495 9676 36912 9704
rect 36495 9673 36507 9676
rect 36449 9667 36507 9673
rect 36906 9664 36912 9676
rect 36964 9664 36970 9716
rect 36998 9664 37004 9716
rect 37056 9704 37062 9716
rect 38930 9704 38936 9716
rect 37056 9676 38936 9704
rect 37056 9664 37062 9676
rect 38930 9664 38936 9676
rect 38988 9664 38994 9716
rect 39022 9664 39028 9716
rect 39080 9664 39086 9716
rect 40678 9664 40684 9716
rect 40736 9704 40742 9716
rect 40865 9707 40923 9713
rect 40865 9704 40877 9707
rect 40736 9676 40877 9704
rect 40736 9664 40742 9676
rect 40865 9673 40877 9676
rect 40911 9673 40923 9707
rect 40865 9667 40923 9673
rect 34146 9636 34152 9648
rect 32355 9608 32904 9636
rect 32968 9608 34152 9636
rect 32355 9605 32367 9608
rect 32309 9599 32367 9605
rect 31389 9571 31447 9577
rect 31389 9568 31401 9571
rect 30484 9540 31401 9568
rect 28169 9531 28227 9537
rect 31389 9537 31401 9540
rect 31435 9537 31447 9571
rect 31389 9531 31447 9537
rect 31478 9528 31484 9580
rect 31536 9528 31542 9580
rect 32968 9577 32996 9608
rect 32953 9571 33011 9577
rect 32953 9537 32965 9571
rect 32999 9537 33011 9571
rect 32953 9531 33011 9537
rect 33134 9528 33140 9580
rect 33192 9528 33198 9580
rect 33226 9528 33232 9580
rect 33284 9528 33290 9580
rect 33318 9528 33324 9580
rect 33376 9528 33382 9580
rect 33980 9577 34008 9608
rect 34146 9596 34152 9608
rect 34204 9596 34210 9648
rect 34241 9639 34299 9645
rect 34241 9605 34253 9639
rect 34287 9636 34299 9639
rect 34330 9636 34336 9648
rect 34287 9608 34336 9636
rect 34287 9605 34299 9608
rect 34241 9599 34299 9605
rect 33965 9571 34023 9577
rect 33965 9537 33977 9571
rect 34011 9537 34023 9571
rect 33965 9531 34023 9537
rect 34054 9528 34060 9580
rect 34112 9568 34118 9580
rect 34256 9568 34284 9599
rect 34330 9596 34336 9608
rect 34388 9596 34394 9648
rect 34698 9596 34704 9648
rect 34756 9596 34762 9648
rect 37550 9596 37556 9648
rect 37608 9596 37614 9648
rect 39298 9636 39304 9648
rect 38778 9608 39304 9636
rect 39298 9596 39304 9608
rect 39356 9596 39362 9648
rect 39390 9596 39396 9648
rect 39448 9596 39454 9648
rect 39850 9596 39856 9648
rect 39908 9596 39914 9648
rect 34790 9568 34796 9580
rect 34112 9540 34284 9568
rect 34440 9540 34796 9568
rect 34112 9528 34118 9540
rect 26234 9460 26240 9512
rect 26292 9460 26298 9512
rect 26328 9503 26386 9509
rect 26328 9469 26340 9503
rect 26374 9469 26386 9503
rect 26328 9463 26386 9469
rect 26421 9503 26479 9509
rect 26421 9469 26433 9503
rect 26467 9469 26479 9503
rect 26878 9500 26884 9512
rect 26421 9463 26479 9469
rect 26712 9472 26884 9500
rect 26344 9432 26372 9463
rect 26160 9404 26372 9432
rect 26436 9432 26464 9463
rect 26712 9432 26740 9472
rect 26878 9460 26884 9472
rect 26936 9460 26942 9512
rect 27062 9460 27068 9512
rect 27120 9460 27126 9512
rect 28074 9460 28080 9512
rect 28132 9460 28138 9512
rect 28534 9460 28540 9512
rect 28592 9460 28598 9512
rect 28626 9460 28632 9512
rect 28684 9460 28690 9512
rect 29270 9500 29276 9512
rect 28736 9472 29276 9500
rect 26436 9404 26740 9432
rect 28552 9432 28580 9460
rect 28736 9432 28764 9472
rect 29270 9460 29276 9472
rect 29328 9500 29334 9512
rect 29546 9500 29552 9512
rect 29328 9472 29552 9500
rect 29328 9460 29334 9472
rect 29546 9460 29552 9472
rect 29604 9460 29610 9512
rect 30466 9460 30472 9512
rect 30524 9500 30530 9512
rect 31202 9500 31208 9512
rect 30524 9472 31208 9500
rect 30524 9460 30530 9472
rect 31202 9460 31208 9472
rect 31260 9460 31266 9512
rect 31294 9460 31300 9512
rect 31352 9500 31358 9512
rect 31849 9503 31907 9509
rect 31849 9500 31861 9503
rect 31352 9472 31861 9500
rect 31352 9460 31358 9472
rect 31849 9469 31861 9472
rect 31895 9469 31907 9503
rect 31849 9463 31907 9469
rect 32490 9460 32496 9512
rect 32548 9500 32554 9512
rect 32548 9472 33456 9500
rect 32548 9460 32554 9472
rect 33134 9432 33140 9444
rect 28552 9404 28764 9432
rect 29932 9404 33140 9432
rect 10744 9336 11560 9364
rect 10744 9324 10750 9336
rect 22370 9324 22376 9376
rect 22428 9364 22434 9376
rect 22465 9367 22523 9373
rect 22465 9364 22477 9367
rect 22428 9336 22477 9364
rect 22428 9324 22434 9336
rect 22465 9333 22477 9336
rect 22511 9333 22523 9367
rect 22465 9327 22523 9333
rect 22830 9324 22836 9376
rect 22888 9364 22894 9376
rect 23017 9367 23075 9373
rect 23017 9364 23029 9367
rect 22888 9336 23029 9364
rect 22888 9324 22894 9336
rect 23017 9333 23029 9336
rect 23063 9333 23075 9367
rect 23017 9327 23075 9333
rect 24026 9324 24032 9376
rect 24084 9364 24090 9376
rect 24670 9364 24676 9376
rect 24084 9336 24676 9364
rect 24084 9324 24090 9336
rect 24670 9324 24676 9336
rect 24728 9324 24734 9376
rect 26694 9324 26700 9376
rect 26752 9324 26758 9376
rect 27525 9367 27583 9373
rect 27525 9333 27537 9367
rect 27571 9364 27583 9367
rect 27614 9364 27620 9376
rect 27571 9336 27620 9364
rect 27571 9333 27583 9336
rect 27525 9327 27583 9333
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 28994 9324 29000 9376
rect 29052 9364 29058 9376
rect 29932 9364 29960 9404
rect 33134 9392 33140 9404
rect 33192 9392 33198 9444
rect 29052 9336 29960 9364
rect 29052 9324 29058 9336
rect 30374 9324 30380 9376
rect 30432 9364 30438 9376
rect 31294 9364 31300 9376
rect 30432 9336 31300 9364
rect 30432 9324 30438 9336
rect 31294 9324 31300 9336
rect 31352 9324 31358 9376
rect 31846 9324 31852 9376
rect 31904 9364 31910 9376
rect 32493 9367 32551 9373
rect 32493 9364 32505 9367
rect 31904 9336 32505 9364
rect 31904 9324 31910 9336
rect 32493 9333 32505 9336
rect 32539 9333 32551 9367
rect 33428 9364 33456 9472
rect 33870 9460 33876 9512
rect 33928 9460 33934 9512
rect 33505 9435 33563 9441
rect 33505 9401 33517 9435
rect 33551 9432 33563 9435
rect 34440 9432 34468 9540
rect 34790 9528 34796 9540
rect 34848 9528 34854 9580
rect 34885 9571 34943 9577
rect 34885 9537 34897 9571
rect 34931 9537 34943 9571
rect 34885 9531 34943 9537
rect 34900 9500 34928 9531
rect 35526 9528 35532 9580
rect 35584 9528 35590 9580
rect 36265 9571 36323 9577
rect 36265 9568 36277 9571
rect 35636 9540 36277 9568
rect 35636 9509 35664 9540
rect 36265 9537 36277 9540
rect 36311 9537 36323 9571
rect 36265 9531 36323 9537
rect 37274 9528 37280 9580
rect 37332 9528 37338 9580
rect 35621 9503 35679 9509
rect 35621 9500 35633 9503
rect 34624 9472 35633 9500
rect 34624 9441 34652 9472
rect 35621 9469 35633 9472
rect 35667 9469 35679 9503
rect 35621 9463 35679 9469
rect 35710 9460 35716 9512
rect 35768 9500 35774 9512
rect 36081 9503 36139 9509
rect 36081 9500 36093 9503
rect 35768 9472 36093 9500
rect 35768 9460 35774 9472
rect 36081 9469 36093 9472
rect 36127 9469 36139 9503
rect 39117 9503 39175 9509
rect 39117 9500 39129 9503
rect 36081 9463 36139 9469
rect 38580 9472 39129 9500
rect 33551 9404 34468 9432
rect 34609 9435 34667 9441
rect 33551 9401 33563 9404
rect 33505 9395 33563 9401
rect 34609 9401 34621 9435
rect 34655 9401 34667 9435
rect 34609 9395 34667 9401
rect 35342 9392 35348 9444
rect 35400 9432 35406 9444
rect 35400 9404 37412 9432
rect 35400 9392 35406 9404
rect 33689 9367 33747 9373
rect 33689 9364 33701 9367
rect 33428 9336 33701 9364
rect 32493 9327 32551 9333
rect 33689 9333 33701 9336
rect 33735 9333 33747 9367
rect 33689 9327 33747 9333
rect 34146 9324 34152 9376
rect 34204 9364 34210 9376
rect 34425 9367 34483 9373
rect 34425 9364 34437 9367
rect 34204 9336 34437 9364
rect 34204 9324 34210 9336
rect 34425 9333 34437 9336
rect 34471 9333 34483 9367
rect 34425 9327 34483 9333
rect 34514 9324 34520 9376
rect 34572 9364 34578 9376
rect 35069 9367 35127 9373
rect 35069 9364 35081 9367
rect 34572 9336 35081 9364
rect 34572 9324 34578 9336
rect 35069 9333 35081 9336
rect 35115 9333 35127 9367
rect 37384 9364 37412 9404
rect 38580 9364 38608 9472
rect 39117 9469 39129 9472
rect 39163 9469 39175 9503
rect 39117 9463 39175 9469
rect 37384 9336 38608 9364
rect 35069 9327 35127 9333
rect 1104 9274 42504 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 42504 9274
rect 1104 9200 42504 9222
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 5442 9160 5448 9172
rect 3936 9132 5448 9160
rect 3936 9120 3942 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5629 9163 5687 9169
rect 5629 9129 5641 9163
rect 5675 9160 5687 9163
rect 5994 9160 6000 9172
rect 5675 9132 6000 9160
rect 5675 9129 5687 9132
rect 5629 9123 5687 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6089 9163 6147 9169
rect 6089 9129 6101 9163
rect 6135 9160 6147 9163
rect 6178 9160 6184 9172
rect 6135 9132 6184 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11020 9132 11161 9160
rect 11020 9120 11026 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 11425 9163 11483 9169
rect 11425 9129 11437 9163
rect 11471 9160 11483 9163
rect 11790 9160 11796 9172
rect 11471 9132 11796 9160
rect 11471 9129 11483 9132
rect 11425 9123 11483 9129
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 20898 9120 20904 9172
rect 20956 9120 20962 9172
rect 22925 9163 22983 9169
rect 22925 9160 22937 9163
rect 21100 9132 22937 9160
rect 20254 9092 20260 9104
rect 19352 9064 20260 9092
rect 3234 8984 3240 9036
rect 3292 9024 3298 9036
rect 7466 9024 7472 9036
rect 3292 8996 7472 9024
rect 3292 8984 3298 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 9024 9459 9027
rect 10686 9024 10692 9036
rect 9447 8996 10692 9024
rect 9447 8993 9459 8996
rect 9401 8987 9459 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 4120 8928 4353 8956
rect 4120 8916 4126 8928
rect 4341 8925 4353 8928
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4614 8916 4620 8968
rect 4672 8916 4678 8968
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5994 8916 6000 8968
rect 6052 8916 6058 8968
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8956 6239 8959
rect 7098 8956 7104 8968
rect 6227 8928 7104 8956
rect 6227 8925 6239 8928
rect 6181 8919 6239 8925
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 11204 8928 11253 8956
rect 11204 8916 11210 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11388 8928 11437 8956
rect 11388 8916 11394 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 5552 8888 5580 8916
rect 5813 8891 5871 8897
rect 5813 8888 5825 8891
rect 5552 8860 5825 8888
rect 5813 8857 5825 8860
rect 5859 8857 5871 8891
rect 5813 8851 5871 8857
rect 9674 8848 9680 8900
rect 9732 8848 9738 8900
rect 10226 8848 10232 8900
rect 10284 8848 10290 8900
rect 19352 8888 19380 9064
rect 20254 9052 20260 9064
rect 20312 9092 20318 9104
rect 20990 9092 20996 9104
rect 20312 9064 20996 9092
rect 20312 9052 20318 9064
rect 20990 9052 20996 9064
rect 21048 9052 21054 9104
rect 19518 8984 19524 9036
rect 19576 8984 19582 9036
rect 20806 8984 20812 9036
rect 20864 9024 20870 9036
rect 21100 9024 21128 9132
rect 22925 9129 22937 9132
rect 22971 9129 22983 9163
rect 22925 9123 22983 9129
rect 23569 9163 23627 9169
rect 23569 9129 23581 9163
rect 23615 9160 23627 9163
rect 23658 9160 23664 9172
rect 23615 9132 23664 9160
rect 23615 9129 23627 9132
rect 23569 9123 23627 9129
rect 23658 9120 23664 9132
rect 23716 9120 23722 9172
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 24489 9163 24547 9169
rect 24489 9160 24501 9163
rect 24176 9132 24501 9160
rect 24176 9120 24182 9132
rect 24489 9129 24501 9132
rect 24535 9129 24547 9163
rect 24489 9123 24547 9129
rect 24670 9120 24676 9172
rect 24728 9160 24734 9172
rect 28534 9160 28540 9172
rect 24728 9132 28540 9160
rect 24728 9120 24734 9132
rect 28534 9120 28540 9132
rect 28592 9120 28598 9172
rect 31754 9120 31760 9172
rect 31812 9160 31818 9172
rect 32493 9163 32551 9169
rect 32493 9160 32505 9163
rect 31812 9132 32505 9160
rect 31812 9120 31818 9132
rect 32493 9129 32505 9132
rect 32539 9129 32551 9163
rect 32493 9123 32551 9129
rect 24394 9052 24400 9104
rect 24452 9092 24458 9104
rect 26878 9092 26884 9104
rect 24452 9064 26884 9092
rect 24452 9052 24458 9064
rect 26878 9052 26884 9064
rect 26936 9052 26942 9104
rect 30466 9092 30472 9104
rect 28828 9064 30472 9092
rect 20864 8996 21128 9024
rect 20864 8984 20870 8996
rect 22370 8984 22376 9036
rect 22428 8984 22434 9036
rect 23750 8984 23756 9036
rect 23808 9024 23814 9036
rect 23937 9027 23995 9033
rect 23937 9024 23949 9027
rect 23808 8996 23949 9024
rect 23808 8984 23814 8996
rect 23937 8993 23949 8996
rect 23983 9024 23995 9027
rect 27614 9024 27620 9036
rect 23983 8996 24624 9024
rect 23983 8993 23995 8996
rect 23937 8987 23995 8993
rect 19426 8916 19432 8968
rect 19484 8916 19490 8968
rect 19536 8956 19564 8984
rect 19797 8959 19855 8965
rect 19797 8956 19809 8959
rect 19536 8928 19809 8956
rect 19797 8925 19809 8928
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 23845 8959 23903 8965
rect 22756 8928 22968 8956
rect 19521 8891 19579 8897
rect 19521 8888 19533 8891
rect 19352 8860 19533 8888
rect 19521 8857 19533 8860
rect 19567 8857 19579 8891
rect 19521 8851 19579 8857
rect 19610 8848 19616 8900
rect 19668 8848 19674 8900
rect 22756 8888 22784 8928
rect 21942 8860 22784 8888
rect 22833 8891 22891 8897
rect 22833 8857 22845 8891
rect 22879 8857 22891 8891
rect 22940 8888 22968 8928
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24394 8956 24400 8968
rect 23891 8928 24400 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 24394 8916 24400 8928
rect 24452 8916 24458 8968
rect 24596 8965 24624 8996
rect 26896 8996 27620 9024
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 26602 8956 26608 8968
rect 24627 8928 26608 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 26602 8916 26608 8928
rect 26660 8916 26666 8968
rect 26694 8916 26700 8968
rect 26752 8965 26758 8968
rect 26896 8965 26924 8996
rect 27614 8984 27620 8996
rect 27672 8984 27678 9036
rect 26752 8959 26785 8965
rect 26773 8925 26785 8959
rect 26752 8919 26785 8925
rect 26881 8959 26939 8965
rect 26881 8925 26893 8959
rect 26927 8925 26939 8959
rect 26881 8919 26939 8925
rect 26752 8916 26758 8919
rect 27522 8916 27528 8968
rect 27580 8916 27586 8968
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8956 28411 8959
rect 28442 8956 28448 8968
rect 28399 8928 28448 8956
rect 28399 8925 28411 8928
rect 28353 8919 28411 8925
rect 28442 8916 28448 8928
rect 28500 8916 28506 8968
rect 28828 8965 28856 9064
rect 30466 9052 30472 9064
rect 30524 9052 30530 9104
rect 32508 9092 32536 9123
rect 33134 9120 33140 9172
rect 33192 9160 33198 9172
rect 33318 9160 33324 9172
rect 33192 9132 33324 9160
rect 33192 9120 33198 9132
rect 33318 9120 33324 9132
rect 33376 9160 33382 9172
rect 33689 9163 33747 9169
rect 33376 9132 33456 9160
rect 33376 9120 33382 9132
rect 32950 9092 32956 9104
rect 32508 9064 32956 9092
rect 32950 9052 32956 9064
rect 33008 9092 33014 9104
rect 33008 9064 33364 9092
rect 33008 9052 33014 9064
rect 30742 9024 30748 9036
rect 30484 8996 30748 9024
rect 28813 8959 28871 8965
rect 28813 8925 28825 8959
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 28994 8916 29000 8968
rect 29052 8916 29058 8968
rect 29086 8916 29092 8968
rect 29144 8916 29150 8968
rect 29178 8916 29184 8968
rect 29236 8916 29242 8968
rect 30484 8965 30512 8996
rect 30742 8984 30748 8996
rect 30800 8984 30806 9036
rect 31021 9027 31079 9033
rect 31021 8993 31033 9027
rect 31067 9024 31079 9027
rect 32585 9027 32643 9033
rect 32585 9024 32597 9027
rect 31067 8996 32597 9024
rect 31067 8993 31079 8996
rect 31021 8987 31079 8993
rect 32585 8993 32597 8996
rect 32631 8993 32643 9027
rect 33042 9024 33048 9036
rect 32585 8987 32643 8993
rect 32784 8996 33048 9024
rect 30469 8959 30527 8965
rect 30469 8925 30481 8959
rect 30515 8925 30527 8959
rect 30469 8919 30527 8925
rect 32122 8916 32128 8968
rect 32180 8956 32186 8968
rect 32784 8956 32812 8996
rect 33042 8984 33048 8996
rect 33100 8984 33106 9036
rect 33336 9033 33364 9064
rect 33321 9027 33379 9033
rect 33321 8993 33333 9027
rect 33367 8993 33379 9027
rect 33428 9024 33456 9132
rect 33689 9129 33701 9163
rect 33735 9160 33747 9163
rect 33870 9160 33876 9172
rect 33735 9132 33876 9160
rect 33735 9129 33747 9132
rect 33689 9123 33747 9129
rect 33870 9120 33876 9132
rect 33928 9120 33934 9172
rect 33962 9120 33968 9172
rect 34020 9160 34026 9172
rect 34606 9160 34612 9172
rect 34020 9132 34612 9160
rect 34020 9120 34026 9132
rect 34606 9120 34612 9132
rect 34664 9120 34670 9172
rect 35250 9120 35256 9172
rect 35308 9160 35314 9172
rect 35526 9160 35532 9172
rect 35308 9132 35532 9160
rect 35308 9120 35314 9132
rect 35526 9120 35532 9132
rect 35584 9120 35590 9172
rect 37366 9120 37372 9172
rect 37424 9160 37430 9172
rect 38470 9160 38476 9172
rect 37424 9132 38476 9160
rect 37424 9120 37430 9132
rect 38470 9120 38476 9132
rect 38528 9120 38534 9172
rect 33594 9052 33600 9104
rect 33652 9092 33658 9104
rect 33652 9064 37504 9092
rect 33652 9052 33658 9064
rect 33428 8996 34192 9024
rect 33321 8987 33379 8993
rect 32180 8928 32812 8956
rect 32180 8916 32186 8928
rect 32858 8916 32864 8968
rect 32916 8956 32922 8968
rect 33137 8959 33195 8965
rect 33137 8956 33149 8959
rect 32916 8928 33149 8956
rect 32916 8916 32922 8928
rect 33137 8925 33149 8928
rect 33183 8925 33195 8959
rect 33137 8919 33195 8925
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8925 33563 8959
rect 33505 8919 33563 8925
rect 33965 8959 34023 8965
rect 33965 8925 33977 8959
rect 34011 8956 34023 8959
rect 34011 8928 34100 8956
rect 34011 8925 34023 8928
rect 33965 8919 34023 8925
rect 24118 8888 24124 8900
rect 22940 8860 24124 8888
rect 22833 8851 22891 8857
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3660 8792 3801 8820
rect 3660 8780 3666 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 4798 8780 4804 8832
rect 4856 8820 4862 8832
rect 4893 8823 4951 8829
rect 4893 8820 4905 8823
rect 4856 8792 4905 8820
rect 4856 8780 4862 8792
rect 4893 8789 4905 8792
rect 4939 8789 4951 8823
rect 4893 8783 4951 8789
rect 5613 8823 5671 8829
rect 5613 8789 5625 8823
rect 5659 8820 5671 8823
rect 5718 8820 5724 8832
rect 5659 8792 5724 8820
rect 5659 8789 5671 8792
rect 5613 8783 5671 8789
rect 5718 8780 5724 8792
rect 5776 8820 5782 8832
rect 6454 8820 6460 8832
rect 5776 8792 6460 8820
rect 5776 8780 5782 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 19245 8823 19303 8829
rect 19245 8789 19257 8823
rect 19291 8820 19303 8823
rect 20346 8820 20352 8832
rect 19291 8792 20352 8820
rect 19291 8789 19303 8792
rect 19245 8783 19303 8789
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 22094 8780 22100 8832
rect 22152 8820 22158 8832
rect 22848 8820 22876 8851
rect 24118 8848 24124 8860
rect 24176 8848 24182 8900
rect 28074 8888 28080 8900
rect 24228 8860 28080 8888
rect 22152 8792 22876 8820
rect 22152 8780 22158 8792
rect 23842 8780 23848 8832
rect 23900 8820 23906 8832
rect 24228 8820 24256 8860
rect 28074 8848 28080 8860
rect 28132 8848 28138 8900
rect 28721 8891 28779 8897
rect 28721 8857 28733 8891
rect 28767 8888 28779 8891
rect 29012 8888 29040 8916
rect 33520 8888 33548 8919
rect 28767 8860 29040 8888
rect 32416 8860 33548 8888
rect 28767 8857 28779 8860
rect 28721 8851 28779 8857
rect 23900 8792 24256 8820
rect 26513 8823 26571 8829
rect 23900 8780 23906 8792
rect 26513 8789 26525 8823
rect 26559 8820 26571 8823
rect 27154 8820 27160 8832
rect 26559 8792 27160 8820
rect 26559 8789 26571 8792
rect 26513 8783 26571 8789
rect 27154 8780 27160 8792
rect 27212 8820 27218 8832
rect 27430 8820 27436 8832
rect 27212 8792 27436 8820
rect 27212 8780 27218 8792
rect 27430 8780 27436 8792
rect 27488 8780 27494 8832
rect 28166 8780 28172 8832
rect 28224 8780 28230 8832
rect 28350 8780 28356 8832
rect 28408 8820 28414 8832
rect 29270 8820 29276 8832
rect 28408 8792 29276 8820
rect 28408 8780 28414 8792
rect 29270 8780 29276 8792
rect 29328 8780 29334 8832
rect 29365 8823 29423 8829
rect 29365 8789 29377 8823
rect 29411 8820 29423 8823
rect 29454 8820 29460 8832
rect 29411 8792 29460 8820
rect 29411 8789 29423 8792
rect 29365 8783 29423 8789
rect 29454 8780 29460 8792
rect 29512 8780 29518 8832
rect 31662 8780 31668 8832
rect 31720 8820 31726 8832
rect 32416 8820 32444 8860
rect 31720 8792 32444 8820
rect 34072 8820 34100 8928
rect 34164 8897 34192 8996
rect 34256 8965 34284 9064
rect 35268 8996 35664 9024
rect 34241 8959 34299 8965
rect 34241 8925 34253 8959
rect 34287 8925 34299 8959
rect 34241 8919 34299 8925
rect 34330 8916 34336 8968
rect 34388 8916 34394 8968
rect 35268 8956 35296 8996
rect 34532 8928 35296 8956
rect 34149 8891 34207 8897
rect 34149 8857 34161 8891
rect 34195 8888 34207 8891
rect 34532 8888 34560 8928
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 35437 8959 35495 8965
rect 35437 8956 35449 8959
rect 35400 8928 35449 8956
rect 35400 8916 35406 8928
rect 35437 8925 35449 8928
rect 35483 8925 35495 8959
rect 35636 8956 35664 8996
rect 35710 8984 35716 9036
rect 35768 9024 35774 9036
rect 36449 9027 36507 9033
rect 36449 9024 36461 9027
rect 35768 8996 36461 9024
rect 35768 8984 35774 8996
rect 36449 8993 36461 8996
rect 36495 8993 36507 9027
rect 37366 9024 37372 9036
rect 36449 8987 36507 8993
rect 36556 8996 37372 9024
rect 36556 8956 36584 8996
rect 37366 8984 37372 8996
rect 37424 8984 37430 9036
rect 35636 8928 36584 8956
rect 37093 8959 37151 8965
rect 35437 8919 35495 8925
rect 37093 8925 37105 8959
rect 37139 8956 37151 8959
rect 37185 8959 37243 8965
rect 37185 8956 37197 8959
rect 37139 8928 37197 8956
rect 37139 8925 37151 8928
rect 37093 8919 37151 8925
rect 37185 8925 37197 8928
rect 37231 8925 37243 8959
rect 37185 8919 37243 8925
rect 34195 8860 34560 8888
rect 34195 8857 34207 8860
rect 34149 8851 34207 8857
rect 34606 8848 34612 8900
rect 34664 8888 34670 8900
rect 37274 8888 37280 8900
rect 34664 8860 37280 8888
rect 34664 8848 34670 8860
rect 37274 8848 37280 8860
rect 37332 8848 37338 8900
rect 37384 8897 37412 8984
rect 37476 8897 37504 9064
rect 37553 8959 37611 8965
rect 37553 8925 37565 8959
rect 37599 8956 37611 8959
rect 37826 8956 37832 8968
rect 37599 8928 37832 8956
rect 37599 8925 37611 8928
rect 37553 8919 37611 8925
rect 37826 8916 37832 8928
rect 37884 8916 37890 8968
rect 37369 8891 37427 8897
rect 37369 8857 37381 8891
rect 37415 8857 37427 8891
rect 37369 8851 37427 8857
rect 37461 8891 37519 8897
rect 37461 8857 37473 8891
rect 37507 8888 37519 8891
rect 37918 8888 37924 8900
rect 37507 8860 37924 8888
rect 37507 8857 37519 8860
rect 37461 8851 37519 8857
rect 37918 8848 37924 8860
rect 37976 8848 37982 8900
rect 34422 8820 34428 8832
rect 34072 8792 34428 8820
rect 31720 8780 31726 8792
rect 34422 8780 34428 8792
rect 34480 8780 34486 8832
rect 34517 8823 34575 8829
rect 34517 8789 34529 8823
rect 34563 8820 34575 8823
rect 34698 8820 34704 8832
rect 34563 8792 34704 8820
rect 34563 8789 34575 8792
rect 34517 8783 34575 8789
rect 34698 8780 34704 8792
rect 34756 8780 34762 8832
rect 35158 8780 35164 8832
rect 35216 8820 35222 8832
rect 37642 8820 37648 8832
rect 35216 8792 37648 8820
rect 35216 8780 35222 8792
rect 37642 8780 37648 8792
rect 37700 8780 37706 8832
rect 37734 8780 37740 8832
rect 37792 8780 37798 8832
rect 1104 8730 42504 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 42504 8730
rect 1104 8656 42504 8678
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 1688 8588 3893 8616
rect 1688 8557 1716 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 4433 8619 4491 8625
rect 3881 8579 3939 8585
rect 4080 8588 4384 8616
rect 1673 8551 1731 8557
rect 1673 8517 1685 8551
rect 1719 8517 1731 8551
rect 3234 8548 3240 8560
rect 2898 8520 3240 8548
rect 1673 8511 1731 8517
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 4080 8557 4108 8588
rect 4065 8551 4123 8557
rect 4065 8548 4077 8551
rect 4028 8520 4077 8548
rect 4028 8508 4034 8520
rect 4065 8517 4077 8520
rect 4111 8517 4123 8551
rect 4265 8551 4323 8557
rect 4265 8548 4277 8551
rect 4065 8511 4123 8517
rect 4172 8520 4277 8548
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4172 8480 4200 8520
rect 4265 8517 4277 8520
rect 4311 8517 4323 8551
rect 4356 8548 4384 8588
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 5461 8619 5519 8625
rect 5461 8616 5473 8619
rect 4479 8588 5473 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 5461 8585 5473 8588
rect 5507 8585 5519 8619
rect 5461 8579 5519 8585
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 5813 8619 5871 8625
rect 5813 8585 5825 8619
rect 5859 8616 5871 8619
rect 6638 8616 6644 8628
rect 5859 8588 6644 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 8849 8619 8907 8625
rect 8849 8616 8861 8619
rect 6972 8588 8861 8616
rect 6972 8576 6978 8588
rect 8849 8585 8861 8588
rect 8895 8585 8907 8619
rect 8849 8579 8907 8585
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 19518 8616 19524 8628
rect 18923 8588 19524 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 21358 8576 21364 8628
rect 21416 8616 21422 8628
rect 26418 8616 26424 8628
rect 21416 8588 26424 8616
rect 21416 8576 21422 8588
rect 5261 8551 5319 8557
rect 4356 8520 4844 8548
rect 4265 8511 4323 8517
rect 4816 8489 4844 8520
rect 5261 8517 5273 8551
rect 5307 8517 5319 8551
rect 5261 8511 5319 8517
rect 6549 8551 6607 8557
rect 6549 8517 6561 8551
rect 6595 8548 6607 8551
rect 6822 8548 6828 8560
rect 6595 8520 6828 8548
rect 6595 8517 6607 8520
rect 6549 8511 6607 8517
rect 3844 8452 4200 8480
rect 4525 8483 4583 8489
rect 3844 8440 3850 8452
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4801 8483 4859 8489
rect 4571 8452 4752 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2740 8384 3249 8412
rect 2740 8372 2746 8384
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3694 8372 3700 8424
rect 3752 8372 3758 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8381 4675 8415
rect 4724 8412 4752 8452
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 5276 8480 5304 8511
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 8021 8551 8079 8557
rect 7064 8520 7328 8548
rect 7064 8508 7070 8520
rect 4801 8443 4859 8449
rect 4908 8452 5304 8480
rect 4908 8424 4936 8452
rect 5718 8440 5724 8492
rect 5776 8440 5782 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 4890 8412 4896 8424
rect 4724 8384 4896 8412
rect 4617 8375 4675 8381
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 3786 8344 3792 8356
rect 3191 8316 3792 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 3786 8304 3792 8316
rect 3844 8344 3850 8356
rect 4062 8344 4068 8356
rect 3844 8316 4068 8344
rect 3844 8304 3850 8316
rect 4062 8304 4068 8316
rect 4120 8344 4126 8356
rect 4632 8344 4660 8375
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5920 8412 5948 8443
rect 6454 8440 6460 8492
rect 6512 8440 6518 8492
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8480 6791 8483
rect 7190 8480 7196 8492
rect 6779 8452 7196 8480
rect 6779 8449 6791 8452
rect 6733 8443 6791 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7300 8489 7328 8520
rect 8021 8517 8033 8551
rect 8067 8548 8079 8551
rect 8662 8548 8668 8560
rect 8067 8520 8668 8548
rect 8067 8517 8079 8520
rect 8021 8511 8079 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 20346 8508 20352 8560
rect 20404 8508 20410 8560
rect 20714 8508 20720 8560
rect 20772 8508 20778 8560
rect 23658 8508 23664 8560
rect 23716 8508 23722 8560
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 5000 8384 5948 8412
rect 6472 8412 6500 8440
rect 6914 8412 6920 8424
rect 6472 8384 6920 8412
rect 5000 8353 5028 8384
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 4120 8316 4660 8344
rect 4985 8347 5043 8353
rect 4120 8304 4126 8316
rect 4985 8313 4997 8347
rect 5031 8313 5043 8347
rect 5534 8344 5540 8356
rect 4985 8307 5043 8313
rect 5092 8316 5540 8344
rect 4249 8279 4307 8285
rect 4249 8245 4261 8279
rect 4295 8276 4307 8279
rect 4801 8279 4859 8285
rect 4801 8276 4813 8279
rect 4295 8248 4813 8276
rect 4295 8245 4307 8248
rect 4249 8239 4307 8245
rect 4801 8245 4813 8248
rect 4847 8276 4859 8279
rect 5092 8276 5120 8316
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 7006 8344 7012 8356
rect 5684 8316 7012 8344
rect 5684 8304 5690 8316
rect 7006 8304 7012 8316
rect 7064 8344 7070 8356
rect 7101 8347 7159 8353
rect 7101 8344 7113 8347
rect 7064 8316 7113 8344
rect 7064 8304 7070 8316
rect 7101 8313 7113 8316
rect 7147 8313 7159 8347
rect 7300 8344 7328 8443
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8941 8483 8999 8489
rect 8941 8480 8953 8483
rect 8352 8452 8953 8480
rect 8352 8440 8358 8452
rect 8941 8449 8953 8452
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16908 8452 16957 8480
rect 16908 8440 16914 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 21545 8483 21603 8489
rect 18380 8452 19274 8480
rect 18380 8440 18386 8452
rect 21545 8449 21557 8483
rect 21591 8480 21603 8483
rect 22370 8480 22376 8492
rect 21591 8452 22376 8480
rect 21591 8449 21603 8452
rect 21545 8443 21603 8449
rect 8202 8372 8208 8424
rect 8260 8372 8266 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8496 8384 8585 8412
rect 8496 8353 8524 8384
rect 8573 8381 8585 8384
rect 8619 8412 8631 8415
rect 8754 8412 8760 8424
rect 8619 8384 8760 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 17221 8415 17279 8421
rect 17221 8381 17233 8415
rect 17267 8412 17279 8415
rect 19150 8412 19156 8424
rect 17267 8384 19156 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 20625 8415 20683 8421
rect 20625 8381 20637 8415
rect 20671 8412 20683 8415
rect 21560 8412 21588 8443
rect 22370 8440 22376 8452
rect 22428 8480 22434 8492
rect 22646 8480 22652 8492
rect 22428 8452 22652 8480
rect 22428 8440 22434 8452
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 23676 8480 23704 8508
rect 23753 8483 23811 8489
rect 23753 8480 23765 8483
rect 23676 8452 23765 8480
rect 23753 8449 23765 8452
rect 23799 8449 23811 8483
rect 23952 8480 23980 8588
rect 26418 8576 26424 8588
rect 26476 8576 26482 8628
rect 26789 8619 26847 8625
rect 26789 8585 26801 8619
rect 26835 8616 26847 8619
rect 28902 8616 28908 8628
rect 26835 8588 28908 8616
rect 26835 8585 26847 8588
rect 26789 8579 26847 8585
rect 28902 8576 28908 8588
rect 28960 8576 28966 8628
rect 30374 8616 30380 8628
rect 29380 8588 30380 8616
rect 24029 8551 24087 8557
rect 24029 8517 24041 8551
rect 24075 8548 24087 8551
rect 26510 8548 26516 8560
rect 24075 8520 24808 8548
rect 24075 8517 24087 8520
rect 24029 8511 24087 8517
rect 23952 8452 24348 8480
rect 23753 8443 23811 8449
rect 20671 8384 21588 8412
rect 23661 8415 23719 8421
rect 20671 8381 20683 8384
rect 20625 8375 20683 8381
rect 23661 8381 23673 8415
rect 23707 8412 23719 8415
rect 23842 8412 23848 8424
rect 23707 8384 23848 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 24026 8372 24032 8424
rect 24084 8412 24090 8424
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 24084 8384 24133 8412
rect 24084 8372 24090 8384
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24320 8412 24348 8452
rect 24394 8440 24400 8492
rect 24452 8440 24458 8492
rect 24780 8489 24808 8520
rect 26160 8520 26516 8548
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 24765 8483 24823 8489
rect 24765 8449 24777 8483
rect 24811 8480 24823 8483
rect 25222 8480 25228 8492
rect 24811 8452 25228 8480
rect 24811 8449 24823 8452
rect 24765 8443 24823 8449
rect 24596 8412 24624 8443
rect 24320 8384 24624 8412
rect 24688 8412 24716 8443
rect 25222 8440 25228 8452
rect 25280 8440 25286 8492
rect 26160 8412 26188 8520
rect 26510 8508 26516 8520
rect 26568 8508 26574 8560
rect 28166 8548 28172 8560
rect 26620 8520 28172 8548
rect 26237 8483 26295 8489
rect 26237 8449 26249 8483
rect 26283 8449 26295 8483
rect 26237 8443 26295 8449
rect 24688 8384 26188 8412
rect 26252 8412 26280 8443
rect 26418 8440 26424 8492
rect 26476 8440 26482 8492
rect 26620 8489 26648 8520
rect 28166 8508 28172 8520
rect 28224 8548 28230 8560
rect 28261 8551 28319 8557
rect 28261 8548 28273 8551
rect 28224 8520 28273 8548
rect 28224 8508 28230 8520
rect 28261 8517 28273 8520
rect 28307 8517 28319 8551
rect 28261 8511 28319 8517
rect 28350 8508 28356 8560
rect 28408 8508 28414 8560
rect 26605 8483 26663 8489
rect 26605 8449 26617 8483
rect 26651 8449 26663 8483
rect 26605 8443 26663 8449
rect 27062 8440 27068 8492
rect 27120 8480 27126 8492
rect 27430 8480 27436 8492
rect 27120 8452 27436 8480
rect 27120 8440 27126 8452
rect 27430 8440 27436 8452
rect 27488 8480 27494 8492
rect 27525 8483 27583 8489
rect 27525 8480 27537 8483
rect 27488 8452 27537 8480
rect 27488 8440 27494 8452
rect 27525 8449 27537 8452
rect 27571 8449 27583 8483
rect 27985 8483 28043 8489
rect 27985 8480 27997 8483
rect 27525 8443 27583 8449
rect 27632 8452 27997 8480
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26252 8384 26985 8412
rect 24121 8375 24179 8381
rect 8481 8347 8539 8353
rect 7300 8316 8432 8344
rect 7101 8307 7159 8313
rect 4847 8248 5120 8276
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 5442 8236 5448 8288
rect 5500 8236 5506 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 6733 8279 6791 8285
rect 6733 8276 6745 8279
rect 6696 8248 6745 8276
rect 6696 8236 6702 8248
rect 6733 8245 6745 8248
rect 6779 8245 6791 8279
rect 6733 8239 6791 8245
rect 8202 8236 8208 8288
rect 8260 8236 8266 8288
rect 8404 8276 8432 8316
rect 8481 8313 8493 8347
rect 8527 8313 8539 8347
rect 10318 8344 10324 8356
rect 8481 8307 8539 8313
rect 8588 8316 10324 8344
rect 8588 8276 8616 8316
rect 10318 8304 10324 8316
rect 10376 8344 10382 8356
rect 11146 8344 11152 8356
rect 10376 8316 11152 8344
rect 10376 8304 10382 8316
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 18693 8347 18751 8353
rect 18693 8313 18705 8347
rect 18739 8344 18751 8347
rect 19334 8344 19340 8356
rect 18739 8316 19340 8344
rect 18739 8313 18751 8316
rect 18693 8307 18751 8313
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 20990 8304 20996 8356
rect 21048 8344 21054 8356
rect 21358 8344 21364 8356
rect 21048 8316 21364 8344
rect 21048 8304 21054 8316
rect 21358 8304 21364 8316
rect 21416 8344 21422 8356
rect 24688 8344 24716 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 27154 8372 27160 8424
rect 27212 8412 27218 8424
rect 27632 8412 27660 8452
rect 27985 8449 27997 8452
rect 28031 8449 28043 8483
rect 27985 8443 28043 8449
rect 28905 8483 28963 8489
rect 28905 8449 28917 8483
rect 28951 8480 28963 8483
rect 29380 8480 29408 8588
rect 30374 8576 30380 8588
rect 30432 8576 30438 8628
rect 32858 8576 32864 8628
rect 32916 8576 32922 8628
rect 34241 8619 34299 8625
rect 34241 8585 34253 8619
rect 34287 8616 34299 8619
rect 34330 8616 34336 8628
rect 34287 8588 34336 8616
rect 34287 8585 34299 8588
rect 34241 8579 34299 8585
rect 30742 8548 30748 8560
rect 30208 8520 30748 8548
rect 28951 8452 29408 8480
rect 28951 8449 28963 8452
rect 28905 8443 28963 8449
rect 29454 8440 29460 8492
rect 29512 8440 29518 8492
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 30208 8489 30236 8520
rect 30742 8508 30748 8520
rect 30800 8508 30806 8560
rect 32950 8508 32956 8560
rect 33008 8548 33014 8560
rect 33962 8548 33968 8560
rect 33008 8520 33456 8548
rect 33008 8508 33014 8520
rect 30193 8483 30251 8489
rect 30193 8480 30205 8483
rect 29604 8452 30205 8480
rect 29604 8440 29610 8452
rect 30193 8449 30205 8452
rect 30239 8449 30251 8483
rect 30193 8443 30251 8449
rect 31570 8440 31576 8492
rect 31628 8440 31634 8492
rect 33045 8483 33103 8489
rect 33045 8480 33057 8483
rect 32784 8452 33057 8480
rect 27212 8384 27660 8412
rect 27893 8415 27951 8421
rect 27212 8372 27218 8384
rect 27893 8381 27905 8415
rect 27939 8381 27951 8415
rect 27893 8375 27951 8381
rect 28813 8415 28871 8421
rect 28813 8381 28825 8415
rect 28859 8381 28871 8415
rect 28813 8375 28871 8381
rect 21416 8316 24716 8344
rect 21416 8304 21422 8316
rect 26326 8304 26332 8356
rect 26384 8344 26390 8356
rect 27709 8347 27767 8353
rect 27709 8344 27721 8347
rect 26384 8316 27721 8344
rect 26384 8304 26390 8316
rect 27709 8313 27721 8316
rect 27755 8313 27767 8347
rect 27908 8344 27936 8375
rect 28074 8344 28080 8356
rect 27908 8316 28080 8344
rect 27709 8307 27767 8313
rect 28074 8304 28080 8316
rect 28132 8344 28138 8356
rect 28828 8344 28856 8375
rect 29178 8372 29184 8424
rect 29236 8372 29242 8424
rect 29270 8372 29276 8424
rect 29328 8372 29334 8424
rect 30466 8372 30472 8424
rect 30524 8372 30530 8424
rect 31941 8415 31999 8421
rect 31941 8381 31953 8415
rect 31987 8412 31999 8415
rect 32125 8415 32183 8421
rect 32125 8412 32137 8415
rect 31987 8384 32137 8412
rect 31987 8381 31999 8384
rect 31941 8375 31999 8381
rect 32125 8381 32137 8384
rect 32171 8381 32183 8415
rect 32125 8375 32183 8381
rect 28132 8316 30328 8344
rect 28132 8304 28138 8316
rect 8404 8248 8616 8276
rect 23474 8236 23480 8288
rect 23532 8236 23538 8288
rect 24949 8279 25007 8285
rect 24949 8245 24961 8279
rect 24995 8276 25007 8279
rect 25406 8276 25412 8288
rect 24995 8248 25412 8276
rect 24995 8245 25007 8248
rect 24949 8239 25007 8245
rect 25406 8236 25412 8248
rect 25464 8236 25470 8288
rect 28258 8236 28264 8288
rect 28316 8276 28322 8288
rect 28629 8279 28687 8285
rect 28629 8276 28641 8279
rect 28316 8248 28641 8276
rect 28316 8236 28322 8248
rect 28629 8245 28641 8248
rect 28675 8245 28687 8279
rect 28629 8239 28687 8245
rect 29822 8236 29828 8288
rect 29880 8276 29886 8288
rect 30101 8279 30159 8285
rect 30101 8276 30113 8279
rect 29880 8248 30113 8276
rect 29880 8236 29886 8248
rect 30101 8245 30113 8248
rect 30147 8245 30159 8279
rect 30300 8276 30328 8316
rect 30558 8276 30564 8288
rect 30300 8248 30564 8276
rect 30101 8239 30159 8245
rect 30558 8236 30564 8248
rect 30616 8236 30622 8288
rect 31938 8236 31944 8288
rect 31996 8276 32002 8288
rect 32784 8285 32812 8452
rect 33045 8449 33057 8452
rect 33091 8449 33103 8483
rect 33045 8443 33103 8449
rect 33134 8440 33140 8492
rect 33192 8440 33198 8492
rect 33229 8483 33287 8489
rect 33229 8449 33241 8483
rect 33275 8480 33287 8483
rect 33318 8480 33324 8492
rect 33275 8452 33324 8480
rect 33275 8449 33287 8452
rect 33229 8443 33287 8449
rect 33318 8440 33324 8452
rect 33376 8440 33382 8492
rect 33428 8489 33456 8520
rect 33612 8520 33968 8548
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8449 33471 8483
rect 33612 8480 33640 8520
rect 33962 8508 33968 8520
rect 34020 8508 34026 8560
rect 34057 8551 34115 8557
rect 34057 8517 34069 8551
rect 34103 8548 34115 8551
rect 34256 8548 34284 8579
rect 34330 8576 34336 8588
rect 34388 8576 34394 8628
rect 34422 8576 34428 8628
rect 34480 8616 34486 8628
rect 36265 8619 36323 8625
rect 36265 8616 36277 8619
rect 34480 8588 36277 8616
rect 34480 8576 34486 8588
rect 36265 8585 36277 8588
rect 36311 8585 36323 8619
rect 36265 8579 36323 8585
rect 34103 8520 34284 8548
rect 34103 8517 34115 8520
rect 34057 8511 34115 8517
rect 35434 8508 35440 8560
rect 35492 8548 35498 8560
rect 36173 8551 36231 8557
rect 36173 8548 36185 8551
rect 35492 8520 36185 8548
rect 35492 8508 35498 8520
rect 36173 8517 36185 8520
rect 36219 8517 36231 8551
rect 36173 8511 36231 8517
rect 37826 8508 37832 8560
rect 37884 8508 37890 8560
rect 33674 8483 33732 8489
rect 33674 8480 33686 8483
rect 33612 8452 33686 8480
rect 33413 8443 33471 8449
rect 33674 8449 33686 8452
rect 33720 8449 33732 8483
rect 33674 8443 33732 8449
rect 33781 8483 33839 8489
rect 33781 8449 33793 8483
rect 33827 8480 33839 8483
rect 34238 8480 34244 8492
rect 33827 8452 34244 8480
rect 33827 8449 33839 8452
rect 33781 8443 33839 8449
rect 34238 8440 34244 8452
rect 34296 8440 34302 8492
rect 35158 8480 35164 8492
rect 34716 8452 35164 8480
rect 32950 8372 32956 8424
rect 33008 8412 33014 8424
rect 34149 8415 34207 8421
rect 34149 8412 34161 8415
rect 33008 8384 34161 8412
rect 33008 8372 33014 8384
rect 34149 8381 34161 8384
rect 34195 8412 34207 8415
rect 34716 8412 34744 8452
rect 35158 8440 35164 8452
rect 35216 8440 35222 8492
rect 36262 8440 36268 8492
rect 36320 8480 36326 8492
rect 37553 8483 37611 8489
rect 37553 8480 37565 8483
rect 36320 8452 37565 8480
rect 36320 8440 36326 8452
rect 37553 8449 37565 8452
rect 37599 8449 37611 8483
rect 37553 8443 37611 8449
rect 37642 8440 37648 8492
rect 37700 8480 37706 8492
rect 37921 8483 37979 8489
rect 37921 8480 37933 8483
rect 37700 8452 37933 8480
rect 37700 8440 37706 8452
rect 37921 8449 37933 8452
rect 37967 8449 37979 8483
rect 37921 8443 37979 8449
rect 34195 8384 34744 8412
rect 34195 8381 34207 8384
rect 34149 8375 34207 8381
rect 34790 8372 34796 8424
rect 34848 8372 34854 8424
rect 35434 8372 35440 8424
rect 35492 8372 35498 8424
rect 36817 8415 36875 8421
rect 36817 8412 36829 8415
rect 35544 8384 36829 8412
rect 34054 8304 34060 8356
rect 34112 8344 34118 8356
rect 35544 8344 35572 8384
rect 36817 8381 36829 8384
rect 36863 8381 36875 8415
rect 36817 8375 36875 8381
rect 37458 8372 37464 8424
rect 37516 8372 37522 8424
rect 34112 8316 35572 8344
rect 34112 8304 34118 8316
rect 35894 8304 35900 8356
rect 35952 8344 35958 8356
rect 37277 8347 37335 8353
rect 37277 8344 37289 8347
rect 35952 8316 37289 8344
rect 35952 8304 35958 8316
rect 37277 8313 37289 8316
rect 37323 8313 37335 8347
rect 37277 8307 37335 8313
rect 32769 8279 32827 8285
rect 32769 8276 32781 8279
rect 31996 8248 32781 8276
rect 31996 8236 32002 8248
rect 32769 8245 32781 8248
rect 32815 8245 32827 8279
rect 32769 8239 32827 8245
rect 33226 8236 33232 8288
rect 33284 8276 33290 8288
rect 33505 8279 33563 8285
rect 33505 8276 33517 8279
rect 33284 8248 33517 8276
rect 33284 8236 33290 8248
rect 33505 8245 33517 8248
rect 33551 8245 33563 8279
rect 33505 8239 33563 8245
rect 1104 8186 42504 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 42504 8186
rect 1104 8112 42504 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 2372 8044 3893 8072
rect 2372 8032 2378 8044
rect 3881 8041 3893 8044
rect 3927 8041 3939 8075
rect 3881 8035 3939 8041
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4488 8044 5028 8072
rect 4488 8032 4494 8044
rect 4525 8007 4583 8013
rect 4525 8004 4537 8007
rect 2746 7976 4537 8004
rect 1394 7896 1400 7948
rect 1452 7896 1458 7948
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2746 7936 2774 7976
rect 4525 7973 4537 7976
rect 4571 7973 4583 8007
rect 4525 7967 4583 7973
rect 1719 7908 2774 7936
rect 3145 7939 3203 7945
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 3145 7905 3157 7939
rect 3191 7905 3203 7939
rect 3145 7899 3203 7905
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 4614 7936 4620 7948
rect 3283 7908 4620 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3160 7868 3188 7899
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 4856 7908 4936 7936
rect 4856 7896 4862 7908
rect 3421 7871 3479 7877
rect 3421 7868 3433 7871
rect 3160 7840 3433 7868
rect 3421 7837 3433 7840
rect 3467 7868 3479 7871
rect 3467 7840 3740 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 2958 7800 2964 7812
rect 2898 7772 2964 7800
rect 2958 7760 2964 7772
rect 3016 7760 3022 7812
rect 3602 7800 3608 7812
rect 3528 7772 3608 7800
rect 3528 7732 3556 7772
rect 3602 7760 3608 7772
rect 3660 7760 3666 7812
rect 3712 7800 3740 7840
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 4120 7840 4261 7868
rect 4120 7828 4126 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4522 7828 4528 7880
rect 4580 7868 4586 7880
rect 4908 7877 4936 7908
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4580 7840 4721 7868
rect 4580 7828 4586 7840
rect 4709 7837 4721 7840
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 5000 7868 5028 8044
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 6144 8044 6469 8072
rect 6144 8032 6150 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 7101 8075 7159 8081
rect 7101 8072 7113 8075
rect 6880 8044 7113 8072
rect 6880 8032 6886 8044
rect 7101 8041 7113 8044
rect 7147 8041 7159 8075
rect 8018 8072 8024 8084
rect 7101 8035 7159 8041
rect 7760 8044 8024 8072
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7760 8013 7788 8044
rect 8018 8032 8024 8044
rect 8076 8072 8082 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 8076 8044 8125 8072
rect 8076 8032 8082 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 7745 8007 7803 8013
rect 7745 8004 7757 8007
rect 7432 7976 7757 8004
rect 7432 7964 7438 7976
rect 7745 7973 7757 7976
rect 7791 7973 7803 8007
rect 7745 7967 7803 7973
rect 7834 7964 7840 8016
rect 7892 7964 7898 8016
rect 8128 8004 8156 8035
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 8757 8075 8815 8081
rect 8757 8072 8769 8075
rect 8720 8044 8769 8072
rect 8720 8032 8726 8044
rect 8757 8041 8769 8044
rect 8803 8041 8815 8075
rect 8757 8035 8815 8041
rect 8772 8004 8800 8035
rect 9030 8032 9036 8084
rect 9088 8072 9094 8084
rect 9493 8075 9551 8081
rect 9493 8072 9505 8075
rect 9088 8044 9505 8072
rect 9088 8032 9094 8044
rect 9493 8041 9505 8044
rect 9539 8041 9551 8075
rect 9493 8035 9551 8041
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19886 8072 19892 8084
rect 19484 8044 19892 8072
rect 19484 8032 19490 8044
rect 19886 8032 19892 8044
rect 19944 8072 19950 8084
rect 19981 8075 20039 8081
rect 19981 8072 19993 8075
rect 19944 8044 19993 8072
rect 19944 8032 19950 8044
rect 19981 8041 19993 8044
rect 20027 8041 20039 8075
rect 19981 8035 20039 8041
rect 25222 8032 25228 8084
rect 25280 8032 25286 8084
rect 27433 8075 27491 8081
rect 27433 8041 27445 8075
rect 27479 8072 27491 8075
rect 27522 8072 27528 8084
rect 27479 8044 27528 8072
rect 27479 8041 27491 8044
rect 27433 8035 27491 8041
rect 27522 8032 27528 8044
rect 27580 8032 27586 8084
rect 28626 8032 28632 8084
rect 28684 8072 28690 8084
rect 28684 8044 29316 8072
rect 28684 8032 28690 8044
rect 8128 7976 8616 8004
rect 8772 7976 9168 8004
rect 5736 7908 6224 7936
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 5000 7840 5089 7868
rect 4893 7831 4951 7837
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 5736 7877 5764 7908
rect 5721 7871 5779 7877
rect 5721 7868 5733 7871
rect 5684 7840 5733 7868
rect 5684 7828 5690 7840
rect 5721 7837 5733 7840
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6086 7868 6092 7880
rect 5951 7840 6092 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6196 7868 6224 7908
rect 6638 7896 6644 7948
rect 6696 7896 6702 7948
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8251 7908 8432 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 6417 7871 6475 7877
rect 6417 7868 6429 7871
rect 6196 7840 6429 7868
rect 6417 7837 6429 7840
rect 6463 7837 6475 7871
rect 6417 7831 6475 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6779 7840 6837 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 6825 7837 6837 7840
rect 6871 7868 6883 7871
rect 7374 7868 7380 7880
rect 6871 7840 7380 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7834 7828 7840 7880
rect 7892 7828 7898 7880
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8404 7877 8432 7908
rect 8588 7877 8616 7976
rect 9030 7896 9036 7948
rect 9088 7896 9094 7948
rect 9140 7945 9168 7976
rect 9125 7939 9183 7945
rect 9125 7905 9137 7939
rect 9171 7905 9183 7939
rect 11425 7939 11483 7945
rect 11425 7936 11437 7939
rect 9125 7899 9183 7905
rect 10704 7908 11437 7936
rect 10704 7880 10732 7908
rect 11425 7905 11437 7908
rect 11471 7905 11483 7939
rect 11425 7899 11483 7905
rect 19334 7896 19340 7948
rect 19392 7896 19398 7948
rect 22370 7896 22376 7948
rect 22428 7896 22434 7948
rect 22465 7939 22523 7945
rect 22465 7905 22477 7939
rect 22511 7936 22523 7939
rect 23382 7936 23388 7948
rect 22511 7908 23388 7936
rect 22511 7905 22523 7908
rect 22465 7899 22523 7905
rect 23382 7896 23388 7908
rect 23440 7936 23446 7948
rect 25682 7936 25688 7948
rect 23440 7908 25688 7936
rect 23440 7896 23446 7908
rect 25682 7896 25688 7908
rect 25740 7896 25746 7948
rect 25961 7939 26019 7945
rect 25961 7905 25973 7939
rect 26007 7936 26019 7939
rect 26326 7936 26332 7948
rect 26007 7908 26332 7936
rect 26007 7905 26019 7908
rect 25961 7899 26019 7905
rect 26326 7896 26332 7908
rect 26384 7896 26390 7948
rect 27430 7896 27436 7948
rect 27488 7936 27494 7948
rect 27525 7939 27583 7945
rect 27525 7936 27537 7939
rect 27488 7908 27537 7936
rect 27488 7896 27494 7908
rect 27525 7905 27537 7908
rect 27571 7905 27583 7939
rect 27525 7899 27583 7905
rect 28902 7896 28908 7948
rect 28960 7936 28966 7948
rect 29288 7945 29316 8044
rect 30466 8032 30472 8084
rect 30524 8072 30530 8084
rect 31389 8075 31447 8081
rect 31389 8072 31401 8075
rect 30524 8044 31401 8072
rect 30524 8032 30530 8044
rect 31389 8041 31401 8044
rect 31435 8041 31447 8075
rect 32950 8072 32956 8084
rect 31389 8035 31447 8041
rect 32048 8044 32956 8072
rect 31202 7964 31208 8016
rect 31260 8004 31266 8016
rect 31297 8007 31355 8013
rect 31297 8004 31309 8007
rect 31260 7976 31309 8004
rect 31260 7964 31266 7976
rect 31297 7973 31309 7976
rect 31343 7973 31355 8007
rect 31297 7967 31355 7973
rect 28997 7939 29055 7945
rect 28997 7936 29009 7939
rect 28960 7908 29009 7936
rect 28960 7896 28966 7908
rect 28997 7905 29009 7908
rect 29043 7905 29055 7939
rect 28997 7899 29055 7905
rect 29273 7939 29331 7945
rect 29273 7905 29285 7939
rect 29319 7936 29331 7939
rect 29546 7936 29552 7948
rect 29319 7908 29552 7936
rect 29319 7905 29331 7908
rect 29273 7899 29331 7905
rect 29546 7896 29552 7908
rect 29604 7896 29610 7948
rect 29822 7896 29828 7948
rect 29880 7896 29886 7948
rect 30558 7896 30564 7948
rect 30616 7936 30622 7948
rect 31573 7939 31631 7945
rect 31573 7936 31585 7939
rect 30616 7908 31585 7936
rect 30616 7896 30622 7908
rect 31573 7905 31585 7908
rect 31619 7905 31631 7939
rect 31846 7936 31852 7948
rect 31573 7899 31631 7905
rect 31772 7908 31852 7936
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 3970 7800 3976 7812
rect 3712 7772 3976 7800
rect 3970 7760 3976 7772
rect 4028 7800 4034 7812
rect 4433 7803 4491 7809
rect 4433 7800 4445 7803
rect 4028 7772 4445 7800
rect 4028 7760 4034 7772
rect 4433 7769 4445 7772
rect 4479 7800 4491 7803
rect 4801 7803 4859 7809
rect 4801 7800 4813 7803
rect 4479 7772 4813 7800
rect 4479 7769 4491 7772
rect 4433 7763 4491 7769
rect 4801 7769 4813 7772
rect 4847 7769 4859 7803
rect 4801 7763 4859 7769
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7101 7803 7159 7809
rect 7101 7800 7113 7803
rect 6972 7772 7113 7800
rect 6972 7760 6978 7772
rect 7101 7769 7113 7772
rect 7147 7769 7159 7803
rect 7101 7763 7159 7769
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 7248 7772 7297 7800
rect 7248 7760 7254 7772
rect 7285 7769 7297 7772
rect 7331 7800 7343 7803
rect 7561 7803 7619 7809
rect 7561 7800 7573 7803
rect 7331 7772 7573 7800
rect 7331 7769 7343 7772
rect 7285 7763 7343 7769
rect 7561 7769 7573 7772
rect 7607 7800 7619 7803
rect 7607 7772 8064 7800
rect 7607 7769 7619 7772
rect 7561 7763 7619 7769
rect 3786 7732 3792 7744
rect 3528 7704 3792 7732
rect 3786 7692 3792 7704
rect 3844 7732 3850 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3844 7704 4077 7732
rect 3844 7692 3850 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4614 7732 4620 7744
rect 4212 7704 4620 7732
rect 4212 7692 4218 7704
rect 4614 7692 4620 7704
rect 4672 7732 4678 7744
rect 4890 7732 4896 7744
rect 4672 7704 4896 7732
rect 4672 7692 4678 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 5316 7704 5825 7732
rect 5316 7692 5322 7704
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6546 7732 6552 7744
rect 6319 7704 6552 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 7929 7735 7987 7741
rect 7929 7732 7941 7735
rect 7708 7704 7941 7732
rect 7708 7692 7714 7704
rect 7929 7701 7941 7704
rect 7975 7701 7987 7735
rect 8036 7732 8064 7772
rect 8110 7732 8116 7744
rect 8036 7704 8116 7732
rect 7929 7695 7987 7701
rect 8110 7692 8116 7704
rect 8168 7732 8174 7744
rect 8404 7732 8432 7831
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9306 7828 9312 7880
rect 9364 7828 9370 7880
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24228 7840 24593 7868
rect 12253 7803 12311 7809
rect 12253 7769 12265 7803
rect 12299 7769 12311 7803
rect 12253 7763 12311 7769
rect 8168 7704 8432 7732
rect 8168 7692 8174 7704
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 11606 7732 11612 7744
rect 9640 7704 11612 7732
rect 9640 7692 9646 7704
rect 11606 7692 11612 7704
rect 11664 7732 11670 7744
rect 12268 7732 12296 7763
rect 20806 7760 20812 7812
rect 20864 7800 20870 7812
rect 20864 7772 20930 7800
rect 20864 7760 20870 7772
rect 22094 7760 22100 7812
rect 22152 7760 22158 7812
rect 22741 7803 22799 7809
rect 22741 7769 22753 7803
rect 22787 7769 22799 7803
rect 24118 7800 24124 7812
rect 23966 7772 24124 7800
rect 22741 7763 22799 7769
rect 11664 7704 12296 7732
rect 11664 7692 11670 7704
rect 20622 7692 20628 7744
rect 20680 7692 20686 7744
rect 22756 7732 22784 7763
rect 24118 7760 24124 7772
rect 24176 7760 24182 7812
rect 23474 7732 23480 7744
rect 22756 7704 23480 7732
rect 23474 7692 23480 7704
rect 23532 7692 23538 7744
rect 24228 7741 24256 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 31665 7871 31723 7877
rect 31665 7837 31677 7871
rect 31711 7868 31723 7871
rect 31772 7868 31800 7908
rect 31846 7896 31852 7908
rect 31904 7896 31910 7948
rect 31938 7896 31944 7948
rect 31996 7896 32002 7948
rect 32048 7945 32076 8044
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 34425 8075 34483 8081
rect 34425 8041 34437 8075
rect 34471 8072 34483 8075
rect 34790 8072 34796 8084
rect 34471 8044 34796 8072
rect 34471 8041 34483 8044
rect 34425 8035 34483 8041
rect 34790 8032 34796 8044
rect 34848 8032 34854 8084
rect 35424 8075 35482 8081
rect 35424 8041 35436 8075
rect 35470 8072 35482 8075
rect 35894 8072 35900 8084
rect 35470 8044 35900 8072
rect 35470 8041 35482 8044
rect 35424 8035 35482 8041
rect 35894 8032 35900 8044
rect 35952 8032 35958 8084
rect 37645 8075 37703 8081
rect 37645 8041 37657 8075
rect 37691 8072 37703 8075
rect 37826 8072 37832 8084
rect 37691 8044 37832 8072
rect 37691 8041 37703 8044
rect 37645 8035 37703 8041
rect 37826 8032 37832 8044
rect 37884 8032 37890 8084
rect 32033 7939 32091 7945
rect 32033 7905 32045 7939
rect 32079 7905 32091 7939
rect 32033 7899 32091 7905
rect 32582 7896 32588 7948
rect 32640 7936 32646 7948
rect 32677 7939 32735 7945
rect 32677 7936 32689 7939
rect 32640 7908 32689 7936
rect 32640 7896 32646 7908
rect 32677 7905 32689 7908
rect 32723 7936 32735 7939
rect 34974 7936 34980 7948
rect 32723 7908 34980 7936
rect 32723 7905 32735 7908
rect 32677 7899 32735 7905
rect 34974 7896 34980 7908
rect 35032 7936 35038 7948
rect 35161 7939 35219 7945
rect 35161 7936 35173 7939
rect 35032 7908 35173 7936
rect 35032 7896 35038 7908
rect 35161 7905 35173 7908
rect 35207 7936 35219 7939
rect 35434 7936 35440 7948
rect 35207 7908 35440 7936
rect 35207 7905 35219 7908
rect 35161 7899 35219 7905
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 36909 7939 36967 7945
rect 36909 7905 36921 7939
rect 36955 7936 36967 7939
rect 37001 7939 37059 7945
rect 37001 7936 37013 7939
rect 36955 7908 37013 7936
rect 36955 7905 36967 7908
rect 36909 7899 36967 7905
rect 37001 7905 37013 7908
rect 37047 7905 37059 7939
rect 37001 7899 37059 7905
rect 32125 7871 32183 7877
rect 32125 7868 32137 7871
rect 31711 7840 31800 7868
rect 31864 7840 32137 7868
rect 31711 7837 31723 7840
rect 31665 7831 31723 7837
rect 27338 7800 27344 7812
rect 27186 7772 27344 7800
rect 27338 7760 27344 7772
rect 27396 7800 27402 7812
rect 27396 7772 27830 7800
rect 27396 7760 27402 7772
rect 29362 7760 29368 7812
rect 29420 7800 29426 7812
rect 31864 7800 31892 7840
rect 32125 7837 32137 7840
rect 32171 7837 32183 7871
rect 32125 7831 32183 7837
rect 29420 7772 30314 7800
rect 31726 7772 31892 7800
rect 29420 7760 29426 7772
rect 24213 7735 24271 7741
rect 24213 7701 24225 7735
rect 24259 7701 24271 7735
rect 30208 7732 30236 7772
rect 31570 7732 31576 7744
rect 30208 7704 31576 7732
rect 24213 7695 24271 7701
rect 31570 7692 31576 7704
rect 31628 7732 31634 7744
rect 31726 7732 31754 7772
rect 32490 7760 32496 7812
rect 32548 7760 32554 7812
rect 32953 7803 33011 7809
rect 32953 7769 32965 7803
rect 32999 7800 33011 7803
rect 33226 7800 33232 7812
rect 32999 7772 33232 7800
rect 32999 7769 33011 7772
rect 32953 7763 33011 7769
rect 33226 7760 33232 7772
rect 33284 7760 33290 7812
rect 35894 7800 35900 7812
rect 33336 7772 33442 7800
rect 35176 7772 35900 7800
rect 31628 7704 31754 7732
rect 31628 7692 31634 7704
rect 33134 7692 33140 7744
rect 33192 7732 33198 7744
rect 33336 7732 33364 7772
rect 35176 7732 35204 7772
rect 35894 7760 35900 7772
rect 35952 7760 35958 7812
rect 33192 7704 35204 7732
rect 33192 7692 33198 7704
rect 1104 7642 42504 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 42504 7642
rect 1104 7568 42504 7590
rect 2682 7488 2688 7540
rect 2740 7488 2746 7540
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3375 7500 4384 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 4154 7460 4160 7472
rect 3712 7432 4160 7460
rect 2314 7352 2320 7404
rect 2372 7352 2378 7404
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 2682 7392 2688 7404
rect 2547 7364 2688 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2424 7256 2452 7355
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 3712 7401 3740 7432
rect 4154 7420 4160 7432
rect 4212 7420 4218 7472
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3007 7364 3709 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3786 7352 3792 7404
rect 3844 7352 3850 7404
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 3970 7392 3976 7404
rect 3927 7364 3976 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 3053 7327 3111 7333
rect 3053 7293 3065 7327
rect 3099 7324 3111 7327
rect 3099 7296 3556 7324
rect 3099 7293 3111 7296
rect 3053 7287 3111 7293
rect 3421 7259 3479 7265
rect 3421 7256 3433 7259
rect 2424 7228 3433 7256
rect 3421 7225 3433 7228
rect 3467 7225 3479 7259
rect 3528 7256 3556 7296
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 4080 7324 4108 7355
rect 4246 7352 4252 7404
rect 4304 7352 4310 7404
rect 4356 7401 4384 7500
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4580 7500 4752 7528
rect 4580 7488 4586 7500
rect 4614 7420 4620 7472
rect 4672 7420 4678 7472
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 4724 7401 4752 7500
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8297 7531 8355 7537
rect 8297 7528 8309 7531
rect 8260 7500 8309 7528
rect 8260 7488 8266 7500
rect 8297 7497 8309 7500
rect 8343 7497 8355 7531
rect 8297 7491 8355 7497
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 19208 7500 19257 7528
rect 19208 7488 19214 7500
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 19245 7491 19303 7497
rect 21637 7531 21695 7537
rect 21637 7497 21649 7531
rect 21683 7528 21695 7531
rect 21818 7528 21824 7540
rect 21683 7500 21824 7528
rect 21683 7497 21695 7500
rect 21637 7491 21695 7497
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 22094 7488 22100 7540
rect 22152 7528 22158 7540
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 22152 7500 22569 7528
rect 22152 7488 22158 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 22557 7491 22615 7497
rect 23937 7531 23995 7537
rect 23937 7497 23949 7531
rect 23983 7528 23995 7531
rect 24394 7528 24400 7540
rect 23983 7500 24400 7528
rect 23983 7497 23995 7500
rect 23937 7491 23995 7497
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 24486 7488 24492 7540
rect 24544 7528 24550 7540
rect 27338 7528 27344 7540
rect 24544 7500 27344 7528
rect 24544 7488 24550 7500
rect 7190 7420 7196 7472
rect 7248 7420 7254 7472
rect 8128 7460 8156 7488
rect 8846 7460 8852 7472
rect 8128 7432 8432 7460
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 3660 7296 4108 7324
rect 4724 7324 4752 7355
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5316 7364 6316 7392
rect 5316 7352 5322 7364
rect 5626 7324 5632 7336
rect 4724 7296 5632 7324
rect 3660 7284 3666 7296
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 4706 7256 4712 7268
rect 3528 7228 4108 7256
rect 3421 7219 3479 7225
rect 4080 7188 4108 7228
rect 4264 7228 4712 7256
rect 4157 7191 4215 7197
rect 4157 7188 4169 7191
rect 4080 7160 4169 7188
rect 4157 7157 4169 7160
rect 4203 7188 4215 7191
rect 4264 7188 4292 7228
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 4816 7228 5120 7256
rect 4203 7160 4292 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4816 7188 4844 7228
rect 4580 7160 4844 7188
rect 4580 7148 4586 7160
rect 4890 7148 4896 7200
rect 4948 7148 4954 7200
rect 5092 7197 5120 7228
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5258 7188 5264 7200
rect 5123 7160 5264 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 6288 7188 6316 7364
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8404 7401 8432 7432
rect 8496 7432 8852 7460
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8076 7364 8217 7392
rect 8076 7352 8082 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8389 7395 8447 7401
rect 8389 7361 8401 7395
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 6362 7284 6368 7336
rect 6420 7284 6426 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7190 7324 7196 7336
rect 6687 7296 7196 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 8496 7324 8524 7432
rect 8846 7420 8852 7432
rect 8904 7460 8910 7472
rect 9277 7463 9335 7469
rect 9277 7460 9289 7463
rect 8904 7432 9289 7460
rect 8904 7420 8910 7432
rect 9277 7429 9289 7432
rect 9323 7429 9335 7463
rect 9277 7423 9335 7429
rect 9490 7420 9496 7472
rect 9548 7420 9554 7472
rect 11146 7420 11152 7472
rect 11204 7420 11210 7472
rect 19794 7420 19800 7472
rect 19852 7420 19858 7472
rect 19886 7420 19892 7472
rect 19944 7420 19950 7472
rect 21266 7420 21272 7472
rect 21324 7420 21330 7472
rect 21358 7420 21364 7472
rect 21416 7420 21422 7472
rect 22465 7463 22523 7469
rect 22465 7460 22477 7463
rect 22066 7432 22477 7460
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11664 7364 11713 7392
rect 11664 7352 11670 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 12124 7364 12265 7392
rect 12124 7352 12130 7364
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7392 19579 7395
rect 19702 7392 19708 7404
rect 19567 7364 19708 7392
rect 19567 7361 19579 7364
rect 19521 7355 19579 7361
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 20956 7364 21097 7392
rect 20956 7352 20962 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 22066 7392 22094 7432
rect 22465 7429 22477 7432
rect 22511 7460 22523 7463
rect 23109 7463 23167 7469
rect 23109 7460 23121 7463
rect 22511 7432 23121 7460
rect 22511 7429 22523 7432
rect 22465 7423 22523 7429
rect 23109 7429 23121 7432
rect 23155 7429 23167 7463
rect 23109 7423 23167 7429
rect 23198 7420 23204 7472
rect 23256 7460 23262 7472
rect 24026 7460 24032 7472
rect 23256 7432 24032 7460
rect 23256 7420 23262 7432
rect 24026 7420 24032 7432
rect 24084 7420 24090 7472
rect 25056 7460 25084 7500
rect 27338 7488 27344 7500
rect 27396 7488 27402 7540
rect 28626 7488 28632 7540
rect 28684 7488 28690 7540
rect 29178 7488 29184 7540
rect 29236 7528 29242 7540
rect 29825 7531 29883 7537
rect 29825 7528 29837 7531
rect 29236 7500 29837 7528
rect 29236 7488 29242 7500
rect 29825 7497 29837 7500
rect 29871 7497 29883 7531
rect 29825 7491 29883 7497
rect 33229 7531 33287 7537
rect 33229 7497 33241 7531
rect 33275 7528 33287 7531
rect 34054 7528 34060 7540
rect 33275 7500 34060 7528
rect 33275 7497 33287 7500
rect 33229 7491 33287 7497
rect 34054 7488 34060 7500
rect 34112 7488 34118 7540
rect 35342 7488 35348 7540
rect 35400 7488 35406 7540
rect 35434 7488 35440 7540
rect 35492 7528 35498 7540
rect 35492 7500 37044 7528
rect 35492 7488 35498 7500
rect 24978 7432 25084 7460
rect 25406 7420 25412 7472
rect 25464 7420 25470 7472
rect 28644 7460 28672 7488
rect 28000 7432 28672 7460
rect 21499 7364 22094 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 22830 7352 22836 7404
rect 22888 7352 22894 7404
rect 23842 7392 23848 7404
rect 23124 7364 23848 7392
rect 11885 7327 11943 7333
rect 11885 7324 11897 7327
rect 7432 7296 8524 7324
rect 9140 7296 11897 7324
rect 7432 7284 7438 7296
rect 9140 7200 9168 7296
rect 11716 7268 11744 7296
rect 11885 7293 11897 7296
rect 11931 7293 11943 7327
rect 11885 7287 11943 7293
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12342 7324 12348 7336
rect 12023 7296 12348 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 20622 7284 20628 7336
rect 20680 7324 20686 7336
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 20680 7296 21833 7324
rect 20680 7284 20686 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 23124 7324 23152 7364
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 25682 7352 25688 7404
rect 25740 7352 25746 7404
rect 28000 7401 28028 7432
rect 33134 7420 33140 7472
rect 33192 7460 33198 7472
rect 33192 7432 33534 7460
rect 33192 7420 33198 7432
rect 34698 7420 34704 7472
rect 34756 7420 34762 7472
rect 36078 7420 36084 7472
rect 36136 7420 36142 7472
rect 37016 7460 37044 7500
rect 37016 7432 37136 7460
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7361 27491 7395
rect 27433 7355 27491 7361
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 22787 7296 23152 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11517 7259 11575 7265
rect 11517 7256 11529 7259
rect 11112 7228 11529 7256
rect 11112 7216 11118 7228
rect 11517 7225 11529 7228
rect 11563 7225 11575 7259
rect 11517 7219 11575 7225
rect 11698 7216 11704 7268
rect 11756 7216 11762 7268
rect 8662 7188 8668 7200
rect 6288 7160 8668 7188
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 9122 7148 9128 7200
rect 9180 7148 9186 7200
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 9272 7160 9321 7188
rect 9272 7148 9278 7160
rect 9309 7157 9321 7160
rect 9355 7157 9367 7191
rect 9309 7151 9367 7157
rect 11238 7148 11244 7200
rect 11296 7148 11302 7200
rect 12158 7148 12164 7200
rect 12216 7148 12222 7200
rect 19702 7148 19708 7200
rect 19760 7188 19766 7200
rect 22756 7188 22784 7287
rect 19760 7160 22784 7188
rect 27448 7188 27476 7355
rect 29362 7352 29368 7404
rect 29420 7352 29426 7404
rect 34974 7352 34980 7404
rect 35032 7352 35038 7404
rect 37108 7401 37136 7432
rect 37093 7395 37151 7401
rect 37093 7361 37105 7395
rect 37139 7361 37151 7395
rect 37093 7355 37151 7361
rect 28258 7284 28264 7336
rect 28316 7284 28322 7336
rect 29733 7327 29791 7333
rect 29733 7293 29745 7327
rect 29779 7324 29791 7327
rect 30377 7327 30435 7333
rect 30377 7324 30389 7327
rect 29779 7296 30389 7324
rect 29779 7293 29791 7296
rect 29733 7287 29791 7293
rect 30377 7293 30389 7296
rect 30423 7293 30435 7327
rect 30377 7287 30435 7293
rect 36817 7327 36875 7333
rect 36817 7293 36829 7327
rect 36863 7324 36875 7327
rect 37734 7324 37740 7336
rect 36863 7296 37740 7324
rect 36863 7293 36875 7296
rect 36817 7287 36875 7293
rect 37734 7284 37740 7296
rect 37792 7284 37798 7336
rect 29748 7228 31754 7256
rect 29748 7188 29776 7228
rect 27448 7160 29776 7188
rect 31726 7188 31754 7228
rect 32490 7188 32496 7200
rect 31726 7160 32496 7188
rect 19760 7148 19766 7160
rect 32490 7148 32496 7160
rect 32548 7148 32554 7200
rect 1104 7098 42504 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 42504 7098
rect 1104 7024 42504 7046
rect 4157 6987 4215 6993
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4614 6984 4620 6996
rect 4203 6956 4620 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 4890 6944 4896 6996
rect 4948 6984 4954 6996
rect 5641 6987 5699 6993
rect 5641 6984 5653 6987
rect 4948 6956 5653 6984
rect 4948 6944 4954 6956
rect 5641 6953 5653 6956
rect 5687 6953 5699 6987
rect 5641 6947 5699 6953
rect 9217 6987 9275 6993
rect 9217 6953 9229 6987
rect 9263 6984 9275 6987
rect 9306 6984 9312 6996
rect 9263 6956 9312 6984
rect 9263 6953 9275 6956
rect 9217 6947 9275 6953
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9401 6987 9459 6993
rect 9401 6953 9413 6987
rect 9447 6984 9459 6987
rect 9858 6984 9864 6996
rect 9447 6956 9864 6984
rect 9447 6953 9459 6956
rect 9401 6947 9459 6953
rect 9858 6944 9864 6956
rect 9916 6984 9922 6996
rect 12066 6984 12072 6996
rect 9916 6956 12072 6984
rect 9916 6944 9922 6956
rect 12066 6944 12072 6956
rect 12124 6984 12130 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 12124 6956 12449 6984
rect 12124 6944 12130 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 7282 6916 7288 6928
rect 6144 6888 7288 6916
rect 6144 6876 6150 6888
rect 7282 6876 7288 6888
rect 7340 6876 7346 6928
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 9582 6848 9588 6860
rect 6052 6820 9588 6848
rect 6052 6808 6058 6820
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 11756 6820 12434 6848
rect 11756 6808 11762 6820
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 6362 6780 6368 6792
rect 5951 6752 6368 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6362 6740 6368 6752
rect 6420 6780 6426 6792
rect 6822 6780 6828 6792
rect 6420 6752 6828 6780
rect 6420 6740 6426 6752
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6749 6975 6783
rect 6917 6743 6975 6749
rect 6086 6712 6092 6724
rect 5198 6684 6092 6712
rect 2958 6604 2964 6656
rect 3016 6644 3022 6656
rect 3510 6644 3516 6656
rect 3016 6616 3516 6644
rect 3016 6604 3022 6616
rect 3510 6604 3516 6616
rect 3568 6644 3574 6656
rect 5276 6644 5304 6684
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 6546 6672 6552 6724
rect 6604 6672 6610 6724
rect 6932 6712 6960 6743
rect 7006 6740 7012 6792
rect 7064 6740 7070 6792
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9677 6783 9735 6789
rect 9677 6780 9689 6783
rect 9600 6752 9689 6780
rect 9600 6724 9628 6752
rect 9677 6749 9689 6752
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 12406 6780 12434 6820
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12406 6752 12541 6780
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12986 6740 12992 6792
rect 13044 6740 13050 6792
rect 7098 6712 7104 6724
rect 6932 6684 7104 6712
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 9582 6672 9588 6724
rect 9640 6672 9646 6724
rect 10226 6672 10232 6724
rect 10284 6712 10290 6724
rect 10284 6684 10548 6712
rect 10284 6672 10290 6684
rect 3568 6616 5304 6644
rect 3568 6604 3574 6616
rect 9030 6604 9036 6656
rect 9088 6604 9094 6656
rect 9385 6647 9443 6653
rect 9385 6613 9397 6647
rect 9431 6644 9443 6647
rect 9674 6644 9680 6656
rect 9431 6616 9680 6644
rect 9431 6613 9443 6616
rect 9385 6607 9443 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 9824 6616 10333 6644
rect 9824 6604 9830 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10520 6644 10548 6684
rect 10594 6672 10600 6724
rect 10652 6712 10658 6724
rect 10965 6715 11023 6721
rect 10965 6712 10977 6715
rect 10652 6684 10977 6712
rect 10652 6672 10658 6684
rect 10965 6681 10977 6684
rect 11011 6681 11023 6715
rect 11422 6712 11428 6724
rect 10965 6675 11023 6681
rect 11072 6684 11428 6712
rect 11072 6644 11100 6684
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 12268 6684 12756 6712
rect 10520 6616 11100 6644
rect 10321 6607 10379 6613
rect 11606 6604 11612 6656
rect 11664 6644 11670 6656
rect 12268 6644 12296 6684
rect 11664 6616 12296 6644
rect 11664 6604 11670 6616
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12728 6653 12756 6684
rect 12621 6647 12679 6653
rect 12621 6644 12633 6647
rect 12400 6616 12633 6644
rect 12400 6604 12406 6616
rect 12621 6613 12633 6616
rect 12667 6613 12679 6647
rect 12621 6607 12679 6613
rect 12713 6647 12771 6653
rect 12713 6613 12725 6647
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 1104 6554 42504 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 42504 6554
rect 1104 6480 42504 6502
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 8352 6412 9505 6440
rect 8352 6400 8358 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 11149 6443 11207 6449
rect 11149 6440 11161 6443
rect 9732 6412 11161 6440
rect 9732 6400 9738 6412
rect 11149 6409 11161 6412
rect 11195 6440 11207 6443
rect 11882 6440 11888 6452
rect 11195 6412 11888 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11882 6400 11888 6412
rect 11940 6440 11946 6452
rect 12342 6440 12348 6452
rect 11940 6412 12348 6440
rect 11940 6400 11946 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 9692 6372 9720 6400
rect 10226 6372 10232 6384
rect 9692 6344 9812 6372
rect 9062 6276 9628 6304
rect 6822 6196 6828 6248
rect 6880 6236 6886 6248
rect 7653 6239 7711 6245
rect 7653 6236 7665 6239
rect 6880 6208 7665 6236
rect 6880 6196 6886 6208
rect 7653 6205 7665 6208
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 9490 6236 9496 6248
rect 7975 6208 9496 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 9490 6196 9496 6208
rect 9548 6196 9554 6248
rect 9600 6236 9628 6276
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 9784 6313 9812 6344
rect 9876 6344 10232 6372
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 9876 6236 9904 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 12158 6372 12164 6384
rect 10428 6344 12164 6372
rect 9950 6264 9956 6316
rect 10008 6264 10014 6316
rect 10428 6313 10456 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 9600 6208 9904 6236
rect 10152 6236 10180 6267
rect 10594 6264 10600 6316
rect 10652 6264 10658 6316
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11054 6304 11060 6316
rect 11011 6276 11060 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 11238 6264 11244 6316
rect 11296 6264 11302 6316
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 11882 6264 11888 6316
rect 11940 6264 11946 6316
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12066 6304 12072 6316
rect 12023 6276 12072 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 10152 6208 11529 6236
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 11848 6208 12434 6236
rect 11848 6196 11854 6208
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 10042 6168 10048 6180
rect 9088 6140 10048 6168
rect 9088 6128 9094 6140
rect 10042 6128 10048 6140
rect 10100 6128 10106 6180
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 9401 6103 9459 6109
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 9582 6100 9588 6112
rect 9447 6072 9588 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9858 6060 9864 6112
rect 9916 6060 9922 6112
rect 10244 6100 10272 6131
rect 10318 6128 10324 6180
rect 10376 6128 10382 6180
rect 11606 6168 11612 6180
rect 10704 6140 11612 6168
rect 10704 6100 10732 6140
rect 11606 6128 11612 6140
rect 11664 6128 11670 6180
rect 12406 6168 12434 6208
rect 12986 6168 12992 6180
rect 12406 6140 12992 6168
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 10244 6072 10732 6100
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 10870 6100 10876 6112
rect 10827 6072 10876 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 1104 6010 42504 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 42504 6010
rect 1104 5936 42504 5958
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 4801 5899 4859 5905
rect 4801 5896 4813 5899
rect 4488 5868 4813 5896
rect 4488 5856 4494 5868
rect 4801 5865 4813 5868
rect 4847 5896 4859 5899
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4847 5868 5089 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 5077 5859 5135 5865
rect 5537 5899 5595 5905
rect 5537 5865 5549 5899
rect 5583 5896 5595 5899
rect 5718 5896 5724 5908
rect 5583 5868 5724 5896
rect 5583 5865 5595 5868
rect 5537 5859 5595 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9217 5899 9275 5905
rect 9217 5896 9229 5899
rect 8996 5868 9229 5896
rect 8996 5856 9002 5868
rect 9217 5865 9229 5868
rect 9263 5865 9275 5899
rect 9217 5859 9275 5865
rect 9490 5856 9496 5908
rect 9548 5856 9554 5908
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 9858 5896 9864 5908
rect 9640 5868 9864 5896
rect 9640 5856 9646 5868
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 11238 5896 11244 5908
rect 10376 5868 11244 5896
rect 10376 5856 10382 5868
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 12342 5856 12348 5908
rect 12400 5856 12406 5908
rect 2314 5828 2320 5840
rect 2240 5800 2320 5828
rect 2240 5769 2268 5800
rect 2314 5788 2320 5800
rect 2372 5828 2378 5840
rect 2372 5800 2774 5828
rect 2372 5788 2378 5800
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5729 2283 5763
rect 2225 5723 2283 5729
rect 2501 5763 2559 5769
rect 2501 5729 2513 5763
rect 2547 5760 2559 5763
rect 2746 5760 2774 5800
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 5316 5800 5488 5828
rect 5316 5788 5322 5800
rect 2547 5732 2636 5760
rect 2746 5732 4568 5760
rect 2547 5729 2559 5732
rect 2501 5723 2559 5729
rect 2130 5652 2136 5704
rect 2188 5652 2194 5704
rect 2608 5701 2636 5732
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5661 2651 5695
rect 2593 5655 2651 5661
rect 2682 5652 2688 5704
rect 2740 5652 2746 5704
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2832 5664 2881 5692
rect 2832 5652 2838 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4338 5692 4344 5704
rect 4295 5664 4344 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4338 5652 4344 5664
rect 4396 5652 4402 5704
rect 4540 5701 4568 5732
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 2148 5624 2176 5652
rect 4430 5624 4436 5636
rect 2148 5596 4436 5624
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 4540 5624 4568 5655
rect 4890 5652 4896 5704
rect 4948 5692 4954 5704
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 4948 5664 5089 5692
rect 4948 5652 4954 5664
rect 5077 5661 5089 5664
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 4769 5627 4827 5633
rect 4769 5624 4781 5627
rect 4540 5596 4781 5624
rect 4769 5593 4781 5596
rect 4815 5593 4827 5627
rect 4769 5587 4827 5593
rect 4982 5584 4988 5636
rect 5040 5624 5046 5636
rect 5368 5624 5396 5655
rect 5040 5596 5396 5624
rect 5460 5624 5488 5800
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 6748 5732 7113 5760
rect 6748 5701 6776 5732
rect 7101 5729 7113 5732
rect 7147 5729 7159 5763
rect 9214 5760 9220 5772
rect 7101 5723 7159 5729
rect 9048 5732 9220 5760
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7300 5624 7328 5655
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9048 5701 9076 5732
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 10336 5760 10364 5856
rect 9692 5732 10364 5760
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8904 5664 8953 5692
rect 8904 5652 8910 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9490 5692 9496 5704
rect 9033 5655 9091 5661
rect 9140 5664 9496 5692
rect 9140 5624 9168 5664
rect 9490 5652 9496 5664
rect 9548 5692 9554 5704
rect 9692 5701 9720 5732
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9548 5664 9689 5692
rect 9548 5652 9554 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 10594 5652 10600 5704
rect 10652 5652 10658 5704
rect 5460 5596 6960 5624
rect 7300 5596 9168 5624
rect 9217 5627 9275 5633
rect 5040 5584 5046 5596
rect 6932 5568 6960 5596
rect 9217 5593 9229 5627
rect 9263 5624 9275 5627
rect 9398 5624 9404 5636
rect 9263 5596 9404 5624
rect 9263 5593 9275 5596
rect 9217 5587 9275 5593
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 9861 5627 9919 5633
rect 9861 5593 9873 5627
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 2958 5516 2964 5568
rect 3016 5556 3022 5568
rect 3053 5559 3111 5565
rect 3053 5556 3065 5559
rect 3016 5528 3065 5556
rect 3016 5516 3022 5528
rect 3053 5525 3065 5528
rect 3099 5525 3111 5559
rect 3053 5519 3111 5525
rect 4065 5559 4123 5565
rect 4065 5525 4077 5559
rect 4111 5556 4123 5559
rect 4154 5556 4160 5568
rect 4111 5528 4160 5556
rect 4111 5525 4123 5528
rect 4065 5519 4123 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4617 5559 4675 5565
rect 4617 5556 4629 5559
rect 4304 5528 4629 5556
rect 4304 5516 4310 5528
rect 4617 5525 4629 5528
rect 4663 5525 4675 5559
rect 4617 5519 4675 5525
rect 6546 5516 6552 5568
rect 6604 5516 6610 5568
rect 6914 5516 6920 5568
rect 6972 5516 6978 5568
rect 8662 5516 8668 5568
rect 8720 5556 8726 5568
rect 9876 5556 9904 5587
rect 10870 5584 10876 5636
rect 10928 5584 10934 5636
rect 11422 5584 11428 5636
rect 11480 5584 11486 5636
rect 11514 5556 11520 5568
rect 8720 5528 11520 5556
rect 8720 5516 8726 5528
rect 11514 5516 11520 5528
rect 11572 5556 11578 5568
rect 11790 5556 11796 5568
rect 11572 5528 11796 5556
rect 11572 5516 11578 5528
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 1104 5466 42504 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 42504 5466
rect 1104 5392 42504 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 4338 5352 4344 5364
rect 2547 5324 4344 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 9309 5355 9367 5361
rect 9309 5321 9321 5355
rect 9355 5352 9367 5355
rect 9398 5352 9404 5364
rect 9355 5324 9404 5352
rect 9355 5321 9367 5324
rect 9309 5315 9367 5321
rect 9398 5312 9404 5324
rect 9456 5352 9462 5364
rect 9858 5352 9864 5364
rect 9456 5324 9864 5352
rect 9456 5312 9462 5324
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10137 5355 10195 5361
rect 10137 5352 10149 5355
rect 10008 5324 10149 5352
rect 10008 5312 10014 5324
rect 10137 5321 10149 5324
rect 10183 5321 10195 5355
rect 10137 5315 10195 5321
rect 3510 5244 3516 5296
rect 3568 5244 3574 5296
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 3936 5256 4292 5284
rect 3936 5244 3942 5256
rect 2222 5176 2228 5228
rect 2280 5176 2286 5228
rect 4264 5225 4292 5256
rect 5994 5244 6000 5296
rect 6052 5244 6058 5296
rect 6546 5244 6552 5296
rect 6604 5284 6610 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 6604 5256 6653 5284
rect 6604 5244 6610 5256
rect 6641 5253 6653 5256
rect 6687 5253 6699 5287
rect 6641 5247 6699 5253
rect 7282 5244 7288 5296
rect 7340 5244 7346 5296
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 11885 5287 11943 5293
rect 8904 5256 10548 5284
rect 8904 5244 8910 5256
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5216 4307 5219
rect 4295 5188 5304 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 2041 5151 2099 5157
rect 2041 5148 2053 5151
rect 1452 5120 2053 5148
rect 1452 5108 1458 5120
rect 2041 5117 2053 5120
rect 2087 5148 2099 5151
rect 2130 5148 2136 5160
rect 2087 5120 2136 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2774 5148 2780 5160
rect 2455 5120 2780 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3973 5151 4031 5157
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4019 5120 4292 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 4264 5080 4292 5120
rect 4338 5108 4344 5160
rect 4396 5148 4402 5160
rect 4706 5148 4712 5160
rect 4396 5120 4712 5148
rect 4396 5108 4402 5120
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5276 5157 5304 5188
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 9180 5188 9229 5216
rect 9180 5176 9186 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 9217 5179 9275 5185
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 9582 5216 9588 5228
rect 9447 5188 9588 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 9766 5216 9772 5228
rect 9723 5188 9772 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 9858 5176 9864 5228
rect 9916 5176 9922 5228
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5534 5148 5540 5160
rect 5307 5120 5540 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5534 5108 5540 5120
rect 5592 5148 5598 5160
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 5592 5120 6377 5148
rect 5592 5108 5598 5120
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 9968 5148 9996 5179
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10520 5225 10548 5256
rect 11885 5253 11897 5287
rect 11931 5284 11943 5287
rect 11974 5284 11980 5296
rect 11931 5256 11980 5284
rect 11931 5253 11943 5256
rect 11885 5247 11943 5253
rect 11974 5244 11980 5256
rect 12032 5244 12038 5296
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10100 5188 10241 5216
rect 10100 5176 10106 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 6365 5111 6423 5117
rect 9416 5120 9996 5148
rect 4614 5080 4620 5092
rect 4264 5052 4620 5080
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 4246 5012 4252 5024
rect 3844 4984 4252 5012
rect 3844 4972 3850 4984
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 4890 5012 4896 5024
rect 4488 4984 4896 5012
rect 4488 4972 4494 4984
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 4985 5015 5043 5021
rect 4985 4981 4997 5015
rect 5031 5012 5043 5015
rect 5350 5012 5356 5024
rect 5031 4984 5356 5012
rect 5031 4981 5043 4984
rect 4985 4975 5043 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 6380 5012 6408 5111
rect 9033 5083 9091 5089
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9416 5080 9444 5120
rect 10428 5080 10456 5179
rect 9079 5052 9444 5080
rect 9784 5052 10456 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 6822 5012 6828 5024
rect 6380 4984 6828 5012
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 7432 4984 8125 5012
rect 7432 4972 7438 4984
rect 8113 4981 8125 4984
rect 8159 5012 8171 5015
rect 9048 5012 9076 5043
rect 9214 5012 9220 5024
rect 8159 4984 9220 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 9585 5015 9643 5021
rect 9585 5012 9597 5015
rect 9364 4984 9597 5012
rect 9364 4972 9370 4984
rect 9585 4981 9597 4984
rect 9631 5012 9643 5015
rect 9784 5012 9812 5052
rect 9631 4984 9812 5012
rect 9631 4981 9643 4984
rect 9585 4975 9643 4981
rect 9858 4972 9864 5024
rect 9916 4972 9922 5024
rect 10226 4972 10232 5024
rect 10284 4972 10290 5024
rect 10778 4972 10784 5024
rect 10836 5012 10842 5024
rect 11793 5015 11851 5021
rect 11793 5012 11805 5015
rect 10836 4984 11805 5012
rect 10836 4972 10842 4984
rect 11793 4981 11805 4984
rect 11839 5012 11851 5015
rect 12434 5012 12440 5024
rect 11839 4984 12440 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 1104 4922 42504 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 42504 4922
rect 1104 4848 42504 4870
rect 1394 4768 1400 4820
rect 1452 4768 1458 4820
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 3510 4808 3516 4820
rect 2464 4780 3516 4808
rect 2464 4768 2470 4780
rect 3510 4768 3516 4780
rect 3568 4768 3574 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4120 4780 4169 4808
rect 4120 4768 4126 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5442 4808 5448 4820
rect 5031 4780 5448 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 7006 4768 7012 4820
rect 7064 4768 7070 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 9125 4811 9183 4817
rect 7524 4780 9076 4808
rect 7524 4768 7530 4780
rect 4433 4743 4491 4749
rect 4433 4709 4445 4743
rect 4479 4740 4491 4743
rect 4706 4740 4712 4752
rect 4479 4712 4712 4740
rect 4479 4709 4491 4712
rect 4433 4703 4491 4709
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 7282 4740 7288 4752
rect 5960 4712 7288 4740
rect 5960 4700 5966 4712
rect 7282 4700 7288 4712
rect 7340 4700 7346 4752
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8665 4743 8723 4749
rect 8665 4740 8677 4743
rect 8352 4712 8677 4740
rect 8352 4700 8358 4712
rect 8665 4709 8677 4712
rect 8711 4709 8723 4743
rect 9048 4740 9076 4780
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9398 4808 9404 4820
rect 9171 4780 9404 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10042 4808 10048 4820
rect 9999 4780 10048 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10778 4740 10784 4752
rect 9048 4712 10784 4740
rect 8665 4703 8723 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 3878 4672 3884 4684
rect 3191 4644 3884 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 4890 4672 4896 4684
rect 4632 4644 4896 4672
rect 3786 4564 3792 4616
rect 3844 4604 3850 4616
rect 4246 4604 4252 4616
rect 3844 4576 4252 4604
rect 3844 4564 3850 4576
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 4632 4613 4660 4644
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 6733 4675 6791 4681
rect 6733 4641 6745 4675
rect 6779 4672 6791 4675
rect 8846 4672 8852 4684
rect 6779 4644 8852 4672
rect 6779 4641 6791 4644
rect 6733 4635 6791 4641
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 7374 4604 7380 4616
rect 6687 4576 7380 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 7374 4564 7380 4576
rect 7432 4604 7438 4616
rect 8404 4613 8432 4644
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9784 4644 10333 4672
rect 8389 4607 8447 4613
rect 7432 4576 8340 4604
rect 7432 4564 7438 4576
rect 2406 4496 2412 4548
rect 2464 4496 2470 4548
rect 2869 4539 2927 4545
rect 2869 4505 2881 4539
rect 2915 4536 2927 4539
rect 2958 4536 2964 4548
rect 2915 4508 2964 4536
rect 2915 4505 2927 4508
rect 2869 4499 2927 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 4157 4539 4215 4545
rect 4157 4505 4169 4539
rect 4203 4536 4215 4539
rect 4430 4536 4436 4548
rect 4203 4508 4436 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 4172 4468 4200 4499
rect 4430 4496 4436 4508
rect 4488 4496 4494 4548
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4536 4767 4539
rect 5276 4536 5304 4564
rect 4755 4508 5304 4536
rect 4755 4505 4767 4508
rect 4709 4499 4767 4505
rect 4816 4480 4844 4508
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 8312 4536 8340 4576
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 8665 4607 8723 4613
rect 8435 4576 8469 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9398 4604 9404 4616
rect 8711 4576 9404 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9784 4613 9812 4644
rect 10321 4641 10333 4644
rect 10367 4672 10379 4675
rect 10410 4672 10416 4684
rect 10367 4644 10416 4672
rect 10367 4641 10379 4644
rect 10321 4635 10379 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 10594 4632 10600 4684
rect 10652 4672 10658 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 10652 4644 12081 4672
rect 10652 4632 10658 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9732 4576 9781 4604
rect 9732 4564 9738 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 9950 4564 9956 4616
rect 10008 4564 10014 4616
rect 10045 4607 10103 4613
rect 10045 4573 10057 4607
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4604 10287 4607
rect 10502 4604 10508 4616
rect 10275 4576 10508 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 8481 4539 8539 4545
rect 8481 4536 8493 4539
rect 8312 4508 8493 4536
rect 8481 4505 8493 4508
rect 8527 4505 8539 4539
rect 8481 4499 8539 4505
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 9093 4539 9151 4545
rect 9093 4536 9105 4539
rect 8904 4508 9105 4536
rect 8904 4496 8910 4508
rect 9093 4505 9105 4508
rect 9139 4505 9151 4539
rect 9093 4499 9151 4505
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 9272 4508 9321 4536
rect 9272 4496 9278 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9309 4499 9367 4505
rect 9582 4496 9588 4548
rect 9640 4536 9646 4548
rect 10060 4536 10088 4567
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12492 4576 12541 4604
rect 12492 4564 12498 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 9640 4508 10088 4536
rect 10137 4539 10195 4545
rect 9640 4496 9646 4508
rect 10137 4505 10149 4539
rect 10183 4536 10195 4539
rect 10183 4508 10548 4536
rect 10183 4505 10195 4508
rect 10137 4499 10195 4505
rect 2740 4440 4200 4468
rect 2740 4428 2746 4440
rect 4338 4428 4344 4480
rect 4396 4428 4402 4480
rect 4798 4428 4804 4480
rect 4856 4428 4862 4480
rect 8570 4428 8576 4480
rect 8628 4468 8634 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8628 4440 8953 4468
rect 8628 4428 8634 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 10520 4468 10548 4508
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11388 4508 11468 4536
rect 11388 4496 11394 4508
rect 11146 4468 11152 4480
rect 10520 4440 11152 4468
rect 8941 4431 8999 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11440 4468 11468 4508
rect 11790 4496 11796 4548
rect 11848 4496 11854 4548
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 11440 4440 12265 4468
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12253 4431 12311 4437
rect 1104 4378 42504 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 42504 4378
rect 1104 4304 42504 4326
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 4985 4267 5043 4273
rect 4985 4264 4997 4267
rect 4672 4236 4997 4264
rect 4672 4224 4678 4236
rect 4985 4233 4997 4236
rect 5031 4233 5043 4267
rect 4985 4227 5043 4233
rect 5350 4224 5356 4276
rect 5408 4224 5414 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 9858 4264 9864 4276
rect 9180 4236 9864 4264
rect 9180 4224 9186 4236
rect 9858 4224 9864 4236
rect 9916 4264 9922 4276
rect 9916 4236 10180 4264
rect 9916 4224 9922 4236
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 5258 4196 5264 4208
rect 4764 4168 5264 4196
rect 4764 4156 4770 4168
rect 5258 4156 5264 4168
rect 5316 4196 5322 4208
rect 5721 4199 5779 4205
rect 5721 4196 5733 4199
rect 5316 4168 5733 4196
rect 5316 4156 5322 4168
rect 5721 4165 5733 4168
rect 5767 4165 5779 4199
rect 9582 4196 9588 4208
rect 5721 4159 5779 4165
rect 8588 4168 9588 4196
rect 8588 4140 8616 4168
rect 9582 4156 9588 4168
rect 9640 4196 9646 4208
rect 10152 4196 10180 4236
rect 10318 4224 10324 4276
rect 10376 4264 10382 4276
rect 11330 4264 11336 4276
rect 10376 4236 11336 4264
rect 10376 4224 10382 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 10502 4196 10508 4208
rect 9640 4168 10088 4196
rect 9640 4156 9646 4168
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4264 4060 4292 4091
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4396 4100 5181 4128
rect 4396 4088 4402 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5552 4100 5917 4128
rect 4264 4032 4476 4060
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 4341 3995 4399 4001
rect 4341 3992 4353 3995
rect 3568 3964 4353 3992
rect 3568 3952 3574 3964
rect 4341 3961 4353 3964
rect 4387 3961 4399 3995
rect 4448 3992 4476 4032
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 4614 4020 4620 4072
rect 4672 4020 4678 4072
rect 4706 4020 4712 4072
rect 4764 4020 4770 4072
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5460 4060 5488 4088
rect 4948 4032 5488 4060
rect 4948 4020 4954 4032
rect 4816 3992 4844 4020
rect 5442 3992 5448 4004
rect 4448 3964 4844 3992
rect 5276 3964 5448 3992
rect 4341 3955 4399 3961
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 3292 3896 4169 3924
rect 3292 3884 3298 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4157 3887 4215 3893
rect 4522 3884 4528 3936
rect 4580 3924 4586 3936
rect 5276 3924 5304 3964
rect 5442 3952 5448 3964
rect 5500 3992 5506 4004
rect 5552 3992 5580 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8294 4128 8300 4140
rect 8251 4100 8300 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8570 4128 8576 4140
rect 8435 4100 8576 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8662 4088 8668 4140
rect 8720 4088 8726 4140
rect 8757 4131 8815 4137
rect 8757 4097 8769 4131
rect 8803 4097 8815 4131
rect 8757 4091 8815 4097
rect 8772 4060 8800 4091
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 10060 4137 10088 4168
rect 10152 4168 10508 4196
rect 10152 4140 10180 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 10045 4131 10103 4137
rect 9079 4100 9260 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8772 4032 9137 4060
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 5500 3964 5580 3992
rect 5500 3952 5506 3964
rect 7926 3952 7932 4004
rect 7984 3992 7990 4004
rect 8481 3995 8539 4001
rect 8481 3992 8493 3995
rect 7984 3964 8493 3992
rect 7984 3952 7990 3964
rect 8481 3961 8493 3964
rect 8527 3961 8539 3995
rect 8481 3955 8539 3961
rect 4580 3896 5304 3924
rect 4580 3884 4586 3896
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5408 3896 5549 3924
rect 5408 3884 5414 3896
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 9232 3924 9260 4100
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10134 4088 10140 4140
rect 10192 4088 10198 4140
rect 10410 4088 10416 4140
rect 10468 4088 10474 4140
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9456 4032 9689 4060
rect 9456 4020 9462 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 9861 3995 9919 4001
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 9950 3992 9956 4004
rect 9907 3964 9956 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 9950 3952 9956 3964
rect 10008 3992 10014 4004
rect 11238 3992 11244 4004
rect 10008 3964 11244 3992
rect 10008 3952 10014 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 8435 3896 9260 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10560 3896 11069 3924
rect 10560 3884 10566 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 1104 3834 42504 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 42504 3834
rect 1104 3760 42504 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 4706 3720 4712 3732
rect 2280 3692 4712 3720
rect 2280 3680 2286 3692
rect 3344 3661 3372 3692
rect 4706 3680 4712 3692
rect 4764 3720 4770 3732
rect 4890 3720 4896 3732
rect 4764 3692 4896 3720
rect 4764 3680 4770 3692
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 5629 3723 5687 3729
rect 5629 3720 5641 3723
rect 5316 3692 5641 3720
rect 5316 3680 5322 3692
rect 5629 3689 5641 3692
rect 5675 3720 5687 3723
rect 10781 3723 10839 3729
rect 5675 3692 6132 3720
rect 5675 3689 5687 3692
rect 5629 3683 5687 3689
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3621 3387 3655
rect 3329 3615 3387 3621
rect 3421 3655 3479 3661
rect 3421 3621 3433 3655
rect 3467 3652 3479 3655
rect 3467 3624 4016 3652
rect 3467 3621 3479 3624
rect 3421 3615 3479 3621
rect 3142 3544 3148 3596
rect 3200 3584 3206 3596
rect 3878 3584 3884 3596
rect 3200 3556 3884 3584
rect 3200 3544 3206 3556
rect 3878 3544 3884 3556
rect 3936 3544 3942 3596
rect 3988 3584 4016 3624
rect 5534 3584 5540 3596
rect 3988 3556 5540 3584
rect 5534 3544 5540 3556
rect 5592 3584 5598 3596
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5592 3556 6009 3584
rect 5592 3544 5598 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 3234 3476 3240 3528
rect 3292 3476 3298 3528
rect 3510 3476 3516 3528
rect 3568 3476 3574 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5500 3488 5733 3516
rect 5500 3476 5506 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 5721 3479 5779 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 6104 3516 6132 3692
rect 10781 3689 10793 3723
rect 10827 3720 10839 3723
rect 10827 3692 11008 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 10873 3655 10931 3661
rect 10873 3652 10885 3655
rect 8128 3624 10885 3652
rect 8128 3593 8156 3624
rect 10873 3621 10885 3624
rect 10919 3621 10931 3655
rect 10980 3652 11008 3692
rect 11238 3680 11244 3732
rect 11296 3680 11302 3732
rect 11790 3652 11796 3664
rect 10980 3624 11796 3652
rect 10873 3615 10931 3621
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 9401 3587 9459 3593
rect 9401 3584 9413 3587
rect 8527 3556 9413 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 9401 3553 9413 3556
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9548 3556 10640 3584
rect 9548 3544 9554 3556
rect 5859 3488 6132 3516
rect 6181 3519 6239 3525
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 6181 3485 6193 3519
rect 6227 3485 6239 3519
rect 6181 3479 6239 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8662 3516 8668 3528
rect 8619 3488 8668 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 4154 3408 4160 3460
rect 4212 3408 4218 3460
rect 5902 3448 5908 3460
rect 5382 3420 5908 3448
rect 5902 3408 5908 3420
rect 5960 3408 5966 3460
rect 6196 3448 6224 3479
rect 8662 3476 8668 3488
rect 8720 3516 8726 3528
rect 9508 3516 9536 3544
rect 8720 3488 9536 3516
rect 10045 3519 10103 3525
rect 8720 3476 8726 3488
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 10134 3516 10140 3528
rect 10091 3488 10140 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3476 10290 3528
rect 10502 3476 10508 3528
rect 10560 3476 10566 3528
rect 10612 3525 10640 3556
rect 11146 3544 11152 3596
rect 11204 3544 11210 3596
rect 41874 3544 41880 3596
rect 41932 3544 41938 3596
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 11514 3516 11520 3528
rect 11471 3488 11520 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 42150 3476 42156 3528
rect 42208 3476 42214 3528
rect 6914 3448 6920 3460
rect 6196 3420 6920 3448
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 3418 3380 3424 3392
rect 3099 3352 3424 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 6196 3380 6224 3420
rect 6914 3408 6920 3420
rect 6972 3448 6978 3460
rect 8846 3448 8852 3460
rect 6972 3420 8852 3448
rect 6972 3408 6978 3420
rect 8846 3408 8852 3420
rect 8904 3448 8910 3460
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 8904 3420 10425 3448
rect 8904 3408 8910 3420
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 10413 3411 10471 3417
rect 4580 3352 6224 3380
rect 8757 3383 8815 3389
rect 4580 3340 4586 3352
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 9766 3380 9772 3392
rect 8803 3352 9772 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 1104 3290 42504 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 42504 3290
rect 1104 3216 42504 3238
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4985 3179 5043 3185
rect 4985 3176 4997 3179
rect 4212 3148 4997 3176
rect 4212 3136 4218 3148
rect 4985 3145 4997 3148
rect 5031 3145 5043 3179
rect 5902 3176 5908 3188
rect 4985 3139 5043 3145
rect 5092 3148 5908 3176
rect 3418 3068 3424 3120
rect 3476 3068 3482 3120
rect 5092 3108 5120 3148
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 9398 3136 9404 3188
rect 9456 3136 9462 3188
rect 10594 3176 10600 3188
rect 9508 3148 10600 3176
rect 4646 3080 5120 3108
rect 5258 3068 5264 3120
rect 5316 3068 5322 3120
rect 5350 3068 5356 3120
rect 5408 3068 5414 3120
rect 7926 3068 7932 3120
rect 7984 3068 7990 3120
rect 3142 3000 3148 3052
rect 3200 3000 3206 3052
rect 4706 3000 4712 3052
rect 4764 3040 4770 3052
rect 5169 3043 5227 3049
rect 5169 3040 5181 3043
rect 4764 3012 5181 3040
rect 4764 3000 4770 3012
rect 5169 3009 5181 3012
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5534 3000 5540 3052
rect 5592 3000 5598 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 9508 3049 9536 3148
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 9766 3068 9772 3120
rect 9824 3068 9830 3120
rect 10318 3068 10324 3120
rect 10376 3068 10382 3120
rect 7653 3043 7711 3049
rect 7653 3040 7665 3043
rect 6880 3012 7665 3040
rect 6880 3000 6886 3012
rect 7653 3009 7665 3012
rect 7699 3009 7711 3043
rect 9493 3043 9551 3049
rect 7653 3003 7711 3009
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4856 2944 4905 2972
rect 4856 2932 4862 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 4893 2935 4951 2941
rect 9048 2836 9076 3026
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 10134 2932 10140 2984
rect 10192 2972 10198 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 10192 2944 11253 2972
rect 10192 2932 10198 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 10318 2836 10324 2848
rect 9048 2808 10324 2836
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 1104 2746 42504 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 42504 2746
rect 1104 2672 42504 2694
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 8812 2400 11713 2428
rect 8812 2388 8818 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2261 11943 2295
rect 11885 2255 11943 2261
rect 1104 2202 42504 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 42504 2202
rect 1104 2128 42504 2150
<< via1 >>
rect 4874 43494 4926 43546
rect 4938 43494 4990 43546
rect 5002 43494 5054 43546
rect 5066 43494 5118 43546
rect 5130 43494 5182 43546
rect 35594 43494 35646 43546
rect 35658 43494 35710 43546
rect 35722 43494 35774 43546
rect 35786 43494 35838 43546
rect 35850 43494 35902 43546
rect 17684 43435 17736 43444
rect 17684 43401 17693 43435
rect 17693 43401 17727 43435
rect 17727 43401 17736 43435
rect 17684 43392 17736 43401
rect 19524 43435 19576 43444
rect 19524 43401 19533 43435
rect 19533 43401 19567 43435
rect 19567 43401 19576 43435
rect 19524 43392 19576 43401
rect 20260 43435 20312 43444
rect 20260 43401 20269 43435
rect 20269 43401 20303 43435
rect 20303 43401 20312 43435
rect 20260 43392 20312 43401
rect 20536 43392 20588 43444
rect 22836 43435 22888 43444
rect 22836 43401 22845 43435
rect 22845 43401 22879 43435
rect 22879 43401 22888 43435
rect 22836 43392 22888 43401
rect 23388 43435 23440 43444
rect 23388 43401 23397 43435
rect 23397 43401 23431 43435
rect 23431 43401 23440 43435
rect 23388 43392 23440 43401
rect 25320 43435 25372 43444
rect 25320 43401 25329 43435
rect 25329 43401 25363 43435
rect 25363 43401 25372 43435
rect 25320 43392 25372 43401
rect 29184 43435 29236 43444
rect 29184 43401 29193 43435
rect 29193 43401 29227 43435
rect 29227 43401 29236 43435
rect 29184 43392 29236 43401
rect 24400 43324 24452 43376
rect 28448 43324 28500 43376
rect 17500 43299 17552 43308
rect 17500 43265 17509 43299
rect 17509 43265 17543 43299
rect 17543 43265 17552 43299
rect 17500 43256 17552 43265
rect 19800 43256 19852 43308
rect 19340 43188 19392 43240
rect 20996 43299 21048 43308
rect 20996 43265 21005 43299
rect 21005 43265 21039 43299
rect 21039 43265 21048 43299
rect 20996 43256 21048 43265
rect 22744 43256 22796 43308
rect 23020 43256 23072 43308
rect 24584 43299 24636 43308
rect 24584 43265 24593 43299
rect 24593 43265 24627 43299
rect 24627 43265 24636 43299
rect 24584 43256 24636 43265
rect 24676 43188 24728 43240
rect 26148 43256 26200 43308
rect 28356 43299 28408 43308
rect 28356 43265 28365 43299
rect 28365 43265 28399 43299
rect 28399 43265 28408 43299
rect 28356 43256 28408 43265
rect 29552 43256 29604 43308
rect 24032 43052 24084 43104
rect 28080 43052 28132 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 17500 42848 17552 42900
rect 26148 42891 26200 42900
rect 26148 42857 26157 42891
rect 26157 42857 26191 42891
rect 26191 42857 26200 42891
rect 26148 42848 26200 42857
rect 28356 42848 28408 42900
rect 24768 42712 24820 42764
rect 27620 42712 27672 42764
rect 15660 42687 15712 42696
rect 15660 42653 15669 42687
rect 15669 42653 15703 42687
rect 15703 42653 15712 42687
rect 15660 42644 15712 42653
rect 19064 42644 19116 42696
rect 16212 42576 16264 42628
rect 16396 42576 16448 42628
rect 18144 42508 18196 42560
rect 19524 42619 19576 42628
rect 19524 42585 19533 42619
rect 19533 42585 19567 42619
rect 19567 42585 19576 42619
rect 19524 42576 19576 42585
rect 19800 42687 19852 42696
rect 19800 42653 19809 42687
rect 19809 42653 19843 42687
rect 19843 42653 19852 42687
rect 19800 42644 19852 42653
rect 19892 42644 19944 42696
rect 24032 42687 24084 42696
rect 24032 42653 24041 42687
rect 24041 42653 24075 42687
rect 24075 42653 24084 42687
rect 24032 42644 24084 42653
rect 25688 42644 25740 42696
rect 29644 42712 29696 42764
rect 37280 42712 37332 42764
rect 19432 42508 19484 42560
rect 20812 42576 20864 42628
rect 21548 42576 21600 42628
rect 22192 42508 22244 42560
rect 22744 42551 22796 42560
rect 22744 42517 22753 42551
rect 22753 42517 22787 42551
rect 22787 42517 22796 42551
rect 22744 42508 22796 42517
rect 23664 42576 23716 42628
rect 24032 42508 24084 42560
rect 27896 42644 27948 42696
rect 29552 42644 29604 42696
rect 26608 42619 26660 42628
rect 26608 42585 26617 42619
rect 26617 42585 26651 42619
rect 26651 42585 26660 42619
rect 26608 42576 26660 42585
rect 28540 42576 28592 42628
rect 28264 42508 28316 42560
rect 28816 42619 28868 42628
rect 28816 42585 28825 42619
rect 28825 42585 28859 42619
rect 28859 42585 28868 42619
rect 28816 42576 28868 42585
rect 35440 42619 35492 42628
rect 35440 42585 35449 42619
rect 35449 42585 35483 42619
rect 35483 42585 35492 42619
rect 35440 42576 35492 42585
rect 36820 42576 36872 42628
rect 37004 42508 37056 42560
rect 4874 42406 4926 42458
rect 4938 42406 4990 42458
rect 5002 42406 5054 42458
rect 5066 42406 5118 42458
rect 5130 42406 5182 42458
rect 35594 42406 35646 42458
rect 35658 42406 35710 42458
rect 35722 42406 35774 42458
rect 35786 42406 35838 42458
rect 35850 42406 35902 42458
rect 16580 42236 16632 42288
rect 15936 42168 15988 42220
rect 16212 42168 16264 42220
rect 17500 42168 17552 42220
rect 18788 42304 18840 42356
rect 19892 42304 19944 42356
rect 22008 42304 22060 42356
rect 24584 42304 24636 42356
rect 24676 42304 24728 42356
rect 18144 42279 18196 42288
rect 18144 42245 18153 42279
rect 18153 42245 18187 42279
rect 18187 42245 18196 42279
rect 18144 42236 18196 42245
rect 19156 42236 19208 42288
rect 20720 42236 20772 42288
rect 26608 42304 26660 42356
rect 28264 42304 28316 42356
rect 29552 42347 29604 42356
rect 29552 42313 29561 42347
rect 29561 42313 29595 42347
rect 29595 42313 29604 42347
rect 29552 42304 29604 42313
rect 35440 42304 35492 42356
rect 19892 42211 19944 42220
rect 19892 42177 19901 42211
rect 19901 42177 19935 42211
rect 19935 42177 19944 42211
rect 19892 42168 19944 42177
rect 24032 42168 24084 42220
rect 25596 42168 25648 42220
rect 27436 42168 27488 42220
rect 28080 42279 28132 42288
rect 28080 42245 28089 42279
rect 28089 42245 28123 42279
rect 28123 42245 28132 42279
rect 28080 42236 28132 42245
rect 28540 42236 28592 42288
rect 29644 42236 29696 42288
rect 19432 42100 19484 42152
rect 19800 42100 19852 42152
rect 20168 42143 20220 42152
rect 20168 42109 20177 42143
rect 20177 42109 20211 42143
rect 20211 42109 20220 42143
rect 20168 42100 20220 42109
rect 22652 42143 22704 42152
rect 22652 42109 22661 42143
rect 22661 42109 22695 42143
rect 22695 42109 22704 42143
rect 22652 42100 22704 42109
rect 23296 42100 23348 42152
rect 27344 42100 27396 42152
rect 20812 41964 20864 42016
rect 21732 41964 21784 42016
rect 21824 42007 21876 42016
rect 21824 41973 21833 42007
rect 21833 41973 21867 42007
rect 21867 41973 21876 42007
rect 21824 41964 21876 41973
rect 24400 42007 24452 42016
rect 24400 41973 24409 42007
rect 24409 41973 24443 42007
rect 24443 41973 24452 42007
rect 24400 41964 24452 41973
rect 25320 41964 25372 42016
rect 26884 41964 26936 42016
rect 34796 42168 34848 42220
rect 35624 42211 35676 42220
rect 35624 42177 35633 42211
rect 35633 42177 35667 42211
rect 35667 42177 35676 42211
rect 35624 42168 35676 42177
rect 36452 42168 36504 42220
rect 36820 42236 36872 42288
rect 37280 42211 37332 42220
rect 37280 42177 37289 42211
rect 37289 42177 37323 42211
rect 37323 42177 37332 42211
rect 37280 42168 37332 42177
rect 27712 42100 27764 42152
rect 28724 42100 28776 42152
rect 28816 42100 28868 42152
rect 30840 42100 30892 42152
rect 30932 42100 30984 42152
rect 31576 42032 31628 42084
rect 32036 42100 32088 42152
rect 35348 42100 35400 42152
rect 30932 41964 30984 42016
rect 31208 41964 31260 42016
rect 32956 41964 33008 42016
rect 36544 42143 36596 42152
rect 36544 42109 36553 42143
rect 36553 42109 36587 42143
rect 36587 42109 36596 42143
rect 36544 42100 36596 42109
rect 36636 42143 36688 42152
rect 36636 42109 36645 42143
rect 36645 42109 36679 42143
rect 36679 42109 36688 42143
rect 36636 42100 36688 42109
rect 37004 42032 37056 42084
rect 36084 42007 36136 42016
rect 36084 41973 36093 42007
rect 36093 41973 36127 42007
rect 36127 41973 36136 42007
rect 36084 41964 36136 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 20168 41760 20220 41812
rect 21548 41760 21600 41812
rect 23296 41803 23348 41812
rect 23296 41769 23305 41803
rect 23305 41769 23339 41803
rect 23339 41769 23348 41803
rect 23296 41760 23348 41769
rect 27344 41803 27396 41812
rect 27344 41769 27353 41803
rect 27353 41769 27387 41803
rect 27387 41769 27396 41803
rect 27344 41760 27396 41769
rect 27436 41760 27488 41812
rect 28540 41760 28592 41812
rect 15660 41624 15712 41676
rect 18788 41624 18840 41676
rect 20076 41667 20128 41676
rect 20076 41633 20085 41667
rect 20085 41633 20119 41667
rect 20119 41633 20128 41667
rect 20076 41624 20128 41633
rect 21088 41667 21140 41676
rect 21088 41633 21097 41667
rect 21097 41633 21131 41667
rect 21131 41633 21140 41667
rect 21088 41624 21140 41633
rect 21732 41624 21784 41676
rect 16396 41556 16448 41608
rect 19984 41599 20036 41608
rect 19984 41565 19993 41599
rect 19993 41565 20027 41599
rect 20027 41565 20036 41599
rect 19984 41556 20036 41565
rect 15384 41488 15436 41540
rect 17408 41531 17460 41540
rect 17408 41497 17417 41531
rect 17417 41497 17451 41531
rect 17451 41497 17460 41531
rect 17408 41488 17460 41497
rect 20720 41556 20772 41608
rect 21824 41556 21876 41608
rect 22008 41599 22060 41608
rect 22008 41565 22017 41599
rect 22017 41565 22051 41599
rect 22051 41565 22060 41599
rect 22008 41556 22060 41565
rect 24032 41624 24084 41676
rect 26884 41667 26936 41676
rect 22744 41556 22796 41608
rect 24400 41556 24452 41608
rect 25872 41599 25924 41608
rect 25872 41565 25881 41599
rect 25881 41565 25915 41599
rect 25915 41565 25924 41599
rect 25872 41556 25924 41565
rect 25964 41599 26016 41608
rect 25964 41565 25973 41599
rect 25973 41565 26007 41599
rect 26007 41565 26016 41599
rect 25964 41556 26016 41565
rect 26056 41599 26108 41608
rect 26056 41565 26065 41599
rect 26065 41565 26099 41599
rect 26099 41565 26108 41599
rect 26056 41556 26108 41565
rect 16580 41463 16632 41472
rect 16580 41429 16589 41463
rect 16589 41429 16623 41463
rect 16623 41429 16632 41463
rect 16580 41420 16632 41429
rect 18328 41420 18380 41472
rect 19432 41420 19484 41472
rect 21364 41531 21416 41540
rect 21364 41497 21373 41531
rect 21373 41497 21407 41531
rect 21407 41497 21416 41531
rect 21364 41488 21416 41497
rect 22192 41531 22244 41540
rect 22192 41497 22201 41531
rect 22201 41497 22235 41531
rect 22235 41497 22244 41531
rect 22192 41488 22244 41497
rect 22836 41488 22888 41540
rect 24676 41488 24728 41540
rect 25504 41488 25556 41540
rect 26884 41633 26893 41667
rect 26893 41633 26927 41667
rect 26927 41633 26936 41667
rect 26884 41624 26936 41633
rect 23756 41463 23808 41472
rect 23756 41429 23765 41463
rect 23765 41429 23799 41463
rect 23799 41429 23808 41463
rect 23756 41420 23808 41429
rect 25688 41463 25740 41472
rect 25688 41429 25697 41463
rect 25697 41429 25731 41463
rect 25731 41429 25740 41463
rect 25688 41420 25740 41429
rect 27068 41599 27120 41608
rect 27068 41565 27077 41599
rect 27077 41565 27111 41599
rect 27111 41565 27120 41599
rect 27068 41556 27120 41565
rect 28724 41692 28776 41744
rect 27344 41624 27396 41676
rect 27620 41667 27672 41676
rect 27620 41633 27629 41667
rect 27629 41633 27663 41667
rect 27663 41633 27672 41667
rect 27620 41624 27672 41633
rect 28172 41556 28224 41608
rect 28724 41599 28776 41608
rect 28724 41565 28733 41599
rect 28733 41565 28767 41599
rect 28767 41565 28776 41599
rect 28724 41556 28776 41565
rect 27804 41488 27856 41540
rect 28540 41488 28592 41540
rect 30472 41599 30524 41608
rect 30472 41565 30481 41599
rect 30481 41565 30515 41599
rect 30515 41565 30524 41599
rect 30472 41556 30524 41565
rect 30840 41803 30892 41812
rect 30840 41769 30849 41803
rect 30849 41769 30883 41803
rect 30883 41769 30892 41803
rect 30840 41760 30892 41769
rect 30932 41760 30984 41812
rect 32220 41760 32272 41812
rect 32864 41760 32916 41812
rect 33048 41760 33100 41812
rect 31116 41692 31168 41744
rect 34796 41803 34848 41812
rect 34796 41769 34805 41803
rect 34805 41769 34839 41803
rect 34839 41769 34848 41803
rect 34796 41760 34848 41769
rect 35348 41803 35400 41812
rect 35348 41769 35357 41803
rect 35357 41769 35391 41803
rect 35391 41769 35400 41803
rect 35348 41760 35400 41769
rect 32128 41624 32180 41676
rect 30932 41556 30984 41608
rect 30748 41531 30800 41540
rect 30748 41497 30757 41531
rect 30757 41497 30791 41531
rect 30791 41497 30800 41531
rect 30748 41488 30800 41497
rect 29092 41463 29144 41472
rect 29092 41429 29101 41463
rect 29101 41429 29135 41463
rect 29135 41429 29144 41463
rect 29092 41420 29144 41429
rect 31116 41599 31168 41608
rect 31116 41565 31125 41599
rect 31125 41565 31159 41599
rect 31159 41565 31168 41599
rect 31116 41556 31168 41565
rect 31208 41556 31260 41608
rect 31576 41556 31628 41608
rect 31668 41488 31720 41540
rect 31852 41599 31904 41608
rect 31852 41565 31861 41599
rect 31861 41565 31895 41599
rect 31895 41565 31904 41599
rect 31852 41556 31904 41565
rect 31944 41599 31996 41608
rect 31944 41565 31953 41599
rect 31953 41565 31987 41599
rect 31987 41565 31996 41599
rect 31944 41556 31996 41565
rect 32036 41599 32088 41608
rect 32036 41565 32045 41599
rect 32045 41565 32079 41599
rect 32079 41565 32088 41599
rect 32036 41556 32088 41565
rect 35624 41692 35676 41744
rect 36360 41760 36412 41812
rect 36636 41760 36688 41812
rect 32404 41556 32456 41608
rect 32772 41599 32824 41608
rect 32772 41565 32781 41599
rect 32781 41565 32815 41599
rect 32815 41565 32824 41599
rect 32772 41556 32824 41565
rect 32864 41599 32916 41608
rect 32864 41565 32873 41599
rect 32873 41565 32907 41599
rect 32907 41565 32916 41599
rect 32864 41556 32916 41565
rect 32956 41599 33008 41608
rect 32956 41565 32965 41599
rect 32965 41565 32999 41599
rect 32999 41565 33008 41599
rect 32956 41556 33008 41565
rect 34520 41556 34572 41608
rect 31852 41420 31904 41472
rect 32680 41420 32732 41472
rect 35716 41599 35768 41608
rect 35716 41565 35725 41599
rect 35725 41565 35759 41599
rect 35759 41565 35768 41599
rect 35716 41556 35768 41565
rect 35900 41556 35952 41608
rect 36268 41667 36320 41676
rect 36268 41633 36277 41667
rect 36277 41633 36311 41667
rect 36311 41633 36320 41667
rect 36268 41624 36320 41633
rect 36820 41599 36872 41608
rect 36820 41565 36829 41599
rect 36829 41565 36863 41599
rect 36863 41565 36872 41599
rect 36820 41556 36872 41565
rect 36912 41599 36964 41608
rect 36912 41565 36921 41599
rect 36921 41565 36955 41599
rect 36955 41565 36964 41599
rect 36912 41556 36964 41565
rect 35072 41463 35124 41472
rect 35072 41429 35081 41463
rect 35081 41429 35115 41463
rect 35115 41429 35124 41463
rect 35072 41420 35124 41429
rect 35440 41420 35492 41472
rect 36820 41420 36872 41472
rect 4874 41318 4926 41370
rect 4938 41318 4990 41370
rect 5002 41318 5054 41370
rect 5066 41318 5118 41370
rect 5130 41318 5182 41370
rect 35594 41318 35646 41370
rect 35658 41318 35710 41370
rect 35722 41318 35774 41370
rect 35786 41318 35838 41370
rect 35850 41318 35902 41370
rect 15384 41216 15436 41268
rect 17040 41148 17092 41200
rect 17592 41191 17644 41200
rect 17592 41157 17617 41191
rect 17617 41157 17644 41191
rect 17592 41148 17644 41157
rect 17960 41123 18012 41132
rect 17960 41089 17969 41123
rect 17969 41089 18003 41123
rect 18003 41089 18012 41123
rect 17960 41080 18012 41089
rect 19432 41216 19484 41268
rect 19984 41259 20036 41268
rect 19984 41225 19993 41259
rect 19993 41225 20027 41259
rect 20027 41225 20036 41259
rect 19984 41216 20036 41225
rect 23756 41216 23808 41268
rect 25872 41216 25924 41268
rect 24032 41148 24084 41200
rect 27344 41259 27396 41268
rect 27344 41225 27353 41259
rect 27353 41225 27387 41259
rect 27387 41225 27396 41259
rect 27344 41216 27396 41225
rect 27620 41148 27672 41200
rect 16580 41012 16632 41064
rect 18144 41012 18196 41064
rect 18788 41012 18840 41064
rect 18052 40944 18104 40996
rect 19248 41012 19300 41064
rect 19984 41012 20036 41064
rect 20904 41080 20956 41132
rect 22560 41080 22612 41132
rect 22928 41080 22980 41132
rect 20996 41012 21048 41064
rect 23388 41080 23440 41132
rect 23756 41123 23808 41132
rect 23756 41089 23765 41123
rect 23765 41089 23799 41123
rect 23799 41089 23808 41123
rect 23756 41080 23808 41089
rect 24768 41123 24820 41132
rect 24768 41089 24777 41123
rect 24777 41089 24811 41123
rect 24811 41089 24820 41123
rect 24768 41080 24820 41089
rect 28908 41148 28960 41200
rect 29644 41148 29696 41200
rect 25044 41055 25096 41064
rect 25044 41021 25053 41055
rect 25053 41021 25087 41055
rect 25087 41021 25096 41055
rect 25044 41012 25096 41021
rect 25596 41012 25648 41064
rect 25780 41012 25832 41064
rect 17500 40876 17552 40928
rect 17776 40919 17828 40928
rect 17776 40885 17785 40919
rect 17785 40885 17819 40919
rect 17819 40885 17828 40919
rect 17776 40876 17828 40885
rect 17868 40876 17920 40928
rect 19800 40987 19852 40996
rect 19800 40953 19809 40987
rect 19809 40953 19843 40987
rect 19843 40953 19852 40987
rect 19800 40944 19852 40953
rect 21088 40876 21140 40928
rect 26148 40876 26200 40928
rect 26240 40876 26292 40928
rect 28172 41012 28224 41064
rect 28356 41055 28408 41064
rect 28356 41021 28365 41055
rect 28365 41021 28399 41055
rect 28399 41021 28408 41055
rect 28356 41012 28408 41021
rect 28908 41055 28960 41064
rect 28908 41021 28917 41055
rect 28917 41021 28951 41055
rect 28951 41021 28960 41055
rect 28908 41012 28960 41021
rect 30748 41080 30800 41132
rect 31116 41080 31168 41132
rect 31668 41148 31720 41200
rect 30564 41012 30616 41064
rect 31852 41148 31904 41200
rect 32772 41148 32824 41200
rect 33232 41148 33284 41200
rect 32220 41123 32272 41132
rect 32220 41089 32229 41123
rect 32229 41089 32263 41123
rect 32263 41089 32272 41123
rect 32220 41080 32272 41089
rect 32404 41123 32456 41132
rect 32404 41089 32413 41123
rect 32413 41089 32447 41123
rect 32447 41089 32456 41123
rect 32404 41080 32456 41089
rect 34152 41148 34204 41200
rect 36176 41148 36228 41200
rect 36728 41148 36780 41200
rect 32496 41055 32548 41064
rect 32496 41021 32505 41055
rect 32505 41021 32539 41055
rect 32539 41021 32548 41055
rect 32496 41012 32548 41021
rect 32864 41012 32916 41064
rect 33140 41012 33192 41064
rect 34704 41012 34756 41064
rect 35072 41012 35124 41064
rect 36268 41080 36320 41132
rect 37188 41080 37240 41132
rect 37280 41080 37332 41132
rect 38200 41123 38252 41132
rect 38200 41089 38209 41123
rect 38209 41089 38243 41123
rect 38243 41089 38252 41123
rect 38200 41080 38252 41089
rect 36360 41012 36412 41064
rect 36912 41012 36964 41064
rect 36544 40944 36596 40996
rect 37372 40944 37424 40996
rect 30564 40876 30616 40928
rect 32772 40876 32824 40928
rect 33324 40876 33376 40928
rect 35348 40876 35400 40928
rect 36820 40876 36872 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 1308 40672 1360 40724
rect 17132 40672 17184 40724
rect 17408 40672 17460 40724
rect 17500 40672 17552 40724
rect 19984 40672 20036 40724
rect 20076 40672 20128 40724
rect 20904 40715 20956 40724
rect 20904 40681 20913 40715
rect 20913 40681 20947 40715
rect 20947 40681 20956 40715
rect 20904 40672 20956 40681
rect 21088 40672 21140 40724
rect 25044 40672 25096 40724
rect 25872 40672 25924 40724
rect 28356 40672 28408 40724
rect 32864 40672 32916 40724
rect 33232 40672 33284 40724
rect 34152 40672 34204 40724
rect 17776 40604 17828 40656
rect 20812 40604 20864 40656
rect 17408 40536 17460 40588
rect 19800 40536 19852 40588
rect 17040 40511 17092 40520
rect 17040 40477 17049 40511
rect 17049 40477 17083 40511
rect 17083 40477 17092 40511
rect 17040 40468 17092 40477
rect 17592 40400 17644 40452
rect 17868 40468 17920 40520
rect 18144 40511 18196 40520
rect 18144 40477 18153 40511
rect 18153 40477 18187 40511
rect 18187 40477 18196 40511
rect 18144 40468 18196 40477
rect 22100 40579 22152 40588
rect 22100 40545 22109 40579
rect 22109 40545 22143 40579
rect 22143 40545 22152 40579
rect 22100 40536 22152 40545
rect 22928 40536 22980 40588
rect 25688 40536 25740 40588
rect 25964 40579 26016 40588
rect 25964 40545 25973 40579
rect 25973 40545 26007 40579
rect 26007 40545 26016 40579
rect 25964 40536 26016 40545
rect 18788 40400 18840 40452
rect 20076 40443 20128 40452
rect 20076 40409 20085 40443
rect 20085 40409 20119 40443
rect 20119 40409 20128 40443
rect 20076 40400 20128 40409
rect 21272 40511 21324 40520
rect 21272 40477 21281 40511
rect 21281 40477 21315 40511
rect 21315 40477 21324 40511
rect 21272 40468 21324 40477
rect 20628 40400 20680 40452
rect 21824 40400 21876 40452
rect 30472 40604 30524 40656
rect 31116 40647 31168 40656
rect 31116 40613 31125 40647
rect 31125 40613 31159 40647
rect 31159 40613 31168 40647
rect 31116 40604 31168 40613
rect 34796 40604 34848 40656
rect 27804 40536 27856 40588
rect 29092 40536 29144 40588
rect 30656 40579 30708 40588
rect 30656 40545 30665 40579
rect 30665 40545 30699 40579
rect 30699 40545 30708 40579
rect 30656 40536 30708 40545
rect 32680 40579 32732 40588
rect 32680 40545 32689 40579
rect 32689 40545 32723 40579
rect 32723 40545 32732 40579
rect 32680 40536 32732 40545
rect 32956 40536 33008 40588
rect 26148 40468 26200 40520
rect 28172 40511 28224 40520
rect 28172 40477 28181 40511
rect 28181 40477 28215 40511
rect 28215 40477 28224 40511
rect 28172 40468 28224 40477
rect 30748 40511 30800 40520
rect 30748 40477 30757 40511
rect 30757 40477 30791 40511
rect 30791 40477 30800 40511
rect 30748 40468 30800 40477
rect 32772 40511 32824 40520
rect 32772 40477 32781 40511
rect 32781 40477 32815 40511
rect 32815 40477 32824 40511
rect 32772 40468 32824 40477
rect 34704 40468 34756 40520
rect 36820 40604 36872 40656
rect 35256 40511 35308 40520
rect 35256 40477 35265 40511
rect 35265 40477 35299 40511
rect 35299 40477 35308 40511
rect 35256 40468 35308 40477
rect 35348 40511 35400 40520
rect 35348 40477 35357 40511
rect 35357 40477 35391 40511
rect 35391 40477 35400 40511
rect 35348 40468 35400 40477
rect 25504 40400 25556 40452
rect 26056 40443 26108 40452
rect 26056 40409 26065 40443
rect 26065 40409 26099 40443
rect 26099 40409 26108 40443
rect 26056 40400 26108 40409
rect 33324 40400 33376 40452
rect 35440 40400 35492 40452
rect 37832 40511 37884 40520
rect 37832 40477 37841 40511
rect 37841 40477 37875 40511
rect 37875 40477 37884 40511
rect 37832 40468 37884 40477
rect 38200 40536 38252 40588
rect 39304 40468 39356 40520
rect 42156 40511 42208 40520
rect 42156 40477 42165 40511
rect 42165 40477 42199 40511
rect 42199 40477 42208 40511
rect 42156 40468 42208 40477
rect 38108 40443 38160 40452
rect 38108 40409 38117 40443
rect 38117 40409 38151 40443
rect 38151 40409 38160 40443
rect 38108 40400 38160 40409
rect 26240 40375 26292 40384
rect 26240 40341 26249 40375
rect 26249 40341 26283 40375
rect 26283 40341 26292 40375
rect 26240 40332 26292 40341
rect 31944 40332 31996 40384
rect 34428 40332 34480 40384
rect 35992 40332 36044 40384
rect 41052 40332 41104 40384
rect 4874 40230 4926 40282
rect 4938 40230 4990 40282
rect 5002 40230 5054 40282
rect 5066 40230 5118 40282
rect 5130 40230 5182 40282
rect 35594 40230 35646 40282
rect 35658 40230 35710 40282
rect 35722 40230 35774 40282
rect 35786 40230 35838 40282
rect 35850 40230 35902 40282
rect 17592 40128 17644 40180
rect 20076 40128 20128 40180
rect 20628 40128 20680 40180
rect 14556 39992 14608 40044
rect 16028 40035 16080 40044
rect 16028 40001 16037 40035
rect 16037 40001 16071 40035
rect 16071 40001 16080 40035
rect 16028 39992 16080 40001
rect 20812 40060 20864 40112
rect 21272 40128 21324 40180
rect 23388 40128 23440 40180
rect 26056 40128 26108 40180
rect 30748 40171 30800 40180
rect 30748 40137 30757 40171
rect 30757 40137 30791 40171
rect 30791 40137 30800 40171
rect 30748 40128 30800 40137
rect 32404 40128 32456 40180
rect 26240 40060 26292 40112
rect 35348 40128 35400 40180
rect 37832 40128 37884 40180
rect 36176 40060 36228 40112
rect 38200 40060 38252 40112
rect 16304 39992 16356 40044
rect 17132 40035 17184 40044
rect 17132 40001 17141 40035
rect 17141 40001 17175 40035
rect 17175 40001 17184 40035
rect 17132 39992 17184 40001
rect 18604 39992 18656 40044
rect 20996 39992 21048 40044
rect 22100 39992 22152 40044
rect 23112 40035 23164 40044
rect 23112 40001 23121 40035
rect 23121 40001 23155 40035
rect 23155 40001 23164 40035
rect 23112 39992 23164 40001
rect 25044 40035 25096 40044
rect 25044 40001 25053 40035
rect 25053 40001 25087 40035
rect 25087 40001 25096 40035
rect 25044 39992 25096 40001
rect 26516 39992 26568 40044
rect 30288 39992 30340 40044
rect 31392 39992 31444 40044
rect 32036 39992 32088 40044
rect 35348 39992 35400 40044
rect 35992 40035 36044 40044
rect 35992 40001 36001 40035
rect 36001 40001 36035 40035
rect 36035 40001 36044 40035
rect 35992 39992 36044 40001
rect 12900 39924 12952 39976
rect 13544 39967 13596 39976
rect 13544 39933 13553 39967
rect 13553 39933 13587 39967
rect 13587 39933 13596 39967
rect 13544 39924 13596 39933
rect 14832 39788 14884 39840
rect 17040 39924 17092 39976
rect 17316 39924 17368 39976
rect 18696 39924 18748 39976
rect 23204 39967 23256 39976
rect 23204 39933 23213 39967
rect 23213 39933 23247 39967
rect 23247 39933 23256 39967
rect 23204 39924 23256 39933
rect 25136 39967 25188 39976
rect 25136 39933 25145 39967
rect 25145 39933 25179 39967
rect 25179 39933 25188 39967
rect 25136 39924 25188 39933
rect 26792 39924 26844 39976
rect 32220 39967 32272 39976
rect 32220 39933 32229 39967
rect 32229 39933 32263 39967
rect 32263 39933 32272 39967
rect 32220 39924 32272 39933
rect 32404 39924 32456 39976
rect 34704 39924 34756 39976
rect 35440 39924 35492 39976
rect 36084 39967 36136 39976
rect 36084 39933 36093 39967
rect 36093 39933 36127 39967
rect 36127 39933 36136 39967
rect 36084 39924 36136 39933
rect 27804 39856 27856 39908
rect 35992 39856 36044 39908
rect 37004 39856 37056 39908
rect 15108 39831 15160 39840
rect 15108 39797 15117 39831
rect 15117 39797 15151 39831
rect 15151 39797 15160 39831
rect 15108 39788 15160 39797
rect 20720 39788 20772 39840
rect 21548 39788 21600 39840
rect 35532 39831 35584 39840
rect 35532 39797 35541 39831
rect 35541 39797 35575 39831
rect 35575 39797 35584 39831
rect 35532 39788 35584 39797
rect 35624 39831 35676 39840
rect 35624 39797 35633 39831
rect 35633 39797 35667 39831
rect 35667 39797 35676 39831
rect 35624 39788 35676 39797
rect 35716 39788 35768 39840
rect 37188 39992 37240 40044
rect 37280 39967 37332 39976
rect 37280 39933 37289 39967
rect 37289 39933 37323 39967
rect 37323 39933 37332 39967
rect 37280 39924 37332 39933
rect 38476 39967 38528 39976
rect 38476 39933 38485 39967
rect 38485 39933 38519 39967
rect 38519 39933 38528 39967
rect 38476 39924 38528 39933
rect 39580 40035 39632 40044
rect 39580 40001 39588 40035
rect 39588 40001 39622 40035
rect 39622 40001 39632 40035
rect 39580 39992 39632 40001
rect 39672 40035 39724 40044
rect 39672 40001 39681 40035
rect 39681 40001 39715 40035
rect 39715 40001 39724 40035
rect 39672 39992 39724 40001
rect 41420 39992 41472 40044
rect 38936 39899 38988 39908
rect 38936 39865 38945 39899
rect 38945 39865 38979 39899
rect 38979 39865 38988 39899
rect 38936 39856 38988 39865
rect 39028 39899 39080 39908
rect 39028 39865 39037 39899
rect 39037 39865 39071 39899
rect 39071 39865 39080 39899
rect 39028 39856 39080 39865
rect 39304 39967 39356 39976
rect 39304 39933 39313 39967
rect 39313 39933 39347 39967
rect 39347 39933 39356 39967
rect 39304 39924 39356 39933
rect 40316 39967 40368 39976
rect 40316 39933 40325 39967
rect 40325 39933 40359 39967
rect 40359 39933 40368 39967
rect 40316 39924 40368 39933
rect 39672 39856 39724 39908
rect 37740 39788 37792 39840
rect 37924 39831 37976 39840
rect 37924 39797 37933 39831
rect 37933 39797 37967 39831
rect 37967 39797 37976 39831
rect 37924 39788 37976 39797
rect 41788 39831 41840 39840
rect 41788 39797 41797 39831
rect 41797 39797 41831 39831
rect 41831 39797 41840 39831
rect 41788 39788 41840 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 13544 39584 13596 39636
rect 14740 39448 14792 39500
rect 14832 39491 14884 39500
rect 14832 39457 14841 39491
rect 14841 39457 14875 39491
rect 14875 39457 14884 39491
rect 14832 39448 14884 39457
rect 18144 39584 18196 39636
rect 17316 39559 17368 39568
rect 17316 39525 17325 39559
rect 17325 39525 17359 39559
rect 17359 39525 17368 39559
rect 17316 39516 17368 39525
rect 17132 39448 17184 39500
rect 17592 39491 17644 39500
rect 17592 39457 17601 39491
rect 17601 39457 17635 39491
rect 17635 39457 17644 39491
rect 17592 39448 17644 39457
rect 15108 39380 15160 39432
rect 18604 39559 18656 39568
rect 18604 39525 18613 39559
rect 18613 39525 18647 39559
rect 18647 39525 18656 39559
rect 18604 39516 18656 39525
rect 18696 39559 18748 39568
rect 18696 39525 18705 39559
rect 18705 39525 18739 39559
rect 18739 39525 18748 39559
rect 18696 39516 18748 39525
rect 20628 39516 20680 39568
rect 15200 39312 15252 39364
rect 15752 39355 15804 39364
rect 15752 39321 15761 39355
rect 15761 39321 15795 39355
rect 15795 39321 15804 39355
rect 15752 39312 15804 39321
rect 16304 39312 16356 39364
rect 14004 39244 14056 39296
rect 15108 39244 15160 39296
rect 17132 39244 17184 39296
rect 17500 39312 17552 39364
rect 18420 39423 18472 39432
rect 18420 39389 18429 39423
rect 18429 39389 18463 39423
rect 18463 39389 18472 39423
rect 18420 39380 18472 39389
rect 19248 39448 19300 39500
rect 20260 39491 20312 39500
rect 20260 39457 20269 39491
rect 20269 39457 20303 39491
rect 20303 39457 20312 39491
rect 20260 39448 20312 39457
rect 23112 39627 23164 39636
rect 23112 39593 23121 39627
rect 23121 39593 23155 39627
rect 23155 39593 23164 39627
rect 23112 39584 23164 39593
rect 23204 39559 23256 39568
rect 23204 39525 23213 39559
rect 23213 39525 23247 39559
rect 23247 39525 23256 39559
rect 23204 39516 23256 39525
rect 21088 39491 21140 39500
rect 21088 39457 21097 39491
rect 21097 39457 21131 39491
rect 21131 39457 21140 39491
rect 21088 39448 21140 39457
rect 21824 39448 21876 39500
rect 23848 39559 23900 39568
rect 19432 39423 19484 39432
rect 19432 39389 19441 39423
rect 19441 39389 19475 39423
rect 19475 39389 19484 39423
rect 19432 39380 19484 39389
rect 19524 39423 19576 39432
rect 19524 39389 19533 39423
rect 19533 39389 19567 39423
rect 19567 39389 19576 39423
rect 19524 39380 19576 39389
rect 19708 39423 19760 39432
rect 19708 39389 19717 39423
rect 19717 39389 19751 39423
rect 19751 39389 19760 39423
rect 19708 39380 19760 39389
rect 20168 39423 20220 39432
rect 20168 39389 20177 39423
rect 20177 39389 20211 39423
rect 20211 39389 20220 39423
rect 20168 39380 20220 39389
rect 22928 39423 22980 39432
rect 22928 39389 22937 39423
rect 22937 39389 22971 39423
rect 22971 39389 22980 39423
rect 22928 39380 22980 39389
rect 23848 39525 23857 39559
rect 23857 39525 23891 39559
rect 23891 39525 23900 39559
rect 23848 39516 23900 39525
rect 25044 39584 25096 39636
rect 25136 39627 25188 39636
rect 25136 39593 25145 39627
rect 25145 39593 25179 39627
rect 25179 39593 25188 39627
rect 25136 39584 25188 39593
rect 26516 39627 26568 39636
rect 26516 39593 26525 39627
rect 26525 39593 26559 39627
rect 26559 39593 26568 39627
rect 26516 39584 26568 39593
rect 26792 39627 26844 39636
rect 26792 39593 26801 39627
rect 26801 39593 26835 39627
rect 26835 39593 26844 39627
rect 26792 39584 26844 39593
rect 28172 39627 28224 39636
rect 28172 39593 28181 39627
rect 28181 39593 28215 39627
rect 28215 39593 28224 39627
rect 28172 39584 28224 39593
rect 30656 39584 30708 39636
rect 31024 39584 31076 39636
rect 31944 39584 31996 39636
rect 32036 39584 32088 39636
rect 32220 39627 32272 39636
rect 32220 39593 32229 39627
rect 32229 39593 32263 39627
rect 32263 39593 32272 39627
rect 32220 39584 32272 39593
rect 34704 39627 34756 39636
rect 34704 39593 34713 39627
rect 34713 39593 34747 39627
rect 34747 39593 34756 39627
rect 34704 39584 34756 39593
rect 24676 39516 24728 39568
rect 25228 39559 25280 39568
rect 25228 39525 25237 39559
rect 25237 39525 25271 39559
rect 25271 39525 25280 39559
rect 25228 39516 25280 39525
rect 27252 39559 27304 39568
rect 24308 39448 24360 39500
rect 27252 39525 27261 39559
rect 27261 39525 27295 39559
rect 27295 39525 27304 39559
rect 27252 39516 27304 39525
rect 28540 39559 28592 39568
rect 28540 39525 28549 39559
rect 28549 39525 28583 39559
rect 28583 39525 28592 39559
rect 28540 39516 28592 39525
rect 29184 39516 29236 39568
rect 30288 39516 30340 39568
rect 32312 39559 32364 39568
rect 32312 39525 32321 39559
rect 32321 39525 32355 39559
rect 32355 39525 32364 39559
rect 32312 39516 32364 39525
rect 35992 39584 36044 39636
rect 36084 39584 36136 39636
rect 37004 39584 37056 39636
rect 38936 39584 38988 39636
rect 39580 39627 39632 39636
rect 39580 39593 39589 39627
rect 39589 39593 39623 39627
rect 39623 39593 39632 39627
rect 39580 39584 39632 39593
rect 42156 39627 42208 39636
rect 20996 39312 21048 39364
rect 21548 39312 21600 39364
rect 23756 39423 23808 39432
rect 23756 39389 23765 39423
rect 23765 39389 23799 39423
rect 23799 39389 23808 39423
rect 23756 39380 23808 39389
rect 24032 39423 24084 39432
rect 24032 39389 24041 39423
rect 24041 39389 24075 39423
rect 24075 39389 24084 39423
rect 24032 39380 24084 39389
rect 24584 39423 24636 39432
rect 24584 39389 24593 39423
rect 24593 39389 24627 39423
rect 24627 39389 24636 39423
rect 24584 39380 24636 39389
rect 24124 39312 24176 39364
rect 23572 39244 23624 39296
rect 24032 39244 24084 39296
rect 25964 39312 26016 39364
rect 30840 39491 30892 39500
rect 30840 39457 30849 39491
rect 30849 39457 30883 39491
rect 30883 39457 30892 39491
rect 30840 39448 30892 39457
rect 31392 39448 31444 39500
rect 27160 39423 27212 39432
rect 27160 39389 27169 39423
rect 27169 39389 27203 39423
rect 27203 39389 27212 39423
rect 27160 39380 27212 39389
rect 27528 39380 27580 39432
rect 31024 39423 31076 39432
rect 29184 39312 29236 39364
rect 27160 39244 27212 39296
rect 31024 39389 31033 39423
rect 31033 39389 31067 39423
rect 31067 39389 31076 39423
rect 31024 39380 31076 39389
rect 32496 39448 32548 39500
rect 34796 39448 34848 39500
rect 31668 39423 31720 39432
rect 31668 39389 31677 39423
rect 31677 39389 31711 39423
rect 31711 39389 31720 39423
rect 31668 39380 31720 39389
rect 31760 39423 31812 39432
rect 31760 39389 31769 39423
rect 31769 39389 31803 39423
rect 31803 39389 31812 39423
rect 31760 39380 31812 39389
rect 31944 39423 31996 39432
rect 31944 39389 31953 39423
rect 31953 39389 31987 39423
rect 31987 39389 31996 39423
rect 31944 39380 31996 39389
rect 36084 39448 36136 39500
rect 37740 39448 37792 39500
rect 38200 39448 38252 39500
rect 39028 39516 39080 39568
rect 42156 39593 42165 39627
rect 42165 39593 42199 39627
rect 42199 39593 42208 39627
rect 42156 39584 42208 39593
rect 35624 39380 35676 39432
rect 35992 39380 36044 39432
rect 36176 39380 36228 39432
rect 31668 39244 31720 39296
rect 32772 39244 32824 39296
rect 34612 39244 34664 39296
rect 35532 39312 35584 39364
rect 37464 39312 37516 39364
rect 38936 39423 38988 39432
rect 38936 39389 38945 39423
rect 38945 39389 38979 39423
rect 38979 39389 38988 39423
rect 38936 39380 38988 39389
rect 39396 39423 39448 39432
rect 39396 39389 39405 39423
rect 39405 39389 39439 39423
rect 39439 39389 39448 39423
rect 39396 39380 39448 39389
rect 39948 39423 40000 39432
rect 39948 39389 39957 39423
rect 39957 39389 39991 39423
rect 39991 39389 40000 39423
rect 39948 39380 40000 39389
rect 40224 39380 40276 39432
rect 40776 39448 40828 39500
rect 39580 39312 39632 39364
rect 40040 39312 40092 39364
rect 40132 39355 40184 39364
rect 40132 39321 40141 39355
rect 40141 39321 40175 39355
rect 40175 39321 40184 39355
rect 40132 39312 40184 39321
rect 40684 39355 40736 39364
rect 40684 39321 40693 39355
rect 40693 39321 40727 39355
rect 40727 39321 40736 39355
rect 40684 39312 40736 39321
rect 41420 39312 41472 39364
rect 36176 39287 36228 39296
rect 36176 39253 36185 39287
rect 36185 39253 36219 39287
rect 36219 39253 36228 39287
rect 36176 39244 36228 39253
rect 37096 39244 37148 39296
rect 38292 39287 38344 39296
rect 38292 39253 38301 39287
rect 38301 39253 38335 39287
rect 38335 39253 38344 39287
rect 38292 39244 38344 39253
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 15752 39040 15804 39092
rect 18420 39040 18472 39092
rect 19524 39040 19576 39092
rect 20168 39040 20220 39092
rect 20260 39040 20312 39092
rect 23756 39040 23808 39092
rect 24584 39040 24636 39092
rect 25228 39083 25280 39092
rect 25228 39049 25237 39083
rect 25237 39049 25271 39083
rect 25271 39049 25280 39083
rect 25228 39040 25280 39049
rect 32312 39040 32364 39092
rect 32496 39083 32548 39092
rect 32496 39049 32505 39083
rect 32505 39049 32539 39083
rect 32539 39049 32548 39083
rect 32496 39040 32548 39049
rect 32772 39083 32824 39092
rect 32772 39049 32781 39083
rect 32781 39049 32815 39083
rect 32815 39049 32824 39083
rect 32772 39040 32824 39049
rect 35348 39040 35400 39092
rect 35808 39083 35860 39092
rect 35808 39049 35817 39083
rect 35817 39049 35851 39083
rect 35851 39049 35860 39083
rect 35808 39040 35860 39049
rect 35992 39040 36044 39092
rect 36176 39040 36228 39092
rect 3608 38947 3660 38956
rect 3608 38913 3617 38947
rect 3617 38913 3651 38947
rect 3651 38913 3660 38947
rect 3608 38904 3660 38913
rect 14556 38904 14608 38956
rect 12900 38836 12952 38888
rect 14096 38836 14148 38888
rect 15200 38904 15252 38956
rect 16028 38904 16080 38956
rect 17500 38947 17552 38956
rect 17500 38913 17509 38947
rect 17509 38913 17543 38947
rect 17543 38913 17552 38947
rect 17500 38904 17552 38913
rect 17684 38947 17736 38956
rect 17684 38913 17693 38947
rect 17693 38913 17727 38947
rect 17727 38913 17736 38947
rect 17684 38904 17736 38913
rect 17132 38879 17184 38888
rect 17132 38845 17141 38879
rect 17141 38845 17175 38879
rect 17175 38845 17184 38879
rect 17132 38836 17184 38845
rect 19248 38947 19300 38956
rect 19248 38913 19257 38947
rect 19257 38913 19291 38947
rect 19291 38913 19300 38947
rect 19248 38904 19300 38913
rect 27160 38972 27212 39024
rect 19524 38904 19576 38956
rect 20996 38947 21048 38956
rect 20996 38913 21035 38947
rect 21035 38913 21048 38947
rect 20996 38904 21048 38913
rect 22100 38904 22152 38956
rect 22928 38904 22980 38956
rect 14740 38768 14792 38820
rect 19708 38836 19760 38888
rect 23756 38947 23808 38956
rect 23756 38913 23765 38947
rect 23765 38913 23799 38947
rect 23799 38913 23808 38947
rect 23756 38904 23808 38913
rect 23940 38947 23992 38956
rect 23940 38913 23949 38947
rect 23949 38913 23983 38947
rect 23983 38913 23992 38947
rect 23940 38904 23992 38913
rect 24124 38836 24176 38888
rect 25136 38947 25188 38956
rect 25136 38913 25145 38947
rect 25145 38913 25179 38947
rect 25179 38913 25188 38947
rect 25136 38904 25188 38913
rect 25228 38947 25280 38956
rect 25228 38913 25237 38947
rect 25237 38913 25271 38947
rect 25271 38913 25280 38947
rect 25228 38904 25280 38913
rect 25688 38904 25740 38956
rect 27528 38904 27580 38956
rect 37464 39040 37516 39092
rect 37924 39040 37976 39092
rect 38476 39040 38528 39092
rect 39948 39083 40000 39092
rect 39948 39049 39957 39083
rect 39957 39049 39991 39083
rect 39991 39049 40000 39083
rect 39948 39040 40000 39049
rect 40040 39040 40092 39092
rect 40684 39083 40736 39092
rect 40684 39049 40693 39083
rect 40693 39049 40727 39083
rect 40727 39049 40736 39083
rect 40684 39040 40736 39049
rect 41052 39083 41104 39092
rect 41052 39049 41061 39083
rect 41061 39049 41095 39083
rect 41095 39049 41104 39083
rect 41052 39040 41104 39049
rect 25964 38836 26016 38888
rect 28540 38904 28592 38956
rect 30196 38904 30248 38956
rect 30564 38904 30616 38956
rect 30748 38947 30800 38956
rect 30748 38913 30757 38947
rect 30757 38913 30791 38947
rect 30791 38913 30800 38947
rect 30748 38904 30800 38913
rect 31024 38947 31076 38956
rect 31024 38913 31033 38947
rect 31033 38913 31067 38947
rect 31067 38913 31076 38947
rect 31024 38904 31076 38913
rect 27988 38836 28040 38888
rect 17500 38768 17552 38820
rect 23572 38811 23624 38820
rect 23572 38777 23581 38811
rect 23581 38777 23615 38811
rect 23615 38777 23624 38811
rect 23572 38768 23624 38777
rect 27252 38768 27304 38820
rect 30932 38768 30984 38820
rect 31944 38904 31996 38956
rect 32496 38947 32548 38956
rect 32496 38913 32505 38947
rect 32505 38913 32539 38947
rect 32539 38913 32548 38947
rect 32496 38904 32548 38913
rect 32772 38937 32824 38946
rect 32772 38903 32781 38937
rect 32781 38903 32815 38937
rect 32815 38903 32824 38937
rect 32772 38894 32824 38903
rect 33048 38947 33100 38956
rect 33048 38913 33057 38947
rect 33057 38913 33091 38947
rect 33091 38913 33100 38947
rect 33048 38904 33100 38913
rect 34428 38904 34480 38956
rect 35348 38947 35400 38956
rect 35348 38913 35357 38947
rect 35357 38913 35391 38947
rect 35391 38913 35400 38947
rect 35348 38904 35400 38913
rect 32680 38879 32732 38888
rect 32680 38845 32689 38879
rect 32689 38845 32723 38879
rect 32723 38845 32732 38879
rect 32680 38836 32732 38845
rect 35992 38904 36044 38956
rect 39396 38904 39448 38956
rect 35900 38879 35952 38888
rect 35900 38845 35909 38879
rect 35909 38845 35943 38879
rect 35943 38845 35952 38879
rect 35900 38836 35952 38845
rect 37372 38836 37424 38888
rect 39120 38879 39172 38888
rect 39120 38845 39129 38879
rect 39129 38845 39163 38879
rect 39163 38845 39172 38879
rect 39120 38836 39172 38845
rect 40132 38947 40184 38956
rect 40132 38913 40141 38947
rect 40141 38913 40175 38947
rect 40175 38913 40184 38947
rect 40132 38904 40184 38913
rect 40224 38904 40276 38956
rect 41788 38904 41840 38956
rect 41144 38879 41196 38888
rect 41144 38845 41153 38879
rect 41153 38845 41187 38879
rect 41187 38845 41196 38879
rect 41144 38836 41196 38845
rect 3240 38700 3292 38752
rect 15016 38743 15068 38752
rect 15016 38709 15025 38743
rect 15025 38709 15059 38743
rect 15059 38709 15068 38743
rect 15016 38700 15068 38709
rect 31392 38700 31444 38752
rect 35532 38811 35584 38820
rect 35532 38777 35541 38811
rect 35541 38777 35575 38811
rect 35575 38777 35584 38811
rect 35532 38768 35584 38777
rect 32680 38700 32732 38752
rect 32956 38700 33008 38752
rect 35348 38700 35400 38752
rect 35900 38700 35952 38752
rect 36084 38743 36136 38752
rect 36084 38709 36093 38743
rect 36093 38709 36127 38743
rect 36127 38709 36136 38743
rect 36084 38700 36136 38709
rect 37372 38700 37424 38752
rect 38936 38768 38988 38820
rect 39672 38768 39724 38820
rect 41052 38768 41104 38820
rect 40500 38700 40552 38752
rect 40868 38700 40920 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1400 38360 1452 38412
rect 3792 38360 3844 38412
rect 3424 38292 3476 38344
rect 5264 38360 5316 38412
rect 6092 38335 6144 38344
rect 6092 38301 6101 38335
rect 6101 38301 6135 38335
rect 6135 38301 6144 38335
rect 6092 38292 6144 38301
rect 7288 38496 7340 38548
rect 14096 38539 14148 38548
rect 14096 38505 14105 38539
rect 14105 38505 14139 38539
rect 14139 38505 14148 38539
rect 14096 38496 14148 38505
rect 19524 38539 19576 38548
rect 19524 38505 19533 38539
rect 19533 38505 19567 38539
rect 19567 38505 19576 38539
rect 19524 38496 19576 38505
rect 19708 38539 19760 38548
rect 19708 38505 19717 38539
rect 19717 38505 19751 38539
rect 19751 38505 19760 38539
rect 19708 38496 19760 38505
rect 20996 38496 21048 38548
rect 21272 38496 21324 38548
rect 13820 38428 13872 38480
rect 19616 38428 19668 38480
rect 7104 38360 7156 38412
rect 8300 38360 8352 38412
rect 14740 38403 14792 38412
rect 14740 38369 14749 38403
rect 14749 38369 14783 38403
rect 14783 38369 14792 38403
rect 14740 38360 14792 38369
rect 19524 38360 19576 38412
rect 22100 38496 22152 38548
rect 23756 38496 23808 38548
rect 23940 38496 23992 38548
rect 25228 38539 25280 38548
rect 25228 38505 25237 38539
rect 25237 38505 25271 38539
rect 25271 38505 25280 38539
rect 25228 38496 25280 38505
rect 25596 38496 25648 38548
rect 25688 38496 25740 38548
rect 28540 38539 28592 38548
rect 28540 38505 28549 38539
rect 28549 38505 28583 38539
rect 28583 38505 28592 38539
rect 28540 38496 28592 38505
rect 29184 38539 29236 38548
rect 29184 38505 29193 38539
rect 29193 38505 29227 38539
rect 29227 38505 29236 38539
rect 29184 38496 29236 38505
rect 31024 38496 31076 38548
rect 22284 38428 22336 38480
rect 6828 38335 6880 38344
rect 6828 38301 6837 38335
rect 6837 38301 6871 38335
rect 6871 38301 6880 38335
rect 6828 38292 6880 38301
rect 11612 38292 11664 38344
rect 15016 38292 15068 38344
rect 19248 38335 19300 38344
rect 19248 38301 19257 38335
rect 19257 38301 19291 38335
rect 19291 38301 19300 38335
rect 19248 38292 19300 38301
rect 19432 38292 19484 38344
rect 19892 38335 19944 38344
rect 19892 38301 19901 38335
rect 19901 38301 19935 38335
rect 19935 38301 19944 38335
rect 19892 38292 19944 38301
rect 20996 38292 21048 38344
rect 21272 38335 21324 38344
rect 21272 38301 21281 38335
rect 21281 38301 21315 38335
rect 21315 38301 21324 38335
rect 21272 38292 21324 38301
rect 21640 38292 21692 38344
rect 22284 38335 22336 38344
rect 22284 38301 22293 38335
rect 22293 38301 22327 38335
rect 22327 38301 22336 38335
rect 22284 38292 22336 38301
rect 22376 38335 22428 38344
rect 22376 38301 22385 38335
rect 22385 38301 22419 38335
rect 22419 38301 22428 38335
rect 22376 38292 22428 38301
rect 25596 38360 25648 38412
rect 25964 38471 26016 38480
rect 25964 38437 25973 38471
rect 25973 38437 26007 38471
rect 26007 38437 26016 38471
rect 25964 38428 26016 38437
rect 28908 38428 28960 38480
rect 1952 38267 2004 38276
rect 1952 38233 1961 38267
rect 1961 38233 1995 38267
rect 1995 38233 2004 38267
rect 1952 38224 2004 38233
rect 2964 38224 3016 38276
rect 2596 38156 2648 38208
rect 3424 38199 3476 38208
rect 3424 38165 3433 38199
rect 3433 38165 3467 38199
rect 3467 38165 3476 38199
rect 3424 38156 3476 38165
rect 3516 38156 3568 38208
rect 4712 38156 4764 38208
rect 4804 38156 4856 38208
rect 5448 38267 5500 38276
rect 5448 38233 5457 38267
rect 5457 38233 5491 38267
rect 5491 38233 5500 38267
rect 5448 38224 5500 38233
rect 5908 38199 5960 38208
rect 5908 38165 5917 38199
rect 5917 38165 5951 38199
rect 5951 38165 5960 38199
rect 5908 38156 5960 38165
rect 6460 38224 6512 38276
rect 7012 38224 7064 38276
rect 9680 38224 9732 38276
rect 12072 38267 12124 38276
rect 12072 38233 12081 38267
rect 12081 38233 12115 38267
rect 12115 38233 12124 38267
rect 12072 38224 12124 38233
rect 14372 38224 14424 38276
rect 19524 38267 19576 38276
rect 19524 38233 19533 38267
rect 19533 38233 19567 38267
rect 19567 38233 19576 38267
rect 19524 38224 19576 38233
rect 7932 38156 7984 38208
rect 8944 38199 8996 38208
rect 8944 38165 8953 38199
rect 8953 38165 8987 38199
rect 8987 38165 8996 38199
rect 8944 38156 8996 38165
rect 14648 38156 14700 38208
rect 19248 38156 19300 38208
rect 21364 38224 21416 38276
rect 23940 38267 23992 38276
rect 23940 38233 23949 38267
rect 23949 38233 23983 38267
rect 23983 38233 23992 38267
rect 25412 38335 25464 38344
rect 25412 38301 25421 38335
rect 25421 38301 25455 38335
rect 25455 38301 25464 38335
rect 25412 38292 25464 38301
rect 25688 38335 25740 38344
rect 25688 38301 25697 38335
rect 25697 38301 25731 38335
rect 25731 38301 25740 38335
rect 25688 38292 25740 38301
rect 23940 38224 23992 38233
rect 26148 38292 26200 38344
rect 36912 38496 36964 38548
rect 37556 38496 37608 38548
rect 40316 38496 40368 38548
rect 32772 38360 32824 38412
rect 34796 38360 34848 38412
rect 37372 38403 37424 38412
rect 37372 38369 37381 38403
rect 37381 38369 37415 38403
rect 37415 38369 37424 38403
rect 37372 38360 37424 38369
rect 28172 38292 28224 38344
rect 28632 38267 28684 38276
rect 28632 38233 28641 38267
rect 28641 38233 28675 38267
rect 28675 38233 28684 38267
rect 28632 38224 28684 38233
rect 28908 38335 28960 38344
rect 28908 38301 28917 38335
rect 28917 38301 28951 38335
rect 28951 38301 28960 38335
rect 28908 38292 28960 38301
rect 32404 38335 32456 38344
rect 32404 38301 32413 38335
rect 32413 38301 32447 38335
rect 32447 38301 32456 38335
rect 32404 38292 32456 38301
rect 29184 38267 29236 38276
rect 29184 38233 29193 38267
rect 29193 38233 29227 38267
rect 29227 38233 29236 38267
rect 29184 38224 29236 38233
rect 29552 38224 29604 38276
rect 32312 38224 32364 38276
rect 32680 38267 32732 38276
rect 32680 38233 32689 38267
rect 32689 38233 32723 38267
rect 32723 38233 32732 38267
rect 32680 38224 32732 38233
rect 33232 38224 33284 38276
rect 21824 38156 21876 38208
rect 22560 38156 22612 38208
rect 25136 38156 25188 38208
rect 26056 38156 26108 38208
rect 31392 38199 31444 38208
rect 31392 38165 31401 38199
rect 31401 38165 31435 38199
rect 31435 38165 31444 38199
rect 31392 38156 31444 38165
rect 33692 38156 33744 38208
rect 35808 38335 35860 38344
rect 35808 38301 35817 38335
rect 35817 38301 35851 38335
rect 35851 38301 35860 38335
rect 35808 38292 35860 38301
rect 37924 38335 37976 38344
rect 37924 38301 37933 38335
rect 37933 38301 37967 38335
rect 37967 38301 37976 38335
rect 37924 38292 37976 38301
rect 41052 38403 41104 38412
rect 41052 38369 41061 38403
rect 41061 38369 41095 38403
rect 41095 38369 41104 38403
rect 41052 38360 41104 38369
rect 38292 38292 38344 38344
rect 39120 38292 39172 38344
rect 39396 38292 39448 38344
rect 40868 38335 40920 38344
rect 40868 38301 40877 38335
rect 40877 38301 40911 38335
rect 40911 38301 40920 38335
rect 40868 38292 40920 38301
rect 41880 38335 41932 38344
rect 41880 38301 41889 38335
rect 41889 38301 41923 38335
rect 41923 38301 41932 38335
rect 41880 38292 41932 38301
rect 40592 38224 40644 38276
rect 34704 38199 34756 38208
rect 34704 38165 34713 38199
rect 34713 38165 34747 38199
rect 34747 38165 34756 38199
rect 34704 38156 34756 38165
rect 35440 38199 35492 38208
rect 35440 38165 35449 38199
rect 35449 38165 35483 38199
rect 35483 38165 35492 38199
rect 35440 38156 35492 38165
rect 40960 38199 41012 38208
rect 40960 38165 40969 38199
rect 40969 38165 41003 38199
rect 41003 38165 41012 38199
rect 40960 38156 41012 38165
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 1952 37952 2004 38004
rect 5816 37952 5868 38004
rect 6092 37952 6144 38004
rect 7012 37995 7064 38004
rect 7012 37961 7021 37995
rect 7021 37961 7055 37995
rect 7055 37961 7064 37995
rect 7012 37952 7064 37961
rect 6460 37884 6512 37936
rect 7472 37952 7524 38004
rect 15108 37952 15160 38004
rect 1860 37859 1912 37868
rect 1860 37825 1869 37859
rect 1869 37825 1903 37859
rect 1903 37825 1912 37859
rect 1860 37816 1912 37825
rect 2044 37859 2096 37868
rect 2044 37825 2053 37859
rect 2053 37825 2087 37859
rect 2087 37825 2096 37859
rect 2044 37816 2096 37825
rect 2596 37859 2648 37868
rect 2596 37825 2605 37859
rect 2605 37825 2639 37859
rect 2639 37825 2648 37859
rect 2596 37816 2648 37825
rect 3516 37816 3568 37868
rect 5540 37816 5592 37868
rect 6920 37816 6972 37868
rect 3332 37748 3384 37800
rect 3700 37791 3752 37800
rect 3700 37757 3709 37791
rect 3709 37757 3743 37791
rect 3743 37757 3752 37791
rect 3700 37748 3752 37757
rect 3792 37791 3844 37800
rect 3792 37757 3801 37791
rect 3801 37757 3835 37791
rect 3835 37757 3844 37791
rect 3792 37748 3844 37757
rect 4620 37748 4672 37800
rect 5172 37680 5224 37732
rect 5448 37680 5500 37732
rect 6644 37791 6696 37800
rect 6644 37757 6653 37791
rect 6653 37757 6687 37791
rect 6687 37757 6696 37791
rect 6644 37748 6696 37757
rect 7012 37748 7064 37800
rect 7288 37859 7340 37868
rect 7288 37825 7297 37859
rect 7297 37825 7331 37859
rect 7331 37825 7340 37859
rect 7288 37816 7340 37825
rect 7380 37859 7432 37868
rect 7380 37825 7389 37859
rect 7389 37825 7423 37859
rect 7423 37825 7432 37859
rect 7380 37816 7432 37825
rect 7472 37859 7524 37868
rect 7472 37825 7507 37859
rect 7507 37825 7524 37859
rect 7472 37816 7524 37825
rect 8944 37884 8996 37936
rect 8024 37816 8076 37868
rect 2872 37612 2924 37664
rect 3148 37612 3200 37664
rect 4804 37612 4856 37664
rect 8024 37680 8076 37732
rect 8116 37680 8168 37732
rect 14464 37816 14516 37868
rect 12900 37748 12952 37800
rect 14096 37748 14148 37800
rect 8576 37680 8628 37732
rect 16856 37859 16908 37868
rect 16856 37825 16865 37859
rect 16865 37825 16899 37859
rect 16899 37825 16908 37859
rect 16856 37816 16908 37825
rect 19248 37952 19300 38004
rect 19432 37952 19484 38004
rect 19616 37952 19668 38004
rect 20076 37884 20128 37936
rect 22376 37884 22428 37936
rect 17684 37748 17736 37800
rect 21364 37816 21416 37868
rect 22652 37816 22704 37868
rect 24124 37859 24176 37868
rect 24124 37825 24133 37859
rect 24133 37825 24167 37859
rect 24167 37825 24176 37859
rect 24124 37816 24176 37825
rect 27068 37859 27120 37868
rect 27068 37825 27077 37859
rect 27077 37825 27111 37859
rect 27111 37825 27120 37859
rect 27068 37816 27120 37825
rect 19892 37748 19944 37800
rect 20996 37791 21048 37800
rect 20996 37757 21005 37791
rect 21005 37757 21039 37791
rect 21039 37757 21048 37791
rect 20996 37748 21048 37757
rect 22468 37791 22520 37800
rect 22468 37757 22477 37791
rect 22477 37757 22511 37791
rect 22511 37757 22520 37791
rect 22468 37748 22520 37757
rect 25412 37680 25464 37732
rect 8392 37612 8444 37664
rect 18972 37612 19024 37664
rect 19616 37612 19668 37664
rect 22100 37612 22152 37664
rect 23572 37655 23624 37664
rect 23572 37621 23581 37655
rect 23581 37621 23615 37655
rect 23615 37621 23624 37655
rect 23572 37612 23624 37621
rect 27620 37995 27672 38004
rect 27620 37961 27635 37995
rect 27635 37961 27669 37995
rect 27669 37961 27672 37995
rect 27620 37952 27672 37961
rect 27988 37995 28040 38004
rect 27988 37961 27997 37995
rect 27997 37961 28031 37995
rect 28031 37961 28040 37995
rect 27988 37952 28040 37961
rect 28632 37995 28684 38004
rect 28632 37961 28641 37995
rect 28641 37961 28675 37995
rect 28675 37961 28684 37995
rect 28632 37952 28684 37961
rect 28908 37952 28960 38004
rect 29552 37995 29604 38004
rect 29552 37961 29561 37995
rect 29561 37961 29595 37995
rect 29595 37961 29604 37995
rect 29552 37952 29604 37961
rect 31392 37952 31444 38004
rect 32680 37952 32732 38004
rect 34704 37952 34756 38004
rect 34796 37995 34848 38004
rect 34796 37961 34805 37995
rect 34805 37961 34839 37995
rect 34839 37961 34848 37995
rect 34796 37952 34848 37961
rect 35992 37995 36044 38004
rect 35992 37961 36001 37995
rect 36001 37961 36035 37995
rect 36035 37961 36044 37995
rect 35992 37952 36044 37961
rect 37924 37952 37976 38004
rect 40500 37995 40552 38004
rect 40500 37961 40509 37995
rect 40509 37961 40543 37995
rect 40543 37961 40552 37995
rect 40500 37952 40552 37961
rect 30748 37884 30800 37936
rect 27896 37859 27948 37868
rect 27896 37825 27905 37859
rect 27905 37825 27939 37859
rect 27939 37825 27948 37859
rect 27896 37816 27948 37825
rect 27988 37748 28040 37800
rect 28908 37816 28960 37868
rect 29276 37859 29328 37868
rect 29276 37825 29285 37859
rect 29285 37825 29319 37859
rect 29319 37825 29328 37859
rect 29276 37816 29328 37825
rect 30196 37816 30248 37868
rect 30564 37859 30616 37868
rect 30564 37825 30573 37859
rect 30573 37825 30607 37859
rect 30607 37825 30616 37859
rect 30564 37816 30616 37825
rect 31300 37816 31352 37868
rect 32404 37884 32456 37936
rect 32956 37884 33008 37936
rect 35440 37884 35492 37936
rect 39856 37884 39908 37936
rect 32128 37859 32180 37868
rect 32128 37825 32137 37859
rect 32137 37825 32171 37859
rect 32171 37825 32180 37859
rect 32128 37816 32180 37825
rect 33140 37859 33192 37868
rect 33140 37825 33149 37859
rect 33149 37825 33183 37859
rect 33183 37825 33192 37859
rect 33140 37816 33192 37825
rect 30012 37791 30064 37800
rect 30012 37757 30021 37791
rect 30021 37757 30055 37791
rect 30055 37757 30064 37791
rect 30012 37748 30064 37757
rect 30104 37791 30156 37800
rect 30104 37757 30113 37791
rect 30113 37757 30147 37791
rect 30147 37757 30156 37791
rect 30104 37748 30156 37757
rect 33416 37816 33468 37868
rect 34244 37748 34296 37800
rect 35440 37748 35492 37800
rect 36452 37791 36504 37800
rect 36452 37757 36461 37791
rect 36461 37757 36495 37791
rect 36495 37757 36504 37791
rect 36452 37748 36504 37757
rect 37648 37816 37700 37868
rect 38476 37816 38528 37868
rect 39948 37859 40000 37868
rect 39948 37825 39957 37859
rect 39957 37825 39991 37859
rect 39991 37825 40000 37859
rect 39948 37816 40000 37825
rect 40040 37816 40092 37868
rect 40316 37816 40368 37868
rect 40684 37859 40736 37868
rect 40684 37825 40693 37859
rect 40693 37825 40727 37859
rect 40727 37825 40736 37859
rect 40684 37816 40736 37825
rect 40776 37816 40828 37868
rect 41696 37816 41748 37868
rect 28908 37612 28960 37664
rect 34520 37680 34572 37732
rect 37372 37680 37424 37732
rect 37464 37612 37516 37664
rect 37740 37723 37792 37732
rect 37740 37689 37749 37723
rect 37749 37689 37783 37723
rect 37783 37689 37792 37723
rect 37740 37680 37792 37689
rect 38292 37680 38344 37732
rect 41512 37680 41564 37732
rect 39396 37612 39448 37664
rect 40316 37655 40368 37664
rect 40316 37621 40325 37655
rect 40325 37621 40359 37655
rect 40359 37621 40368 37655
rect 40316 37612 40368 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1860 37408 1912 37460
rect 3424 37451 3476 37460
rect 3424 37417 3433 37451
rect 3433 37417 3467 37451
rect 3467 37417 3476 37451
rect 3424 37408 3476 37417
rect 5908 37408 5960 37460
rect 7012 37451 7064 37460
rect 7012 37417 7021 37451
rect 7021 37417 7055 37451
rect 7055 37417 7064 37451
rect 7012 37408 7064 37417
rect 7288 37408 7340 37460
rect 12072 37451 12124 37460
rect 12072 37417 12081 37451
rect 12081 37417 12115 37451
rect 12115 37417 12124 37451
rect 12072 37408 12124 37417
rect 1400 37315 1452 37324
rect 1400 37281 1409 37315
rect 1409 37281 1443 37315
rect 1443 37281 1452 37315
rect 1400 37272 1452 37281
rect 2044 37272 2096 37324
rect 3700 37340 3752 37392
rect 4068 37340 4120 37392
rect 4160 37340 4212 37392
rect 5172 37340 5224 37392
rect 3792 37272 3844 37324
rect 2780 37204 2832 37256
rect 2964 37204 3016 37256
rect 1676 37179 1728 37188
rect 1676 37145 1685 37179
rect 1685 37145 1719 37179
rect 1719 37145 1728 37179
rect 1676 37136 1728 37145
rect 4804 37136 4856 37188
rect 5172 37247 5224 37256
rect 5172 37213 5181 37247
rect 5181 37213 5215 37247
rect 5215 37213 5224 37247
rect 5172 37204 5224 37213
rect 6828 37272 6880 37324
rect 7932 37340 7984 37392
rect 14096 37451 14148 37460
rect 14096 37417 14105 37451
rect 14105 37417 14139 37451
rect 14139 37417 14148 37451
rect 14096 37408 14148 37417
rect 14464 37408 14516 37460
rect 15108 37408 15160 37460
rect 20996 37408 21048 37460
rect 24124 37408 24176 37460
rect 26056 37408 26108 37460
rect 26332 37408 26384 37460
rect 27988 37451 28040 37460
rect 27988 37417 27997 37451
rect 27997 37417 28031 37451
rect 28031 37417 28040 37451
rect 27988 37408 28040 37417
rect 34244 37451 34296 37460
rect 34244 37417 34253 37451
rect 34253 37417 34287 37451
rect 34287 37417 34296 37451
rect 34244 37408 34296 37417
rect 36452 37451 36504 37460
rect 36452 37417 36461 37451
rect 36461 37417 36495 37451
rect 36495 37417 36504 37451
rect 36452 37408 36504 37417
rect 39396 37451 39448 37460
rect 39396 37417 39405 37451
rect 39405 37417 39439 37451
rect 39439 37417 39448 37451
rect 39396 37408 39448 37417
rect 39856 37408 39908 37460
rect 14556 37340 14608 37392
rect 14740 37340 14792 37392
rect 7104 37247 7156 37256
rect 7104 37213 7113 37247
rect 7113 37213 7147 37247
rect 7147 37213 7156 37247
rect 7104 37204 7156 37213
rect 8300 37204 8352 37256
rect 4160 37068 4212 37120
rect 4436 37068 4488 37120
rect 5356 37068 5408 37120
rect 5540 37068 5592 37120
rect 6368 37068 6420 37120
rect 6920 37136 6972 37188
rect 8576 37247 8628 37256
rect 8576 37213 8585 37247
rect 8585 37213 8619 37247
rect 8619 37213 8628 37247
rect 8576 37204 8628 37213
rect 9680 37272 9732 37324
rect 7472 37068 7524 37120
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 8116 37068 8168 37120
rect 8392 37111 8444 37120
rect 8392 37077 8401 37111
rect 8401 37077 8435 37111
rect 8435 37077 8444 37111
rect 12256 37247 12308 37256
rect 12256 37213 12265 37247
rect 12265 37213 12299 37247
rect 12299 37213 12308 37247
rect 12256 37204 12308 37213
rect 12532 37204 12584 37256
rect 14372 37204 14424 37256
rect 15016 37272 15068 37324
rect 14556 37247 14608 37256
rect 14556 37213 14565 37247
rect 14565 37213 14599 37247
rect 14599 37213 14608 37247
rect 14556 37204 14608 37213
rect 12164 37136 12216 37188
rect 12900 37136 12952 37188
rect 17316 37272 17368 37324
rect 17684 37272 17736 37324
rect 19708 37272 19760 37324
rect 22100 37315 22152 37324
rect 22100 37281 22109 37315
rect 22109 37281 22143 37315
rect 22143 37281 22152 37315
rect 22100 37272 22152 37281
rect 25044 37272 25096 37324
rect 28908 37340 28960 37392
rect 30564 37340 30616 37392
rect 35348 37340 35400 37392
rect 30104 37272 30156 37324
rect 17592 37204 17644 37256
rect 17776 37204 17828 37256
rect 18788 37247 18840 37256
rect 18788 37213 18797 37247
rect 18797 37213 18831 37247
rect 18831 37213 18840 37247
rect 18788 37204 18840 37213
rect 18972 37247 19024 37256
rect 18972 37213 18981 37247
rect 18981 37213 19015 37247
rect 19015 37213 19024 37247
rect 18972 37204 19024 37213
rect 16212 37136 16264 37188
rect 19616 37247 19668 37256
rect 19616 37213 19625 37247
rect 19625 37213 19659 37247
rect 19659 37213 19668 37247
rect 19616 37204 19668 37213
rect 8392 37068 8444 37077
rect 14556 37068 14608 37120
rect 15384 37068 15436 37120
rect 21548 37136 21600 37188
rect 22192 37136 22244 37188
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 25780 37204 25832 37256
rect 22652 37136 22704 37188
rect 22744 37179 22796 37188
rect 22744 37145 22753 37179
rect 22753 37145 22787 37179
rect 22787 37145 22796 37179
rect 22744 37136 22796 37145
rect 25136 37136 25188 37188
rect 17776 37111 17828 37120
rect 17776 37077 17785 37111
rect 17785 37077 17819 37111
rect 17819 37077 17828 37111
rect 17776 37068 17828 37077
rect 17868 37111 17920 37120
rect 17868 37077 17877 37111
rect 17877 37077 17911 37111
rect 17911 37077 17920 37111
rect 17868 37068 17920 37077
rect 19248 37111 19300 37120
rect 19248 37077 19257 37111
rect 19257 37077 19291 37111
rect 19291 37077 19300 37111
rect 19248 37068 19300 37077
rect 19800 37068 19852 37120
rect 24400 37068 24452 37120
rect 29460 37204 29512 37256
rect 29552 37204 29604 37256
rect 30196 37247 30248 37256
rect 30196 37213 30205 37247
rect 30205 37213 30239 37247
rect 30239 37213 30248 37247
rect 30196 37204 30248 37213
rect 31852 37204 31904 37256
rect 31944 37204 31996 37256
rect 32772 37204 32824 37256
rect 33140 37247 33192 37256
rect 33140 37213 33149 37247
rect 33149 37213 33183 37247
rect 33183 37213 33192 37247
rect 33140 37204 33192 37213
rect 33968 37247 34020 37256
rect 33968 37213 33977 37247
rect 33977 37213 34011 37247
rect 34011 37213 34020 37247
rect 33968 37204 34020 37213
rect 34152 37247 34204 37256
rect 34152 37213 34161 37247
rect 34161 37213 34195 37247
rect 34195 37213 34204 37247
rect 36912 37340 36964 37392
rect 37464 37383 37516 37392
rect 37464 37349 37473 37383
rect 37473 37349 37507 37383
rect 37507 37349 37516 37383
rect 37464 37340 37516 37349
rect 37740 37340 37792 37392
rect 34152 37204 34204 37213
rect 26516 37179 26568 37188
rect 26516 37145 26525 37179
rect 26525 37145 26559 37179
rect 26559 37145 26568 37179
rect 26516 37136 26568 37145
rect 28172 37136 28224 37188
rect 31392 37136 31444 37188
rect 28080 37111 28132 37120
rect 28080 37077 28089 37111
rect 28089 37077 28123 37111
rect 28123 37077 28132 37111
rect 28080 37068 28132 37077
rect 29644 37111 29696 37120
rect 29644 37077 29653 37111
rect 29653 37077 29687 37111
rect 29687 37077 29696 37111
rect 29644 37068 29696 37077
rect 30472 37068 30524 37120
rect 31668 37111 31720 37120
rect 31668 37077 31677 37111
rect 31677 37077 31711 37111
rect 31711 37077 31720 37111
rect 31668 37068 31720 37077
rect 32496 37068 32548 37120
rect 34520 37136 34572 37188
rect 35256 37247 35308 37256
rect 35256 37213 35265 37247
rect 35265 37213 35299 37247
rect 35299 37213 35308 37247
rect 35256 37204 35308 37213
rect 35348 37247 35400 37256
rect 35348 37213 35357 37247
rect 35357 37213 35391 37247
rect 35391 37213 35400 37247
rect 35348 37204 35400 37213
rect 35440 37247 35492 37256
rect 35440 37213 35449 37247
rect 35449 37213 35483 37247
rect 35483 37213 35492 37247
rect 35440 37204 35492 37213
rect 37372 37247 37424 37256
rect 37372 37213 37381 37247
rect 37381 37213 37415 37247
rect 37415 37213 37424 37247
rect 37372 37204 37424 37213
rect 37648 37247 37700 37256
rect 37648 37213 37657 37247
rect 37657 37213 37691 37247
rect 37691 37213 37700 37247
rect 37648 37204 37700 37213
rect 40776 37272 40828 37324
rect 35992 37179 36044 37188
rect 33416 37068 33468 37120
rect 35992 37145 36001 37179
rect 36001 37145 36035 37179
rect 36035 37145 36044 37179
rect 35992 37136 36044 37145
rect 36912 37136 36964 37188
rect 39948 37204 40000 37256
rect 40040 37247 40092 37256
rect 40040 37213 40049 37247
rect 40049 37213 40083 37247
rect 40083 37213 40092 37247
rect 40040 37204 40092 37213
rect 36268 37068 36320 37120
rect 40316 37136 40368 37188
rect 40408 37179 40460 37188
rect 40408 37145 40417 37179
rect 40417 37145 40451 37179
rect 40451 37145 40460 37179
rect 40408 37136 40460 37145
rect 40500 37136 40552 37188
rect 40684 37068 40736 37120
rect 41880 37111 41932 37120
rect 41880 37077 41889 37111
rect 41889 37077 41923 37111
rect 41923 37077 41932 37111
rect 41880 37068 41932 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 1676 36864 1728 36916
rect 2872 36864 2924 36916
rect 4620 36864 4672 36916
rect 5172 36907 5224 36916
rect 5172 36873 5181 36907
rect 5181 36873 5215 36907
rect 5215 36873 5224 36907
rect 5172 36864 5224 36873
rect 5356 36907 5408 36916
rect 5356 36873 5365 36907
rect 5365 36873 5399 36907
rect 5399 36873 5408 36907
rect 5356 36864 5408 36873
rect 6920 36864 6972 36916
rect 8116 36864 8168 36916
rect 2872 36771 2924 36780
rect 2872 36737 2881 36771
rect 2881 36737 2915 36771
rect 2915 36737 2924 36771
rect 2872 36728 2924 36737
rect 3148 36771 3200 36780
rect 3148 36737 3157 36771
rect 3157 36737 3191 36771
rect 3191 36737 3200 36771
rect 3148 36728 3200 36737
rect 3792 36796 3844 36848
rect 6644 36796 6696 36848
rect 12532 36864 12584 36916
rect 14188 36864 14240 36916
rect 3516 36728 3568 36780
rect 4436 36771 4488 36780
rect 4436 36737 4445 36771
rect 4445 36737 4479 36771
rect 4479 36737 4488 36771
rect 4436 36728 4488 36737
rect 4528 36771 4580 36780
rect 4528 36737 4537 36771
rect 4537 36737 4571 36771
rect 4571 36737 4580 36771
rect 4528 36728 4580 36737
rect 3240 36660 3292 36712
rect 3332 36660 3384 36712
rect 4344 36660 4396 36712
rect 4988 36728 5040 36780
rect 4804 36592 4856 36644
rect 4068 36524 4120 36576
rect 6552 36771 6604 36780
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 6828 36703 6880 36712
rect 6828 36669 6837 36703
rect 6837 36669 6871 36703
rect 6871 36669 6880 36703
rect 6828 36660 6880 36669
rect 7196 36660 7248 36712
rect 7472 36660 7524 36712
rect 13176 36839 13228 36848
rect 13176 36805 13185 36839
rect 13185 36805 13219 36839
rect 13219 36805 13228 36839
rect 13176 36796 13228 36805
rect 15384 36864 15436 36916
rect 16856 36864 16908 36916
rect 17316 36864 17368 36916
rect 17592 36864 17644 36916
rect 15108 36796 15160 36848
rect 10048 36660 10100 36712
rect 5632 36524 5684 36576
rect 7104 36524 7156 36576
rect 9864 36524 9916 36576
rect 10508 36524 10560 36576
rect 11980 36728 12032 36780
rect 12624 36771 12676 36780
rect 12624 36737 12633 36771
rect 12633 36737 12667 36771
rect 12667 36737 12676 36771
rect 12624 36728 12676 36737
rect 17408 36728 17460 36780
rect 17684 36771 17736 36780
rect 17684 36737 17693 36771
rect 17693 36737 17727 36771
rect 17727 36737 17736 36771
rect 17684 36728 17736 36737
rect 11336 36703 11388 36712
rect 11336 36669 11345 36703
rect 11345 36669 11379 36703
rect 11379 36669 11388 36703
rect 11336 36660 11388 36669
rect 12072 36703 12124 36712
rect 12072 36669 12081 36703
rect 12081 36669 12115 36703
rect 12115 36669 12124 36703
rect 12072 36660 12124 36669
rect 12900 36703 12952 36712
rect 12900 36669 12909 36703
rect 12909 36669 12943 36703
rect 12943 36669 12952 36703
rect 14740 36703 14792 36712
rect 12900 36660 12952 36669
rect 14740 36669 14749 36703
rect 14749 36669 14783 36703
rect 14783 36669 14792 36703
rect 14740 36660 14792 36669
rect 15752 36660 15804 36712
rect 16304 36660 16356 36712
rect 11612 36592 11664 36644
rect 16212 36592 16264 36644
rect 17868 36703 17920 36712
rect 17868 36669 17877 36703
rect 17877 36669 17911 36703
rect 17911 36669 17920 36703
rect 17868 36660 17920 36669
rect 19248 36864 19300 36916
rect 19892 36907 19944 36916
rect 19892 36873 19901 36907
rect 19901 36873 19935 36907
rect 19935 36873 19944 36907
rect 19892 36864 19944 36873
rect 22744 36864 22796 36916
rect 23572 36864 23624 36916
rect 25044 36864 25096 36916
rect 26516 36864 26568 36916
rect 27896 36907 27948 36916
rect 27896 36873 27905 36907
rect 27905 36873 27939 36907
rect 27939 36873 27948 36907
rect 27896 36864 27948 36873
rect 18144 36771 18196 36780
rect 18144 36737 18153 36771
rect 18153 36737 18187 36771
rect 18187 36737 18196 36771
rect 18144 36728 18196 36737
rect 21548 36796 21600 36848
rect 22652 36796 22704 36848
rect 23204 36796 23256 36848
rect 24400 36796 24452 36848
rect 26056 36796 26108 36848
rect 28080 36796 28132 36848
rect 21916 36771 21968 36780
rect 21916 36737 21925 36771
rect 21925 36737 21959 36771
rect 21959 36737 21968 36771
rect 21916 36728 21968 36737
rect 22468 36728 22520 36780
rect 24492 36728 24544 36780
rect 26332 36771 26384 36780
rect 26332 36737 26341 36771
rect 26341 36737 26375 36771
rect 26375 36737 26384 36771
rect 26332 36728 26384 36737
rect 27620 36728 27672 36780
rect 27712 36728 27764 36780
rect 28908 36728 28960 36780
rect 29184 36728 29236 36780
rect 31300 36864 31352 36916
rect 31392 36864 31444 36916
rect 30472 36839 30524 36848
rect 30472 36805 30481 36839
rect 30481 36805 30515 36839
rect 30515 36805 30524 36839
rect 30472 36796 30524 36805
rect 31944 36907 31996 36916
rect 31944 36873 31953 36907
rect 31953 36873 31987 36907
rect 31987 36873 31996 36907
rect 31944 36864 31996 36873
rect 32312 36796 32364 36848
rect 32496 36796 32548 36848
rect 36912 36907 36964 36916
rect 36912 36873 36921 36907
rect 36921 36873 36955 36907
rect 36955 36873 36964 36907
rect 36912 36864 36964 36873
rect 37648 36864 37700 36916
rect 38476 36864 38528 36916
rect 39948 36864 40000 36916
rect 40776 36864 40828 36916
rect 41328 36864 41380 36916
rect 31576 36728 31628 36780
rect 20076 36660 20128 36712
rect 11060 36524 11112 36576
rect 12256 36567 12308 36576
rect 12256 36533 12265 36567
rect 12265 36533 12299 36567
rect 12299 36533 12308 36567
rect 12256 36524 12308 36533
rect 16672 36567 16724 36576
rect 16672 36533 16681 36567
rect 16681 36533 16715 36567
rect 16715 36533 16724 36567
rect 16672 36524 16724 36533
rect 18052 36592 18104 36644
rect 19524 36592 19576 36644
rect 23112 36703 23164 36712
rect 23112 36669 23121 36703
rect 23121 36669 23155 36703
rect 23155 36669 23164 36703
rect 23112 36660 23164 36669
rect 25596 36660 25648 36712
rect 27344 36660 27396 36712
rect 29736 36660 29788 36712
rect 23480 36592 23532 36644
rect 25780 36592 25832 36644
rect 34336 36771 34388 36780
rect 34336 36737 34345 36771
rect 34345 36737 34379 36771
rect 34379 36737 34388 36771
rect 34336 36728 34388 36737
rect 34428 36728 34480 36780
rect 35716 36728 35768 36780
rect 36268 36728 36320 36780
rect 36544 36728 36596 36780
rect 36820 36771 36872 36780
rect 36820 36737 36829 36771
rect 36829 36737 36863 36771
rect 36863 36737 36872 36771
rect 36820 36728 36872 36737
rect 36912 36660 36964 36712
rect 37004 36660 37056 36712
rect 38200 36728 38252 36780
rect 38292 36771 38344 36780
rect 38292 36737 38301 36771
rect 38301 36737 38335 36771
rect 38335 36737 38344 36771
rect 38292 36728 38344 36737
rect 38936 36728 38988 36780
rect 39120 36771 39172 36780
rect 39120 36737 39129 36771
rect 39129 36737 39163 36771
rect 39163 36737 39172 36771
rect 39120 36728 39172 36737
rect 40500 36728 40552 36780
rect 19156 36524 19208 36576
rect 19616 36524 19668 36576
rect 19984 36567 20036 36576
rect 19984 36533 19993 36567
rect 19993 36533 20027 36567
rect 20027 36533 20036 36567
rect 19984 36524 20036 36533
rect 29092 36567 29144 36576
rect 29092 36533 29101 36567
rect 29101 36533 29135 36567
rect 29135 36533 29144 36567
rect 29092 36524 29144 36533
rect 34152 36635 34204 36644
rect 34152 36601 34161 36635
rect 34161 36601 34195 36635
rect 34195 36601 34204 36635
rect 34152 36592 34204 36601
rect 34520 36635 34572 36644
rect 34520 36601 34529 36635
rect 34529 36601 34563 36635
rect 34563 36601 34572 36635
rect 34520 36592 34572 36601
rect 35992 36592 36044 36644
rect 36544 36592 36596 36644
rect 31576 36524 31628 36576
rect 34336 36524 34388 36576
rect 35624 36524 35676 36576
rect 39212 36660 39264 36712
rect 39396 36592 39448 36644
rect 39856 36592 39908 36644
rect 38200 36524 38252 36576
rect 38936 36524 38988 36576
rect 39028 36524 39080 36576
rect 41512 36660 41564 36712
rect 41604 36703 41656 36712
rect 41604 36669 41613 36703
rect 41613 36669 41647 36703
rect 41647 36669 41656 36703
rect 41604 36660 41656 36669
rect 40040 36567 40092 36576
rect 40040 36533 40049 36567
rect 40049 36533 40083 36567
rect 40083 36533 40092 36567
rect 40040 36524 40092 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4988 36320 5040 36372
rect 5448 36320 5500 36372
rect 7196 36320 7248 36372
rect 11336 36363 11388 36372
rect 11336 36329 11345 36363
rect 11345 36329 11379 36363
rect 11379 36329 11388 36363
rect 11336 36320 11388 36329
rect 13176 36320 13228 36372
rect 15752 36363 15804 36372
rect 15752 36329 15761 36363
rect 15761 36329 15795 36363
rect 15795 36329 15804 36363
rect 15752 36320 15804 36329
rect 2872 36116 2924 36168
rect 2964 36159 3016 36168
rect 2964 36125 2973 36159
rect 2973 36125 3007 36159
rect 3007 36125 3016 36159
rect 2964 36116 3016 36125
rect 3792 36184 3844 36236
rect 3976 36252 4028 36304
rect 6552 36252 6604 36304
rect 7012 36252 7064 36304
rect 8024 36252 8076 36304
rect 6092 36184 6144 36236
rect 3884 36159 3936 36168
rect 3884 36125 3893 36159
rect 3893 36125 3927 36159
rect 3927 36125 3936 36159
rect 3884 36116 3936 36125
rect 4068 36116 4120 36168
rect 5172 36116 5224 36168
rect 7104 36159 7156 36168
rect 7104 36125 7113 36159
rect 7113 36125 7147 36159
rect 7147 36125 7156 36159
rect 7104 36116 7156 36125
rect 7380 36184 7432 36236
rect 8116 36184 8168 36236
rect 12348 36252 12400 36304
rect 21916 36320 21968 36372
rect 9864 36227 9916 36236
rect 9864 36193 9873 36227
rect 9873 36193 9907 36227
rect 9907 36193 9916 36227
rect 9864 36184 9916 36193
rect 10508 36184 10560 36236
rect 9588 36159 9640 36168
rect 9588 36125 9597 36159
rect 9597 36125 9631 36159
rect 9631 36125 9640 36159
rect 9588 36116 9640 36125
rect 12256 36227 12308 36236
rect 12256 36193 12265 36227
rect 12265 36193 12299 36227
rect 12299 36193 12308 36227
rect 12256 36184 12308 36193
rect 14556 36227 14608 36236
rect 14556 36193 14565 36227
rect 14565 36193 14599 36227
rect 14599 36193 14608 36227
rect 14556 36184 14608 36193
rect 13268 36116 13320 36168
rect 13820 36159 13872 36168
rect 13820 36125 13829 36159
rect 13829 36125 13863 36159
rect 13863 36125 13872 36159
rect 13820 36116 13872 36125
rect 14280 36116 14332 36168
rect 16304 36184 16356 36236
rect 2872 35980 2924 36032
rect 3516 36048 3568 36100
rect 3700 36048 3752 36100
rect 6368 36048 6420 36100
rect 4068 35980 4120 36032
rect 5356 35980 5408 36032
rect 7564 36048 7616 36100
rect 9772 36048 9824 36100
rect 12624 36048 12676 36100
rect 16672 36116 16724 36168
rect 16856 36184 16908 36236
rect 17500 36184 17552 36236
rect 19708 36184 19760 36236
rect 19892 36184 19944 36236
rect 22192 36227 22244 36236
rect 22192 36193 22201 36227
rect 22201 36193 22235 36227
rect 22235 36193 22244 36227
rect 22192 36184 22244 36193
rect 19984 36116 20036 36168
rect 25136 36252 25188 36304
rect 23940 36227 23992 36236
rect 23940 36193 23949 36227
rect 23949 36193 23983 36227
rect 23983 36193 23992 36227
rect 23940 36184 23992 36193
rect 29184 36320 29236 36372
rect 29552 36363 29604 36372
rect 29552 36329 29561 36363
rect 29561 36329 29595 36363
rect 29595 36329 29604 36363
rect 29552 36320 29604 36329
rect 34336 36320 34388 36372
rect 27344 36252 27396 36304
rect 31300 36227 31352 36236
rect 31300 36193 31309 36227
rect 31309 36193 31343 36227
rect 31343 36193 31352 36227
rect 31300 36184 31352 36193
rect 31484 36184 31536 36236
rect 31944 36227 31996 36236
rect 31944 36193 31953 36227
rect 31953 36193 31987 36227
rect 31987 36193 31996 36227
rect 31944 36184 31996 36193
rect 35716 36184 35768 36236
rect 11704 36023 11756 36032
rect 11704 35989 11713 36023
rect 11713 35989 11747 36023
rect 11747 35989 11756 36023
rect 11704 35980 11756 35989
rect 13084 35980 13136 36032
rect 15660 36048 15712 36100
rect 14464 36023 14516 36032
rect 14464 35989 14473 36023
rect 14473 35989 14507 36023
rect 14507 35989 14516 36023
rect 14464 35980 14516 35989
rect 15292 35980 15344 36032
rect 16856 36048 16908 36100
rect 20904 36048 20956 36100
rect 21640 36048 21692 36100
rect 22468 36091 22520 36100
rect 22468 36057 22477 36091
rect 22477 36057 22511 36091
rect 22511 36057 22520 36091
rect 22468 36048 22520 36057
rect 27436 36116 27488 36168
rect 32772 36159 32824 36168
rect 32772 36125 32781 36159
rect 32781 36125 32815 36159
rect 32815 36125 32824 36159
rect 32772 36116 32824 36125
rect 16948 36023 17000 36032
rect 16948 35989 16957 36023
rect 16957 35989 16991 36023
rect 16991 35989 17000 36023
rect 16948 35980 17000 35989
rect 17040 36023 17092 36032
rect 17040 35989 17049 36023
rect 17049 35989 17083 36023
rect 17083 35989 17092 36023
rect 17040 35980 17092 35989
rect 18236 35980 18288 36032
rect 19708 36023 19760 36032
rect 19708 35989 19717 36023
rect 19717 35989 19751 36023
rect 19751 35989 19760 36023
rect 19708 35980 19760 35989
rect 22560 35980 22612 36032
rect 27068 36048 27120 36100
rect 27896 36091 27948 36100
rect 27896 36057 27905 36091
rect 27905 36057 27939 36091
rect 27939 36057 27948 36091
rect 27896 36048 27948 36057
rect 29276 36048 29328 36100
rect 29736 36048 29788 36100
rect 31024 36091 31076 36100
rect 31024 36057 31033 36091
rect 31033 36057 31067 36091
rect 31067 36057 31076 36091
rect 31024 36048 31076 36057
rect 34060 36048 34112 36100
rect 24032 35980 24084 36032
rect 24584 35980 24636 36032
rect 27528 36023 27580 36032
rect 27528 35989 27537 36023
rect 27537 35989 27571 36023
rect 27571 35989 27580 36023
rect 27528 35980 27580 35989
rect 27712 35980 27764 36032
rect 30748 35980 30800 36032
rect 32680 35980 32732 36032
rect 33416 36023 33468 36032
rect 33416 35989 33425 36023
rect 33425 35989 33459 36023
rect 33459 35989 33468 36023
rect 33416 35980 33468 35989
rect 33784 36023 33836 36032
rect 33784 35989 33793 36023
rect 33793 35989 33827 36023
rect 33827 35989 33836 36023
rect 33784 35980 33836 35989
rect 34244 36023 34296 36032
rect 34244 35989 34253 36023
rect 34253 35989 34287 36023
rect 34287 35989 34296 36023
rect 34244 35980 34296 35989
rect 34428 35980 34480 36032
rect 35440 36116 35492 36168
rect 36820 36363 36872 36372
rect 36820 36329 36829 36363
rect 36829 36329 36863 36363
rect 36863 36329 36872 36363
rect 36820 36320 36872 36329
rect 38292 36320 38344 36372
rect 39120 36320 39172 36372
rect 41604 36320 41656 36372
rect 36452 36184 36504 36236
rect 38108 36184 38160 36236
rect 35624 36091 35676 36100
rect 35624 36057 35633 36091
rect 35633 36057 35667 36091
rect 35667 36057 35676 36091
rect 36912 36159 36964 36168
rect 36912 36125 36921 36159
rect 36921 36125 36955 36159
rect 36955 36125 36964 36159
rect 36912 36116 36964 36125
rect 37372 36159 37424 36168
rect 37372 36125 37381 36159
rect 37381 36125 37415 36159
rect 37415 36125 37424 36159
rect 37372 36116 37424 36125
rect 38752 36116 38804 36168
rect 39028 36116 39080 36168
rect 35624 36048 35676 36057
rect 36452 36048 36504 36100
rect 37648 36091 37700 36100
rect 37648 36057 37657 36091
rect 37657 36057 37691 36091
rect 37691 36057 37700 36091
rect 37648 36048 37700 36057
rect 40132 36227 40184 36236
rect 40132 36193 40141 36227
rect 40141 36193 40175 36227
rect 40175 36193 40184 36227
rect 40132 36184 40184 36193
rect 41328 36184 41380 36236
rect 39212 36159 39264 36168
rect 39212 36125 39221 36159
rect 39221 36125 39255 36159
rect 39255 36125 39264 36159
rect 39212 36116 39264 36125
rect 39396 36159 39448 36168
rect 39396 36125 39405 36159
rect 39405 36125 39439 36159
rect 39439 36125 39448 36159
rect 39396 36116 39448 36125
rect 40040 36048 40092 36100
rect 36084 35980 36136 36032
rect 36544 36023 36596 36032
rect 36544 35989 36553 36023
rect 36553 35989 36587 36023
rect 36587 35989 36596 36023
rect 36544 35980 36596 35989
rect 38936 35980 38988 36032
rect 39304 35980 39356 36032
rect 41236 35980 41288 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 3608 35776 3660 35828
rect 5632 35776 5684 35828
rect 6092 35819 6144 35828
rect 6092 35785 6101 35819
rect 6101 35785 6135 35819
rect 6135 35785 6144 35819
rect 6092 35776 6144 35785
rect 9680 35776 9732 35828
rect 2780 35640 2832 35692
rect 3700 35640 3752 35692
rect 3884 35640 3936 35692
rect 1400 35615 1452 35624
rect 1400 35581 1409 35615
rect 1409 35581 1443 35615
rect 1443 35581 1452 35615
rect 1400 35572 1452 35581
rect 2872 35572 2924 35624
rect 3424 35572 3476 35624
rect 3516 35572 3568 35624
rect 12072 35776 12124 35828
rect 14280 35776 14332 35828
rect 14648 35819 14700 35828
rect 14648 35785 14657 35819
rect 14657 35785 14691 35819
rect 14691 35785 14700 35819
rect 14648 35776 14700 35785
rect 16948 35819 17000 35828
rect 16948 35785 16957 35819
rect 16957 35785 16991 35819
rect 16991 35785 17000 35819
rect 16948 35776 17000 35785
rect 17132 35776 17184 35828
rect 20904 35776 20956 35828
rect 22468 35776 22520 35828
rect 24584 35776 24636 35828
rect 27528 35776 27580 35828
rect 27896 35776 27948 35828
rect 29092 35776 29144 35828
rect 29644 35776 29696 35828
rect 11704 35708 11756 35760
rect 14188 35708 14240 35760
rect 18236 35751 18288 35760
rect 18236 35717 18245 35751
rect 18245 35717 18279 35751
rect 18279 35717 18288 35751
rect 18236 35708 18288 35717
rect 19524 35708 19576 35760
rect 22836 35708 22888 35760
rect 23204 35708 23256 35760
rect 4620 35640 4672 35692
rect 5264 35683 5316 35692
rect 5264 35649 5273 35683
rect 5273 35649 5307 35683
rect 5307 35649 5316 35683
rect 5264 35640 5316 35649
rect 4896 35615 4948 35624
rect 4896 35581 4905 35615
rect 4905 35581 4939 35615
rect 4939 35581 4948 35615
rect 4896 35572 4948 35581
rect 2136 35436 2188 35488
rect 5448 35640 5500 35692
rect 5632 35615 5684 35624
rect 5632 35581 5641 35615
rect 5641 35581 5675 35615
rect 5675 35581 5684 35615
rect 5632 35572 5684 35581
rect 5908 35683 5960 35692
rect 5908 35649 5917 35683
rect 5917 35649 5951 35683
rect 5951 35649 5960 35683
rect 5908 35640 5960 35649
rect 7656 35640 7708 35692
rect 8208 35640 8260 35692
rect 6276 35572 6328 35624
rect 9496 35572 9548 35624
rect 9864 35572 9916 35624
rect 11520 35615 11572 35624
rect 11520 35581 11529 35615
rect 11529 35581 11563 35615
rect 11563 35581 11572 35615
rect 11520 35572 11572 35581
rect 14280 35640 14332 35692
rect 15200 35640 15252 35692
rect 15476 35683 15528 35692
rect 15476 35649 15485 35683
rect 15485 35649 15519 35683
rect 15519 35649 15528 35683
rect 15476 35640 15528 35649
rect 17040 35683 17092 35692
rect 17040 35649 17049 35683
rect 17049 35649 17083 35683
rect 17083 35649 17092 35683
rect 17040 35640 17092 35649
rect 14372 35572 14424 35624
rect 15108 35615 15160 35624
rect 15108 35581 15117 35615
rect 15117 35581 15151 35615
rect 15151 35581 15160 35615
rect 15108 35572 15160 35581
rect 15292 35615 15344 35624
rect 15292 35581 15301 35615
rect 15301 35581 15335 35615
rect 15335 35581 15344 35615
rect 15292 35572 15344 35581
rect 16580 35572 16632 35624
rect 16856 35615 16908 35624
rect 16856 35581 16865 35615
rect 16865 35581 16899 35615
rect 16899 35581 16908 35615
rect 16856 35572 16908 35581
rect 3976 35436 4028 35488
rect 4068 35436 4120 35488
rect 5448 35504 5500 35556
rect 7840 35436 7892 35488
rect 13268 35479 13320 35488
rect 13268 35445 13277 35479
rect 13277 35445 13311 35479
rect 13311 35445 13320 35479
rect 13268 35436 13320 35445
rect 15660 35479 15712 35488
rect 15660 35445 15669 35479
rect 15669 35445 15703 35479
rect 15703 35445 15712 35479
rect 15660 35436 15712 35445
rect 16028 35436 16080 35488
rect 17316 35572 17368 35624
rect 19892 35640 19944 35692
rect 20168 35683 20220 35692
rect 20168 35649 20177 35683
rect 20177 35649 20211 35683
rect 20211 35649 20220 35683
rect 20168 35640 20220 35649
rect 20536 35640 20588 35692
rect 20076 35572 20128 35624
rect 20444 35615 20496 35624
rect 20444 35581 20453 35615
rect 20453 35581 20487 35615
rect 20487 35581 20496 35615
rect 20444 35572 20496 35581
rect 19800 35547 19852 35556
rect 19800 35513 19809 35547
rect 19809 35513 19843 35547
rect 19843 35513 19852 35547
rect 19800 35504 19852 35513
rect 23296 35640 23348 35692
rect 25780 35708 25832 35760
rect 31208 35776 31260 35828
rect 32772 35776 32824 35828
rect 34428 35776 34480 35828
rect 37648 35776 37700 35828
rect 22284 35615 22336 35624
rect 22284 35581 22293 35615
rect 22293 35581 22327 35615
rect 22327 35581 22336 35615
rect 22284 35572 22336 35581
rect 23112 35572 23164 35624
rect 24768 35572 24820 35624
rect 26148 35572 26200 35624
rect 26976 35572 27028 35624
rect 24032 35504 24084 35556
rect 25412 35504 25464 35556
rect 27344 35504 27396 35556
rect 28724 35615 28776 35624
rect 28724 35581 28733 35615
rect 28733 35581 28767 35615
rect 28767 35581 28776 35615
rect 28724 35572 28776 35581
rect 29000 35572 29052 35624
rect 30104 35640 30156 35692
rect 30748 35708 30800 35760
rect 34060 35708 34112 35760
rect 39120 35708 39172 35760
rect 40408 35776 40460 35828
rect 40592 35819 40644 35828
rect 40592 35785 40601 35819
rect 40601 35785 40635 35819
rect 40635 35785 40644 35819
rect 40592 35776 40644 35785
rect 41144 35776 41196 35828
rect 41696 35708 41748 35760
rect 31576 35640 31628 35692
rect 33876 35640 33928 35692
rect 36912 35683 36964 35692
rect 36912 35649 36921 35683
rect 36921 35649 36955 35683
rect 36955 35649 36964 35683
rect 36912 35640 36964 35649
rect 39304 35683 39356 35692
rect 39304 35649 39313 35683
rect 39313 35649 39347 35683
rect 39347 35649 39356 35683
rect 39304 35640 39356 35649
rect 41420 35683 41472 35692
rect 41420 35649 41429 35683
rect 41429 35649 41463 35683
rect 41463 35649 41472 35683
rect 41420 35640 41472 35649
rect 30840 35572 30892 35624
rect 31208 35572 31260 35624
rect 32404 35572 32456 35624
rect 33784 35572 33836 35624
rect 34704 35572 34756 35624
rect 35440 35572 35492 35624
rect 35992 35615 36044 35624
rect 35992 35581 36001 35615
rect 36001 35581 36035 35615
rect 36035 35581 36044 35615
rect 35992 35572 36044 35581
rect 36084 35615 36136 35624
rect 36084 35581 36093 35615
rect 36093 35581 36127 35615
rect 36127 35581 36136 35615
rect 36084 35572 36136 35581
rect 36544 35572 36596 35624
rect 38476 35615 38528 35624
rect 38476 35581 38485 35615
rect 38485 35581 38519 35615
rect 38519 35581 38528 35615
rect 38476 35572 38528 35581
rect 40132 35572 40184 35624
rect 40408 35572 40460 35624
rect 41052 35572 41104 35624
rect 41512 35615 41564 35624
rect 41512 35581 41521 35615
rect 41521 35581 41555 35615
rect 41555 35581 41564 35615
rect 41512 35572 41564 35581
rect 41144 35504 41196 35556
rect 20444 35436 20496 35488
rect 26148 35436 26200 35488
rect 31024 35436 31076 35488
rect 33232 35436 33284 35488
rect 33876 35436 33928 35488
rect 35532 35479 35584 35488
rect 35532 35445 35541 35479
rect 35541 35445 35575 35479
rect 35575 35445 35584 35479
rect 35532 35436 35584 35445
rect 36360 35436 36412 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3884 35232 3936 35284
rect 5264 35232 5316 35284
rect 9864 35275 9916 35284
rect 9864 35241 9873 35275
rect 9873 35241 9907 35275
rect 9907 35241 9916 35275
rect 9864 35232 9916 35241
rect 9680 35164 9732 35216
rect 1400 35096 1452 35148
rect 2136 35139 2188 35148
rect 2136 35105 2145 35139
rect 2145 35105 2179 35139
rect 2179 35105 2188 35139
rect 2136 35096 2188 35105
rect 2688 35096 2740 35148
rect 6828 35096 6880 35148
rect 7288 35096 7340 35148
rect 9588 35096 9640 35148
rect 11520 35096 11572 35148
rect 3608 35028 3660 35080
rect 3884 35028 3936 35080
rect 10048 35071 10100 35080
rect 10048 35037 10057 35071
rect 10057 35037 10091 35071
rect 10091 35037 10100 35071
rect 10048 35028 10100 35037
rect 3700 34960 3752 35012
rect 3976 34960 4028 35012
rect 4344 35003 4396 35012
rect 4344 34969 4353 35003
rect 4353 34969 4387 35003
rect 4387 34969 4396 35003
rect 4344 34960 4396 34969
rect 4068 34892 4120 34944
rect 4712 34935 4764 34944
rect 4712 34901 4721 34935
rect 4721 34901 4755 34935
rect 4755 34901 4764 34935
rect 4712 34892 4764 34901
rect 6368 34960 6420 35012
rect 7564 34960 7616 35012
rect 9128 34960 9180 35012
rect 9680 34960 9732 35012
rect 5264 34892 5316 34944
rect 6460 34892 6512 34944
rect 8576 34892 8628 34944
rect 10508 35071 10560 35080
rect 10508 35037 10517 35071
rect 10517 35037 10551 35071
rect 10551 35037 10560 35071
rect 10508 35028 10560 35037
rect 12256 35232 12308 35284
rect 15476 35232 15528 35284
rect 16580 35232 16632 35284
rect 16948 35232 17000 35284
rect 17868 35232 17920 35284
rect 14004 35164 14056 35216
rect 15292 35139 15344 35148
rect 15292 35105 15301 35139
rect 15301 35105 15335 35139
rect 15335 35105 15344 35139
rect 15292 35096 15344 35105
rect 19708 35232 19760 35284
rect 22284 35232 22336 35284
rect 23296 35232 23348 35284
rect 24768 35275 24820 35284
rect 24768 35241 24777 35275
rect 24777 35241 24811 35275
rect 24811 35241 24820 35275
rect 24768 35232 24820 35241
rect 27712 35232 27764 35284
rect 31668 35232 31720 35284
rect 36912 35232 36964 35284
rect 40408 35275 40460 35284
rect 40408 35241 40417 35275
rect 40417 35241 40451 35275
rect 40451 35241 40460 35275
rect 40408 35232 40460 35241
rect 41236 35275 41288 35284
rect 41236 35241 41245 35275
rect 41245 35241 41279 35275
rect 41279 35241 41288 35275
rect 41236 35232 41288 35241
rect 20444 35164 20496 35216
rect 20168 35096 20220 35148
rect 22376 35207 22428 35216
rect 22376 35173 22385 35207
rect 22385 35173 22419 35207
rect 22419 35173 22428 35207
rect 22376 35164 22428 35173
rect 36452 35164 36504 35216
rect 23388 35096 23440 35148
rect 13544 35071 13596 35080
rect 13544 35037 13553 35071
rect 13553 35037 13587 35071
rect 13587 35037 13596 35071
rect 13544 35028 13596 35037
rect 14004 35028 14056 35080
rect 14280 35071 14332 35080
rect 14280 35037 14289 35071
rect 14289 35037 14323 35071
rect 14323 35037 14332 35071
rect 14280 35028 14332 35037
rect 15108 35028 15160 35080
rect 15660 35028 15712 35080
rect 10968 34960 11020 35012
rect 16488 34960 16540 35012
rect 17316 35071 17368 35080
rect 17316 35037 17325 35071
rect 17325 35037 17359 35071
rect 17359 35037 17368 35071
rect 17316 35028 17368 35037
rect 24032 35096 24084 35148
rect 25596 35096 25648 35148
rect 27436 35096 27488 35148
rect 29000 35096 29052 35148
rect 25412 35028 25464 35080
rect 29276 35096 29328 35148
rect 31944 35139 31996 35148
rect 31944 35105 31953 35139
rect 31953 35105 31987 35139
rect 31987 35105 31996 35139
rect 31944 35096 31996 35105
rect 34796 35096 34848 35148
rect 37280 35096 37332 35148
rect 38476 35139 38528 35148
rect 38476 35105 38485 35139
rect 38485 35105 38519 35139
rect 38519 35105 38528 35139
rect 38476 35096 38528 35105
rect 39212 35096 39264 35148
rect 40040 35096 40092 35148
rect 41144 35096 41196 35148
rect 29184 35028 29236 35080
rect 36360 35028 36412 35080
rect 22284 34960 22336 35012
rect 23204 34960 23256 35012
rect 26148 35003 26200 35012
rect 26148 34969 26157 35003
rect 26157 34969 26191 35003
rect 26191 34969 26200 35003
rect 26148 34960 26200 34969
rect 32220 35003 32272 35012
rect 32220 34969 32229 35003
rect 32229 34969 32263 35003
rect 32263 34969 32272 35003
rect 32220 34960 32272 34969
rect 35532 34960 35584 35012
rect 11060 34892 11112 34944
rect 13912 34935 13964 34944
rect 13912 34901 13921 34935
rect 13921 34901 13955 34935
rect 13955 34901 13964 34935
rect 13912 34892 13964 34901
rect 15200 34892 15252 34944
rect 15660 34892 15712 34944
rect 17592 34892 17644 34944
rect 20536 34892 20588 34944
rect 20628 34892 20680 34944
rect 22744 34892 22796 34944
rect 23848 34935 23900 34944
rect 23848 34901 23857 34935
rect 23857 34901 23891 34935
rect 23891 34901 23900 34935
rect 23848 34892 23900 34901
rect 23940 34935 23992 34944
rect 23940 34901 23949 34935
rect 23949 34901 23983 34935
rect 23983 34901 23992 34935
rect 23940 34892 23992 34901
rect 25228 34935 25280 34944
rect 25228 34901 25237 34935
rect 25237 34901 25271 34935
rect 25271 34901 25280 34935
rect 25228 34892 25280 34901
rect 27712 34892 27764 34944
rect 29460 34892 29512 34944
rect 31760 34935 31812 34944
rect 31760 34901 31769 34935
rect 31769 34901 31803 34935
rect 31803 34901 31812 34935
rect 31760 34892 31812 34901
rect 32036 34892 32088 34944
rect 32128 34892 32180 34944
rect 33048 34892 33100 34944
rect 38108 34960 38160 35012
rect 38936 34960 38988 35012
rect 40776 35003 40828 35012
rect 40776 34969 40785 35003
rect 40785 34969 40819 35003
rect 40819 34969 40828 35003
rect 40776 34960 40828 34969
rect 36820 34935 36872 34944
rect 36820 34901 36829 34935
rect 36829 34901 36863 34935
rect 36863 34901 36872 34935
rect 36820 34892 36872 34901
rect 37924 34935 37976 34944
rect 37924 34901 37933 34935
rect 37933 34901 37967 34935
rect 37967 34901 37976 34935
rect 37924 34892 37976 34901
rect 38384 34935 38436 34944
rect 38384 34901 38393 34935
rect 38393 34901 38427 34935
rect 38427 34901 38436 34935
rect 38384 34892 38436 34901
rect 40040 34935 40092 34944
rect 40040 34901 40049 34935
rect 40049 34901 40083 34935
rect 40083 34901 40092 34935
rect 40040 34892 40092 34901
rect 41236 34892 41288 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 2964 34688 3016 34740
rect 4620 34688 4672 34740
rect 5540 34688 5592 34740
rect 3976 34620 4028 34672
rect 3608 34595 3660 34604
rect 3608 34561 3617 34595
rect 3617 34561 3651 34595
rect 3651 34561 3660 34595
rect 3608 34552 3660 34561
rect 4068 34552 4120 34604
rect 4712 34552 4764 34604
rect 5632 34620 5684 34672
rect 6184 34620 6236 34672
rect 6644 34663 6696 34672
rect 6644 34629 6653 34663
rect 6653 34629 6687 34663
rect 6687 34629 6696 34663
rect 6644 34620 6696 34629
rect 8208 34620 8260 34672
rect 9404 34620 9456 34672
rect 10968 34663 11020 34672
rect 10968 34629 10977 34663
rect 10977 34629 11011 34663
rect 11011 34629 11020 34663
rect 10968 34620 11020 34629
rect 11612 34688 11664 34740
rect 14464 34688 14516 34740
rect 16028 34731 16080 34740
rect 16028 34697 16037 34731
rect 16037 34697 16071 34731
rect 16071 34697 16080 34731
rect 16028 34688 16080 34697
rect 16488 34731 16540 34740
rect 16488 34697 16497 34731
rect 16497 34697 16531 34731
rect 16531 34697 16540 34731
rect 16488 34688 16540 34697
rect 12164 34620 12216 34672
rect 12624 34620 12676 34672
rect 5172 34552 5224 34604
rect 6092 34552 6144 34604
rect 6276 34552 6328 34604
rect 7288 34484 7340 34536
rect 7564 34484 7616 34536
rect 7840 34595 7892 34604
rect 7840 34561 7849 34595
rect 7849 34561 7883 34595
rect 7883 34561 7892 34595
rect 7840 34552 7892 34561
rect 7932 34595 7984 34604
rect 7932 34561 7941 34595
rect 7941 34561 7975 34595
rect 7975 34561 7984 34595
rect 7932 34552 7984 34561
rect 10048 34552 10100 34604
rect 10324 34552 10376 34604
rect 11060 34552 11112 34604
rect 12900 34595 12952 34604
rect 12900 34561 12909 34595
rect 12909 34561 12943 34595
rect 12943 34561 12952 34595
rect 12900 34552 12952 34561
rect 15568 34620 15620 34672
rect 14924 34552 14976 34604
rect 17316 34620 17368 34672
rect 17868 34688 17920 34740
rect 20076 34731 20128 34740
rect 20076 34697 20085 34731
rect 20085 34697 20119 34731
rect 20119 34697 20128 34731
rect 20076 34688 20128 34697
rect 18236 34620 18288 34672
rect 20628 34731 20680 34740
rect 20628 34697 20637 34731
rect 20637 34697 20671 34731
rect 20671 34697 20680 34731
rect 20628 34688 20680 34697
rect 23480 34731 23532 34740
rect 23480 34697 23489 34731
rect 23489 34697 23523 34731
rect 23523 34697 23532 34731
rect 23480 34688 23532 34697
rect 23940 34688 23992 34740
rect 25228 34731 25280 34740
rect 25228 34697 25237 34731
rect 25237 34697 25271 34731
rect 25271 34697 25280 34731
rect 25228 34688 25280 34697
rect 26056 34731 26108 34740
rect 26056 34697 26065 34731
rect 26065 34697 26099 34731
rect 26099 34697 26108 34731
rect 26056 34688 26108 34697
rect 29184 34731 29236 34740
rect 29184 34697 29193 34731
rect 29193 34697 29227 34731
rect 29227 34697 29236 34731
rect 29184 34688 29236 34697
rect 30012 34731 30064 34740
rect 30012 34697 30021 34731
rect 30021 34697 30055 34731
rect 30055 34697 30064 34731
rect 30012 34688 30064 34697
rect 23296 34620 23348 34672
rect 16948 34595 17000 34604
rect 16948 34561 16982 34595
rect 16982 34561 17000 34595
rect 16948 34552 17000 34561
rect 20444 34552 20496 34604
rect 23204 34595 23256 34604
rect 23204 34561 23213 34595
rect 23213 34561 23247 34595
rect 23247 34561 23256 34595
rect 23204 34552 23256 34561
rect 26148 34620 26200 34672
rect 27712 34663 27764 34672
rect 27712 34629 27721 34663
rect 27721 34629 27755 34663
rect 27755 34629 27764 34663
rect 27712 34620 27764 34629
rect 29276 34620 29328 34672
rect 29184 34552 29236 34604
rect 30932 34620 30984 34672
rect 32680 34663 32732 34672
rect 32680 34629 32689 34663
rect 32689 34629 32723 34663
rect 32723 34629 32732 34663
rect 32680 34620 32732 34629
rect 34704 34688 34756 34740
rect 38936 34688 38988 34740
rect 39212 34688 39264 34740
rect 40776 34731 40828 34740
rect 40776 34697 40785 34731
rect 40785 34697 40819 34731
rect 40819 34697 40828 34731
rect 40776 34688 40828 34697
rect 40960 34731 41012 34740
rect 40960 34697 40969 34731
rect 40969 34697 41003 34731
rect 41003 34697 41012 34731
rect 40960 34688 41012 34697
rect 41328 34688 41380 34740
rect 41420 34731 41472 34740
rect 41420 34697 41429 34731
rect 41429 34697 41463 34731
rect 41463 34697 41472 34731
rect 41420 34688 41472 34697
rect 31576 34552 31628 34604
rect 32404 34595 32456 34604
rect 32404 34561 32413 34595
rect 32413 34561 32447 34595
rect 32447 34561 32456 34595
rect 32404 34552 32456 34561
rect 6460 34416 6512 34468
rect 7748 34416 7800 34468
rect 12992 34527 13044 34536
rect 12992 34493 13001 34527
rect 13001 34493 13035 34527
rect 13035 34493 13044 34527
rect 12992 34484 13044 34493
rect 13176 34527 13228 34536
rect 13176 34493 13185 34527
rect 13185 34493 13219 34527
rect 13219 34493 13228 34527
rect 13176 34484 13228 34493
rect 14004 34484 14056 34536
rect 15476 34484 15528 34536
rect 22376 34527 22428 34536
rect 22376 34493 22385 34527
rect 22385 34493 22419 34527
rect 22419 34493 22428 34527
rect 22376 34484 22428 34493
rect 23848 34484 23900 34536
rect 24032 34527 24084 34536
rect 24032 34493 24041 34527
rect 24041 34493 24075 34527
rect 24075 34493 24084 34527
rect 24032 34484 24084 34493
rect 25688 34527 25740 34536
rect 25688 34493 25697 34527
rect 25697 34493 25731 34527
rect 25731 34493 25740 34527
rect 25688 34484 25740 34493
rect 23388 34416 23440 34468
rect 27436 34527 27488 34536
rect 27436 34493 27445 34527
rect 27445 34493 27479 34527
rect 27479 34493 27488 34527
rect 27436 34484 27488 34493
rect 34796 34595 34848 34604
rect 34796 34561 34805 34595
rect 34805 34561 34839 34595
rect 34839 34561 34848 34595
rect 34796 34552 34848 34561
rect 30196 34416 30248 34468
rect 33876 34484 33928 34536
rect 36360 34620 36412 34672
rect 37924 34620 37976 34672
rect 38752 34552 38804 34604
rect 41512 34620 41564 34672
rect 39948 34552 40000 34604
rect 40408 34552 40460 34604
rect 41972 34552 42024 34604
rect 36452 34484 36504 34536
rect 37372 34527 37424 34536
rect 37372 34493 37381 34527
rect 37381 34493 37415 34527
rect 37415 34493 37424 34527
rect 37372 34484 37424 34493
rect 41144 34484 41196 34536
rect 31944 34416 31996 34468
rect 32128 34416 32180 34468
rect 5908 34348 5960 34400
rect 6368 34348 6420 34400
rect 8116 34348 8168 34400
rect 8392 34391 8444 34400
rect 8392 34357 8401 34391
rect 8401 34357 8435 34391
rect 8435 34357 8444 34391
rect 8392 34348 8444 34357
rect 8576 34391 8628 34400
rect 8576 34357 8585 34391
rect 8585 34357 8619 34391
rect 8619 34357 8628 34391
rect 8576 34348 8628 34357
rect 15660 34348 15712 34400
rect 16028 34348 16080 34400
rect 21180 34348 21232 34400
rect 24308 34391 24360 34400
rect 24308 34357 24317 34391
rect 24317 34357 24351 34391
rect 24351 34357 24360 34391
rect 24308 34348 24360 34357
rect 30840 34391 30892 34400
rect 30840 34357 30849 34391
rect 30849 34357 30883 34391
rect 30883 34357 30892 34391
rect 30840 34348 30892 34357
rect 34796 34348 34848 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 5264 34187 5316 34196
rect 5264 34153 5273 34187
rect 5273 34153 5307 34187
rect 5307 34153 5316 34187
rect 5264 34144 5316 34153
rect 7932 34144 7984 34196
rect 8116 34187 8168 34196
rect 8116 34153 8125 34187
rect 8125 34153 8159 34187
rect 8159 34153 8168 34187
rect 8116 34144 8168 34153
rect 12992 34144 13044 34196
rect 14280 34144 14332 34196
rect 14924 34187 14976 34196
rect 14924 34153 14933 34187
rect 14933 34153 14967 34187
rect 14967 34153 14976 34187
rect 14924 34144 14976 34153
rect 17868 34144 17920 34196
rect 5724 34008 5776 34060
rect 5816 34051 5868 34060
rect 5816 34017 5825 34051
rect 5825 34017 5859 34051
rect 5859 34017 5868 34051
rect 5816 34008 5868 34017
rect 5908 34051 5960 34060
rect 5908 34017 5917 34051
rect 5917 34017 5951 34051
rect 5951 34017 5960 34051
rect 5908 34008 5960 34017
rect 5540 33983 5592 33992
rect 5540 33949 5549 33983
rect 5549 33949 5583 33983
rect 5583 33949 5592 33983
rect 5540 33940 5592 33949
rect 6644 34076 6696 34128
rect 6460 33983 6512 33992
rect 6460 33949 6469 33983
rect 6469 33949 6503 33983
rect 6503 33949 6512 33983
rect 6460 33940 6512 33949
rect 7288 33983 7340 33992
rect 7288 33949 7297 33983
rect 7297 33949 7331 33983
rect 7331 33949 7340 33983
rect 7288 33940 7340 33949
rect 7380 33940 7432 33992
rect 7656 34008 7708 34060
rect 7748 33983 7800 33992
rect 6368 33872 6420 33924
rect 6920 33872 6972 33924
rect 7748 33949 7757 33983
rect 7757 33949 7791 33983
rect 7791 33949 7800 33983
rect 7748 33940 7800 33949
rect 7840 33983 7892 33992
rect 7840 33949 7849 33983
rect 7849 33949 7883 33983
rect 7883 33949 7892 33983
rect 7840 33940 7892 33949
rect 8024 33940 8076 33992
rect 8576 33983 8628 33992
rect 8576 33949 8585 33983
rect 8585 33949 8619 33983
rect 8619 33949 8628 33983
rect 8576 33940 8628 33949
rect 9404 33940 9456 33992
rect 11612 34008 11664 34060
rect 12624 34008 12676 34060
rect 17960 34076 18012 34128
rect 13912 34008 13964 34060
rect 15476 34051 15528 34060
rect 15476 34017 15485 34051
rect 15485 34017 15519 34051
rect 15519 34017 15528 34051
rect 15476 34008 15528 34017
rect 22284 34187 22336 34196
rect 22284 34153 22293 34187
rect 22293 34153 22327 34187
rect 22327 34153 22336 34187
rect 22284 34144 22336 34153
rect 23940 34144 23992 34196
rect 6092 33804 6144 33856
rect 7932 33872 7984 33924
rect 13820 33983 13872 33992
rect 13820 33949 13829 33983
rect 13829 33949 13863 33983
rect 13863 33949 13872 33983
rect 13820 33940 13872 33949
rect 15108 33940 15160 33992
rect 16028 33940 16080 33992
rect 17316 33940 17368 33992
rect 17868 33940 17920 33992
rect 18512 33983 18564 33992
rect 18512 33949 18521 33983
rect 18521 33949 18555 33983
rect 18555 33949 18564 33983
rect 18512 33940 18564 33949
rect 22836 34051 22888 34060
rect 22836 34017 22845 34051
rect 22845 34017 22879 34051
rect 22879 34017 22888 34051
rect 22836 34008 22888 34017
rect 27436 34144 27488 34196
rect 27620 34144 27672 34196
rect 28724 34144 28776 34196
rect 29460 34144 29512 34196
rect 31484 34187 31536 34196
rect 31484 34153 31493 34187
rect 31493 34153 31527 34187
rect 31527 34153 31536 34187
rect 31484 34144 31536 34153
rect 34244 34144 34296 34196
rect 34796 34144 34848 34196
rect 35992 34144 36044 34196
rect 38384 34144 38436 34196
rect 25688 34076 25740 34128
rect 26976 34119 27028 34128
rect 26976 34085 26985 34119
rect 26985 34085 27019 34119
rect 27019 34085 27028 34119
rect 26976 34076 27028 34085
rect 21180 33983 21232 33992
rect 8484 33804 8536 33856
rect 11152 33804 11204 33856
rect 15292 33847 15344 33856
rect 15292 33813 15301 33847
rect 15301 33813 15335 33847
rect 15335 33813 15344 33847
rect 15292 33804 15344 33813
rect 21180 33949 21214 33983
rect 21214 33949 21232 33983
rect 21180 33940 21232 33949
rect 23112 33915 23164 33924
rect 23112 33881 23146 33915
rect 23146 33881 23164 33915
rect 16120 33804 16172 33856
rect 23112 33872 23164 33881
rect 23204 33872 23256 33924
rect 25044 33872 25096 33924
rect 27528 34051 27580 34060
rect 27528 34017 27537 34051
rect 27537 34017 27571 34051
rect 27571 34017 27580 34051
rect 27528 34008 27580 34017
rect 29184 34008 29236 34060
rect 30196 34051 30248 34060
rect 30196 34017 30205 34051
rect 30205 34017 30239 34051
rect 30239 34017 30248 34051
rect 30196 34008 30248 34017
rect 31760 34008 31812 34060
rect 28632 33940 28684 33992
rect 30012 33940 30064 33992
rect 32128 34051 32180 34060
rect 32128 34017 32137 34051
rect 32137 34017 32171 34051
rect 32171 34017 32180 34051
rect 32128 34008 32180 34017
rect 32312 33940 32364 33992
rect 32220 33872 32272 33924
rect 36084 34008 36136 34060
rect 33784 33940 33836 33992
rect 36820 34076 36872 34128
rect 33968 33872 34020 33924
rect 40408 34008 40460 34060
rect 40776 34144 40828 34196
rect 41972 34187 42024 34196
rect 41972 34153 41981 34187
rect 41981 34153 42015 34187
rect 42015 34153 42024 34187
rect 41972 34144 42024 34153
rect 40040 33940 40092 33992
rect 41328 33940 41380 33992
rect 17960 33804 18012 33856
rect 18144 33804 18196 33856
rect 20628 33847 20680 33856
rect 20628 33813 20637 33847
rect 20637 33813 20671 33847
rect 20671 33813 20680 33847
rect 20628 33804 20680 33813
rect 22744 33804 22796 33856
rect 23388 33804 23440 33856
rect 26056 33847 26108 33856
rect 26056 33813 26065 33847
rect 26065 33813 26099 33847
rect 26099 33813 26108 33847
rect 26056 33804 26108 33813
rect 28172 33847 28224 33856
rect 28172 33813 28181 33847
rect 28181 33813 28215 33847
rect 28215 33813 28224 33847
rect 28172 33804 28224 33813
rect 28632 33804 28684 33856
rect 29920 33847 29972 33856
rect 29920 33813 29929 33847
rect 29929 33813 29963 33847
rect 29963 33813 29972 33847
rect 29920 33804 29972 33813
rect 30012 33847 30064 33856
rect 30012 33813 30021 33847
rect 30021 33813 30055 33847
rect 30055 33813 30064 33847
rect 30012 33804 30064 33813
rect 32036 33804 32088 33856
rect 32588 33804 32640 33856
rect 34060 33804 34112 33856
rect 36176 33847 36228 33856
rect 36176 33813 36185 33847
rect 36185 33813 36219 33847
rect 36219 33813 36228 33847
rect 36176 33804 36228 33813
rect 36452 33804 36504 33856
rect 38936 33872 38988 33924
rect 39580 33872 39632 33924
rect 40868 33915 40920 33924
rect 40868 33881 40902 33915
rect 40902 33881 40920 33915
rect 40868 33872 40920 33881
rect 36820 33804 36872 33856
rect 38660 33847 38712 33856
rect 38660 33813 38669 33847
rect 38669 33813 38703 33847
rect 38703 33813 38712 33847
rect 38660 33804 38712 33813
rect 39672 33847 39724 33856
rect 39672 33813 39681 33847
rect 39681 33813 39715 33847
rect 39715 33813 39724 33847
rect 39672 33804 39724 33813
rect 40408 33804 40460 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 1676 33600 1728 33652
rect 2688 33600 2740 33652
rect 3516 33600 3568 33652
rect 4804 33600 4856 33652
rect 5724 33600 5776 33652
rect 6736 33600 6788 33652
rect 3608 33532 3660 33584
rect 6460 33532 6512 33584
rect 7104 33600 7156 33652
rect 9404 33600 9456 33652
rect 13544 33600 13596 33652
rect 15108 33600 15160 33652
rect 2780 33464 2832 33516
rect 4068 33464 4120 33516
rect 4804 33464 4856 33516
rect 5448 33464 5500 33516
rect 5632 33464 5684 33516
rect 7840 33532 7892 33584
rect 9128 33532 9180 33584
rect 7196 33464 7248 33516
rect 7932 33464 7984 33516
rect 10232 33507 10284 33516
rect 10232 33473 10266 33507
rect 10266 33473 10284 33507
rect 10232 33464 10284 33473
rect 11520 33464 11572 33516
rect 12808 33464 12860 33516
rect 16120 33643 16172 33652
rect 16120 33609 16129 33643
rect 16129 33609 16163 33643
rect 16163 33609 16172 33643
rect 16120 33600 16172 33609
rect 16948 33600 17000 33652
rect 17592 33643 17644 33652
rect 17592 33609 17601 33643
rect 17601 33609 17635 33643
rect 17635 33609 17644 33643
rect 17592 33600 17644 33609
rect 18512 33600 18564 33652
rect 23112 33600 23164 33652
rect 24308 33600 24360 33652
rect 25044 33643 25096 33652
rect 25044 33609 25053 33643
rect 25053 33609 25087 33643
rect 25087 33609 25096 33643
rect 25044 33600 25096 33609
rect 26056 33600 26108 33652
rect 30932 33600 30984 33652
rect 32588 33643 32640 33652
rect 32588 33609 32597 33643
rect 32597 33609 32631 33643
rect 32631 33609 32640 33643
rect 32588 33600 32640 33609
rect 33416 33643 33468 33652
rect 33416 33609 33425 33643
rect 33425 33609 33459 33643
rect 33459 33609 33468 33643
rect 33416 33600 33468 33609
rect 36176 33600 36228 33652
rect 36820 33600 36872 33652
rect 38752 33600 38804 33652
rect 39580 33643 39632 33652
rect 39580 33609 39589 33643
rect 39589 33609 39623 33643
rect 39623 33609 39632 33643
rect 39580 33600 39632 33609
rect 39948 33643 40000 33652
rect 39948 33609 39957 33643
rect 39957 33609 39991 33643
rect 39991 33609 40000 33643
rect 39948 33600 40000 33609
rect 40408 33643 40460 33652
rect 40408 33609 40417 33643
rect 40417 33609 40451 33643
rect 40451 33609 40460 33643
rect 40408 33600 40460 33609
rect 40868 33600 40920 33652
rect 18052 33532 18104 33584
rect 20536 33532 20588 33584
rect 20628 33532 20680 33584
rect 15476 33464 15528 33516
rect 2136 33396 2188 33448
rect 3516 33439 3568 33448
rect 3516 33405 3525 33439
rect 3525 33405 3559 33439
rect 3559 33405 3568 33439
rect 3516 33396 3568 33405
rect 3608 33439 3660 33448
rect 3608 33405 3617 33439
rect 3617 33405 3651 33439
rect 3651 33405 3660 33439
rect 3608 33396 3660 33405
rect 6920 33396 6972 33448
rect 7380 33439 7432 33448
rect 7380 33405 7389 33439
rect 7389 33405 7423 33439
rect 7423 33405 7432 33439
rect 7380 33396 7432 33405
rect 7472 33396 7524 33448
rect 8024 33396 8076 33448
rect 9956 33439 10008 33448
rect 7288 33328 7340 33380
rect 3148 33303 3200 33312
rect 3148 33269 3157 33303
rect 3157 33269 3191 33303
rect 3191 33269 3200 33303
rect 3148 33260 3200 33269
rect 3240 33303 3292 33312
rect 3240 33269 3249 33303
rect 3249 33269 3283 33303
rect 3283 33269 3292 33303
rect 3240 33260 3292 33269
rect 3792 33260 3844 33312
rect 6828 33303 6880 33312
rect 6828 33269 6837 33303
rect 6837 33269 6871 33303
rect 6871 33269 6880 33303
rect 6828 33260 6880 33269
rect 7104 33303 7156 33312
rect 7104 33269 7113 33303
rect 7113 33269 7147 33303
rect 7147 33269 7156 33303
rect 7104 33260 7156 33269
rect 9956 33405 9965 33439
rect 9965 33405 9999 33439
rect 9999 33405 10008 33439
rect 9956 33396 10008 33405
rect 15568 33439 15620 33448
rect 15568 33405 15577 33439
rect 15577 33405 15611 33439
rect 15611 33405 15620 33439
rect 15568 33396 15620 33405
rect 16488 33464 16540 33516
rect 17868 33464 17920 33516
rect 19524 33464 19576 33516
rect 22836 33532 22888 33584
rect 23940 33532 23992 33584
rect 22100 33507 22152 33516
rect 22100 33473 22134 33507
rect 22134 33473 22152 33507
rect 22100 33464 22152 33473
rect 22376 33464 22428 33516
rect 11060 33260 11112 33312
rect 13452 33303 13504 33312
rect 13452 33269 13461 33303
rect 13461 33269 13495 33303
rect 13495 33269 13504 33303
rect 13452 33260 13504 33269
rect 15292 33260 15344 33312
rect 17040 33260 17092 33312
rect 18420 33439 18472 33448
rect 18420 33405 18429 33439
rect 18429 33405 18463 33439
rect 18463 33405 18472 33439
rect 18420 33396 18472 33405
rect 19432 33396 19484 33448
rect 20076 33396 20128 33448
rect 20628 33439 20680 33448
rect 20628 33405 20637 33439
rect 20637 33405 20671 33439
rect 20671 33405 20680 33439
rect 20628 33396 20680 33405
rect 24032 33396 24084 33448
rect 25872 33464 25924 33516
rect 28356 33464 28408 33516
rect 29736 33507 29788 33516
rect 29736 33473 29770 33507
rect 29770 33473 29788 33507
rect 29736 33464 29788 33473
rect 36544 33532 36596 33584
rect 39304 33532 39356 33584
rect 39672 33532 39724 33584
rect 32588 33464 32640 33516
rect 33784 33507 33836 33516
rect 33784 33473 33793 33507
rect 33793 33473 33827 33507
rect 33827 33473 33836 33507
rect 33784 33464 33836 33473
rect 34060 33464 34112 33516
rect 38108 33464 38160 33516
rect 38568 33464 38620 33516
rect 23388 33328 23440 33380
rect 25780 33396 25832 33448
rect 29460 33439 29512 33448
rect 29460 33405 29469 33439
rect 29469 33405 29503 33439
rect 29503 33405 29512 33439
rect 29460 33396 29512 33405
rect 30564 33328 30616 33380
rect 32680 33328 32732 33380
rect 33968 33439 34020 33448
rect 33968 33405 33977 33439
rect 33977 33405 34011 33439
rect 34011 33405 34020 33439
rect 33968 33396 34020 33405
rect 35808 33396 35860 33448
rect 36452 33396 36504 33448
rect 37372 33396 37424 33448
rect 38384 33396 38436 33448
rect 23480 33260 23532 33312
rect 30196 33260 30248 33312
rect 32128 33303 32180 33312
rect 32128 33269 32137 33303
rect 32137 33269 32171 33303
rect 32171 33269 32180 33303
rect 32128 33260 32180 33269
rect 35440 33303 35492 33312
rect 35440 33269 35449 33303
rect 35449 33269 35483 33303
rect 35483 33269 35492 33303
rect 35440 33260 35492 33269
rect 37648 33260 37700 33312
rect 39028 33396 39080 33448
rect 39120 33371 39172 33380
rect 39120 33337 39129 33371
rect 39129 33337 39163 33371
rect 39163 33337 39172 33371
rect 39120 33328 39172 33337
rect 40040 33396 40092 33448
rect 40316 33507 40368 33516
rect 40316 33473 40325 33507
rect 40325 33473 40359 33507
rect 40359 33473 40368 33507
rect 40316 33464 40368 33473
rect 40960 33396 41012 33448
rect 38844 33260 38896 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5356 32988 5408 33040
rect 6828 33056 6880 33108
rect 7380 33099 7432 33108
rect 7380 33065 7389 33099
rect 7389 33065 7423 33099
rect 7423 33065 7432 33099
rect 7380 33056 7432 33065
rect 10232 33099 10284 33108
rect 10232 33065 10241 33099
rect 10241 33065 10275 33099
rect 10275 33065 10284 33099
rect 10232 33056 10284 33065
rect 10324 33099 10376 33108
rect 10324 33065 10333 33099
rect 10333 33065 10367 33099
rect 10367 33065 10376 33099
rect 10324 33056 10376 33065
rect 10876 33056 10928 33108
rect 6368 32988 6420 33040
rect 1676 32963 1728 32972
rect 1676 32929 1685 32963
rect 1685 32929 1719 32963
rect 1719 32929 1728 32963
rect 1676 32920 1728 32929
rect 3516 32920 3568 32972
rect 9956 32988 10008 33040
rect 2964 32784 3016 32836
rect 3608 32852 3660 32904
rect 4068 32852 4120 32904
rect 4712 32784 4764 32836
rect 5356 32895 5408 32904
rect 5356 32861 5365 32895
rect 5365 32861 5399 32895
rect 5399 32861 5408 32895
rect 5356 32852 5408 32861
rect 5632 32852 5684 32904
rect 5908 32852 5960 32904
rect 6736 32852 6788 32904
rect 6920 32895 6972 32904
rect 6920 32861 6929 32895
rect 6929 32861 6963 32895
rect 6963 32861 6972 32895
rect 6920 32852 6972 32861
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 7656 32895 7708 32904
rect 7656 32861 7665 32895
rect 7665 32861 7699 32895
rect 7699 32861 7708 32895
rect 7656 32852 7708 32861
rect 10324 32920 10376 32972
rect 10968 32963 11020 32972
rect 10968 32929 10977 32963
rect 10977 32929 11011 32963
rect 11011 32929 11020 32963
rect 10968 32920 11020 32929
rect 12808 33099 12860 33108
rect 12808 33065 12817 33099
rect 12817 33065 12851 33099
rect 12851 33065 12860 33099
rect 12808 33056 12860 33065
rect 13912 33056 13964 33108
rect 13820 32988 13872 33040
rect 16488 33056 16540 33108
rect 22100 33056 22152 33108
rect 23848 33056 23900 33108
rect 13176 32920 13228 32972
rect 13544 32920 13596 32972
rect 8392 32852 8444 32904
rect 8484 32784 8536 32836
rect 10876 32784 10928 32836
rect 11152 32852 11204 32904
rect 13452 32852 13504 32904
rect 14004 32852 14056 32904
rect 14372 32852 14424 32904
rect 15568 32920 15620 32972
rect 20076 32963 20128 32972
rect 20076 32929 20085 32963
rect 20085 32929 20119 32963
rect 20119 32929 20128 32963
rect 20076 32920 20128 32929
rect 20628 32920 20680 32972
rect 22376 32963 22428 32972
rect 22376 32929 22385 32963
rect 22385 32929 22419 32963
rect 22419 32929 22428 32963
rect 22376 32920 22428 32929
rect 26148 32920 26200 32972
rect 26700 32963 26752 32972
rect 26700 32929 26709 32963
rect 26709 32929 26743 32963
rect 26743 32929 26752 32963
rect 26700 32920 26752 32929
rect 29736 33056 29788 33108
rect 32312 33056 32364 33108
rect 38660 33056 38712 33108
rect 21824 32852 21876 32904
rect 23480 32852 23532 32904
rect 24124 32895 24176 32904
rect 24124 32861 24133 32895
rect 24133 32861 24167 32895
rect 24167 32861 24176 32895
rect 24124 32852 24176 32861
rect 27896 32852 27948 32904
rect 12164 32784 12216 32836
rect 15200 32827 15252 32836
rect 15200 32793 15209 32827
rect 15209 32793 15243 32827
rect 15243 32793 15252 32827
rect 15200 32784 15252 32793
rect 15292 32784 15344 32836
rect 17316 32827 17368 32836
rect 17316 32793 17325 32827
rect 17325 32793 17359 32827
rect 17359 32793 17368 32827
rect 17316 32784 17368 32793
rect 19432 32784 19484 32836
rect 23388 32784 23440 32836
rect 24492 32784 24544 32836
rect 28172 32920 28224 32972
rect 30196 32920 30248 32972
rect 38844 33099 38896 33108
rect 38844 33065 38853 33099
rect 38853 33065 38887 33099
rect 38887 33065 38896 33099
rect 38844 33056 38896 33065
rect 30564 32852 30616 32904
rect 40960 32963 41012 32972
rect 40960 32929 40969 32963
rect 40969 32929 41003 32963
rect 41003 32929 41012 32963
rect 40960 32920 41012 32929
rect 41420 32920 41472 32972
rect 29460 32784 29512 32836
rect 3332 32716 3384 32768
rect 3516 32716 3568 32768
rect 3608 32716 3660 32768
rect 4804 32759 4856 32768
rect 4804 32725 4813 32759
rect 4813 32725 4847 32759
rect 4847 32725 4856 32759
rect 4804 32716 4856 32725
rect 5264 32716 5316 32768
rect 5540 32759 5592 32768
rect 5540 32725 5549 32759
rect 5549 32725 5583 32759
rect 5583 32725 5592 32759
rect 5540 32716 5592 32725
rect 14280 32716 14332 32768
rect 14556 32716 14608 32768
rect 18052 32716 18104 32768
rect 19156 32716 19208 32768
rect 22100 32759 22152 32768
rect 22100 32725 22109 32759
rect 22109 32725 22143 32759
rect 22143 32725 22152 32759
rect 22100 32716 22152 32725
rect 24400 32759 24452 32768
rect 24400 32725 24409 32759
rect 24409 32725 24443 32759
rect 24443 32725 24452 32759
rect 24400 32716 24452 32725
rect 25688 32716 25740 32768
rect 27252 32759 27304 32768
rect 27252 32725 27261 32759
rect 27261 32725 27295 32759
rect 27295 32725 27304 32759
rect 27252 32716 27304 32725
rect 28356 32716 28408 32768
rect 28816 32716 28868 32768
rect 31024 32716 31076 32768
rect 31300 32784 31352 32836
rect 32128 32852 32180 32904
rect 35072 32895 35124 32904
rect 35072 32861 35081 32895
rect 35081 32861 35115 32895
rect 35115 32861 35124 32895
rect 35072 32852 35124 32861
rect 37372 32895 37424 32904
rect 37372 32861 37381 32895
rect 37381 32861 37415 32895
rect 37415 32861 37424 32895
rect 37372 32852 37424 32861
rect 37648 32895 37700 32904
rect 37648 32861 37682 32895
rect 37682 32861 37700 32895
rect 37648 32852 37700 32861
rect 33140 32784 33192 32836
rect 35348 32827 35400 32836
rect 35348 32793 35382 32827
rect 35382 32793 35400 32827
rect 35348 32784 35400 32793
rect 38844 32784 38896 32836
rect 34060 32716 34112 32768
rect 36820 32716 36872 32768
rect 40592 32716 40644 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 2136 32555 2188 32564
rect 2136 32521 2145 32555
rect 2145 32521 2179 32555
rect 2179 32521 2188 32555
rect 2136 32512 2188 32521
rect 2596 32444 2648 32496
rect 3332 32512 3384 32564
rect 3240 32376 3292 32428
rect 3332 32419 3384 32428
rect 3332 32385 3341 32419
rect 3341 32385 3375 32419
rect 3375 32385 3384 32419
rect 3332 32376 3384 32385
rect 3608 32419 3660 32428
rect 3608 32385 3617 32419
rect 3617 32385 3651 32419
rect 3651 32385 3660 32419
rect 3608 32376 3660 32385
rect 3792 32419 3844 32428
rect 3792 32385 3801 32419
rect 3801 32385 3835 32419
rect 3835 32385 3844 32419
rect 3792 32376 3844 32385
rect 5816 32512 5868 32564
rect 14004 32512 14056 32564
rect 6276 32444 6328 32496
rect 7656 32444 7708 32496
rect 13544 32444 13596 32496
rect 14556 32555 14608 32564
rect 14556 32521 14565 32555
rect 14565 32521 14599 32555
rect 14599 32521 14608 32555
rect 14556 32512 14608 32521
rect 17316 32512 17368 32564
rect 18052 32512 18104 32564
rect 18420 32512 18472 32564
rect 22652 32512 22704 32564
rect 23204 32512 23256 32564
rect 23388 32555 23440 32564
rect 23388 32521 23397 32555
rect 23397 32521 23431 32555
rect 23431 32521 23440 32555
rect 23388 32512 23440 32521
rect 24400 32512 24452 32564
rect 26148 32555 26200 32564
rect 26148 32521 26157 32555
rect 26157 32521 26191 32555
rect 26191 32521 26200 32555
rect 26148 32512 26200 32521
rect 28172 32512 28224 32564
rect 33140 32555 33192 32564
rect 33140 32521 33149 32555
rect 33149 32521 33183 32555
rect 33183 32521 33192 32555
rect 33140 32512 33192 32521
rect 36452 32555 36504 32564
rect 36452 32521 36461 32555
rect 36461 32521 36495 32555
rect 36495 32521 36504 32555
rect 36452 32512 36504 32521
rect 38936 32512 38988 32564
rect 41420 32512 41472 32564
rect 19432 32444 19484 32496
rect 19616 32444 19668 32496
rect 20076 32444 20128 32496
rect 24124 32444 24176 32496
rect 3056 32351 3108 32360
rect 3056 32317 3065 32351
rect 3065 32317 3099 32351
rect 3099 32317 3108 32351
rect 6920 32376 6972 32428
rect 7196 32376 7248 32428
rect 8392 32419 8444 32428
rect 8392 32385 8401 32419
rect 8401 32385 8435 32419
rect 8435 32385 8444 32419
rect 8392 32376 8444 32385
rect 3056 32308 3108 32317
rect 3792 32172 3844 32224
rect 4620 32308 4672 32360
rect 7380 32308 7432 32360
rect 8208 32308 8260 32360
rect 9312 32308 9364 32360
rect 12072 32308 12124 32360
rect 14372 32376 14424 32428
rect 14464 32419 14516 32428
rect 14464 32385 14473 32419
rect 14473 32385 14507 32419
rect 14507 32385 14516 32419
rect 14464 32376 14516 32385
rect 18420 32376 18472 32428
rect 19156 32419 19208 32428
rect 15476 32308 15528 32360
rect 18052 32308 18104 32360
rect 7748 32240 7800 32292
rect 16028 32240 16080 32292
rect 18788 32240 18840 32292
rect 4620 32172 4672 32224
rect 5080 32172 5132 32224
rect 5632 32172 5684 32224
rect 5908 32172 5960 32224
rect 7932 32215 7984 32224
rect 7932 32181 7941 32215
rect 7941 32181 7975 32215
rect 7975 32181 7984 32215
rect 7932 32172 7984 32181
rect 8668 32215 8720 32224
rect 8668 32181 8677 32215
rect 8677 32181 8711 32215
rect 8711 32181 8720 32215
rect 8668 32172 8720 32181
rect 10508 32172 10560 32224
rect 17500 32172 17552 32224
rect 17776 32172 17828 32224
rect 19156 32385 19164 32419
rect 19164 32385 19198 32419
rect 19198 32385 19208 32419
rect 19156 32376 19208 32385
rect 19248 32419 19300 32428
rect 19248 32385 19257 32419
rect 19257 32385 19291 32419
rect 19291 32385 19300 32419
rect 19248 32376 19300 32385
rect 27436 32444 27488 32496
rect 25044 32419 25096 32428
rect 25044 32385 25078 32419
rect 25078 32385 25096 32419
rect 25044 32376 25096 32385
rect 26976 32419 27028 32428
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 27252 32419 27304 32428
rect 27252 32385 27286 32419
rect 27286 32385 27304 32419
rect 27252 32376 27304 32385
rect 20168 32351 20220 32360
rect 20168 32317 20177 32351
rect 20177 32317 20211 32351
rect 20211 32317 20220 32351
rect 20168 32308 20220 32317
rect 20536 32308 20588 32360
rect 21916 32308 21968 32360
rect 24032 32351 24084 32360
rect 24032 32317 24041 32351
rect 24041 32317 24075 32351
rect 24075 32317 24084 32351
rect 24032 32308 24084 32317
rect 24124 32308 24176 32360
rect 28816 32444 28868 32496
rect 33416 32444 33468 32496
rect 35440 32444 35492 32496
rect 28540 32376 28592 32428
rect 29644 32376 29696 32428
rect 29920 32419 29972 32428
rect 29920 32385 29929 32419
rect 29929 32385 29963 32419
rect 29963 32385 29972 32419
rect 29920 32376 29972 32385
rect 33508 32419 33560 32428
rect 33508 32385 33517 32419
rect 33517 32385 33551 32419
rect 33551 32385 33560 32419
rect 33508 32376 33560 32385
rect 34060 32376 34112 32428
rect 34704 32376 34756 32428
rect 35072 32419 35124 32428
rect 35072 32385 35081 32419
rect 35081 32385 35115 32419
rect 35115 32385 35124 32419
rect 35072 32376 35124 32385
rect 37648 32419 37700 32428
rect 37648 32385 37682 32419
rect 37682 32385 37700 32419
rect 37648 32376 37700 32385
rect 40592 32487 40644 32496
rect 40592 32453 40626 32487
rect 40626 32453 40644 32487
rect 40592 32444 40644 32453
rect 40408 32376 40460 32428
rect 41972 32376 42024 32428
rect 18972 32240 19024 32292
rect 20904 32172 20956 32224
rect 21824 32172 21876 32224
rect 28356 32172 28408 32224
rect 30012 32308 30064 32360
rect 32128 32351 32180 32360
rect 32128 32317 32137 32351
rect 32137 32317 32171 32351
rect 32171 32317 32180 32351
rect 32128 32308 32180 32317
rect 34244 32308 34296 32360
rect 37372 32351 37424 32360
rect 37372 32317 37381 32351
rect 37381 32317 37415 32351
rect 37415 32317 37424 32351
rect 37372 32308 37424 32317
rect 31300 32240 31352 32292
rect 33048 32240 33100 32292
rect 29460 32172 29512 32224
rect 30564 32215 30616 32224
rect 30564 32181 30573 32215
rect 30573 32181 30607 32215
rect 30607 32181 30616 32215
rect 30564 32172 30616 32181
rect 30656 32215 30708 32224
rect 30656 32181 30665 32215
rect 30665 32181 30699 32215
rect 30699 32181 30708 32215
rect 30656 32172 30708 32181
rect 31024 32172 31076 32224
rect 31392 32172 31444 32224
rect 32772 32215 32824 32224
rect 32772 32181 32781 32215
rect 32781 32181 32815 32215
rect 32815 32181 32824 32215
rect 32772 32172 32824 32181
rect 38292 32172 38344 32224
rect 42064 32215 42116 32224
rect 42064 32181 42073 32215
rect 42073 32181 42107 32215
rect 42107 32181 42116 32215
rect 42064 32172 42116 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 3056 31968 3108 32020
rect 4712 32011 4764 32020
rect 4712 31977 4721 32011
rect 4721 31977 4755 32011
rect 4755 31977 4764 32011
rect 4712 31968 4764 31977
rect 5356 31968 5408 32020
rect 5724 31968 5776 32020
rect 6368 32011 6420 32020
rect 6368 31977 6377 32011
rect 6377 31977 6411 32011
rect 6411 31977 6420 32011
rect 6368 31968 6420 31977
rect 7380 31968 7432 32020
rect 8208 31968 8260 32020
rect 9312 32011 9364 32020
rect 9312 31977 9321 32011
rect 9321 31977 9355 32011
rect 9355 31977 9364 32011
rect 9312 31968 9364 31977
rect 12900 31968 12952 32020
rect 13544 32011 13596 32020
rect 13544 31977 13553 32011
rect 13553 31977 13587 32011
rect 13587 31977 13596 32011
rect 13544 31968 13596 31977
rect 15200 31968 15252 32020
rect 16028 31968 16080 32020
rect 16764 31968 16816 32020
rect 4804 31832 4856 31884
rect 3424 31764 3476 31816
rect 5264 31764 5316 31816
rect 5908 31900 5960 31952
rect 6368 31832 6420 31884
rect 7748 31832 7800 31884
rect 10416 31832 10468 31884
rect 5632 31807 5684 31816
rect 5632 31773 5641 31807
rect 5641 31773 5675 31807
rect 5675 31773 5684 31807
rect 5632 31764 5684 31773
rect 6644 31807 6696 31816
rect 5356 31696 5408 31748
rect 6644 31773 6653 31807
rect 6653 31773 6687 31807
rect 6687 31773 6696 31807
rect 6644 31764 6696 31773
rect 6828 31807 6880 31816
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 6920 31807 6972 31816
rect 6920 31773 6929 31807
rect 6929 31773 6963 31807
rect 6963 31773 6972 31807
rect 6920 31764 6972 31773
rect 6000 31696 6052 31748
rect 7196 31739 7248 31748
rect 7196 31705 7205 31739
rect 7205 31705 7239 31739
rect 7239 31705 7248 31739
rect 7196 31696 7248 31705
rect 3976 31628 4028 31680
rect 8208 31628 8260 31680
rect 10784 31739 10836 31748
rect 10784 31705 10793 31739
rect 10793 31705 10827 31739
rect 10827 31705 10836 31739
rect 10784 31696 10836 31705
rect 10876 31696 10928 31748
rect 11520 31764 11572 31816
rect 12164 31807 12216 31816
rect 12164 31773 12173 31807
rect 12173 31773 12207 31807
rect 12207 31773 12216 31807
rect 12164 31764 12216 31773
rect 13820 31807 13872 31816
rect 13820 31773 13829 31807
rect 13829 31773 13863 31807
rect 13863 31773 13872 31807
rect 13820 31764 13872 31773
rect 15844 31807 15896 31816
rect 15844 31773 15853 31807
rect 15853 31773 15887 31807
rect 15887 31773 15896 31807
rect 15844 31764 15896 31773
rect 16948 31900 17000 31952
rect 18052 32011 18104 32020
rect 18052 31977 18061 32011
rect 18061 31977 18095 32011
rect 18095 31977 18104 32011
rect 18052 31968 18104 31977
rect 18788 31968 18840 32020
rect 21180 31968 21232 32020
rect 20168 31900 20220 31952
rect 16396 31764 16448 31816
rect 16580 31807 16632 31816
rect 16580 31773 16589 31807
rect 16589 31773 16623 31807
rect 16623 31773 16632 31807
rect 16580 31764 16632 31773
rect 16764 31764 16816 31816
rect 16856 31807 16908 31816
rect 16856 31773 16865 31807
rect 16865 31773 16899 31807
rect 16899 31773 16908 31807
rect 16856 31764 16908 31773
rect 12072 31696 12124 31748
rect 17132 31764 17184 31816
rect 17316 31807 17368 31816
rect 17316 31773 17325 31807
rect 17325 31773 17359 31807
rect 17359 31773 17368 31807
rect 17316 31764 17368 31773
rect 17408 31764 17460 31816
rect 18052 31764 18104 31816
rect 18328 31807 18380 31816
rect 18328 31773 18337 31807
rect 18337 31773 18371 31807
rect 18371 31773 18380 31807
rect 18328 31764 18380 31773
rect 10968 31628 11020 31680
rect 13452 31628 13504 31680
rect 16672 31628 16724 31680
rect 17316 31628 17368 31680
rect 17684 31628 17736 31680
rect 18604 31807 18656 31816
rect 18604 31773 18612 31807
rect 18612 31773 18646 31807
rect 18646 31773 18656 31807
rect 18604 31764 18656 31773
rect 18788 31807 18840 31816
rect 18788 31773 18797 31807
rect 18797 31773 18831 31807
rect 18831 31773 18840 31807
rect 18788 31764 18840 31773
rect 19432 31764 19484 31816
rect 20812 31764 20864 31816
rect 19616 31696 19668 31748
rect 20996 31807 21048 31816
rect 20996 31773 21005 31807
rect 21005 31773 21039 31807
rect 21039 31773 21048 31807
rect 20996 31764 21048 31773
rect 21456 31900 21508 31952
rect 25044 31968 25096 32020
rect 26700 31968 26752 32020
rect 27528 31968 27580 32020
rect 28540 32011 28592 32020
rect 28540 31977 28549 32011
rect 28549 31977 28583 32011
rect 28583 31977 28592 32011
rect 28540 31968 28592 31977
rect 28632 31900 28684 31952
rect 25504 31832 25556 31884
rect 25688 31875 25740 31884
rect 25688 31841 25697 31875
rect 25697 31841 25731 31875
rect 25731 31841 25740 31875
rect 25688 31832 25740 31841
rect 25780 31875 25832 31884
rect 25780 31841 25789 31875
rect 25789 31841 25823 31875
rect 25823 31841 25832 31875
rect 25780 31832 25832 31841
rect 30656 31968 30708 32020
rect 32128 31968 32180 32020
rect 35348 31968 35400 32020
rect 37648 31968 37700 32020
rect 33784 31900 33836 31952
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 21640 31807 21692 31816
rect 21640 31773 21649 31807
rect 21649 31773 21683 31807
rect 21683 31773 21692 31807
rect 21640 31764 21692 31773
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 23756 31807 23808 31816
rect 23756 31773 23765 31807
rect 23765 31773 23799 31807
rect 23799 31773 23808 31807
rect 23756 31764 23808 31773
rect 23848 31807 23900 31816
rect 23848 31773 23857 31807
rect 23857 31773 23891 31807
rect 23891 31773 23900 31807
rect 23848 31764 23900 31773
rect 24124 31807 24176 31816
rect 24124 31773 24133 31807
rect 24133 31773 24167 31807
rect 24167 31773 24176 31807
rect 24124 31764 24176 31773
rect 26976 31764 27028 31816
rect 27528 31764 27580 31816
rect 29460 31832 29512 31884
rect 34244 31943 34296 31952
rect 34244 31909 34253 31943
rect 34253 31909 34287 31943
rect 34287 31909 34296 31943
rect 34244 31900 34296 31909
rect 35808 31832 35860 31884
rect 36820 31875 36872 31884
rect 36820 31841 36829 31875
rect 36829 31841 36863 31875
rect 36863 31841 36872 31875
rect 36820 31832 36872 31841
rect 38292 31875 38344 31884
rect 38292 31841 38301 31875
rect 38301 31841 38335 31875
rect 38335 31841 38344 31875
rect 38292 31832 38344 31841
rect 39028 31875 39080 31884
rect 39028 31841 39037 31875
rect 39037 31841 39071 31875
rect 39071 31841 39080 31875
rect 39028 31832 39080 31841
rect 41236 31943 41288 31952
rect 41236 31909 41245 31943
rect 41245 31909 41279 31943
rect 41279 31909 41288 31943
rect 41236 31900 41288 31909
rect 20720 31628 20772 31680
rect 21456 31696 21508 31748
rect 26240 31696 26292 31748
rect 30380 31764 30432 31816
rect 31208 31764 31260 31816
rect 33324 31764 33376 31816
rect 33416 31764 33468 31816
rect 37372 31764 37424 31816
rect 40408 31764 40460 31816
rect 30196 31696 30248 31748
rect 32128 31739 32180 31748
rect 32128 31705 32146 31739
rect 32146 31705 32180 31739
rect 32128 31696 32180 31705
rect 22376 31628 22428 31680
rect 23480 31628 23532 31680
rect 25596 31671 25648 31680
rect 25596 31637 25605 31671
rect 25605 31637 25639 31671
rect 25639 31637 25648 31671
rect 25596 31628 25648 31637
rect 30012 31628 30064 31680
rect 31576 31628 31628 31680
rect 32588 31628 32640 31680
rect 32864 31628 32916 31680
rect 34520 31628 34572 31680
rect 35992 31628 36044 31680
rect 36084 31628 36136 31680
rect 38292 31628 38344 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 2596 31467 2648 31476
rect 2596 31433 2605 31467
rect 2605 31433 2639 31467
rect 2639 31433 2648 31467
rect 2596 31424 2648 31433
rect 3608 31424 3660 31476
rect 4068 31424 4120 31476
rect 5172 31467 5224 31476
rect 5172 31433 5181 31467
rect 5181 31433 5215 31467
rect 5215 31433 5224 31467
rect 5172 31424 5224 31433
rect 5356 31467 5408 31476
rect 5356 31433 5383 31467
rect 5383 31433 5408 31467
rect 5356 31424 5408 31433
rect 2872 31356 2924 31408
rect 3516 31356 3568 31408
rect 5908 31424 5960 31476
rect 7196 31424 7248 31476
rect 6092 31356 6144 31408
rect 3240 31288 3292 31340
rect 3148 31220 3200 31272
rect 3056 31152 3108 31204
rect 5816 31288 5868 31340
rect 6368 31288 6420 31340
rect 4620 31220 4672 31272
rect 7748 31331 7800 31340
rect 7748 31297 7757 31331
rect 7757 31297 7791 31331
rect 7791 31297 7800 31331
rect 7748 31288 7800 31297
rect 8668 31424 8720 31476
rect 13820 31424 13872 31476
rect 8024 31356 8076 31408
rect 10968 31356 11020 31408
rect 15292 31424 15344 31476
rect 15384 31424 15436 31476
rect 15936 31467 15988 31476
rect 15936 31433 15945 31467
rect 15945 31433 15979 31467
rect 15979 31433 15988 31467
rect 15936 31424 15988 31433
rect 17040 31467 17092 31476
rect 17040 31433 17049 31467
rect 17049 31433 17083 31467
rect 17083 31433 17092 31467
rect 17040 31424 17092 31433
rect 17316 31424 17368 31476
rect 19064 31424 19116 31476
rect 19616 31467 19668 31476
rect 19616 31433 19625 31467
rect 19625 31433 19659 31467
rect 19659 31433 19668 31467
rect 19616 31424 19668 31433
rect 21640 31424 21692 31476
rect 23848 31424 23900 31476
rect 7932 31288 7984 31340
rect 11520 31331 11572 31340
rect 6920 31220 6972 31272
rect 10140 31220 10192 31272
rect 11520 31297 11529 31331
rect 11529 31297 11563 31331
rect 11563 31297 11572 31331
rect 11520 31288 11572 31297
rect 12072 31263 12124 31272
rect 12072 31229 12081 31263
rect 12081 31229 12115 31263
rect 12115 31229 12124 31263
rect 12072 31220 12124 31229
rect 4896 31152 4948 31204
rect 1676 31084 1728 31136
rect 2964 31084 3016 31136
rect 3332 31084 3384 31136
rect 4068 31127 4120 31136
rect 4068 31093 4077 31127
rect 4077 31093 4111 31127
rect 4111 31093 4120 31127
rect 4068 31084 4120 31093
rect 6092 31152 6144 31204
rect 13728 31152 13780 31204
rect 15200 31263 15252 31272
rect 15200 31229 15209 31263
rect 15209 31229 15243 31263
rect 15243 31229 15252 31263
rect 15200 31220 15252 31229
rect 16212 31331 16264 31340
rect 16212 31297 16221 31331
rect 16221 31297 16255 31331
rect 16255 31297 16264 31331
rect 16212 31288 16264 31297
rect 16396 31288 16448 31340
rect 16856 31288 16908 31340
rect 17316 31288 17368 31340
rect 17500 31331 17552 31340
rect 17500 31297 17509 31331
rect 17509 31297 17543 31331
rect 17543 31297 17552 31331
rect 17500 31288 17552 31297
rect 15476 31152 15528 31204
rect 5632 31127 5684 31136
rect 5632 31093 5641 31127
rect 5641 31093 5675 31127
rect 5675 31093 5684 31127
rect 5632 31084 5684 31093
rect 5816 31084 5868 31136
rect 8208 31084 8260 31136
rect 11980 31127 12032 31136
rect 11980 31093 11989 31127
rect 11989 31093 12023 31127
rect 12023 31093 12032 31127
rect 11980 31084 12032 31093
rect 12164 31084 12216 31136
rect 14372 31084 14424 31136
rect 15660 31084 15712 31136
rect 15752 31084 15804 31136
rect 17776 31331 17828 31340
rect 17776 31297 17785 31331
rect 17785 31297 17819 31331
rect 17819 31297 17828 31331
rect 17776 31288 17828 31297
rect 17868 31331 17920 31340
rect 17868 31297 17877 31331
rect 17877 31297 17911 31331
rect 17911 31297 17920 31331
rect 17868 31288 17920 31297
rect 18880 31288 18932 31340
rect 19800 31356 19852 31408
rect 19708 31331 19760 31340
rect 19708 31297 19717 31331
rect 19717 31297 19751 31331
rect 19751 31297 19760 31331
rect 19708 31288 19760 31297
rect 16396 31152 16448 31204
rect 19432 31220 19484 31272
rect 20168 31288 20220 31340
rect 20076 31152 20128 31204
rect 20352 31331 20404 31340
rect 20352 31297 20361 31331
rect 20361 31297 20395 31331
rect 20395 31297 20404 31331
rect 20352 31288 20404 31297
rect 20996 31399 21048 31408
rect 20996 31365 21005 31399
rect 21005 31365 21039 31399
rect 21039 31365 21048 31399
rect 20996 31356 21048 31365
rect 21732 31356 21784 31408
rect 23480 31356 23532 31408
rect 25136 31424 25188 31476
rect 25320 31424 25372 31476
rect 26240 31424 26292 31476
rect 29644 31424 29696 31476
rect 27712 31356 27764 31408
rect 30380 31424 30432 31476
rect 32772 31424 32824 31476
rect 33324 31467 33376 31476
rect 33324 31433 33333 31467
rect 33333 31433 33367 31467
rect 33367 31433 33376 31467
rect 33324 31424 33376 31433
rect 34520 31424 34572 31476
rect 35348 31356 35400 31408
rect 20904 31331 20956 31340
rect 20904 31297 20911 31331
rect 20911 31297 20956 31331
rect 20904 31288 20956 31297
rect 21640 31288 21692 31340
rect 24952 31331 25004 31340
rect 24952 31297 24961 31331
rect 24961 31297 24995 31331
rect 24995 31297 25004 31331
rect 24952 31288 25004 31297
rect 25228 31288 25280 31340
rect 22468 31220 22520 31272
rect 22928 31263 22980 31272
rect 22928 31229 22937 31263
rect 22937 31229 22971 31263
rect 22971 31229 22980 31263
rect 22928 31220 22980 31229
rect 16856 31084 16908 31136
rect 17040 31084 17092 31136
rect 18328 31084 18380 31136
rect 19892 31084 19944 31136
rect 20720 31152 20772 31204
rect 21088 31152 21140 31204
rect 23848 31220 23900 31272
rect 24400 31220 24452 31272
rect 28816 31288 28868 31340
rect 29552 31288 29604 31340
rect 30104 31331 30156 31340
rect 30104 31297 30113 31331
rect 30113 31297 30147 31331
rect 30147 31297 30156 31331
rect 30104 31288 30156 31297
rect 30564 31288 30616 31340
rect 30748 31288 30800 31340
rect 32496 31331 32548 31340
rect 32496 31297 32505 31331
rect 32505 31297 32539 31331
rect 32539 31297 32548 31331
rect 32496 31288 32548 31297
rect 34152 31288 34204 31340
rect 34612 31288 34664 31340
rect 24216 31152 24268 31204
rect 24584 31152 24636 31204
rect 27528 31263 27580 31272
rect 27528 31229 27537 31263
rect 27537 31229 27571 31263
rect 27571 31229 27580 31263
rect 27528 31220 27580 31229
rect 30288 31263 30340 31272
rect 30288 31229 30297 31263
rect 30297 31229 30331 31263
rect 30331 31229 30340 31263
rect 30288 31220 30340 31229
rect 31024 31263 31076 31272
rect 31024 31229 31033 31263
rect 31033 31229 31067 31263
rect 31067 31229 31076 31263
rect 31024 31220 31076 31229
rect 32680 31263 32732 31272
rect 32680 31229 32689 31263
rect 32689 31229 32723 31263
rect 32723 31229 32732 31263
rect 32680 31220 32732 31229
rect 34244 31220 34296 31272
rect 34520 31220 34572 31272
rect 34796 31220 34848 31272
rect 35992 31288 36044 31340
rect 36268 31220 36320 31272
rect 36636 31356 36688 31408
rect 37004 31356 37056 31408
rect 37280 31331 37332 31340
rect 37280 31297 37289 31331
rect 37289 31297 37323 31331
rect 37323 31297 37332 31331
rect 37280 31288 37332 31297
rect 37464 31288 37516 31340
rect 37832 31288 37884 31340
rect 40132 31331 40184 31340
rect 40132 31297 40141 31331
rect 40141 31297 40175 31331
rect 40175 31297 40184 31331
rect 40132 31288 40184 31297
rect 41972 31424 42024 31476
rect 40408 31331 40460 31340
rect 40408 31297 40417 31331
rect 40417 31297 40451 31331
rect 40451 31297 40460 31331
rect 40408 31288 40460 31297
rect 41788 31288 41840 31340
rect 41052 31220 41104 31272
rect 34336 31152 34388 31204
rect 37740 31152 37792 31204
rect 20536 31127 20588 31136
rect 20536 31093 20545 31127
rect 20545 31093 20579 31127
rect 20579 31093 20588 31127
rect 20536 31084 20588 31093
rect 20812 31084 20864 31136
rect 24308 31084 24360 31136
rect 32772 31084 32824 31136
rect 34796 31084 34848 31136
rect 37648 31084 37700 31136
rect 40868 31084 40920 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3148 30923 3200 30932
rect 3148 30889 3157 30923
rect 3157 30889 3191 30923
rect 3191 30889 3200 30923
rect 3148 30880 3200 30889
rect 3240 30923 3292 30932
rect 3240 30889 3249 30923
rect 3249 30889 3283 30923
rect 3283 30889 3292 30923
rect 3240 30880 3292 30889
rect 3516 30880 3568 30932
rect 4804 30880 4856 30932
rect 5632 30880 5684 30932
rect 10784 30923 10836 30932
rect 10784 30889 10793 30923
rect 10793 30889 10827 30923
rect 10827 30889 10836 30923
rect 10784 30880 10836 30889
rect 12900 30880 12952 30932
rect 14464 30880 14516 30932
rect 15016 30923 15068 30932
rect 15016 30889 15025 30923
rect 15025 30889 15059 30923
rect 15059 30889 15068 30923
rect 15016 30880 15068 30889
rect 15844 30880 15896 30932
rect 16212 30880 16264 30932
rect 16396 30880 16448 30932
rect 17408 30880 17460 30932
rect 18788 30880 18840 30932
rect 19432 30923 19484 30932
rect 19432 30889 19441 30923
rect 19441 30889 19475 30923
rect 19475 30889 19484 30923
rect 19432 30880 19484 30889
rect 3792 30855 3844 30864
rect 3792 30821 3801 30855
rect 3801 30821 3835 30855
rect 3835 30821 3844 30855
rect 3792 30812 3844 30821
rect 5540 30812 5592 30864
rect 4620 30744 4672 30796
rect 4896 30744 4948 30796
rect 5172 30787 5224 30796
rect 5172 30753 5181 30787
rect 5181 30753 5215 30787
rect 5215 30753 5224 30787
rect 5172 30744 5224 30753
rect 6920 30787 6972 30796
rect 6920 30753 6929 30787
rect 6929 30753 6963 30787
rect 6963 30753 6972 30787
rect 6920 30744 6972 30753
rect 10508 30787 10560 30796
rect 10508 30753 10517 30787
rect 10517 30753 10551 30787
rect 10551 30753 10560 30787
rect 10508 30744 10560 30753
rect 10876 30787 10928 30796
rect 10876 30753 10885 30787
rect 10885 30753 10919 30787
rect 10919 30753 10928 30787
rect 10876 30744 10928 30753
rect 19800 30880 19852 30932
rect 20352 30880 20404 30932
rect 20628 30923 20680 30932
rect 20628 30889 20637 30923
rect 20637 30889 20671 30923
rect 20671 30889 20680 30923
rect 20628 30880 20680 30889
rect 23664 30880 23716 30932
rect 23756 30880 23808 30932
rect 14372 30787 14424 30796
rect 14372 30753 14381 30787
rect 14381 30753 14415 30787
rect 14415 30753 14424 30787
rect 14372 30744 14424 30753
rect 15660 30744 15712 30796
rect 16580 30787 16632 30796
rect 16580 30753 16589 30787
rect 16589 30753 16623 30787
rect 16623 30753 16632 30787
rect 16580 30744 16632 30753
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 3056 30608 3108 30660
rect 3516 30719 3568 30728
rect 3516 30685 3525 30719
rect 3525 30685 3559 30719
rect 3559 30685 3568 30719
rect 3516 30676 3568 30685
rect 4068 30719 4120 30728
rect 4068 30685 4077 30719
rect 4077 30685 4111 30719
rect 4111 30685 4120 30719
rect 4068 30676 4120 30685
rect 4252 30676 4304 30728
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 6000 30676 6052 30728
rect 6092 30719 6144 30728
rect 6092 30685 6101 30719
rect 6101 30685 6135 30719
rect 6135 30685 6144 30719
rect 6092 30676 6144 30685
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 10600 30676 10652 30685
rect 13452 30719 13504 30728
rect 13452 30685 13461 30719
rect 13461 30685 13495 30719
rect 13495 30685 13504 30719
rect 13452 30676 13504 30685
rect 13820 30676 13872 30728
rect 14188 30676 14240 30728
rect 15568 30719 15620 30728
rect 15568 30685 15577 30719
rect 15577 30685 15611 30719
rect 15611 30685 15620 30719
rect 15568 30676 15620 30685
rect 16120 30676 16172 30728
rect 16304 30719 16356 30728
rect 16304 30685 16313 30719
rect 16313 30685 16347 30719
rect 16347 30685 16356 30719
rect 16304 30676 16356 30685
rect 5264 30608 5316 30660
rect 3148 30540 3200 30592
rect 4068 30540 4120 30592
rect 4620 30540 4672 30592
rect 5448 30583 5500 30592
rect 5448 30549 5457 30583
rect 5457 30549 5491 30583
rect 5491 30549 5500 30583
rect 5448 30540 5500 30549
rect 6184 30651 6236 30660
rect 6184 30617 6193 30651
rect 6193 30617 6227 30651
rect 6227 30617 6236 30651
rect 6184 30608 6236 30617
rect 11152 30651 11204 30660
rect 11152 30617 11161 30651
rect 11161 30617 11195 30651
rect 11195 30617 11204 30651
rect 11152 30608 11204 30617
rect 10692 30540 10744 30592
rect 10968 30540 11020 30592
rect 15108 30608 15160 30660
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 18420 30744 18472 30796
rect 18880 30787 18932 30796
rect 18880 30753 18889 30787
rect 18889 30753 18923 30787
rect 18923 30753 18932 30787
rect 18880 30744 18932 30753
rect 17684 30719 17736 30728
rect 17684 30685 17693 30719
rect 17693 30685 17727 30719
rect 17727 30685 17736 30719
rect 17684 30676 17736 30685
rect 17776 30676 17828 30728
rect 18144 30719 18196 30728
rect 18144 30685 18153 30719
rect 18153 30685 18187 30719
rect 18187 30685 18196 30719
rect 18144 30676 18196 30685
rect 18512 30676 18564 30728
rect 12716 30583 12768 30592
rect 12716 30549 12725 30583
rect 12725 30549 12759 30583
rect 12759 30549 12768 30583
rect 12716 30540 12768 30549
rect 13728 30540 13780 30592
rect 15200 30540 15252 30592
rect 17040 30608 17092 30660
rect 17132 30651 17184 30660
rect 17132 30617 17141 30651
rect 17141 30617 17175 30651
rect 17175 30617 17184 30651
rect 17132 30608 17184 30617
rect 16488 30540 16540 30592
rect 17408 30540 17460 30592
rect 18696 30540 18748 30592
rect 19524 30651 19576 30660
rect 19524 30617 19533 30651
rect 19533 30617 19567 30651
rect 19567 30617 19576 30651
rect 19524 30608 19576 30617
rect 21640 30812 21692 30864
rect 24952 30880 25004 30932
rect 24584 30812 24636 30864
rect 20076 30744 20128 30796
rect 20812 30787 20864 30796
rect 19800 30608 19852 30660
rect 19892 30608 19944 30660
rect 20352 30719 20404 30728
rect 20352 30685 20381 30719
rect 20381 30685 20404 30719
rect 20352 30676 20404 30685
rect 20812 30753 20821 30787
rect 20821 30753 20855 30787
rect 20855 30753 20864 30787
rect 20812 30744 20864 30753
rect 21088 30744 21140 30796
rect 21916 30744 21968 30796
rect 24952 30744 25004 30796
rect 20720 30676 20772 30728
rect 22100 30676 22152 30728
rect 23756 30719 23808 30728
rect 23756 30685 23765 30719
rect 23765 30685 23799 30719
rect 23799 30685 23808 30719
rect 23756 30676 23808 30685
rect 24032 30676 24084 30728
rect 24400 30676 24452 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 24676 30719 24728 30728
rect 24676 30685 24685 30719
rect 24685 30685 24719 30719
rect 24719 30685 24728 30719
rect 24676 30676 24728 30685
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 31024 30923 31076 30932
rect 31024 30889 31033 30923
rect 31033 30889 31067 30923
rect 31067 30889 31076 30923
rect 31024 30880 31076 30889
rect 32128 30880 32180 30932
rect 34796 30880 34848 30932
rect 35992 30880 36044 30932
rect 37464 30880 37516 30932
rect 41052 30923 41104 30932
rect 41052 30889 41061 30923
rect 41061 30889 41095 30923
rect 41095 30889 41104 30923
rect 41052 30880 41104 30889
rect 22652 30608 22704 30660
rect 23848 30651 23900 30660
rect 23848 30617 23857 30651
rect 23857 30617 23891 30651
rect 23891 30617 23900 30651
rect 23848 30608 23900 30617
rect 26056 30676 26108 30728
rect 28264 30744 28316 30796
rect 30840 30812 30892 30864
rect 32496 30812 32548 30864
rect 31576 30787 31628 30796
rect 31576 30753 31585 30787
rect 31585 30753 31619 30787
rect 31619 30753 31628 30787
rect 31576 30744 31628 30753
rect 32772 30787 32824 30796
rect 32772 30753 32781 30787
rect 32781 30753 32815 30787
rect 32815 30753 32824 30787
rect 32772 30744 32824 30753
rect 34704 30787 34756 30796
rect 34704 30753 34713 30787
rect 34713 30753 34747 30787
rect 34747 30753 34756 30787
rect 34704 30744 34756 30753
rect 36176 30744 36228 30796
rect 36360 30744 36412 30796
rect 27620 30719 27672 30728
rect 27620 30685 27665 30719
rect 27665 30685 27672 30719
rect 27620 30676 27672 30685
rect 28080 30676 28132 30728
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 25228 30608 25280 30660
rect 20444 30540 20496 30592
rect 21456 30583 21508 30592
rect 21456 30549 21465 30583
rect 21465 30549 21499 30583
rect 21499 30549 21508 30583
rect 21456 30540 21508 30549
rect 21732 30540 21784 30592
rect 21824 30583 21876 30592
rect 21824 30549 21833 30583
rect 21833 30549 21867 30583
rect 21867 30549 21876 30583
rect 21824 30540 21876 30549
rect 22376 30540 22428 30592
rect 24124 30540 24176 30592
rect 25964 30540 26016 30592
rect 27160 30583 27212 30592
rect 27160 30549 27169 30583
rect 27169 30549 27203 30583
rect 27203 30549 27212 30583
rect 27160 30540 27212 30549
rect 28356 30540 28408 30592
rect 29184 30651 29236 30660
rect 29184 30617 29193 30651
rect 29193 30617 29227 30651
rect 29227 30617 29236 30651
rect 29184 30608 29236 30617
rect 29092 30583 29144 30592
rect 29092 30549 29101 30583
rect 29101 30549 29135 30583
rect 29135 30549 29144 30583
rect 29092 30540 29144 30549
rect 29736 30676 29788 30728
rect 30380 30676 30432 30728
rect 30564 30719 30616 30728
rect 30564 30685 30573 30719
rect 30573 30685 30607 30719
rect 30607 30685 30616 30719
rect 30564 30676 30616 30685
rect 33784 30608 33836 30660
rect 34336 30608 34388 30660
rect 31576 30540 31628 30592
rect 36636 30540 36688 30592
rect 37004 30719 37056 30728
rect 37004 30685 37013 30719
rect 37013 30685 37047 30719
rect 37047 30685 37056 30719
rect 37004 30676 37056 30685
rect 37648 30787 37700 30796
rect 37648 30753 37657 30787
rect 37657 30753 37691 30787
rect 37691 30753 37700 30787
rect 37648 30744 37700 30753
rect 40408 30787 40460 30796
rect 40408 30753 40417 30787
rect 40417 30753 40451 30787
rect 40451 30753 40460 30787
rect 40408 30744 40460 30753
rect 37372 30719 37424 30728
rect 37372 30685 37381 30719
rect 37381 30685 37415 30719
rect 37415 30685 37424 30719
rect 37372 30676 37424 30685
rect 36912 30651 36964 30660
rect 36912 30617 36921 30651
rect 36921 30617 36955 30651
rect 36955 30617 36964 30651
rect 36912 30608 36964 30617
rect 38936 30608 38988 30660
rect 37924 30540 37976 30592
rect 38292 30540 38344 30592
rect 40868 30719 40920 30728
rect 40868 30685 40877 30719
rect 40877 30685 40911 30719
rect 40911 30685 40920 30719
rect 40868 30676 40920 30685
rect 40040 30608 40092 30660
rect 39672 30540 39724 30592
rect 40316 30540 40368 30592
rect 40592 30540 40644 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 3148 30336 3200 30388
rect 3240 30379 3292 30388
rect 3240 30345 3249 30379
rect 3249 30345 3283 30379
rect 3283 30345 3292 30379
rect 3240 30336 3292 30345
rect 4068 30336 4120 30388
rect 2872 30311 2924 30320
rect 2872 30277 2881 30311
rect 2881 30277 2915 30311
rect 2915 30277 2924 30311
rect 2872 30268 2924 30277
rect 2964 30200 3016 30252
rect 3332 30200 3384 30252
rect 3792 30311 3844 30320
rect 3792 30277 3801 30311
rect 3801 30277 3835 30311
rect 3835 30277 3844 30311
rect 3792 30268 3844 30277
rect 5632 30336 5684 30388
rect 6092 30336 6144 30388
rect 6920 30336 6972 30388
rect 3700 30064 3752 30116
rect 3792 30039 3844 30048
rect 3792 30005 3801 30039
rect 3801 30005 3835 30039
rect 3835 30005 3844 30039
rect 3792 29996 3844 30005
rect 4068 30200 4120 30252
rect 4252 30243 4304 30252
rect 4252 30209 4261 30243
rect 4261 30209 4295 30243
rect 4295 30209 4304 30243
rect 4252 30200 4304 30209
rect 4436 30243 4488 30252
rect 4436 30209 4445 30243
rect 4445 30209 4479 30243
rect 4479 30209 4488 30243
rect 4436 30200 4488 30209
rect 4528 30243 4580 30252
rect 4528 30209 4537 30243
rect 4537 30209 4571 30243
rect 4571 30209 4580 30243
rect 4528 30200 4580 30209
rect 4712 30243 4764 30252
rect 4712 30209 4721 30243
rect 4721 30209 4755 30243
rect 4755 30209 4764 30243
rect 4712 30200 4764 30209
rect 6276 30268 6328 30320
rect 6552 30268 6604 30320
rect 4896 30243 4948 30252
rect 4896 30209 4905 30243
rect 4905 30209 4939 30243
rect 4939 30209 4948 30243
rect 4896 30200 4948 30209
rect 10140 30311 10192 30320
rect 10140 30277 10149 30311
rect 10149 30277 10183 30311
rect 10183 30277 10192 30311
rect 10140 30268 10192 30277
rect 11152 30336 11204 30388
rect 15292 30336 15344 30388
rect 15660 30336 15712 30388
rect 10416 30243 10468 30252
rect 10416 30209 10425 30243
rect 10425 30209 10459 30243
rect 10459 30209 10468 30243
rect 10416 30200 10468 30209
rect 4252 30064 4304 30116
rect 7840 30175 7892 30184
rect 7840 30141 7849 30175
rect 7849 30141 7883 30175
rect 7883 30141 7892 30175
rect 7840 30132 7892 30141
rect 9036 30132 9088 30184
rect 10692 30200 10744 30252
rect 10968 30200 11020 30252
rect 12716 30268 12768 30320
rect 15752 30268 15804 30320
rect 16488 30268 16540 30320
rect 17776 30336 17828 30388
rect 18696 30379 18748 30388
rect 18696 30345 18705 30379
rect 18705 30345 18739 30379
rect 18739 30345 18748 30379
rect 18696 30336 18748 30345
rect 20168 30336 20220 30388
rect 20536 30336 20588 30388
rect 20720 30336 20772 30388
rect 17040 30268 17092 30320
rect 17408 30268 17460 30320
rect 10600 30132 10652 30184
rect 11152 30132 11204 30184
rect 14832 30243 14884 30252
rect 14832 30209 14841 30243
rect 14841 30209 14875 30243
rect 14875 30209 14884 30243
rect 14832 30200 14884 30209
rect 15016 30243 15068 30252
rect 15016 30209 15025 30243
rect 15025 30209 15059 30243
rect 15059 30209 15068 30243
rect 15016 30200 15068 30209
rect 15200 30243 15252 30252
rect 15200 30209 15209 30243
rect 15209 30209 15243 30243
rect 15243 30209 15252 30243
rect 15200 30200 15252 30209
rect 15292 30243 15344 30252
rect 15292 30209 15301 30243
rect 15301 30209 15335 30243
rect 15335 30209 15344 30243
rect 15292 30200 15344 30209
rect 12256 30132 12308 30184
rect 5632 30064 5684 30116
rect 10876 30064 10928 30116
rect 12992 30175 13044 30184
rect 12992 30141 13001 30175
rect 13001 30141 13035 30175
rect 13035 30141 13044 30175
rect 12992 30132 13044 30141
rect 14924 30132 14976 30184
rect 15476 30175 15528 30184
rect 15476 30141 15485 30175
rect 15485 30141 15519 30175
rect 15519 30141 15528 30175
rect 15476 30132 15528 30141
rect 15936 30243 15988 30252
rect 15936 30209 15945 30243
rect 15945 30209 15979 30243
rect 15979 30209 15988 30243
rect 15936 30200 15988 30209
rect 16120 30243 16172 30252
rect 16120 30209 16129 30243
rect 16129 30209 16163 30243
rect 16163 30209 16172 30243
rect 16120 30200 16172 30209
rect 17040 30132 17092 30184
rect 17408 30132 17460 30184
rect 15568 30064 15620 30116
rect 17960 30268 18012 30320
rect 18236 30243 18288 30252
rect 18236 30209 18245 30243
rect 18245 30209 18279 30243
rect 18279 30209 18288 30243
rect 18236 30200 18288 30209
rect 19616 30268 19668 30320
rect 18512 30132 18564 30184
rect 18972 30175 19024 30184
rect 18972 30141 18981 30175
rect 18981 30141 19015 30175
rect 19015 30141 19024 30175
rect 20628 30200 20680 30252
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 22100 30336 22152 30388
rect 22376 30336 22428 30388
rect 22652 30336 22704 30388
rect 21732 30268 21784 30320
rect 18972 30132 19024 30141
rect 19800 30132 19852 30184
rect 3976 29996 4028 30048
rect 4068 29996 4120 30048
rect 4528 29996 4580 30048
rect 5356 29996 5408 30048
rect 5540 29996 5592 30048
rect 9312 29996 9364 30048
rect 15292 29996 15344 30048
rect 16304 29996 16356 30048
rect 16948 29996 17000 30048
rect 20260 30064 20312 30116
rect 17960 29996 18012 30048
rect 18604 30039 18656 30048
rect 18604 30005 18613 30039
rect 18613 30005 18647 30039
rect 18647 30005 18656 30039
rect 18604 29996 18656 30005
rect 21180 30064 21232 30116
rect 21824 30243 21876 30252
rect 21824 30209 21833 30243
rect 21833 30209 21867 30243
rect 21867 30209 21876 30243
rect 21824 30200 21876 30209
rect 22836 30268 22888 30320
rect 21916 30132 21968 30184
rect 22008 30064 22060 30116
rect 22376 30200 22428 30252
rect 24584 30336 24636 30388
rect 25596 30336 25648 30388
rect 30564 30336 30616 30388
rect 30840 30379 30892 30388
rect 30840 30345 30849 30379
rect 30849 30345 30883 30379
rect 30883 30345 30892 30379
rect 30840 30336 30892 30345
rect 34796 30336 34848 30388
rect 24676 30268 24728 30320
rect 23940 30200 23992 30252
rect 26884 30268 26936 30320
rect 28816 30311 28868 30320
rect 28816 30277 28825 30311
rect 28825 30277 28859 30311
rect 28859 30277 28868 30311
rect 28816 30268 28868 30277
rect 30104 30311 30156 30320
rect 30104 30277 30113 30311
rect 30113 30277 30147 30311
rect 30147 30277 30156 30311
rect 30104 30268 30156 30277
rect 25780 30243 25832 30252
rect 25780 30209 25789 30243
rect 25789 30209 25823 30243
rect 25823 30209 25832 30243
rect 25780 30200 25832 30209
rect 25964 30243 26016 30252
rect 25964 30209 25973 30243
rect 25973 30209 26007 30243
rect 26007 30209 26016 30243
rect 25964 30200 26016 30209
rect 26240 30243 26292 30252
rect 26240 30209 26249 30243
rect 26249 30209 26283 30243
rect 26283 30209 26292 30243
rect 26240 30200 26292 30209
rect 28356 30200 28408 30252
rect 28632 30200 28684 30252
rect 29552 30243 29604 30252
rect 29552 30209 29561 30243
rect 29561 30209 29595 30243
rect 29595 30209 29604 30243
rect 29552 30200 29604 30209
rect 29736 30200 29788 30252
rect 29828 30200 29880 30252
rect 32496 30268 32548 30320
rect 22192 30064 22244 30116
rect 24308 30132 24360 30184
rect 26792 30175 26844 30184
rect 26792 30141 26801 30175
rect 26801 30141 26835 30175
rect 26835 30141 26844 30175
rect 26792 30132 26844 30141
rect 26976 30175 27028 30184
rect 26976 30141 26985 30175
rect 26985 30141 27019 30175
rect 27019 30141 27028 30175
rect 26976 30132 27028 30141
rect 24952 30064 25004 30116
rect 26608 30107 26660 30116
rect 26608 30073 26617 30107
rect 26617 30073 26651 30107
rect 26651 30073 26660 30107
rect 26608 30064 26660 30073
rect 30196 30132 30248 30184
rect 30748 30243 30800 30252
rect 30748 30209 30757 30243
rect 30757 30209 30791 30243
rect 30791 30209 30800 30243
rect 30748 30200 30800 30209
rect 31484 30200 31536 30252
rect 31576 30243 31628 30252
rect 31576 30209 31585 30243
rect 31585 30209 31619 30243
rect 31619 30209 31628 30243
rect 31576 30200 31628 30209
rect 31668 30243 31720 30252
rect 31668 30209 31677 30243
rect 31677 30209 31711 30243
rect 31711 30209 31720 30243
rect 31668 30200 31720 30209
rect 34060 30311 34112 30320
rect 34060 30277 34069 30311
rect 34069 30277 34103 30311
rect 34103 30277 34112 30311
rect 34060 30268 34112 30277
rect 36268 30379 36320 30388
rect 36268 30345 36277 30379
rect 36277 30345 36311 30379
rect 36311 30345 36320 30379
rect 36268 30336 36320 30345
rect 35992 30268 36044 30320
rect 36912 30336 36964 30388
rect 37832 30379 37884 30388
rect 37832 30345 37841 30379
rect 37841 30345 37875 30379
rect 37875 30345 37884 30379
rect 37832 30336 37884 30345
rect 37924 30336 37976 30388
rect 38568 30336 38620 30388
rect 37648 30311 37700 30320
rect 37648 30277 37657 30311
rect 37657 30277 37691 30311
rect 37691 30277 37700 30311
rect 37648 30268 37700 30277
rect 38844 30268 38896 30320
rect 39580 30268 39632 30320
rect 40132 30268 40184 30320
rect 35624 30243 35676 30252
rect 30380 30132 30432 30184
rect 29460 30064 29512 30116
rect 22652 29996 22704 30048
rect 22744 30039 22796 30048
rect 22744 30005 22753 30039
rect 22753 30005 22787 30039
rect 22787 30005 22796 30039
rect 22744 29996 22796 30005
rect 23756 29996 23808 30048
rect 27068 29996 27120 30048
rect 27712 29996 27764 30048
rect 30288 30039 30340 30048
rect 30288 30005 30297 30039
rect 30297 30005 30331 30039
rect 30331 30005 30340 30039
rect 30288 29996 30340 30005
rect 30840 30064 30892 30116
rect 32220 30175 32272 30184
rect 32220 30141 32229 30175
rect 32229 30141 32263 30175
rect 32263 30141 32272 30175
rect 32220 30132 32272 30141
rect 33416 30132 33468 30184
rect 34152 30132 34204 30184
rect 34336 30132 34388 30184
rect 31024 29996 31076 30048
rect 31484 29996 31536 30048
rect 34244 30064 34296 30116
rect 34428 30107 34480 30116
rect 34428 30073 34437 30107
rect 34437 30073 34471 30107
rect 34471 30073 34480 30107
rect 34428 30064 34480 30073
rect 34796 30175 34848 30184
rect 34796 30141 34805 30175
rect 34805 30141 34839 30175
rect 34839 30141 34848 30175
rect 34796 30132 34848 30141
rect 34888 30175 34940 30184
rect 34888 30141 34897 30175
rect 34897 30141 34931 30175
rect 34931 30141 34940 30175
rect 34888 30132 34940 30141
rect 35624 30209 35633 30243
rect 35633 30209 35667 30243
rect 35667 30209 35676 30243
rect 35624 30200 35676 30209
rect 35532 30132 35584 30184
rect 36360 30200 36412 30252
rect 36544 30243 36596 30252
rect 36544 30209 36553 30243
rect 36553 30209 36587 30243
rect 36587 30209 36596 30243
rect 36544 30200 36596 30209
rect 36728 30243 36780 30252
rect 36728 30209 36773 30243
rect 36773 30209 36780 30243
rect 36728 30200 36780 30209
rect 33876 30039 33928 30048
rect 33876 30005 33885 30039
rect 33885 30005 33919 30039
rect 33919 30005 33928 30039
rect 33876 29996 33928 30005
rect 35164 30107 35216 30116
rect 35164 30073 35173 30107
rect 35173 30073 35207 30107
rect 35207 30073 35216 30107
rect 35164 30064 35216 30073
rect 35900 30132 35952 30184
rect 36084 30132 36136 30184
rect 36176 30132 36228 30184
rect 38108 30243 38160 30252
rect 38108 30209 38117 30243
rect 38117 30209 38151 30243
rect 38151 30209 38160 30243
rect 38108 30200 38160 30209
rect 37832 30132 37884 30184
rect 38568 30200 38620 30252
rect 39212 30243 39264 30252
rect 39212 30209 39221 30243
rect 39221 30209 39255 30243
rect 39255 30209 39264 30243
rect 39212 30200 39264 30209
rect 38384 30064 38436 30116
rect 39672 30200 39724 30252
rect 40224 30200 40276 30252
rect 40500 30243 40552 30252
rect 40500 30209 40509 30243
rect 40509 30209 40543 30243
rect 40543 30209 40552 30243
rect 40500 30200 40552 30209
rect 40868 30243 40920 30252
rect 40868 30209 40877 30243
rect 40877 30209 40911 30243
rect 40911 30209 40920 30243
rect 40868 30200 40920 30209
rect 41880 30243 41932 30252
rect 41880 30209 41889 30243
rect 41889 30209 41923 30243
rect 41923 30209 41932 30243
rect 41880 30200 41932 30209
rect 40040 30064 40092 30116
rect 40684 29996 40736 30048
rect 42064 30039 42116 30048
rect 42064 30005 42073 30039
rect 42073 30005 42107 30039
rect 42107 30005 42116 30039
rect 42064 29996 42116 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3424 29792 3476 29844
rect 5540 29835 5592 29844
rect 5540 29801 5549 29835
rect 5549 29801 5583 29835
rect 5583 29801 5592 29835
rect 5540 29792 5592 29801
rect 7840 29792 7892 29844
rect 17408 29792 17460 29844
rect 17684 29792 17736 29844
rect 20260 29792 20312 29844
rect 1768 29588 1820 29640
rect 2688 29631 2740 29640
rect 2688 29597 2697 29631
rect 2697 29597 2731 29631
rect 2731 29597 2740 29631
rect 2688 29588 2740 29597
rect 2872 29631 2924 29640
rect 2872 29597 2881 29631
rect 2881 29597 2915 29631
rect 2915 29597 2924 29631
rect 2872 29588 2924 29597
rect 3516 29724 3568 29776
rect 3976 29724 4028 29776
rect 3240 29631 3292 29640
rect 3240 29597 3249 29631
rect 3249 29597 3283 29631
rect 3283 29597 3292 29631
rect 3240 29588 3292 29597
rect 3792 29656 3844 29708
rect 3608 29631 3660 29640
rect 3608 29597 3617 29631
rect 3617 29597 3651 29631
rect 3651 29597 3660 29631
rect 3608 29588 3660 29597
rect 3976 29631 4028 29640
rect 3976 29597 3985 29631
rect 3985 29597 4019 29631
rect 4019 29597 4028 29631
rect 3976 29588 4028 29597
rect 4068 29631 4120 29640
rect 4068 29597 4077 29631
rect 4077 29597 4111 29631
rect 4111 29597 4120 29631
rect 4068 29588 4120 29597
rect 5080 29656 5132 29708
rect 9588 29699 9640 29708
rect 9588 29665 9597 29699
rect 9597 29665 9631 29699
rect 9631 29665 9640 29699
rect 9588 29656 9640 29665
rect 12900 29656 12952 29708
rect 13176 29656 13228 29708
rect 17776 29656 17828 29708
rect 21180 29656 21232 29708
rect 4344 29631 4396 29640
rect 4344 29597 4353 29631
rect 4353 29597 4387 29631
rect 4387 29597 4396 29631
rect 4344 29588 4396 29597
rect 5356 29631 5408 29640
rect 5356 29597 5365 29631
rect 5365 29597 5399 29631
rect 5399 29597 5408 29631
rect 5356 29588 5408 29597
rect 9312 29631 9364 29640
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 10232 29588 10284 29640
rect 11060 29588 11112 29640
rect 2964 29495 3016 29504
rect 2964 29461 2973 29495
rect 2973 29461 3007 29495
rect 3007 29461 3016 29495
rect 2964 29452 3016 29461
rect 4252 29520 4304 29572
rect 8668 29520 8720 29572
rect 12716 29563 12768 29572
rect 12716 29529 12725 29563
rect 12725 29529 12759 29563
rect 12759 29529 12768 29563
rect 12716 29520 12768 29529
rect 20628 29588 20680 29640
rect 22008 29724 22060 29776
rect 22744 29792 22796 29844
rect 24860 29792 24912 29844
rect 26884 29835 26936 29844
rect 26884 29801 26893 29835
rect 26893 29801 26927 29835
rect 26927 29801 26936 29835
rect 26884 29792 26936 29801
rect 28908 29792 28960 29844
rect 30748 29792 30800 29844
rect 31668 29792 31720 29844
rect 34612 29792 34664 29844
rect 34980 29792 35032 29844
rect 22836 29724 22888 29776
rect 21824 29656 21876 29708
rect 21732 29631 21784 29640
rect 21732 29597 21741 29631
rect 21741 29597 21775 29631
rect 21775 29597 21784 29631
rect 21732 29588 21784 29597
rect 21916 29631 21968 29640
rect 21916 29597 21925 29631
rect 21925 29597 21959 29631
rect 21959 29597 21968 29631
rect 21916 29588 21968 29597
rect 23020 29656 23072 29708
rect 22744 29631 22796 29640
rect 22744 29597 22753 29631
rect 22753 29597 22787 29631
rect 22787 29597 22796 29631
rect 22744 29588 22796 29597
rect 3608 29452 3660 29504
rect 4068 29452 4120 29504
rect 8024 29495 8076 29504
rect 8024 29461 8033 29495
rect 8033 29461 8067 29495
rect 8067 29461 8076 29495
rect 8024 29452 8076 29461
rect 8484 29495 8536 29504
rect 8484 29461 8493 29495
rect 8493 29461 8527 29495
rect 8527 29461 8536 29495
rect 8484 29452 8536 29461
rect 8944 29495 8996 29504
rect 8944 29461 8953 29495
rect 8953 29461 8987 29495
rect 8987 29461 8996 29495
rect 8944 29452 8996 29461
rect 9404 29495 9456 29504
rect 9404 29461 9413 29495
rect 9413 29461 9447 29495
rect 9447 29461 9456 29495
rect 9404 29452 9456 29461
rect 9772 29495 9824 29504
rect 9772 29461 9781 29495
rect 9781 29461 9815 29495
rect 9815 29461 9824 29495
rect 9772 29452 9824 29461
rect 10048 29452 10100 29504
rect 12440 29452 12492 29504
rect 18052 29452 18104 29504
rect 20536 29495 20588 29504
rect 20536 29461 20545 29495
rect 20545 29461 20579 29495
rect 20579 29461 20588 29495
rect 20536 29452 20588 29461
rect 20812 29563 20864 29572
rect 20812 29529 20821 29563
rect 20821 29529 20855 29563
rect 20855 29529 20864 29563
rect 20812 29520 20864 29529
rect 20996 29563 21048 29572
rect 20996 29529 21005 29563
rect 21005 29529 21039 29563
rect 21039 29529 21048 29563
rect 20996 29520 21048 29529
rect 21548 29520 21600 29572
rect 22284 29520 22336 29572
rect 23204 29588 23256 29640
rect 23388 29588 23440 29640
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 24124 29520 24176 29572
rect 24676 29520 24728 29572
rect 25964 29724 26016 29776
rect 27804 29724 27856 29776
rect 27988 29724 28040 29776
rect 25780 29656 25832 29708
rect 26608 29656 26660 29708
rect 29460 29724 29512 29776
rect 25596 29588 25648 29640
rect 27068 29631 27120 29640
rect 27068 29597 27077 29631
rect 27077 29597 27111 29631
rect 27111 29597 27120 29631
rect 27068 29588 27120 29597
rect 27160 29631 27212 29640
rect 27160 29597 27169 29631
rect 27169 29597 27203 29631
rect 27203 29597 27212 29631
rect 27160 29588 27212 29597
rect 21180 29452 21232 29504
rect 23204 29452 23256 29504
rect 24400 29452 24452 29504
rect 25780 29452 25832 29504
rect 26240 29520 26292 29572
rect 27712 29588 27764 29640
rect 29000 29656 29052 29708
rect 29644 29699 29696 29708
rect 29644 29665 29653 29699
rect 29653 29665 29687 29699
rect 29687 29665 29696 29699
rect 29644 29656 29696 29665
rect 29000 29520 29052 29572
rect 29368 29631 29420 29640
rect 29368 29597 29377 29631
rect 29377 29597 29411 29631
rect 29411 29597 29420 29631
rect 29368 29588 29420 29597
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 30196 29588 30248 29640
rect 30288 29631 30340 29640
rect 30288 29597 30297 29631
rect 30297 29597 30331 29631
rect 30331 29597 30340 29631
rect 32496 29724 32548 29776
rect 31484 29699 31536 29708
rect 31484 29665 31493 29699
rect 31493 29665 31527 29699
rect 31527 29665 31536 29699
rect 31484 29656 31536 29665
rect 30288 29588 30340 29597
rect 30656 29588 30708 29640
rect 31116 29588 31168 29640
rect 35348 29724 35400 29776
rect 35532 29792 35584 29844
rect 37280 29792 37332 29844
rect 38108 29792 38160 29844
rect 38292 29792 38344 29844
rect 40408 29792 40460 29844
rect 41880 29792 41932 29844
rect 33416 29656 33468 29708
rect 33600 29631 33652 29640
rect 33600 29597 33608 29631
rect 33608 29597 33642 29631
rect 33642 29597 33652 29631
rect 33600 29588 33652 29597
rect 34888 29656 34940 29708
rect 34704 29588 34756 29640
rect 35072 29631 35124 29640
rect 35072 29597 35081 29631
rect 35081 29597 35115 29631
rect 35115 29597 35124 29631
rect 35072 29588 35124 29597
rect 35532 29656 35584 29708
rect 35808 29588 35860 29640
rect 35992 29656 36044 29708
rect 36544 29724 36596 29776
rect 37096 29724 37148 29776
rect 37648 29699 37700 29708
rect 37648 29665 37657 29699
rect 37657 29665 37691 29699
rect 37691 29665 37700 29699
rect 37648 29656 37700 29665
rect 27712 29452 27764 29504
rect 27896 29495 27948 29504
rect 27896 29461 27905 29495
rect 27905 29461 27939 29495
rect 27939 29461 27948 29495
rect 27896 29452 27948 29461
rect 29460 29452 29512 29504
rect 29736 29452 29788 29504
rect 33048 29520 33100 29572
rect 30564 29452 30616 29504
rect 31024 29452 31076 29504
rect 31760 29452 31812 29504
rect 32956 29452 33008 29504
rect 34152 29520 34204 29572
rect 34888 29520 34940 29572
rect 35992 29520 36044 29572
rect 36452 29588 36504 29640
rect 37280 29588 37332 29640
rect 37832 29631 37884 29640
rect 37832 29597 37841 29631
rect 37841 29597 37875 29631
rect 37875 29597 37884 29631
rect 37832 29588 37884 29597
rect 33232 29452 33284 29504
rect 33600 29452 33652 29504
rect 35440 29452 35492 29504
rect 38200 29631 38252 29640
rect 38200 29597 38209 29631
rect 38209 29597 38243 29631
rect 38243 29597 38252 29631
rect 38200 29588 38252 29597
rect 38384 29631 38436 29640
rect 38384 29597 38393 29631
rect 38393 29597 38427 29631
rect 38427 29597 38436 29631
rect 38384 29588 38436 29597
rect 38660 29656 38712 29708
rect 39304 29656 39356 29708
rect 40684 29699 40736 29708
rect 40684 29665 40693 29699
rect 40693 29665 40727 29699
rect 40727 29665 40736 29699
rect 40684 29656 40736 29665
rect 40224 29588 40276 29640
rect 40408 29631 40460 29640
rect 40408 29597 40417 29631
rect 40417 29597 40451 29631
rect 40451 29597 40460 29631
rect 40408 29588 40460 29597
rect 38844 29520 38896 29572
rect 37188 29452 37240 29504
rect 37924 29452 37976 29504
rect 40040 29563 40092 29572
rect 40040 29529 40049 29563
rect 40049 29529 40083 29563
rect 40083 29529 40092 29563
rect 40040 29520 40092 29529
rect 41420 29520 41472 29572
rect 40224 29495 40276 29504
rect 40224 29461 40233 29495
rect 40233 29461 40267 29495
rect 40267 29461 40276 29495
rect 40224 29452 40276 29461
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 5172 29248 5224 29300
rect 5448 29291 5500 29300
rect 5448 29257 5457 29291
rect 5457 29257 5491 29291
rect 5491 29257 5500 29291
rect 5448 29248 5500 29257
rect 3056 29180 3108 29232
rect 3240 29180 3292 29232
rect 3792 29112 3844 29164
rect 8944 29248 8996 29300
rect 10232 29248 10284 29300
rect 10692 29291 10744 29300
rect 10692 29257 10701 29291
rect 10701 29257 10735 29291
rect 10735 29257 10744 29291
rect 10692 29248 10744 29257
rect 10968 29291 11020 29300
rect 10968 29257 10977 29291
rect 10977 29257 11011 29291
rect 11011 29257 11020 29291
rect 10968 29248 11020 29257
rect 12992 29248 13044 29300
rect 14280 29291 14332 29300
rect 14280 29257 14289 29291
rect 14289 29257 14323 29291
rect 14323 29257 14332 29291
rect 14280 29248 14332 29257
rect 14832 29248 14884 29300
rect 15476 29291 15528 29300
rect 15476 29257 15485 29291
rect 15485 29257 15519 29291
rect 15519 29257 15528 29291
rect 15476 29248 15528 29257
rect 16028 29291 16080 29300
rect 16028 29257 16037 29291
rect 16037 29257 16071 29291
rect 16071 29257 16080 29291
rect 16028 29248 16080 29257
rect 16948 29291 17000 29300
rect 16948 29257 16957 29291
rect 16957 29257 16991 29291
rect 16991 29257 17000 29291
rect 16948 29248 17000 29257
rect 17040 29248 17092 29300
rect 10784 29180 10836 29232
rect 4252 29155 4304 29164
rect 4252 29121 4261 29155
rect 4261 29121 4295 29155
rect 4295 29121 4304 29155
rect 4252 29112 4304 29121
rect 5356 29112 5408 29164
rect 5724 29112 5776 29164
rect 6920 29155 6972 29164
rect 6920 29121 6929 29155
rect 6929 29121 6963 29155
rect 6963 29121 6972 29155
rect 6920 29112 6972 29121
rect 8392 29155 8444 29164
rect 8392 29121 8401 29155
rect 8401 29121 8435 29155
rect 8435 29121 8444 29155
rect 8392 29112 8444 29121
rect 9128 29112 9180 29164
rect 1676 29087 1728 29096
rect 1676 29053 1685 29087
rect 1685 29053 1719 29087
rect 1719 29053 1728 29087
rect 1676 29044 1728 29053
rect 3240 29044 3292 29096
rect 3516 29087 3568 29096
rect 3516 29053 3525 29087
rect 3525 29053 3559 29087
rect 3559 29053 3568 29087
rect 3516 29044 3568 29053
rect 3608 29087 3660 29096
rect 3608 29053 3617 29087
rect 3617 29053 3651 29087
rect 3651 29053 3660 29087
rect 3608 29044 3660 29053
rect 4344 29087 4396 29096
rect 4344 29053 4353 29087
rect 4353 29053 4387 29087
rect 4387 29053 4396 29087
rect 4344 29044 4396 29053
rect 4804 29044 4856 29096
rect 10048 29155 10100 29164
rect 10048 29121 10057 29155
rect 10057 29121 10091 29155
rect 10091 29121 10100 29155
rect 10048 29112 10100 29121
rect 10232 29155 10284 29164
rect 10232 29121 10241 29155
rect 10241 29121 10275 29155
rect 10275 29121 10284 29155
rect 10232 29112 10284 29121
rect 10692 29155 10744 29164
rect 10692 29121 10701 29155
rect 10701 29121 10735 29155
rect 10735 29121 10744 29155
rect 10692 29112 10744 29121
rect 12716 29180 12768 29232
rect 13176 29180 13228 29232
rect 10508 29044 10560 29096
rect 13084 29155 13136 29164
rect 13084 29121 13093 29155
rect 13093 29121 13127 29155
rect 13127 29121 13136 29155
rect 13084 29112 13136 29121
rect 13452 29112 13504 29164
rect 3240 28951 3292 28960
rect 3240 28917 3249 28951
rect 3249 28917 3283 28951
rect 3283 28917 3292 28951
rect 3240 28908 3292 28917
rect 4620 28908 4672 28960
rect 4896 28908 4948 28960
rect 9036 28908 9088 28960
rect 10232 28976 10284 29028
rect 12532 28976 12584 29028
rect 12716 28976 12768 29028
rect 13268 28976 13320 29028
rect 14188 29112 14240 29164
rect 15384 29180 15436 29232
rect 15568 29180 15620 29232
rect 16212 29180 16264 29232
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 17040 29112 17092 29164
rect 17132 29155 17184 29164
rect 17132 29121 17141 29155
rect 17141 29121 17175 29155
rect 17175 29121 17184 29155
rect 17132 29112 17184 29121
rect 17592 29155 17644 29164
rect 17592 29121 17601 29155
rect 17601 29121 17635 29155
rect 17635 29121 17644 29155
rect 17592 29112 17644 29121
rect 15292 29087 15344 29096
rect 15292 29053 15301 29087
rect 15301 29053 15335 29087
rect 15335 29053 15344 29087
rect 15292 29044 15344 29053
rect 15660 29087 15712 29096
rect 15660 29053 15669 29087
rect 15669 29053 15703 29087
rect 15703 29053 15712 29087
rect 15660 29044 15712 29053
rect 17408 29044 17460 29096
rect 17960 29155 18012 29164
rect 17960 29121 17969 29155
rect 17969 29121 18003 29155
rect 18003 29121 18012 29155
rect 17960 29112 18012 29121
rect 18236 29112 18288 29164
rect 19248 29248 19300 29300
rect 23204 29248 23256 29300
rect 21640 29180 21692 29232
rect 22376 29180 22428 29232
rect 22928 29180 22980 29232
rect 24492 29180 24544 29232
rect 20260 29155 20312 29164
rect 20260 29121 20269 29155
rect 20269 29121 20303 29155
rect 20303 29121 20312 29155
rect 20260 29112 20312 29121
rect 20536 29112 20588 29164
rect 21916 29155 21968 29164
rect 21916 29121 21925 29155
rect 21925 29121 21959 29155
rect 21959 29121 21968 29155
rect 21916 29112 21968 29121
rect 18144 29044 18196 29096
rect 18696 29044 18748 29096
rect 18788 29044 18840 29096
rect 23388 29112 23440 29164
rect 24308 29112 24360 29164
rect 25780 29155 25832 29164
rect 25780 29121 25789 29155
rect 25789 29121 25823 29155
rect 25823 29121 25832 29155
rect 25780 29112 25832 29121
rect 26792 29248 26844 29300
rect 28448 29248 28500 29300
rect 32496 29248 32548 29300
rect 32864 29248 32916 29300
rect 29184 29180 29236 29232
rect 30932 29180 30984 29232
rect 26424 29112 26476 29164
rect 27528 29112 27580 29164
rect 23480 29044 23532 29096
rect 21180 28976 21232 29028
rect 24584 28976 24636 29028
rect 24676 28976 24728 29028
rect 10324 28951 10376 28960
rect 10324 28917 10333 28951
rect 10333 28917 10367 28951
rect 10367 28917 10376 28951
rect 10324 28908 10376 28917
rect 10600 28951 10652 28960
rect 10600 28917 10609 28951
rect 10609 28917 10643 28951
rect 10643 28917 10652 28951
rect 10600 28908 10652 28917
rect 13636 28951 13688 28960
rect 13636 28917 13645 28951
rect 13645 28917 13679 28951
rect 13679 28917 13688 28951
rect 13636 28908 13688 28917
rect 13728 28951 13780 28960
rect 13728 28917 13737 28951
rect 13737 28917 13771 28951
rect 13771 28917 13780 28951
rect 13728 28908 13780 28917
rect 13912 28908 13964 28960
rect 16304 28908 16356 28960
rect 16396 28908 16448 28960
rect 16764 28908 16816 28960
rect 18512 28908 18564 28960
rect 21088 28908 21140 28960
rect 22008 28908 22060 28960
rect 25228 28908 25280 28960
rect 25320 28908 25372 28960
rect 27620 28976 27672 29028
rect 27804 29155 27856 29164
rect 27804 29121 27813 29155
rect 27813 29121 27847 29155
rect 27847 29121 27856 29155
rect 27804 29112 27856 29121
rect 29460 29155 29512 29164
rect 29460 29121 29469 29155
rect 29469 29121 29503 29155
rect 29503 29121 29512 29155
rect 29460 29112 29512 29121
rect 29644 29155 29696 29164
rect 29644 29121 29653 29155
rect 29653 29121 29687 29155
rect 29687 29121 29696 29155
rect 29644 29112 29696 29121
rect 30472 29155 30524 29164
rect 30472 29121 30481 29155
rect 30481 29121 30515 29155
rect 30515 29121 30524 29155
rect 30472 29112 30524 29121
rect 31024 29112 31076 29164
rect 31484 29155 31536 29164
rect 31484 29121 31492 29155
rect 31492 29121 31526 29155
rect 31526 29121 31536 29155
rect 31484 29112 31536 29121
rect 31668 29112 31720 29164
rect 32312 29180 32364 29232
rect 32956 29180 33008 29232
rect 32772 29112 32824 29164
rect 34152 29248 34204 29300
rect 34428 29248 34480 29300
rect 34888 29291 34940 29300
rect 34888 29257 34897 29291
rect 34897 29257 34931 29291
rect 34931 29257 34940 29291
rect 34888 29248 34940 29257
rect 36360 29248 36412 29300
rect 36544 29248 36596 29300
rect 33140 29180 33192 29232
rect 33232 29155 33284 29164
rect 33232 29121 33241 29155
rect 33241 29121 33275 29155
rect 33275 29121 33284 29155
rect 33232 29112 33284 29121
rect 27804 28976 27856 29028
rect 27988 28976 28040 29028
rect 29644 28976 29696 29028
rect 30472 28976 30524 29028
rect 30656 28976 30708 29028
rect 31760 29044 31812 29096
rect 33048 29044 33100 29096
rect 34612 29180 34664 29232
rect 33876 29112 33928 29164
rect 34152 29155 34204 29164
rect 34152 29121 34161 29155
rect 34161 29121 34195 29155
rect 34195 29121 34204 29155
rect 34152 29112 34204 29121
rect 34336 29112 34388 29164
rect 34520 29112 34572 29164
rect 35072 29155 35124 29164
rect 35072 29121 35081 29155
rect 35081 29121 35115 29155
rect 35115 29121 35124 29155
rect 35072 29112 35124 29121
rect 35992 29180 36044 29232
rect 29736 28908 29788 28960
rect 31576 28976 31628 29028
rect 33140 29019 33192 29028
rect 33140 28985 33149 29019
rect 33149 28985 33183 29019
rect 33183 28985 33192 29019
rect 33140 28976 33192 28985
rect 33784 29044 33836 29096
rect 30840 28908 30892 28960
rect 32956 28908 33008 28960
rect 33324 28908 33376 28960
rect 33968 28976 34020 29028
rect 34980 29044 35032 29096
rect 35440 29112 35492 29164
rect 38844 29248 38896 29300
rect 40040 29248 40092 29300
rect 37924 29223 37976 29232
rect 37924 29189 37933 29223
rect 37933 29189 37967 29223
rect 37967 29189 37976 29223
rect 37924 29180 37976 29189
rect 39212 29223 39264 29232
rect 37556 29155 37608 29164
rect 37556 29121 37565 29155
rect 37565 29121 37599 29155
rect 37599 29121 37608 29155
rect 37556 29112 37608 29121
rect 38108 29146 38160 29198
rect 34244 28976 34296 29028
rect 37188 29044 37240 29096
rect 37832 29044 37884 29096
rect 36360 28976 36412 29028
rect 37740 28976 37792 29028
rect 38108 29044 38160 29096
rect 39212 29189 39221 29223
rect 39221 29189 39255 29223
rect 39255 29189 39264 29223
rect 39212 29180 39264 29189
rect 39856 29180 39908 29232
rect 40224 29180 40276 29232
rect 41972 29180 42024 29232
rect 39120 29112 39172 29164
rect 39580 29112 39632 29164
rect 39028 28976 39080 29028
rect 34428 28908 34480 28960
rect 35716 28908 35768 28960
rect 36912 28908 36964 28960
rect 37648 28908 37700 28960
rect 39948 29044 40000 29096
rect 42064 29019 42116 29028
rect 42064 28985 42073 29019
rect 42073 28985 42107 29019
rect 42107 28985 42116 29019
rect 42064 28976 42116 28985
rect 40408 28908 40460 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1676 28704 1728 28756
rect 3240 28704 3292 28756
rect 5264 28704 5316 28756
rect 7104 28704 7156 28756
rect 9128 28747 9180 28756
rect 9128 28713 9137 28747
rect 9137 28713 9171 28747
rect 9171 28713 9180 28747
rect 9128 28704 9180 28713
rect 9680 28704 9732 28756
rect 12808 28704 12860 28756
rect 13636 28704 13688 28756
rect 16580 28704 16632 28756
rect 3516 28636 3568 28688
rect 2964 28500 3016 28552
rect 3056 28543 3108 28552
rect 3056 28509 3065 28543
rect 3065 28509 3099 28543
rect 3099 28509 3108 28543
rect 3056 28500 3108 28509
rect 17040 28704 17092 28756
rect 10324 28636 10376 28688
rect 4620 28568 4672 28620
rect 5172 28611 5224 28620
rect 5172 28577 5181 28611
rect 5181 28577 5215 28611
rect 5215 28577 5224 28611
rect 5172 28568 5224 28577
rect 9588 28568 9640 28620
rect 3884 28432 3936 28484
rect 4344 28475 4396 28484
rect 4344 28441 4353 28475
rect 4353 28441 4387 28475
rect 4387 28441 4396 28475
rect 4344 28432 4396 28441
rect 4896 28543 4948 28552
rect 4896 28509 4905 28543
rect 4905 28509 4939 28543
rect 4939 28509 4948 28543
rect 4896 28500 4948 28509
rect 6552 28500 6604 28552
rect 8392 28500 8444 28552
rect 9772 28500 9824 28552
rect 10048 28500 10100 28552
rect 10140 28543 10192 28552
rect 10140 28509 10149 28543
rect 10149 28509 10183 28543
rect 10183 28509 10192 28543
rect 10140 28500 10192 28509
rect 5540 28432 5592 28484
rect 8024 28432 8076 28484
rect 5724 28364 5776 28416
rect 10600 28568 10652 28620
rect 12532 28636 12584 28688
rect 13728 28636 13780 28688
rect 16212 28636 16264 28688
rect 16488 28636 16540 28688
rect 16764 28679 16816 28688
rect 16764 28645 16773 28679
rect 16773 28645 16807 28679
rect 16807 28645 16816 28679
rect 16764 28636 16816 28645
rect 16948 28636 17000 28688
rect 17132 28636 17184 28688
rect 17868 28704 17920 28756
rect 18696 28704 18748 28756
rect 20996 28747 21048 28756
rect 20996 28713 21005 28747
rect 21005 28713 21039 28747
rect 21039 28713 21048 28747
rect 20996 28704 21048 28713
rect 22468 28704 22520 28756
rect 25504 28704 25556 28756
rect 30656 28704 30708 28756
rect 32772 28704 32824 28756
rect 33048 28704 33100 28756
rect 33508 28704 33560 28756
rect 34520 28747 34572 28756
rect 34520 28713 34529 28747
rect 34529 28713 34563 28747
rect 34563 28713 34572 28747
rect 34520 28704 34572 28713
rect 34704 28704 34756 28756
rect 35440 28704 35492 28756
rect 36176 28704 36228 28756
rect 37740 28704 37792 28756
rect 11612 28543 11664 28552
rect 11612 28509 11621 28543
rect 11621 28509 11655 28543
rect 11655 28509 11664 28543
rect 11612 28500 11664 28509
rect 16672 28611 16724 28620
rect 12072 28500 12124 28552
rect 12256 28543 12308 28552
rect 12256 28509 12265 28543
rect 12265 28509 12299 28543
rect 12299 28509 12308 28543
rect 12256 28500 12308 28509
rect 12532 28500 12584 28552
rect 12716 28543 12768 28552
rect 12716 28509 12725 28543
rect 12725 28509 12759 28543
rect 12759 28509 12768 28543
rect 12716 28500 12768 28509
rect 13268 28500 13320 28552
rect 13544 28500 13596 28552
rect 14096 28543 14148 28552
rect 14096 28509 14105 28543
rect 14105 28509 14139 28543
rect 14139 28509 14148 28543
rect 14096 28500 14148 28509
rect 10968 28364 11020 28416
rect 11520 28364 11572 28416
rect 12992 28432 13044 28484
rect 13084 28475 13136 28484
rect 13084 28441 13093 28475
rect 13093 28441 13127 28475
rect 13127 28441 13136 28475
rect 13084 28432 13136 28441
rect 13176 28475 13228 28484
rect 13176 28441 13185 28475
rect 13185 28441 13219 28475
rect 13219 28441 13228 28475
rect 13176 28432 13228 28441
rect 11980 28364 12032 28416
rect 12256 28364 12308 28416
rect 12532 28407 12584 28416
rect 12532 28373 12541 28407
rect 12541 28373 12575 28407
rect 12575 28373 12584 28407
rect 12532 28364 12584 28373
rect 12900 28364 12952 28416
rect 13820 28432 13872 28484
rect 14464 28432 14516 28484
rect 13360 28364 13412 28416
rect 13912 28364 13964 28416
rect 15200 28364 15252 28416
rect 15752 28432 15804 28484
rect 15936 28364 15988 28416
rect 16672 28577 16681 28611
rect 16681 28577 16715 28611
rect 16715 28577 16724 28611
rect 18788 28679 18840 28688
rect 18788 28645 18797 28679
rect 18797 28645 18831 28679
rect 18831 28645 18840 28679
rect 18788 28636 18840 28645
rect 24860 28636 24912 28688
rect 16672 28568 16724 28577
rect 16212 28543 16264 28552
rect 16212 28509 16221 28543
rect 16221 28509 16255 28543
rect 16255 28509 16264 28543
rect 16212 28500 16264 28509
rect 16304 28432 16356 28484
rect 17684 28500 17736 28552
rect 18236 28543 18288 28552
rect 18236 28509 18245 28543
rect 18245 28509 18279 28543
rect 18279 28509 18288 28543
rect 18236 28500 18288 28509
rect 18880 28568 18932 28620
rect 22836 28568 22888 28620
rect 18604 28500 18656 28552
rect 18788 28543 18840 28552
rect 18788 28509 18797 28543
rect 18797 28509 18831 28543
rect 18831 28509 18840 28543
rect 18788 28500 18840 28509
rect 21180 28543 21232 28552
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 21640 28500 21692 28552
rect 21916 28543 21968 28552
rect 21916 28509 21925 28543
rect 21925 28509 21959 28543
rect 21959 28509 21968 28543
rect 21916 28500 21968 28509
rect 22008 28543 22060 28552
rect 22008 28509 22017 28543
rect 22017 28509 22051 28543
rect 22051 28509 22060 28543
rect 22008 28500 22060 28509
rect 17500 28432 17552 28484
rect 18052 28432 18104 28484
rect 19432 28432 19484 28484
rect 19984 28432 20036 28484
rect 22468 28500 22520 28552
rect 25228 28568 25280 28620
rect 24952 28500 25004 28552
rect 25320 28543 25372 28552
rect 25320 28509 25329 28543
rect 25329 28509 25363 28543
rect 25363 28509 25372 28543
rect 25320 28500 25372 28509
rect 22560 28432 22612 28484
rect 24768 28432 24820 28484
rect 25688 28543 25740 28552
rect 25688 28509 25697 28543
rect 25697 28509 25731 28543
rect 25731 28509 25740 28543
rect 25688 28500 25740 28509
rect 25964 28543 26016 28552
rect 25964 28509 25968 28543
rect 25968 28509 26002 28543
rect 26002 28509 26016 28543
rect 25964 28500 26016 28509
rect 26056 28543 26108 28552
rect 26056 28509 26065 28543
rect 26065 28509 26099 28543
rect 26099 28509 26108 28543
rect 26056 28500 26108 28509
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 17592 28364 17644 28373
rect 18512 28364 18564 28416
rect 21916 28364 21968 28416
rect 22284 28364 22336 28416
rect 23020 28364 23072 28416
rect 25228 28364 25280 28416
rect 26332 28543 26384 28552
rect 26332 28509 26340 28543
rect 26340 28509 26374 28543
rect 26374 28509 26384 28543
rect 26332 28500 26384 28509
rect 29368 28679 29420 28688
rect 29368 28645 29377 28679
rect 29377 28645 29411 28679
rect 29411 28645 29420 28679
rect 29368 28636 29420 28645
rect 26976 28568 27028 28620
rect 27344 28500 27396 28552
rect 29736 28543 29788 28552
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 29828 28543 29880 28552
rect 29828 28509 29837 28543
rect 29837 28509 29871 28543
rect 29871 28509 29880 28543
rect 29828 28500 29880 28509
rect 31208 28636 31260 28688
rect 31668 28636 31720 28688
rect 32680 28636 32732 28688
rect 34796 28636 34848 28688
rect 35256 28568 35308 28620
rect 30196 28500 30248 28552
rect 31116 28543 31168 28552
rect 31116 28509 31125 28543
rect 31125 28509 31159 28543
rect 31159 28509 31168 28543
rect 31116 28500 31168 28509
rect 31300 28543 31352 28552
rect 31300 28509 31309 28543
rect 31309 28509 31343 28543
rect 31343 28509 31352 28543
rect 31300 28500 31352 28509
rect 35532 28636 35584 28688
rect 36544 28636 36596 28688
rect 36728 28636 36780 28688
rect 27252 28364 27304 28416
rect 27344 28364 27396 28416
rect 28080 28364 28132 28416
rect 28356 28432 28408 28484
rect 29368 28432 29420 28484
rect 29920 28432 29972 28484
rect 32404 28475 32456 28484
rect 32404 28441 32413 28475
rect 32413 28441 32447 28475
rect 32447 28441 32456 28475
rect 32404 28432 32456 28441
rect 33324 28432 33376 28484
rect 34060 28432 34112 28484
rect 29276 28364 29328 28416
rect 30748 28364 30800 28416
rect 31024 28364 31076 28416
rect 31668 28364 31720 28416
rect 33416 28364 33468 28416
rect 35440 28543 35492 28552
rect 35440 28509 35449 28543
rect 35449 28509 35483 28543
rect 35483 28509 35492 28543
rect 35440 28500 35492 28509
rect 35072 28475 35124 28484
rect 35072 28441 35081 28475
rect 35081 28441 35115 28475
rect 35115 28441 35124 28475
rect 35072 28432 35124 28441
rect 35164 28475 35216 28484
rect 35164 28441 35173 28475
rect 35173 28441 35207 28475
rect 35207 28441 35216 28475
rect 35164 28432 35216 28441
rect 35440 28364 35492 28416
rect 35716 28543 35768 28552
rect 35716 28509 35725 28543
rect 35725 28509 35759 28543
rect 35759 28509 35768 28543
rect 35716 28500 35768 28509
rect 35808 28543 35860 28552
rect 35808 28509 35817 28543
rect 35817 28509 35851 28543
rect 35851 28509 35860 28543
rect 35808 28500 35860 28509
rect 35992 28364 36044 28416
rect 36176 28407 36228 28416
rect 36176 28373 36185 28407
rect 36185 28373 36219 28407
rect 36219 28373 36228 28407
rect 36176 28364 36228 28373
rect 36360 28543 36412 28552
rect 36360 28509 36369 28543
rect 36369 28509 36403 28543
rect 36403 28509 36412 28543
rect 36360 28500 36412 28509
rect 37372 28611 37424 28620
rect 37372 28577 37381 28611
rect 37381 28577 37415 28611
rect 37415 28577 37424 28611
rect 37372 28568 37424 28577
rect 37648 28611 37700 28620
rect 37648 28577 37657 28611
rect 37657 28577 37691 28611
rect 37691 28577 37700 28611
rect 37648 28568 37700 28577
rect 38844 28568 38896 28620
rect 39120 28568 39172 28620
rect 37004 28500 37056 28552
rect 41420 28500 41472 28552
rect 38936 28432 38988 28484
rect 39580 28432 39632 28484
rect 39856 28432 39908 28484
rect 40500 28475 40552 28484
rect 40500 28441 40509 28475
rect 40509 28441 40543 28475
rect 40543 28441 40552 28475
rect 40500 28432 40552 28441
rect 41880 28543 41932 28552
rect 41880 28509 41889 28543
rect 41889 28509 41923 28543
rect 41923 28509 41932 28543
rect 41880 28500 41932 28509
rect 36360 28364 36412 28416
rect 36728 28364 36780 28416
rect 37740 28364 37792 28416
rect 39120 28407 39172 28416
rect 39120 28373 39129 28407
rect 39129 28373 39163 28407
rect 39163 28373 39172 28407
rect 39120 28364 39172 28373
rect 39764 28364 39816 28416
rect 40684 28407 40736 28416
rect 40684 28373 40693 28407
rect 40693 28373 40727 28407
rect 40727 28373 40736 28407
rect 40684 28364 40736 28373
rect 41696 28407 41748 28416
rect 41696 28373 41705 28407
rect 41705 28373 41739 28407
rect 41739 28373 41748 28407
rect 41696 28364 41748 28373
rect 42064 28407 42116 28416
rect 42064 28373 42073 28407
rect 42073 28373 42107 28407
rect 42107 28373 42116 28407
rect 42064 28364 42116 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 3976 28160 4028 28212
rect 4344 28160 4396 28212
rect 5356 28160 5408 28212
rect 5540 28203 5592 28212
rect 5540 28169 5549 28203
rect 5549 28169 5583 28203
rect 5583 28169 5592 28203
rect 5540 28160 5592 28169
rect 8484 28203 8536 28212
rect 8484 28169 8493 28203
rect 8493 28169 8527 28203
rect 8527 28169 8536 28203
rect 8484 28160 8536 28169
rect 8668 28203 8720 28212
rect 8668 28169 8677 28203
rect 8677 28169 8711 28203
rect 8711 28169 8720 28203
rect 8668 28160 8720 28169
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 11612 28160 11664 28212
rect 3056 28092 3108 28144
rect 3884 28024 3936 28076
rect 5448 28092 5500 28144
rect 5632 28092 5684 28144
rect 7104 28024 7156 28076
rect 9680 28024 9732 28076
rect 11980 28067 12032 28076
rect 11980 28033 11989 28067
rect 11989 28033 12023 28067
rect 12023 28033 12032 28067
rect 11980 28024 12032 28033
rect 12072 28067 12124 28076
rect 12072 28033 12081 28067
rect 12081 28033 12115 28067
rect 12115 28033 12124 28067
rect 12072 28024 12124 28033
rect 4896 27999 4948 28008
rect 4896 27965 4905 27999
rect 4905 27965 4939 27999
rect 4939 27965 4948 27999
rect 4896 27956 4948 27965
rect 5264 27999 5316 28008
rect 5264 27965 5273 27999
rect 5273 27965 5307 27999
rect 5307 27965 5316 27999
rect 5264 27956 5316 27965
rect 5172 27888 5224 27940
rect 5724 27956 5776 28008
rect 8116 27956 8168 28008
rect 10140 27956 10192 28008
rect 12532 28160 12584 28212
rect 12808 28203 12860 28212
rect 12808 28169 12817 28203
rect 12817 28169 12851 28203
rect 12851 28169 12860 28203
rect 12808 28160 12860 28169
rect 12992 28160 13044 28212
rect 12348 28092 12400 28144
rect 12900 28092 12952 28144
rect 12992 28067 13044 28076
rect 12992 28033 12996 28067
rect 12996 28033 13030 28067
rect 13030 28033 13044 28067
rect 12992 28024 13044 28033
rect 13176 28067 13228 28076
rect 13176 28033 13185 28067
rect 13185 28033 13219 28067
rect 13219 28033 13228 28067
rect 13176 28024 13228 28033
rect 13544 28024 13596 28076
rect 13636 28024 13688 28076
rect 13912 28024 13964 28076
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 14556 28024 14608 28076
rect 14924 28135 14976 28144
rect 14924 28101 14933 28135
rect 14933 28101 14967 28135
rect 14967 28101 14976 28135
rect 14924 28092 14976 28101
rect 16488 28160 16540 28212
rect 16580 28160 16632 28212
rect 15844 28092 15896 28144
rect 15936 28092 15988 28144
rect 15200 28067 15252 28076
rect 15200 28033 15209 28067
rect 15209 28033 15243 28067
rect 15243 28033 15252 28067
rect 15200 28024 15252 28033
rect 5264 27820 5316 27872
rect 10048 27888 10100 27940
rect 10692 27888 10744 27940
rect 10508 27820 10560 27872
rect 14372 27956 14424 28008
rect 16120 28024 16172 28076
rect 16304 28067 16356 28076
rect 16304 28033 16313 28067
rect 16313 28033 16347 28067
rect 16347 28033 16356 28067
rect 16304 28024 16356 28033
rect 12716 27931 12768 27940
rect 12716 27897 12725 27931
rect 12725 27897 12759 27931
rect 12759 27897 12768 27931
rect 12716 27888 12768 27897
rect 16212 27956 16264 28008
rect 17132 28024 17184 28076
rect 17408 28067 17460 28076
rect 17408 28033 17417 28067
rect 17417 28033 17451 28067
rect 17451 28033 17460 28067
rect 17408 28024 17460 28033
rect 18236 28092 18288 28144
rect 17684 28067 17736 28076
rect 17684 28033 17693 28067
rect 17693 28033 17727 28067
rect 17727 28033 17736 28067
rect 17684 28024 17736 28033
rect 16488 27956 16540 28008
rect 16304 27888 16356 27940
rect 16764 27888 16816 27940
rect 18052 28067 18104 28076
rect 18052 28033 18061 28067
rect 18061 28033 18095 28067
rect 18095 28033 18104 28067
rect 18052 28024 18104 28033
rect 19432 28203 19484 28212
rect 19432 28169 19441 28203
rect 19441 28169 19475 28203
rect 19475 28169 19484 28203
rect 19432 28160 19484 28169
rect 18788 28092 18840 28144
rect 18604 28067 18656 28076
rect 18604 28033 18613 28067
rect 18613 28033 18647 28067
rect 18647 28033 18656 28067
rect 18604 28024 18656 28033
rect 20812 28092 20864 28144
rect 22836 28160 22888 28212
rect 23388 28160 23440 28212
rect 24768 28203 24820 28212
rect 24768 28169 24777 28203
rect 24777 28169 24811 28203
rect 24811 28169 24820 28203
rect 24768 28160 24820 28169
rect 25136 28160 25188 28212
rect 20996 28067 21048 28076
rect 20996 28033 21005 28067
rect 21005 28033 21039 28067
rect 21039 28033 21048 28067
rect 20996 28024 21048 28033
rect 13912 27820 13964 27872
rect 14648 27863 14700 27872
rect 14648 27829 14657 27863
rect 14657 27829 14691 27863
rect 14691 27829 14700 27863
rect 14648 27820 14700 27829
rect 15752 27863 15804 27872
rect 15752 27829 15761 27863
rect 15761 27829 15795 27863
rect 15795 27829 15804 27863
rect 15752 27820 15804 27829
rect 15844 27820 15896 27872
rect 17592 27820 17644 27872
rect 17776 27863 17828 27872
rect 17776 27829 17785 27863
rect 17785 27829 17819 27863
rect 17819 27829 17828 27863
rect 17776 27820 17828 27829
rect 18236 27888 18288 27940
rect 18512 27820 18564 27872
rect 19248 27820 19300 27872
rect 21364 27956 21416 28008
rect 23848 28092 23900 28144
rect 24124 28067 24176 28076
rect 22100 27999 22152 28008
rect 22100 27965 22109 27999
rect 22109 27965 22143 27999
rect 22143 27965 22152 27999
rect 22100 27956 22152 27965
rect 22560 27956 22612 28008
rect 22836 27956 22888 28008
rect 24124 28033 24133 28067
rect 24133 28033 24167 28067
rect 24167 28033 24176 28067
rect 24124 28024 24176 28033
rect 24400 28135 24452 28144
rect 24400 28101 24409 28135
rect 24409 28101 24443 28135
rect 24443 28101 24452 28135
rect 24400 28092 24452 28101
rect 24584 28135 24636 28144
rect 24584 28101 24593 28135
rect 24593 28101 24627 28135
rect 24627 28101 24636 28135
rect 24584 28092 24636 28101
rect 25228 28135 25280 28144
rect 25228 28101 25237 28135
rect 25237 28101 25271 28135
rect 25271 28101 25280 28135
rect 25228 28092 25280 28101
rect 25596 28160 25648 28212
rect 26056 28160 26108 28212
rect 25688 28092 25740 28144
rect 24768 28024 24820 28076
rect 24952 28067 25004 28076
rect 24952 28033 24961 28067
rect 24961 28033 24995 28067
rect 24995 28033 25004 28067
rect 24952 28024 25004 28033
rect 28356 28160 28408 28212
rect 28908 28160 28960 28212
rect 29368 28160 29420 28212
rect 29828 28160 29880 28212
rect 29276 28135 29328 28144
rect 29276 28101 29285 28135
rect 29285 28101 29319 28135
rect 29319 28101 29328 28135
rect 29276 28092 29328 28101
rect 29644 28092 29696 28144
rect 29920 28135 29972 28144
rect 29920 28101 29929 28135
rect 29929 28101 29963 28135
rect 29963 28101 29972 28135
rect 29920 28092 29972 28101
rect 25688 27956 25740 28008
rect 27620 28067 27672 28076
rect 27620 28033 27629 28067
rect 27629 28033 27663 28067
rect 27663 28033 27672 28067
rect 27620 28024 27672 28033
rect 27804 28067 27856 28076
rect 27804 28033 27813 28067
rect 27813 28033 27847 28067
rect 27847 28033 27856 28067
rect 27804 28024 27856 28033
rect 28080 28024 28132 28076
rect 28816 28024 28868 28076
rect 29276 27956 29328 28008
rect 31116 28160 31168 28212
rect 31300 28160 31352 28212
rect 34520 28160 34572 28212
rect 34796 28160 34848 28212
rect 35348 28160 35400 28212
rect 30104 28092 30156 28144
rect 30932 28092 30984 28144
rect 31944 28024 31996 28076
rect 32588 28092 32640 28144
rect 32680 28092 32732 28144
rect 32772 28067 32824 28076
rect 32772 28033 32781 28067
rect 32781 28033 32815 28067
rect 32815 28033 32824 28067
rect 32772 28024 32824 28033
rect 30472 27999 30524 28008
rect 30472 27965 30481 27999
rect 30481 27965 30515 27999
rect 30515 27965 30524 27999
rect 30472 27956 30524 27965
rect 30932 27956 30984 28008
rect 24308 27931 24360 27940
rect 24308 27897 24317 27931
rect 24317 27897 24351 27931
rect 24351 27897 24360 27931
rect 24308 27888 24360 27897
rect 26332 27888 26384 27940
rect 27804 27888 27856 27940
rect 27988 27888 28040 27940
rect 28356 27888 28408 27940
rect 30104 27888 30156 27940
rect 31668 27956 31720 28008
rect 33048 28067 33100 28076
rect 33048 28033 33057 28067
rect 33057 28033 33091 28067
rect 33091 28033 33100 28067
rect 33048 28024 33100 28033
rect 33324 28024 33376 28076
rect 34428 28092 34480 28144
rect 36176 28160 36228 28212
rect 36268 28160 36320 28212
rect 33508 28067 33560 28076
rect 33508 28033 33518 28067
rect 33518 28033 33552 28067
rect 33552 28033 33560 28067
rect 33508 28024 33560 28033
rect 33784 28067 33836 28076
rect 33784 28033 33793 28067
rect 33793 28033 33827 28067
rect 33827 28033 33836 28067
rect 33784 28024 33836 28033
rect 33968 28024 34020 28076
rect 34336 28067 34388 28076
rect 34336 28033 34345 28067
rect 34345 28033 34379 28067
rect 34379 28033 34388 28067
rect 34336 28024 34388 28033
rect 35256 28067 35308 28076
rect 35256 28033 35265 28067
rect 35265 28033 35299 28067
rect 35299 28033 35308 28067
rect 35256 28024 35308 28033
rect 36636 28024 36688 28076
rect 37464 28160 37516 28212
rect 37556 28160 37608 28212
rect 40500 28160 40552 28212
rect 39488 28092 39540 28144
rect 40040 28135 40092 28144
rect 40040 28101 40049 28135
rect 40049 28101 40083 28135
rect 40083 28101 40092 28135
rect 40040 28092 40092 28101
rect 40684 28135 40736 28144
rect 40684 28101 40693 28135
rect 40693 28101 40727 28135
rect 40727 28101 40736 28135
rect 40684 28092 40736 28101
rect 41420 28092 41472 28144
rect 37464 28067 37516 28076
rect 37464 28033 37471 28067
rect 37471 28033 37516 28067
rect 37464 28024 37516 28033
rect 33048 27888 33100 27940
rect 34152 27888 34204 27940
rect 35164 27956 35216 28008
rect 36268 27956 36320 28008
rect 36912 27956 36964 28008
rect 37740 28067 37792 28076
rect 37740 28033 37773 28067
rect 37773 28033 37792 28067
rect 37740 28024 37792 28033
rect 38936 28067 38988 28076
rect 38936 28033 38945 28067
rect 38945 28033 38979 28067
rect 38979 28033 38988 28067
rect 38936 28024 38988 28033
rect 39764 28067 39816 28076
rect 39764 28033 39773 28067
rect 39773 28033 39807 28067
rect 39807 28033 39816 28067
rect 39764 28024 39816 28033
rect 37924 27956 37976 28008
rect 40224 28024 40276 28076
rect 40316 27956 40368 28008
rect 40408 27999 40460 28008
rect 40408 27965 40417 27999
rect 40417 27965 40451 27999
rect 40451 27965 40460 27999
rect 40408 27956 40460 27965
rect 26884 27820 26936 27872
rect 27620 27820 27672 27872
rect 30840 27820 30892 27872
rect 31760 27820 31812 27872
rect 34704 27820 34756 27872
rect 40224 27888 40276 27940
rect 35624 27820 35676 27872
rect 36912 27820 36964 27872
rect 37004 27863 37056 27872
rect 37004 27829 37013 27863
rect 37013 27829 37047 27863
rect 37047 27829 37056 27863
rect 37004 27820 37056 27829
rect 39028 27863 39080 27872
rect 39028 27829 39037 27863
rect 39037 27829 39071 27863
rect 39071 27829 39080 27863
rect 39028 27820 39080 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3976 27616 4028 27668
rect 4344 27616 4396 27668
rect 4896 27616 4948 27668
rect 12072 27616 12124 27668
rect 14924 27616 14976 27668
rect 15844 27616 15896 27668
rect 16948 27616 17000 27668
rect 17776 27616 17828 27668
rect 19340 27616 19392 27668
rect 21180 27616 21232 27668
rect 5172 27591 5224 27600
rect 5172 27557 5181 27591
rect 5181 27557 5215 27591
rect 5215 27557 5224 27591
rect 5172 27548 5224 27557
rect 14004 27548 14056 27600
rect 14188 27548 14240 27600
rect 16028 27548 16080 27600
rect 18696 27548 18748 27600
rect 21272 27548 21324 27600
rect 22100 27616 22152 27668
rect 32404 27616 32456 27668
rect 33048 27616 33100 27668
rect 33968 27616 34020 27668
rect 34796 27616 34848 27668
rect 22744 27548 22796 27600
rect 4804 27480 4856 27532
rect 12256 27523 12308 27532
rect 12256 27489 12265 27523
rect 12265 27489 12299 27523
rect 12299 27489 12308 27523
rect 12256 27480 12308 27489
rect 14096 27480 14148 27532
rect 4068 27455 4120 27464
rect 4068 27421 4077 27455
rect 4077 27421 4111 27455
rect 4111 27421 4120 27455
rect 4068 27412 4120 27421
rect 4712 27412 4764 27464
rect 5264 27455 5316 27464
rect 5264 27421 5273 27455
rect 5273 27421 5307 27455
rect 5307 27421 5316 27455
rect 5264 27412 5316 27421
rect 10784 27412 10836 27464
rect 12624 27412 12676 27464
rect 10416 27344 10468 27396
rect 11428 27387 11480 27396
rect 11428 27353 11437 27387
rect 11437 27353 11471 27387
rect 11471 27353 11480 27387
rect 11428 27344 11480 27353
rect 13268 27412 13320 27464
rect 16212 27480 16264 27532
rect 15476 27412 15528 27464
rect 15752 27412 15804 27464
rect 16120 27455 16172 27464
rect 16120 27421 16129 27455
rect 16129 27421 16163 27455
rect 16163 27421 16172 27455
rect 16120 27412 16172 27421
rect 16396 27455 16448 27464
rect 16396 27421 16405 27455
rect 16405 27421 16439 27455
rect 16439 27421 16448 27455
rect 16396 27412 16448 27421
rect 18144 27480 18196 27532
rect 17132 27412 17184 27464
rect 4528 27276 4580 27328
rect 5448 27276 5500 27328
rect 5724 27276 5776 27328
rect 10600 27276 10652 27328
rect 12348 27276 12400 27328
rect 12808 27276 12860 27328
rect 15936 27344 15988 27396
rect 16488 27344 16540 27396
rect 16672 27344 16724 27396
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 18236 27455 18288 27464
rect 18236 27421 18245 27455
rect 18245 27421 18279 27455
rect 18279 27421 18288 27455
rect 18236 27412 18288 27421
rect 18788 27480 18840 27532
rect 19524 27412 19576 27464
rect 20536 27412 20588 27464
rect 21456 27412 21508 27464
rect 17776 27387 17828 27396
rect 17776 27353 17785 27387
rect 17785 27353 17819 27387
rect 17819 27353 17828 27387
rect 17776 27344 17828 27353
rect 17868 27387 17920 27396
rect 17868 27353 17877 27387
rect 17877 27353 17911 27387
rect 17911 27353 17920 27387
rect 17868 27344 17920 27353
rect 14740 27276 14792 27328
rect 17408 27319 17460 27328
rect 17408 27285 17417 27319
rect 17417 27285 17451 27319
rect 17451 27285 17460 27319
rect 17408 27276 17460 27285
rect 17592 27276 17644 27328
rect 19616 27344 19668 27396
rect 21180 27387 21232 27396
rect 21180 27353 21189 27387
rect 21189 27353 21223 27387
rect 21223 27353 21232 27387
rect 21180 27344 21232 27353
rect 21916 27412 21968 27464
rect 22192 27412 22244 27464
rect 22376 27455 22428 27464
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 24216 27548 24268 27600
rect 23296 27455 23348 27464
rect 23296 27421 23305 27455
rect 23305 27421 23339 27455
rect 23339 27421 23348 27455
rect 23296 27412 23348 27421
rect 24124 27412 24176 27464
rect 26056 27523 26108 27532
rect 26056 27489 26065 27523
rect 26065 27489 26099 27523
rect 26099 27489 26108 27523
rect 26056 27480 26108 27489
rect 28908 27591 28960 27600
rect 28908 27557 28917 27591
rect 28917 27557 28951 27591
rect 28951 27557 28960 27591
rect 28908 27548 28960 27557
rect 29184 27548 29236 27600
rect 29828 27548 29880 27600
rect 24676 27412 24728 27464
rect 24768 27412 24820 27464
rect 26608 27412 26660 27464
rect 26884 27455 26936 27464
rect 26884 27421 26893 27455
rect 26893 27421 26927 27455
rect 26927 27421 26936 27455
rect 26884 27412 26936 27421
rect 20352 27276 20404 27328
rect 21824 27276 21876 27328
rect 23388 27276 23440 27328
rect 24584 27276 24636 27328
rect 25688 27276 25740 27328
rect 25872 27276 25924 27328
rect 26516 27319 26568 27328
rect 26516 27285 26525 27319
rect 26525 27285 26559 27319
rect 26559 27285 26568 27319
rect 26516 27276 26568 27285
rect 26700 27387 26752 27396
rect 26700 27353 26709 27387
rect 26709 27353 26743 27387
rect 26743 27353 26752 27387
rect 26700 27344 26752 27353
rect 27068 27387 27120 27396
rect 27068 27353 27077 27387
rect 27077 27353 27111 27387
rect 27111 27353 27120 27387
rect 27068 27344 27120 27353
rect 27344 27344 27396 27396
rect 27436 27387 27488 27396
rect 27436 27353 27445 27387
rect 27445 27353 27479 27387
rect 27479 27353 27488 27387
rect 27436 27344 27488 27353
rect 27896 27344 27948 27396
rect 30196 27523 30248 27532
rect 30196 27489 30205 27523
rect 30205 27489 30239 27523
rect 30239 27489 30248 27523
rect 30196 27480 30248 27489
rect 29184 27412 29236 27464
rect 30012 27412 30064 27464
rect 30840 27412 30892 27464
rect 31484 27412 31536 27464
rect 32312 27387 32364 27396
rect 32312 27353 32321 27387
rect 32321 27353 32355 27387
rect 32355 27353 32364 27387
rect 32312 27344 32364 27353
rect 35072 27548 35124 27600
rect 33876 27480 33928 27532
rect 34428 27523 34480 27532
rect 34428 27489 34437 27523
rect 34437 27489 34471 27523
rect 34471 27489 34480 27523
rect 34428 27480 34480 27489
rect 35256 27548 35308 27600
rect 39856 27548 39908 27600
rect 33600 27412 33652 27464
rect 34612 27412 34664 27464
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 32956 27344 33008 27396
rect 33508 27344 33560 27396
rect 33968 27344 34020 27396
rect 35164 27455 35216 27464
rect 35164 27421 35178 27455
rect 35178 27421 35212 27455
rect 35212 27421 35216 27455
rect 35440 27480 35492 27532
rect 36084 27480 36136 27532
rect 35164 27412 35216 27421
rect 35992 27455 36044 27464
rect 35992 27421 35999 27455
rect 35999 27421 36044 27455
rect 35992 27412 36044 27421
rect 37004 27480 37056 27532
rect 37280 27480 37332 27532
rect 38292 27480 38344 27532
rect 38936 27480 38988 27532
rect 39120 27480 39172 27532
rect 36268 27455 36320 27464
rect 36268 27421 36282 27455
rect 36282 27421 36316 27455
rect 36316 27421 36320 27455
rect 36268 27412 36320 27421
rect 36452 27412 36504 27464
rect 35624 27344 35676 27396
rect 38108 27344 38160 27396
rect 28080 27276 28132 27328
rect 29920 27276 29972 27328
rect 31300 27319 31352 27328
rect 31300 27285 31309 27319
rect 31309 27285 31343 27319
rect 31343 27285 31352 27319
rect 31300 27276 31352 27285
rect 31392 27276 31444 27328
rect 31760 27319 31812 27328
rect 31760 27285 31769 27319
rect 31769 27285 31803 27319
rect 31803 27285 31812 27319
rect 31760 27276 31812 27285
rect 34060 27276 34112 27328
rect 35440 27276 35492 27328
rect 36360 27276 36412 27328
rect 37832 27276 37884 27328
rect 38016 27276 38068 27328
rect 38476 27276 38528 27328
rect 38752 27276 38804 27328
rect 38936 27276 38988 27328
rect 39212 27387 39264 27396
rect 39212 27353 39221 27387
rect 39221 27353 39255 27387
rect 39255 27353 39264 27387
rect 39212 27344 39264 27353
rect 40316 27387 40368 27396
rect 40316 27353 40325 27387
rect 40325 27353 40359 27387
rect 40359 27353 40368 27387
rect 40316 27344 40368 27353
rect 40776 27455 40828 27464
rect 40776 27421 40785 27455
rect 40785 27421 40819 27455
rect 40819 27421 40828 27455
rect 40776 27412 40828 27421
rect 41604 27412 41656 27464
rect 39396 27319 39448 27328
rect 39396 27285 39405 27319
rect 39405 27285 39439 27319
rect 39439 27285 39448 27319
rect 39396 27276 39448 27285
rect 40224 27276 40276 27328
rect 41052 27344 41104 27396
rect 41144 27319 41196 27328
rect 41144 27285 41153 27319
rect 41153 27285 41187 27319
rect 41187 27285 41196 27319
rect 41144 27276 41196 27285
rect 41512 27319 41564 27328
rect 41512 27285 41521 27319
rect 41521 27285 41555 27319
rect 41555 27285 41564 27319
rect 41512 27276 41564 27285
rect 41880 27319 41932 27328
rect 41880 27285 41889 27319
rect 41889 27285 41923 27319
rect 41923 27285 41932 27319
rect 41880 27276 41932 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 3056 27115 3108 27124
rect 3056 27081 3065 27115
rect 3065 27081 3099 27115
rect 3099 27081 3108 27115
rect 3056 27072 3108 27081
rect 4804 27072 4856 27124
rect 1768 26936 1820 26988
rect 3516 27004 3568 27056
rect 8116 27072 8168 27124
rect 10232 27072 10284 27124
rect 10416 27115 10468 27124
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 10600 27072 10652 27124
rect 12808 27072 12860 27124
rect 13176 27072 13228 27124
rect 8208 27004 8260 27056
rect 3332 26936 3384 26988
rect 3884 26936 3936 26988
rect 2596 26800 2648 26852
rect 4344 26979 4396 26988
rect 4344 26945 4353 26979
rect 4353 26945 4387 26979
rect 4387 26945 4396 26979
rect 4344 26936 4396 26945
rect 4528 26936 4580 26988
rect 4804 26868 4856 26920
rect 5448 26936 5500 26988
rect 9680 26936 9732 26988
rect 10048 26979 10100 26988
rect 10048 26945 10057 26979
rect 10057 26945 10091 26979
rect 10091 26945 10100 26979
rect 10048 26936 10100 26945
rect 10140 26936 10192 26988
rect 4712 26800 4764 26852
rect 6000 26868 6052 26920
rect 7196 26868 7248 26920
rect 8208 26868 8260 26920
rect 8576 26868 8628 26920
rect 10508 26936 10560 26988
rect 12348 26936 12400 26988
rect 13912 27047 13964 27056
rect 13912 27013 13921 27047
rect 13921 27013 13955 27047
rect 13955 27013 13964 27047
rect 13912 27004 13964 27013
rect 13084 26979 13136 26988
rect 10968 26911 11020 26920
rect 10968 26877 10977 26911
rect 10977 26877 11011 26911
rect 11011 26877 11020 26911
rect 10968 26868 11020 26877
rect 11520 26911 11572 26920
rect 11520 26877 11529 26911
rect 11529 26877 11563 26911
rect 11563 26877 11572 26911
rect 11520 26868 11572 26877
rect 848 26732 900 26784
rect 2872 26775 2924 26784
rect 2872 26741 2881 26775
rect 2881 26741 2915 26775
rect 2915 26741 2924 26775
rect 2872 26732 2924 26741
rect 3792 26775 3844 26784
rect 3792 26741 3801 26775
rect 3801 26741 3835 26775
rect 3835 26741 3844 26775
rect 3792 26732 3844 26741
rect 5264 26800 5316 26852
rect 5724 26800 5776 26852
rect 10232 26800 10284 26852
rect 13084 26945 13093 26979
rect 13093 26945 13127 26979
rect 13127 26945 13136 26979
rect 13084 26936 13136 26945
rect 13360 26979 13412 26988
rect 13360 26945 13369 26979
rect 13369 26945 13403 26979
rect 13403 26945 13412 26979
rect 13360 26936 13412 26945
rect 13176 26868 13228 26920
rect 12624 26800 12676 26852
rect 14648 27004 14700 27056
rect 16672 27072 16724 27124
rect 17500 27072 17552 27124
rect 17776 27072 17828 27124
rect 15200 27004 15252 27056
rect 16304 27004 16356 27056
rect 17408 27004 17460 27056
rect 18144 27047 18196 27056
rect 18144 27013 18153 27047
rect 18153 27013 18187 27047
rect 18187 27013 18196 27047
rect 18144 27004 18196 27013
rect 19984 27072 20036 27124
rect 24952 27072 25004 27124
rect 25872 27072 25924 27124
rect 26700 27072 26752 27124
rect 27068 27072 27120 27124
rect 27436 27072 27488 27124
rect 28080 27072 28132 27124
rect 35164 27072 35216 27124
rect 36268 27072 36320 27124
rect 37004 27072 37056 27124
rect 40040 27072 40092 27124
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 18052 26936 18104 26988
rect 21456 27004 21508 27056
rect 22928 27004 22980 27056
rect 24584 27004 24636 27056
rect 26516 27004 26568 27056
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 18696 26936 18748 26945
rect 14096 26868 14148 26920
rect 17776 26868 17828 26920
rect 19432 26868 19484 26920
rect 19524 26911 19576 26920
rect 19524 26877 19533 26911
rect 19533 26877 19567 26911
rect 19567 26877 19576 26911
rect 19524 26868 19576 26877
rect 20444 26868 20496 26920
rect 20996 26911 21048 26920
rect 20996 26877 21005 26911
rect 21005 26877 21039 26911
rect 21039 26877 21048 26911
rect 20996 26868 21048 26877
rect 21364 26868 21416 26920
rect 24308 26911 24360 26920
rect 24308 26877 24317 26911
rect 24317 26877 24351 26911
rect 24351 26877 24360 26911
rect 24308 26868 24360 26877
rect 6552 26732 6604 26784
rect 8392 26732 8444 26784
rect 11244 26732 11296 26784
rect 11704 26775 11756 26784
rect 11704 26741 11713 26775
rect 11713 26741 11747 26775
rect 11747 26741 11756 26775
rect 11704 26732 11756 26741
rect 18604 26800 18656 26852
rect 14924 26732 14976 26784
rect 16764 26732 16816 26784
rect 19156 26732 19208 26784
rect 23296 26800 23348 26852
rect 21548 26732 21600 26784
rect 27252 26979 27304 26988
rect 27252 26945 27261 26979
rect 27261 26945 27295 26979
rect 27295 26945 27304 26979
rect 27252 26936 27304 26945
rect 29828 27047 29880 27056
rect 29828 27013 29837 27047
rect 29837 27013 29871 27047
rect 29871 27013 29880 27047
rect 29828 27004 29880 27013
rect 30748 27004 30800 27056
rect 36452 27004 36504 27056
rect 36636 27004 36688 27056
rect 38660 27004 38712 27056
rect 39396 27004 39448 27056
rect 39580 27004 39632 27056
rect 25872 26868 25924 26920
rect 26608 26868 26660 26920
rect 29276 26936 29328 26988
rect 27988 26868 28040 26920
rect 29920 26979 29972 26988
rect 29920 26945 29929 26979
rect 29929 26945 29963 26979
rect 29963 26945 29972 26979
rect 29920 26936 29972 26945
rect 32312 26936 32364 26988
rect 41236 26979 41288 26988
rect 41236 26945 41245 26979
rect 41245 26945 41279 26979
rect 41279 26945 41288 26979
rect 41236 26936 41288 26945
rect 34428 26868 34480 26920
rect 38292 26868 38344 26920
rect 40408 26868 40460 26920
rect 42156 26911 42208 26920
rect 42156 26877 42165 26911
rect 42165 26877 42199 26911
rect 42199 26877 42208 26911
rect 42156 26868 42208 26877
rect 40224 26800 40276 26852
rect 41052 26800 41104 26852
rect 41696 26800 41748 26852
rect 25964 26775 26016 26784
rect 25964 26741 25973 26775
rect 25973 26741 26007 26775
rect 26007 26741 26016 26775
rect 25964 26732 26016 26741
rect 40776 26732 40828 26784
rect 41512 26775 41564 26784
rect 41512 26741 41521 26775
rect 41521 26741 41555 26775
rect 41555 26741 41564 26775
rect 41512 26732 41564 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4804 26528 4856 26580
rect 3792 26392 3844 26444
rect 6184 26528 6236 26580
rect 8576 26571 8628 26580
rect 8576 26537 8585 26571
rect 8585 26537 8619 26571
rect 8619 26537 8628 26571
rect 8576 26528 8628 26537
rect 7564 26460 7616 26512
rect 10232 26528 10284 26580
rect 10508 26528 10560 26580
rect 10876 26528 10928 26580
rect 3056 26256 3108 26308
rect 4620 26367 4672 26376
rect 4620 26333 4629 26367
rect 4629 26333 4663 26367
rect 4663 26333 4672 26367
rect 4620 26324 4672 26333
rect 4712 26324 4764 26376
rect 5080 26367 5132 26376
rect 5080 26333 5089 26367
rect 5089 26333 5123 26367
rect 5123 26333 5132 26367
rect 5080 26324 5132 26333
rect 5172 26324 5224 26376
rect 5724 26392 5776 26444
rect 11336 26528 11388 26580
rect 12256 26528 12308 26580
rect 12624 26528 12676 26580
rect 13728 26571 13780 26580
rect 13728 26537 13737 26571
rect 13737 26537 13771 26571
rect 13771 26537 13780 26571
rect 13728 26528 13780 26537
rect 14188 26528 14240 26580
rect 12808 26460 12860 26512
rect 8024 26367 8076 26376
rect 8024 26333 8033 26367
rect 8033 26333 8067 26367
rect 8067 26333 8076 26367
rect 8024 26324 8076 26333
rect 8116 26324 8168 26376
rect 8576 26324 8628 26376
rect 9680 26324 9732 26376
rect 11244 26435 11296 26444
rect 11244 26401 11253 26435
rect 11253 26401 11287 26435
rect 11287 26401 11296 26435
rect 11244 26392 11296 26401
rect 12440 26392 12492 26444
rect 13084 26392 13136 26444
rect 13636 26392 13688 26444
rect 5724 26299 5776 26308
rect 5724 26265 5733 26299
rect 5733 26265 5767 26299
rect 5767 26265 5776 26299
rect 5724 26256 5776 26265
rect 6460 26256 6512 26308
rect 7104 26256 7156 26308
rect 8484 26256 8536 26308
rect 13084 26256 13136 26308
rect 14556 26367 14608 26376
rect 14556 26333 14565 26367
rect 14565 26333 14599 26367
rect 14599 26333 14608 26367
rect 14556 26324 14608 26333
rect 14740 26324 14792 26376
rect 16948 26460 17000 26512
rect 17776 26460 17828 26512
rect 18144 26460 18196 26512
rect 18788 26460 18840 26512
rect 19156 26528 19208 26580
rect 19616 26571 19668 26580
rect 19616 26537 19625 26571
rect 19625 26537 19659 26571
rect 19659 26537 19668 26571
rect 19616 26528 19668 26537
rect 20996 26528 21048 26580
rect 21456 26528 21508 26580
rect 21548 26528 21600 26580
rect 15200 26435 15252 26444
rect 15200 26401 15209 26435
rect 15209 26401 15243 26435
rect 15243 26401 15252 26435
rect 15200 26392 15252 26401
rect 15660 26392 15712 26444
rect 17592 26367 17644 26376
rect 17592 26333 17601 26367
rect 17601 26333 17635 26367
rect 17635 26333 17644 26367
rect 17592 26324 17644 26333
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 18236 26392 18288 26444
rect 18512 26392 18564 26444
rect 23204 26460 23256 26512
rect 24308 26528 24360 26580
rect 24676 26528 24728 26580
rect 33324 26528 33376 26580
rect 35440 26528 35492 26580
rect 36636 26528 36688 26580
rect 38936 26528 38988 26580
rect 19432 26392 19484 26444
rect 20352 26392 20404 26444
rect 21364 26392 21416 26444
rect 21456 26392 21508 26444
rect 17868 26256 17920 26308
rect 18604 26324 18656 26376
rect 19248 26367 19300 26376
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 2044 26188 2096 26240
rect 2872 26188 2924 26240
rect 5080 26188 5132 26240
rect 5816 26188 5868 26240
rect 7012 26188 7064 26240
rect 13452 26231 13504 26240
rect 13452 26197 13461 26231
rect 13461 26197 13495 26231
rect 13495 26197 13504 26231
rect 13452 26188 13504 26197
rect 15108 26188 15160 26240
rect 15384 26231 15436 26240
rect 15384 26197 15393 26231
rect 15393 26197 15427 26231
rect 15427 26197 15436 26231
rect 15384 26188 15436 26197
rect 17408 26231 17460 26240
rect 17408 26197 17417 26231
rect 17417 26197 17451 26231
rect 17451 26197 17460 26231
rect 17408 26188 17460 26197
rect 18236 26188 18288 26240
rect 20720 26256 20772 26308
rect 20444 26231 20496 26240
rect 20444 26197 20453 26231
rect 20453 26197 20487 26231
rect 20487 26197 20496 26231
rect 20444 26188 20496 26197
rect 21364 26299 21416 26308
rect 21364 26265 21373 26299
rect 21373 26265 21407 26299
rect 21407 26265 21416 26299
rect 21364 26256 21416 26265
rect 21456 26256 21508 26308
rect 22928 26256 22980 26308
rect 23020 26188 23072 26240
rect 24124 26324 24176 26376
rect 24400 26256 24452 26308
rect 25504 26503 25556 26512
rect 25504 26469 25513 26503
rect 25513 26469 25547 26503
rect 25547 26469 25556 26503
rect 25504 26460 25556 26469
rect 41052 26460 41104 26512
rect 25964 26392 26016 26444
rect 31760 26392 31812 26444
rect 35256 26392 35308 26444
rect 35440 26392 35492 26444
rect 36728 26392 36780 26444
rect 37832 26392 37884 26444
rect 41328 26392 41380 26444
rect 24768 26367 24820 26376
rect 24768 26333 24777 26367
rect 24777 26333 24811 26367
rect 24811 26333 24820 26367
rect 24768 26324 24820 26333
rect 24952 26367 25004 26376
rect 24952 26333 24961 26367
rect 24961 26333 24995 26367
rect 24995 26333 25004 26367
rect 24952 26324 25004 26333
rect 25228 26367 25280 26376
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 25780 26324 25832 26376
rect 26332 26324 26384 26376
rect 27068 26324 27120 26376
rect 29552 26324 29604 26376
rect 33600 26324 33652 26376
rect 35348 26367 35400 26376
rect 35348 26333 35357 26367
rect 35357 26333 35391 26367
rect 35391 26333 35400 26367
rect 35348 26324 35400 26333
rect 36084 26324 36136 26376
rect 37464 26324 37516 26376
rect 38016 26324 38068 26376
rect 38752 26367 38804 26376
rect 38752 26333 38761 26367
rect 38761 26333 38795 26367
rect 38795 26333 38804 26367
rect 38752 26324 38804 26333
rect 26976 26256 27028 26308
rect 28724 26256 28776 26308
rect 35992 26256 36044 26308
rect 36544 26299 36596 26308
rect 36544 26265 36553 26299
rect 36553 26265 36587 26299
rect 36587 26265 36596 26299
rect 36544 26256 36596 26265
rect 38108 26299 38160 26308
rect 38108 26265 38117 26299
rect 38117 26265 38151 26299
rect 38151 26265 38160 26299
rect 38108 26256 38160 26265
rect 38384 26256 38436 26308
rect 40408 26256 40460 26308
rect 26608 26188 26660 26240
rect 27160 26188 27212 26240
rect 31760 26188 31812 26240
rect 32956 26231 33008 26240
rect 32956 26197 32965 26231
rect 32965 26197 32999 26231
rect 32999 26197 33008 26231
rect 32956 26188 33008 26197
rect 33416 26231 33468 26240
rect 33416 26197 33425 26231
rect 33425 26197 33459 26231
rect 33459 26197 33468 26231
rect 33416 26188 33468 26197
rect 36176 26231 36228 26240
rect 36176 26197 36185 26231
rect 36185 26197 36219 26231
rect 36219 26197 36228 26231
rect 36176 26188 36228 26197
rect 36912 26188 36964 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 3884 25984 3936 26036
rect 5724 25984 5776 26036
rect 8024 25984 8076 26036
rect 8484 25984 8536 26036
rect 16672 25984 16724 26036
rect 20720 26027 20772 26036
rect 20720 25993 20729 26027
rect 20729 25993 20763 26027
rect 20763 25993 20772 26027
rect 20720 25984 20772 25993
rect 21364 25984 21416 26036
rect 22836 25984 22888 26036
rect 23204 25984 23256 26036
rect 23296 25984 23348 26036
rect 25044 25984 25096 26036
rect 25228 25984 25280 26036
rect 2044 25891 2096 25900
rect 2044 25857 2053 25891
rect 2053 25857 2087 25891
rect 2087 25857 2096 25891
rect 2044 25848 2096 25857
rect 2596 25891 2648 25900
rect 2596 25857 2605 25891
rect 2605 25857 2639 25891
rect 2639 25857 2648 25891
rect 2596 25848 2648 25857
rect 2872 25891 2924 25900
rect 2872 25857 2881 25891
rect 2881 25857 2915 25891
rect 2915 25857 2924 25891
rect 2872 25848 2924 25857
rect 4068 25916 4120 25968
rect 5632 25916 5684 25968
rect 8392 25916 8444 25968
rect 3332 25891 3384 25900
rect 3332 25857 3341 25891
rect 3341 25857 3375 25891
rect 3375 25857 3384 25891
rect 3332 25848 3384 25857
rect 3516 25891 3568 25900
rect 3516 25857 3525 25891
rect 3525 25857 3559 25891
rect 3559 25857 3568 25891
rect 3516 25848 3568 25857
rect 4620 25848 4672 25900
rect 4804 25848 4856 25900
rect 5264 25891 5316 25900
rect 5264 25857 5272 25891
rect 5272 25857 5306 25891
rect 5306 25857 5316 25891
rect 5264 25848 5316 25857
rect 5356 25891 5408 25900
rect 5356 25857 5365 25891
rect 5365 25857 5399 25891
rect 5399 25857 5408 25891
rect 5356 25848 5408 25857
rect 6552 25891 6604 25900
rect 6552 25857 6561 25891
rect 6561 25857 6595 25891
rect 6595 25857 6604 25891
rect 6552 25848 6604 25857
rect 7012 25891 7064 25900
rect 7012 25857 7021 25891
rect 7021 25857 7055 25891
rect 7055 25857 7064 25891
rect 7012 25848 7064 25857
rect 7656 25891 7708 25900
rect 7656 25857 7665 25891
rect 7665 25857 7699 25891
rect 7699 25857 7708 25891
rect 7656 25848 7708 25857
rect 7840 25891 7892 25900
rect 7840 25857 7849 25891
rect 7849 25857 7883 25891
rect 7883 25857 7892 25891
rect 7840 25848 7892 25857
rect 4068 25644 4120 25696
rect 7104 25780 7156 25832
rect 6644 25712 6696 25764
rect 8300 25891 8352 25900
rect 8300 25857 8309 25891
rect 8309 25857 8343 25891
rect 8343 25857 8352 25891
rect 8300 25848 8352 25857
rect 10048 25916 10100 25968
rect 13452 25959 13504 25968
rect 13452 25925 13461 25959
rect 13461 25925 13495 25959
rect 13495 25925 13504 25959
rect 13452 25916 13504 25925
rect 15016 25916 15068 25968
rect 17408 25959 17460 25968
rect 17408 25925 17417 25959
rect 17417 25925 17451 25959
rect 17451 25925 17460 25959
rect 17408 25916 17460 25925
rect 18052 25916 18104 25968
rect 19156 25916 19208 25968
rect 8208 25780 8260 25832
rect 9680 25891 9732 25900
rect 9680 25857 9689 25891
rect 9689 25857 9723 25891
rect 9723 25857 9732 25891
rect 9680 25848 9732 25857
rect 9772 25848 9824 25900
rect 14740 25848 14792 25900
rect 16672 25848 16724 25900
rect 20904 25916 20956 25968
rect 21272 25916 21324 25968
rect 20260 25848 20312 25900
rect 14096 25780 14148 25832
rect 14464 25780 14516 25832
rect 16396 25780 16448 25832
rect 17132 25823 17184 25832
rect 17132 25789 17141 25823
rect 17141 25789 17175 25823
rect 17175 25789 17184 25823
rect 17132 25780 17184 25789
rect 18420 25780 18472 25832
rect 23388 25848 23440 25900
rect 9312 25712 9364 25764
rect 18788 25712 18840 25764
rect 21548 25780 21600 25832
rect 20352 25712 20404 25764
rect 23480 25780 23532 25832
rect 23572 25780 23624 25832
rect 23848 25823 23900 25832
rect 23848 25789 23857 25823
rect 23857 25789 23891 25823
rect 23891 25789 23900 25823
rect 23848 25780 23900 25789
rect 7472 25644 7524 25696
rect 8852 25687 8904 25696
rect 8852 25653 8861 25687
rect 8861 25653 8895 25687
rect 8895 25653 8904 25687
rect 8852 25644 8904 25653
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 12256 25644 12308 25696
rect 17040 25644 17092 25696
rect 17960 25644 18012 25696
rect 18604 25644 18656 25696
rect 19156 25644 19208 25696
rect 22100 25644 22152 25696
rect 23020 25644 23072 25696
rect 23664 25644 23716 25696
rect 23848 25687 23900 25696
rect 23848 25653 23857 25687
rect 23857 25653 23891 25687
rect 23891 25653 23900 25687
rect 23848 25644 23900 25653
rect 24400 25891 24452 25900
rect 24400 25857 24409 25891
rect 24409 25857 24443 25891
rect 24443 25857 24452 25891
rect 24400 25848 24452 25857
rect 24860 25891 24912 25900
rect 24860 25857 24869 25891
rect 24869 25857 24903 25891
rect 24903 25857 24912 25891
rect 24860 25848 24912 25857
rect 25044 25891 25096 25900
rect 25044 25857 25053 25891
rect 25053 25857 25087 25891
rect 25087 25857 25096 25891
rect 25044 25848 25096 25857
rect 27160 26027 27212 26036
rect 27160 25993 27169 26027
rect 27169 25993 27203 26027
rect 27203 25993 27212 26027
rect 27160 25984 27212 25993
rect 32220 25984 32272 26036
rect 25412 25891 25464 25900
rect 25412 25857 25423 25891
rect 25423 25857 25464 25891
rect 25412 25848 25464 25857
rect 25504 25891 25556 25900
rect 25504 25857 25513 25891
rect 25513 25857 25547 25891
rect 25547 25857 25556 25891
rect 25504 25848 25556 25857
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 25872 25891 25924 25900
rect 25872 25857 25881 25891
rect 25881 25857 25915 25891
rect 25915 25857 25924 25891
rect 25872 25848 25924 25857
rect 25964 25891 26016 25900
rect 25964 25857 25973 25891
rect 25973 25857 26007 25891
rect 26007 25857 26016 25891
rect 25964 25848 26016 25857
rect 26148 25848 26200 25900
rect 26332 25891 26384 25900
rect 26332 25857 26341 25891
rect 26341 25857 26375 25891
rect 26375 25857 26384 25891
rect 26332 25848 26384 25857
rect 25596 25823 25648 25832
rect 25596 25789 25605 25823
rect 25605 25789 25639 25823
rect 25639 25789 25648 25823
rect 25596 25780 25648 25789
rect 25780 25780 25832 25832
rect 26976 25891 27028 25900
rect 26976 25857 26985 25891
rect 26985 25857 27019 25891
rect 27019 25857 27028 25891
rect 26976 25848 27028 25857
rect 28724 25891 28776 25900
rect 28724 25857 28733 25891
rect 28733 25857 28767 25891
rect 28767 25857 28776 25891
rect 28724 25848 28776 25857
rect 28816 25891 28868 25900
rect 28816 25857 28825 25891
rect 28825 25857 28859 25891
rect 28859 25857 28868 25891
rect 28816 25848 28868 25857
rect 28908 25891 28960 25900
rect 28908 25857 28917 25891
rect 28917 25857 28951 25891
rect 28951 25857 28960 25891
rect 28908 25848 28960 25857
rect 24400 25712 24452 25764
rect 24860 25712 24912 25764
rect 24952 25712 25004 25764
rect 25136 25712 25188 25764
rect 26608 25780 26660 25832
rect 30012 25848 30064 25900
rect 29276 25780 29328 25832
rect 29552 25823 29604 25832
rect 29552 25789 29561 25823
rect 29561 25789 29595 25823
rect 29595 25789 29604 25823
rect 29552 25780 29604 25789
rect 29092 25712 29144 25764
rect 24768 25644 24820 25696
rect 25964 25644 26016 25696
rect 26608 25687 26660 25696
rect 26608 25653 26617 25687
rect 26617 25653 26651 25687
rect 26651 25653 26660 25687
rect 26608 25644 26660 25653
rect 28540 25687 28592 25696
rect 28540 25653 28549 25687
rect 28549 25653 28583 25687
rect 28583 25653 28592 25687
rect 28540 25644 28592 25653
rect 28724 25644 28776 25696
rect 30012 25712 30064 25764
rect 29736 25644 29788 25696
rect 30380 25891 30432 25900
rect 30380 25857 30389 25891
rect 30389 25857 30423 25891
rect 30423 25857 30432 25891
rect 30380 25848 30432 25857
rect 31392 25848 31444 25900
rect 32036 25848 32088 25900
rect 32956 25916 33008 25968
rect 34152 25916 34204 25968
rect 34796 25984 34848 26036
rect 35348 25984 35400 26036
rect 36728 25984 36780 26036
rect 31760 25823 31812 25832
rect 31760 25789 31769 25823
rect 31769 25789 31803 25823
rect 31803 25789 31812 25823
rect 31760 25780 31812 25789
rect 33692 25780 33744 25832
rect 34152 25823 34204 25832
rect 34152 25789 34161 25823
rect 34161 25789 34195 25823
rect 34195 25789 34204 25823
rect 34152 25780 34204 25789
rect 30380 25712 30432 25764
rect 31208 25687 31260 25696
rect 31208 25653 31217 25687
rect 31217 25653 31251 25687
rect 31251 25653 31260 25687
rect 31208 25644 31260 25653
rect 32496 25644 32548 25696
rect 32772 25644 32824 25696
rect 34612 25823 34664 25832
rect 34612 25789 34621 25823
rect 34621 25789 34655 25823
rect 34655 25789 34664 25823
rect 34612 25780 34664 25789
rect 39212 25984 39264 26036
rect 41604 25984 41656 26036
rect 39488 25916 39540 25968
rect 41420 25916 41472 25968
rect 36912 25891 36964 25900
rect 36912 25857 36921 25891
rect 36921 25857 36955 25891
rect 36955 25857 36964 25891
rect 36912 25848 36964 25857
rect 37372 25848 37424 25900
rect 37004 25780 37056 25832
rect 37556 25780 37608 25832
rect 38108 25780 38160 25832
rect 38568 25780 38620 25832
rect 39028 25891 39080 25900
rect 39028 25857 39037 25891
rect 39037 25857 39071 25891
rect 39071 25857 39080 25891
rect 39028 25848 39080 25857
rect 40224 25848 40276 25900
rect 40132 25780 40184 25832
rect 38476 25712 38528 25764
rect 36084 25687 36136 25696
rect 36084 25653 36093 25687
rect 36093 25653 36127 25687
rect 36127 25653 36136 25687
rect 36084 25644 36136 25653
rect 36268 25644 36320 25696
rect 37096 25644 37148 25696
rect 37280 25687 37332 25696
rect 37280 25653 37289 25687
rect 37289 25653 37323 25687
rect 37323 25653 37332 25687
rect 37280 25644 37332 25653
rect 40132 25687 40184 25696
rect 40132 25653 40141 25687
rect 40141 25653 40175 25687
rect 40175 25653 40184 25687
rect 40132 25644 40184 25653
rect 40408 25823 40460 25832
rect 40408 25789 40417 25823
rect 40417 25789 40451 25823
rect 40451 25789 40460 25823
rect 40408 25780 40460 25789
rect 41144 25780 41196 25832
rect 42064 25644 42116 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5264 25440 5316 25492
rect 7564 25483 7616 25492
rect 7564 25449 7573 25483
rect 7573 25449 7607 25483
rect 7607 25449 7616 25483
rect 7564 25440 7616 25449
rect 10048 25440 10100 25492
rect 11428 25440 11480 25492
rect 17500 25440 17552 25492
rect 17684 25440 17736 25492
rect 20260 25483 20312 25492
rect 20260 25449 20269 25483
rect 20269 25449 20303 25483
rect 20303 25449 20312 25483
rect 20260 25440 20312 25449
rect 21548 25483 21600 25492
rect 21548 25449 21557 25483
rect 21557 25449 21591 25483
rect 21591 25449 21600 25483
rect 21548 25440 21600 25449
rect 14372 25372 14424 25424
rect 16764 25372 16816 25424
rect 4160 25304 4212 25356
rect 4620 25304 4672 25356
rect 11704 25304 11756 25356
rect 12440 25304 12492 25356
rect 13176 25304 13228 25356
rect 16672 25304 16724 25356
rect 2872 25143 2924 25152
rect 2872 25109 2881 25143
rect 2881 25109 2915 25143
rect 2915 25109 2924 25143
rect 2872 25100 2924 25109
rect 3424 25236 3476 25288
rect 3516 25279 3568 25288
rect 3516 25245 3525 25279
rect 3525 25245 3559 25279
rect 3559 25245 3568 25279
rect 3516 25236 3568 25245
rect 5356 25236 5408 25288
rect 6276 25236 6328 25288
rect 9680 25236 9732 25288
rect 15108 25279 15160 25288
rect 15108 25245 15117 25279
rect 15117 25245 15151 25279
rect 15151 25245 15160 25279
rect 15108 25236 15160 25245
rect 4068 25211 4120 25220
rect 4068 25177 4077 25211
rect 4077 25177 4111 25211
rect 4111 25177 4120 25211
rect 4068 25168 4120 25177
rect 6460 25211 6512 25220
rect 6460 25177 6494 25211
rect 6494 25177 6512 25211
rect 6460 25168 6512 25177
rect 8852 25168 8904 25220
rect 11428 25168 11480 25220
rect 15476 25279 15528 25288
rect 15476 25245 15485 25279
rect 15485 25245 15519 25279
rect 15519 25245 15528 25279
rect 15476 25236 15528 25245
rect 15568 25236 15620 25288
rect 16028 25236 16080 25288
rect 16580 25279 16632 25288
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 17040 25347 17092 25356
rect 17040 25313 17049 25347
rect 17049 25313 17083 25347
rect 17083 25313 17092 25347
rect 17040 25304 17092 25313
rect 17408 25372 17460 25424
rect 17592 25372 17644 25424
rect 17960 25304 18012 25356
rect 16672 25211 16724 25220
rect 16672 25177 16681 25211
rect 16681 25177 16715 25211
rect 16715 25177 16724 25211
rect 16672 25168 16724 25177
rect 16764 25211 16816 25220
rect 16764 25177 16773 25211
rect 16773 25177 16807 25211
rect 16807 25177 16816 25211
rect 16764 25168 16816 25177
rect 3424 25100 3476 25152
rect 3976 25100 4028 25152
rect 5632 25100 5684 25152
rect 11796 25100 11848 25152
rect 13360 25100 13412 25152
rect 14556 25100 14608 25152
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 18236 25304 18288 25356
rect 18328 25347 18380 25356
rect 18328 25313 18337 25347
rect 18337 25313 18371 25347
rect 18371 25313 18380 25347
rect 18328 25304 18380 25313
rect 18512 25304 18564 25356
rect 17684 25168 17736 25220
rect 18144 25279 18196 25288
rect 18144 25245 18153 25279
rect 18153 25245 18187 25279
rect 18187 25245 18196 25279
rect 18144 25236 18196 25245
rect 18420 25279 18472 25288
rect 18420 25245 18429 25279
rect 18429 25245 18463 25279
rect 18463 25245 18472 25279
rect 18420 25236 18472 25245
rect 20260 25279 20312 25288
rect 20260 25245 20269 25279
rect 20269 25245 20303 25279
rect 20303 25245 20312 25279
rect 20260 25236 20312 25245
rect 20996 25236 21048 25288
rect 21732 25279 21784 25288
rect 21732 25245 21741 25279
rect 21741 25245 21775 25279
rect 21775 25245 21784 25279
rect 21732 25236 21784 25245
rect 22100 25440 22152 25492
rect 23848 25440 23900 25492
rect 25872 25440 25924 25492
rect 26148 25440 26200 25492
rect 24400 25372 24452 25424
rect 22652 25304 22704 25356
rect 23480 25304 23532 25356
rect 23848 25304 23900 25356
rect 22284 25236 22336 25288
rect 22468 25279 22520 25288
rect 22468 25245 22477 25279
rect 22477 25245 22511 25279
rect 22511 25245 22520 25279
rect 22468 25236 22520 25245
rect 22836 25279 22888 25288
rect 22836 25245 22845 25279
rect 22845 25245 22879 25279
rect 22879 25245 22888 25279
rect 22836 25236 22888 25245
rect 23020 25279 23072 25288
rect 23020 25245 23029 25279
rect 23029 25245 23063 25279
rect 23063 25245 23072 25279
rect 23020 25236 23072 25245
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 23940 25279 23992 25288
rect 23940 25245 23949 25279
rect 23949 25245 23983 25279
rect 23983 25245 23992 25279
rect 23940 25236 23992 25245
rect 18788 25168 18840 25220
rect 17592 25100 17644 25152
rect 24676 25279 24728 25288
rect 24676 25245 24685 25279
rect 24685 25245 24719 25279
rect 24719 25245 24728 25279
rect 24676 25236 24728 25245
rect 24860 25236 24912 25288
rect 25044 25279 25096 25288
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 25596 25372 25648 25424
rect 28816 25440 28868 25492
rect 30380 25483 30432 25492
rect 30380 25449 30389 25483
rect 30389 25449 30423 25483
rect 30423 25449 30432 25483
rect 30380 25440 30432 25449
rect 31852 25440 31904 25492
rect 32220 25440 32272 25492
rect 32864 25440 32916 25492
rect 33416 25440 33468 25492
rect 35164 25440 35216 25492
rect 36084 25440 36136 25492
rect 36452 25440 36504 25492
rect 36820 25440 36872 25492
rect 39212 25440 39264 25492
rect 29000 25372 29052 25424
rect 29092 25372 29144 25424
rect 25964 25304 26016 25356
rect 25780 25279 25832 25288
rect 25780 25245 25789 25279
rect 25789 25245 25823 25279
rect 25823 25245 25832 25279
rect 25780 25236 25832 25245
rect 25228 25168 25280 25220
rect 27896 25236 27948 25288
rect 28540 25347 28592 25356
rect 28540 25313 28549 25347
rect 28549 25313 28583 25347
rect 28583 25313 28592 25347
rect 28540 25304 28592 25313
rect 28724 25347 28776 25356
rect 28724 25313 28733 25347
rect 28733 25313 28767 25347
rect 28767 25313 28776 25347
rect 28724 25304 28776 25313
rect 28908 25304 28960 25356
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 35348 25372 35400 25424
rect 31116 25304 31168 25356
rect 31668 25304 31720 25356
rect 32680 25347 32732 25356
rect 32680 25313 32689 25347
rect 32689 25313 32723 25347
rect 32723 25313 32732 25347
rect 32680 25304 32732 25313
rect 34796 25347 34848 25356
rect 34796 25313 34805 25347
rect 34805 25313 34839 25347
rect 34839 25313 34848 25347
rect 34796 25304 34848 25313
rect 36176 25304 36228 25356
rect 36452 25304 36504 25356
rect 37648 25372 37700 25424
rect 37740 25372 37792 25424
rect 37280 25304 37332 25356
rect 38384 25304 38436 25356
rect 40500 25440 40552 25492
rect 42156 25483 42208 25492
rect 42156 25449 42165 25483
rect 42165 25449 42199 25483
rect 42199 25449 42208 25483
rect 42156 25440 42208 25449
rect 30748 25279 30800 25288
rect 30748 25245 30757 25279
rect 30757 25245 30791 25279
rect 30791 25245 30800 25279
rect 30748 25236 30800 25245
rect 32772 25236 32824 25288
rect 33416 25236 33468 25288
rect 33784 25279 33836 25288
rect 33784 25245 33793 25279
rect 33793 25245 33827 25279
rect 33827 25245 33836 25279
rect 33784 25236 33836 25245
rect 33876 25279 33928 25288
rect 33876 25245 33885 25279
rect 33885 25245 33919 25279
rect 33919 25245 33928 25279
rect 33876 25236 33928 25245
rect 33968 25236 34020 25288
rect 34520 25236 34572 25288
rect 35992 25279 36044 25288
rect 35992 25245 36001 25279
rect 36001 25245 36035 25279
rect 36035 25245 36044 25279
rect 35992 25236 36044 25245
rect 24032 25100 24084 25152
rect 25780 25100 25832 25152
rect 26424 25211 26476 25220
rect 26424 25177 26433 25211
rect 26433 25177 26467 25211
rect 26467 25177 26476 25211
rect 26424 25168 26476 25177
rect 29184 25168 29236 25220
rect 27344 25100 27396 25152
rect 27804 25100 27856 25152
rect 28080 25143 28132 25152
rect 28080 25109 28089 25143
rect 28089 25109 28123 25143
rect 28123 25109 28132 25143
rect 28080 25100 28132 25109
rect 29000 25100 29052 25152
rect 30840 25168 30892 25220
rect 31208 25168 31260 25220
rect 32496 25168 32548 25220
rect 36084 25168 36136 25220
rect 37556 25236 37608 25288
rect 39304 25236 39356 25288
rect 39580 25236 39632 25288
rect 39948 25236 40000 25288
rect 40408 25279 40460 25288
rect 40408 25245 40417 25279
rect 40417 25245 40451 25279
rect 40451 25245 40460 25279
rect 40408 25236 40460 25245
rect 38292 25168 38344 25220
rect 40684 25211 40736 25220
rect 40684 25177 40693 25211
rect 40693 25177 40727 25211
rect 40727 25177 40736 25211
rect 40684 25168 40736 25177
rect 41420 25168 41472 25220
rect 30196 25100 30248 25152
rect 30564 25143 30616 25152
rect 30564 25109 30573 25143
rect 30573 25109 30607 25143
rect 30607 25109 30616 25143
rect 30564 25100 30616 25109
rect 31024 25100 31076 25152
rect 35256 25100 35308 25152
rect 36820 25100 36872 25152
rect 37280 25143 37332 25152
rect 37280 25109 37289 25143
rect 37289 25109 37323 25143
rect 37323 25109 37332 25143
rect 37280 25100 37332 25109
rect 37740 25100 37792 25152
rect 39580 25100 39632 25152
rect 41604 25100 41656 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 2596 24896 2648 24948
rect 3240 24896 3292 24948
rect 3424 24896 3476 24948
rect 5356 24896 5408 24948
rect 6460 24896 6512 24948
rect 7564 24896 7616 24948
rect 7656 24939 7708 24948
rect 7656 24905 7665 24939
rect 7665 24905 7699 24939
rect 7699 24905 7708 24939
rect 7656 24896 7708 24905
rect 8208 24896 8260 24948
rect 3056 24760 3108 24812
rect 3700 24760 3752 24812
rect 4804 24828 4856 24880
rect 6552 24828 6604 24880
rect 4712 24760 4764 24812
rect 5632 24760 5684 24812
rect 6644 24803 6696 24812
rect 6644 24769 6653 24803
rect 6653 24769 6687 24803
rect 6687 24769 6696 24803
rect 6644 24760 6696 24769
rect 6828 24803 6880 24812
rect 6828 24769 6837 24803
rect 6837 24769 6871 24803
rect 6871 24769 6880 24803
rect 6828 24760 6880 24769
rect 7380 24760 7432 24812
rect 7564 24803 7616 24812
rect 7564 24769 7573 24803
rect 7573 24769 7607 24803
rect 7607 24769 7616 24803
rect 7564 24760 7616 24769
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 1676 24735 1728 24744
rect 1676 24701 1685 24735
rect 1685 24701 1719 24735
rect 1719 24701 1728 24735
rect 1676 24692 1728 24701
rect 3424 24692 3476 24744
rect 4160 24624 4212 24676
rect 5356 24692 5408 24744
rect 7840 24760 7892 24812
rect 8760 24760 8812 24812
rect 9312 24803 9364 24812
rect 9312 24769 9321 24803
rect 9321 24769 9355 24803
rect 9355 24769 9364 24803
rect 9312 24760 9364 24769
rect 9588 24803 9640 24812
rect 9588 24769 9597 24803
rect 9597 24769 9631 24803
rect 9631 24769 9640 24803
rect 9588 24760 9640 24769
rect 11796 24871 11848 24880
rect 11796 24837 11805 24871
rect 11805 24837 11839 24871
rect 11839 24837 11848 24871
rect 11796 24828 11848 24837
rect 13084 24828 13136 24880
rect 14556 24871 14608 24880
rect 14556 24837 14565 24871
rect 14565 24837 14599 24871
rect 14599 24837 14608 24871
rect 14556 24828 14608 24837
rect 16028 24939 16080 24948
rect 16028 24905 16037 24939
rect 16037 24905 16071 24939
rect 16071 24905 16080 24939
rect 16028 24896 16080 24905
rect 16672 24939 16724 24948
rect 16672 24905 16681 24939
rect 16681 24905 16715 24939
rect 16715 24905 16724 24939
rect 16672 24896 16724 24905
rect 17040 24896 17092 24948
rect 17408 24896 17460 24948
rect 18328 24939 18380 24948
rect 18328 24905 18337 24939
rect 18337 24905 18371 24939
rect 18371 24905 18380 24939
rect 18328 24896 18380 24905
rect 18420 24896 18472 24948
rect 15016 24828 15068 24880
rect 17592 24828 17644 24880
rect 10692 24760 10744 24812
rect 11336 24760 11388 24812
rect 6644 24624 6696 24676
rect 6000 24556 6052 24608
rect 7380 24556 7432 24608
rect 11060 24692 11112 24744
rect 8300 24624 8352 24676
rect 9588 24624 9640 24676
rect 16212 24803 16264 24812
rect 16212 24769 16221 24803
rect 16221 24769 16255 24803
rect 16255 24769 16264 24803
rect 16212 24760 16264 24769
rect 17040 24803 17092 24812
rect 17040 24769 17049 24803
rect 17049 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 18880 24896 18932 24948
rect 20076 24896 20128 24948
rect 20260 24896 20312 24948
rect 21732 24896 21784 24948
rect 22468 24939 22520 24948
rect 22468 24905 22477 24939
rect 22477 24905 22511 24939
rect 22511 24905 22520 24939
rect 22468 24896 22520 24905
rect 23940 24896 23992 24948
rect 24768 24896 24820 24948
rect 26424 24896 26476 24948
rect 27620 24896 27672 24948
rect 27896 24896 27948 24948
rect 13728 24692 13780 24744
rect 9772 24556 9824 24608
rect 13360 24556 13412 24608
rect 13544 24599 13596 24608
rect 13544 24565 13553 24599
rect 13553 24565 13587 24599
rect 13587 24565 13596 24599
rect 13544 24556 13596 24565
rect 15752 24556 15804 24608
rect 17960 24556 18012 24608
rect 18696 24760 18748 24812
rect 19524 24803 19576 24812
rect 19524 24769 19533 24803
rect 19533 24769 19567 24803
rect 19567 24769 19576 24803
rect 19524 24760 19576 24769
rect 19708 24803 19760 24812
rect 19708 24769 19717 24803
rect 19717 24769 19751 24803
rect 19751 24769 19760 24803
rect 19708 24760 19760 24769
rect 18972 24692 19024 24744
rect 18512 24624 18564 24676
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 20168 24803 20220 24812
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 20996 24871 21048 24880
rect 20996 24837 21005 24871
rect 21005 24837 21039 24871
rect 21039 24837 21048 24871
rect 20996 24828 21048 24837
rect 21456 24803 21508 24812
rect 21456 24769 21465 24803
rect 21465 24769 21499 24803
rect 21499 24769 21508 24803
rect 23388 24828 23440 24880
rect 21456 24760 21508 24769
rect 21732 24692 21784 24744
rect 23572 24760 23624 24812
rect 24032 24760 24084 24812
rect 24676 24828 24728 24880
rect 24492 24803 24544 24812
rect 24492 24769 24501 24803
rect 24501 24769 24535 24803
rect 24535 24769 24544 24803
rect 24492 24760 24544 24769
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 26608 24760 26660 24812
rect 28080 24828 28132 24880
rect 29736 24871 29788 24880
rect 29736 24837 29745 24871
rect 29745 24837 29779 24871
rect 29779 24837 29788 24871
rect 29736 24828 29788 24837
rect 30564 24896 30616 24948
rect 33876 24939 33928 24948
rect 33876 24905 33885 24939
rect 33885 24905 33919 24939
rect 33919 24905 33928 24939
rect 33876 24896 33928 24905
rect 34612 24896 34664 24948
rect 35164 24939 35216 24948
rect 35164 24905 35173 24939
rect 35173 24905 35207 24939
rect 35207 24905 35216 24939
rect 35164 24896 35216 24905
rect 35256 24939 35308 24948
rect 35256 24905 35265 24939
rect 35265 24905 35299 24939
rect 35299 24905 35308 24939
rect 35256 24896 35308 24905
rect 31024 24828 31076 24880
rect 31944 24828 31996 24880
rect 32588 24871 32640 24880
rect 32588 24837 32623 24871
rect 32623 24837 32640 24871
rect 32588 24828 32640 24837
rect 23480 24692 23532 24744
rect 23848 24692 23900 24744
rect 24400 24692 24452 24744
rect 25780 24692 25832 24744
rect 26056 24692 26108 24744
rect 31852 24760 31904 24812
rect 32036 24760 32088 24812
rect 33416 24828 33468 24880
rect 27528 24735 27580 24744
rect 27528 24701 27537 24735
rect 27537 24701 27571 24735
rect 27571 24701 27580 24735
rect 27528 24692 27580 24701
rect 31392 24692 31444 24744
rect 19616 24556 19668 24608
rect 20168 24556 20220 24608
rect 20444 24556 20496 24608
rect 24584 24624 24636 24676
rect 27160 24624 27212 24676
rect 29184 24624 29236 24676
rect 25320 24556 25372 24608
rect 29828 24556 29880 24608
rect 31760 24735 31812 24744
rect 31760 24701 31769 24735
rect 31769 24701 31803 24735
rect 31803 24701 31812 24735
rect 31760 24692 31812 24701
rect 33048 24803 33100 24812
rect 33048 24769 33057 24803
rect 33057 24769 33091 24803
rect 33091 24769 33100 24803
rect 33048 24760 33100 24769
rect 33692 24828 33744 24880
rect 34704 24828 34756 24880
rect 35624 24828 35676 24880
rect 35992 24896 36044 24948
rect 39580 24896 39632 24948
rect 40684 24896 40736 24948
rect 41052 24896 41104 24948
rect 36268 24828 36320 24880
rect 32680 24692 32732 24744
rect 33232 24692 33284 24744
rect 33416 24692 33468 24744
rect 33784 24599 33836 24608
rect 33784 24565 33793 24599
rect 33793 24565 33827 24599
rect 33827 24565 33836 24599
rect 33784 24556 33836 24565
rect 34152 24803 34204 24812
rect 34152 24769 34161 24803
rect 34161 24769 34195 24803
rect 34195 24769 34204 24803
rect 34152 24760 34204 24769
rect 34520 24803 34572 24812
rect 34520 24769 34529 24803
rect 34529 24769 34563 24803
rect 34563 24769 34572 24803
rect 34520 24760 34572 24769
rect 35164 24760 35216 24812
rect 35440 24760 35492 24812
rect 36544 24760 36596 24812
rect 34888 24692 34940 24744
rect 35348 24735 35400 24744
rect 35348 24701 35357 24735
rect 35357 24701 35391 24735
rect 35391 24701 35400 24735
rect 35348 24692 35400 24701
rect 36084 24692 36136 24744
rect 36360 24735 36412 24744
rect 36360 24701 36369 24735
rect 36369 24701 36403 24735
rect 36403 24701 36412 24735
rect 36360 24692 36412 24701
rect 36176 24624 36228 24676
rect 36636 24624 36688 24676
rect 36820 24760 36872 24812
rect 37740 24828 37792 24880
rect 38568 24828 38620 24880
rect 39304 24828 39356 24880
rect 37372 24692 37424 24744
rect 38292 24760 38344 24812
rect 37648 24735 37700 24744
rect 37648 24701 37657 24735
rect 37657 24701 37691 24735
rect 37691 24701 37700 24735
rect 37648 24692 37700 24701
rect 37832 24735 37884 24744
rect 37832 24701 37841 24735
rect 37841 24701 37875 24735
rect 37875 24701 37884 24735
rect 37832 24692 37884 24701
rect 39028 24692 39080 24744
rect 36728 24556 36780 24608
rect 37280 24556 37332 24608
rect 38476 24556 38528 24608
rect 41420 24828 41472 24880
rect 41512 24760 41564 24812
rect 41972 24760 42024 24812
rect 40592 24599 40644 24608
rect 40592 24565 40601 24599
rect 40601 24565 40635 24599
rect 40635 24565 40644 24599
rect 40592 24556 40644 24565
rect 41512 24624 41564 24676
rect 41696 24556 41748 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1676 24352 1728 24404
rect 3516 24352 3568 24404
rect 6920 24352 6972 24404
rect 1768 24284 1820 24336
rect 2872 24216 2924 24268
rect 2780 24148 2832 24200
rect 2964 24191 3016 24200
rect 2964 24157 2973 24191
rect 2973 24157 3007 24191
rect 3007 24157 3016 24191
rect 2964 24148 3016 24157
rect 7104 24284 7156 24336
rect 6000 24259 6052 24268
rect 6000 24225 6009 24259
rect 6009 24225 6043 24259
rect 6043 24225 6052 24259
rect 6000 24216 6052 24225
rect 6276 24216 6328 24268
rect 7288 24216 7340 24268
rect 7656 24216 7708 24268
rect 8208 24259 8260 24268
rect 8208 24225 8217 24259
rect 8217 24225 8251 24259
rect 8251 24225 8260 24259
rect 8208 24216 8260 24225
rect 8300 24259 8352 24268
rect 8300 24225 8309 24259
rect 8309 24225 8343 24259
rect 8343 24225 8352 24259
rect 8300 24216 8352 24225
rect 9680 24352 9732 24404
rect 10692 24395 10744 24404
rect 10692 24361 10701 24395
rect 10701 24361 10735 24395
rect 10735 24361 10744 24395
rect 10692 24352 10744 24361
rect 15016 24352 15068 24404
rect 18604 24352 18656 24404
rect 11336 24216 11388 24268
rect 3056 24080 3108 24132
rect 3240 24191 3292 24200
rect 3240 24157 3249 24191
rect 3249 24157 3283 24191
rect 3283 24157 3292 24191
rect 3240 24148 3292 24157
rect 3424 24191 3476 24200
rect 3424 24157 3433 24191
rect 3433 24157 3467 24191
rect 3467 24157 3476 24191
rect 3424 24148 3476 24157
rect 4804 24148 4856 24200
rect 5540 24191 5592 24200
rect 5540 24157 5549 24191
rect 5549 24157 5583 24191
rect 5583 24157 5592 24191
rect 5540 24148 5592 24157
rect 5632 24191 5684 24200
rect 5632 24157 5641 24191
rect 5641 24157 5675 24191
rect 5675 24157 5684 24191
rect 5632 24148 5684 24157
rect 6644 24191 6696 24200
rect 6644 24157 6653 24191
rect 6653 24157 6687 24191
rect 6687 24157 6696 24191
rect 6644 24148 6696 24157
rect 5356 24080 5408 24132
rect 2688 24012 2740 24064
rect 2872 24055 2924 24064
rect 2872 24021 2881 24055
rect 2881 24021 2915 24055
rect 2915 24021 2924 24055
rect 2872 24012 2924 24021
rect 7012 24080 7064 24132
rect 7196 24080 7248 24132
rect 7288 24080 7340 24132
rect 7104 24012 7156 24064
rect 7472 24080 7524 24132
rect 8576 24148 8628 24200
rect 16028 24216 16080 24268
rect 16948 24216 17000 24268
rect 13544 24191 13596 24200
rect 13544 24157 13553 24191
rect 13553 24157 13587 24191
rect 13587 24157 13596 24191
rect 13544 24148 13596 24157
rect 15016 24148 15068 24200
rect 15108 24191 15160 24200
rect 15108 24157 15117 24191
rect 15117 24157 15151 24191
rect 15151 24157 15160 24191
rect 15108 24148 15160 24157
rect 16672 24148 16724 24200
rect 17132 24148 17184 24200
rect 17592 24191 17644 24200
rect 17592 24157 17601 24191
rect 17601 24157 17635 24191
rect 17635 24157 17644 24191
rect 17592 24148 17644 24157
rect 7656 24080 7708 24132
rect 9588 24123 9640 24132
rect 9588 24089 9622 24123
rect 9622 24089 9640 24123
rect 9588 24080 9640 24089
rect 11796 24123 11848 24132
rect 11796 24089 11805 24123
rect 11805 24089 11839 24123
rect 11839 24089 11848 24123
rect 11796 24080 11848 24089
rect 13084 24080 13136 24132
rect 16580 24080 16632 24132
rect 17776 24080 17828 24132
rect 9312 24012 9364 24064
rect 11428 24055 11480 24064
rect 11428 24021 11437 24055
rect 11437 24021 11471 24055
rect 11471 24021 11480 24055
rect 11428 24012 11480 24021
rect 13268 24055 13320 24064
rect 13268 24021 13277 24055
rect 13277 24021 13311 24055
rect 13311 24021 13320 24055
rect 13268 24012 13320 24021
rect 14004 24012 14056 24064
rect 16948 24012 17000 24064
rect 18512 24191 18564 24200
rect 18512 24157 18522 24191
rect 18522 24157 18556 24191
rect 18556 24157 18564 24191
rect 18512 24148 18564 24157
rect 19064 24352 19116 24404
rect 19248 24395 19300 24404
rect 19248 24361 19257 24395
rect 19257 24361 19291 24395
rect 19291 24361 19300 24395
rect 19248 24352 19300 24361
rect 20444 24395 20496 24404
rect 20444 24361 20453 24395
rect 20453 24361 20487 24395
rect 20487 24361 20496 24395
rect 20444 24352 20496 24361
rect 21456 24352 21508 24404
rect 21732 24395 21784 24404
rect 21732 24361 21741 24395
rect 21741 24361 21775 24395
rect 21775 24361 21784 24395
rect 21732 24352 21784 24361
rect 29552 24395 29604 24404
rect 29552 24361 29561 24395
rect 29561 24361 29595 24395
rect 29595 24361 29604 24395
rect 29552 24352 29604 24361
rect 33048 24352 33100 24404
rect 18972 24284 19024 24336
rect 26884 24284 26936 24336
rect 31944 24284 31996 24336
rect 32404 24284 32456 24336
rect 19064 24148 19116 24200
rect 19156 24148 19208 24200
rect 19616 24191 19668 24200
rect 19616 24157 19625 24191
rect 19625 24157 19659 24191
rect 19659 24157 19668 24191
rect 19616 24148 19668 24157
rect 19892 24216 19944 24268
rect 20076 24191 20128 24200
rect 18236 24080 18288 24132
rect 18788 24080 18840 24132
rect 19248 24012 19300 24064
rect 19524 24123 19576 24132
rect 19524 24089 19533 24123
rect 19533 24089 19567 24123
rect 19567 24089 19576 24123
rect 19524 24080 19576 24089
rect 19708 24080 19760 24132
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20996 24148 21048 24200
rect 22836 24216 22888 24268
rect 23204 24216 23256 24268
rect 33784 24216 33836 24268
rect 23020 24148 23072 24200
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 25320 24191 25372 24200
rect 25320 24157 25329 24191
rect 25329 24157 25363 24191
rect 25363 24157 25372 24191
rect 25320 24148 25372 24157
rect 25964 24191 26016 24200
rect 25964 24157 25973 24191
rect 25973 24157 26007 24191
rect 26007 24157 26016 24191
rect 25964 24148 26016 24157
rect 26056 24191 26108 24200
rect 26056 24157 26065 24191
rect 26065 24157 26099 24191
rect 26099 24157 26108 24191
rect 26056 24148 26108 24157
rect 26700 24148 26752 24200
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 29000 24148 29052 24200
rect 24400 24080 24452 24132
rect 29828 24191 29880 24200
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 31392 24148 31444 24200
rect 31760 24080 31812 24132
rect 35256 24352 35308 24404
rect 35440 24352 35492 24404
rect 36452 24352 36504 24404
rect 36544 24395 36596 24404
rect 36544 24361 36553 24395
rect 36553 24361 36587 24395
rect 36587 24361 36596 24395
rect 36544 24352 36596 24361
rect 34520 24284 34572 24336
rect 36912 24352 36964 24404
rect 37832 24352 37884 24404
rect 41696 24352 41748 24404
rect 42064 24352 42116 24404
rect 36728 24284 36780 24336
rect 35624 24216 35676 24268
rect 36176 24259 36228 24268
rect 36176 24225 36185 24259
rect 36185 24225 36219 24259
rect 36219 24225 36228 24259
rect 36176 24216 36228 24225
rect 36268 24148 36320 24200
rect 36544 24148 36596 24200
rect 37096 24191 37148 24200
rect 37096 24157 37105 24191
rect 37105 24157 37139 24191
rect 37139 24157 37148 24191
rect 37096 24148 37148 24157
rect 37280 24191 37332 24200
rect 37280 24157 37289 24191
rect 37289 24157 37323 24191
rect 37323 24157 37332 24191
rect 37280 24148 37332 24157
rect 37556 24148 37608 24200
rect 39396 24148 39448 24200
rect 39948 24148 40000 24200
rect 35532 24123 35584 24132
rect 35532 24089 35541 24123
rect 35541 24089 35575 24123
rect 35575 24089 35584 24123
rect 35532 24080 35584 24089
rect 36820 24080 36872 24132
rect 26976 24012 27028 24064
rect 28816 24012 28868 24064
rect 29828 24012 29880 24064
rect 35440 24012 35492 24064
rect 36452 24012 36504 24064
rect 40960 24080 41012 24132
rect 41420 24080 41472 24132
rect 37464 24012 37516 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 2780 23808 2832 23860
rect 3056 23851 3108 23860
rect 3056 23817 3065 23851
rect 3065 23817 3099 23851
rect 3099 23817 3108 23851
rect 3056 23808 3108 23817
rect 6828 23808 6880 23860
rect 6920 23851 6972 23860
rect 6920 23817 6929 23851
rect 6929 23817 6963 23851
rect 6963 23817 6972 23851
rect 6920 23808 6972 23817
rect 7840 23808 7892 23860
rect 3424 23740 3476 23792
rect 2688 23715 2740 23724
rect 2688 23681 2697 23715
rect 2697 23681 2731 23715
rect 2731 23681 2740 23715
rect 2688 23672 2740 23681
rect 3240 23672 3292 23724
rect 6552 23740 6604 23792
rect 5264 23672 5316 23724
rect 6276 23672 6328 23724
rect 7288 23740 7340 23792
rect 6828 23715 6880 23724
rect 6828 23681 6837 23715
rect 6837 23681 6871 23715
rect 6871 23681 6880 23715
rect 6828 23672 6880 23681
rect 7380 23672 7432 23724
rect 7932 23672 7984 23724
rect 9312 23783 9364 23792
rect 9312 23749 9321 23783
rect 9321 23749 9355 23783
rect 9355 23749 9364 23783
rect 9312 23740 9364 23749
rect 9588 23851 9640 23860
rect 9588 23817 9597 23851
rect 9597 23817 9631 23851
rect 9631 23817 9640 23851
rect 9588 23808 9640 23817
rect 11796 23851 11848 23860
rect 11796 23817 11805 23851
rect 11805 23817 11839 23851
rect 11839 23817 11848 23851
rect 11796 23808 11848 23817
rect 13268 23808 13320 23860
rect 11428 23740 11480 23792
rect 15016 23808 15068 23860
rect 18420 23851 18472 23860
rect 18420 23817 18429 23851
rect 18429 23817 18463 23851
rect 18463 23817 18472 23851
rect 18420 23808 18472 23817
rect 18696 23808 18748 23860
rect 18972 23851 19024 23860
rect 18972 23817 18981 23851
rect 18981 23817 19015 23851
rect 19015 23817 19024 23851
rect 18972 23808 19024 23817
rect 3148 23604 3200 23656
rect 3332 23604 3384 23656
rect 3700 23604 3752 23656
rect 2964 23579 3016 23588
rect 2964 23545 2973 23579
rect 2973 23545 3007 23579
rect 3007 23545 3016 23579
rect 2964 23536 3016 23545
rect 3792 23536 3844 23588
rect 5172 23604 5224 23656
rect 6552 23647 6604 23656
rect 6552 23613 6561 23647
rect 6561 23613 6595 23647
rect 6595 23613 6604 23647
rect 6552 23604 6604 23613
rect 7104 23604 7156 23656
rect 7196 23647 7248 23656
rect 7196 23613 7205 23647
rect 7205 23613 7239 23647
rect 7239 23613 7248 23647
rect 7196 23604 7248 23613
rect 9128 23604 9180 23656
rect 9496 23672 9548 23724
rect 9680 23672 9732 23724
rect 9864 23672 9916 23724
rect 11060 23672 11112 23724
rect 13728 23715 13780 23724
rect 13728 23681 13737 23715
rect 13737 23681 13771 23715
rect 13771 23681 13780 23715
rect 13728 23672 13780 23681
rect 14004 23715 14056 23724
rect 14004 23681 14038 23715
rect 14038 23681 14056 23715
rect 14004 23672 14056 23681
rect 9312 23604 9364 23656
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 16948 23783 17000 23792
rect 16948 23749 16957 23783
rect 16957 23749 16991 23783
rect 16991 23749 17000 23783
rect 16948 23740 17000 23749
rect 18236 23740 18288 23792
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 16396 23715 16448 23724
rect 16396 23681 16405 23715
rect 16405 23681 16439 23715
rect 16439 23681 16448 23715
rect 16396 23672 16448 23681
rect 16672 23715 16724 23724
rect 8576 23536 8628 23588
rect 4988 23511 5040 23520
rect 4988 23477 4997 23511
rect 4997 23477 5031 23511
rect 5031 23477 5040 23511
rect 4988 23468 5040 23477
rect 7840 23468 7892 23520
rect 10508 23468 10560 23520
rect 14740 23468 14792 23520
rect 15108 23511 15160 23520
rect 15108 23477 15117 23511
rect 15117 23477 15151 23511
rect 15151 23477 15160 23511
rect 15108 23468 15160 23477
rect 15200 23511 15252 23520
rect 15200 23477 15209 23511
rect 15209 23477 15243 23511
rect 15243 23477 15252 23511
rect 15200 23468 15252 23477
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 15752 23647 15804 23656
rect 15752 23613 15761 23647
rect 15761 23613 15795 23647
rect 15795 23613 15804 23647
rect 15752 23604 15804 23613
rect 15936 23604 15988 23656
rect 16672 23681 16688 23715
rect 16688 23681 16722 23715
rect 16722 23681 16724 23715
rect 16672 23672 16724 23681
rect 18052 23672 18104 23724
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 18696 23672 18748 23724
rect 20076 23783 20128 23792
rect 20076 23749 20085 23783
rect 20085 23749 20119 23783
rect 20119 23749 20128 23783
rect 20076 23740 20128 23749
rect 22376 23851 22428 23860
rect 22376 23817 22385 23851
rect 22385 23817 22419 23851
rect 22419 23817 22428 23851
rect 22376 23808 22428 23817
rect 24492 23808 24544 23860
rect 25964 23808 26016 23860
rect 26792 23808 26844 23860
rect 29000 23808 29052 23860
rect 29920 23808 29972 23860
rect 32312 23808 32364 23860
rect 22928 23740 22980 23792
rect 24584 23740 24636 23792
rect 25320 23740 25372 23792
rect 33784 23740 33836 23792
rect 38200 23808 38252 23860
rect 40960 23851 41012 23860
rect 40960 23817 40969 23851
rect 40969 23817 41003 23851
rect 41003 23817 41012 23851
rect 40960 23808 41012 23817
rect 41328 23851 41380 23860
rect 41328 23817 41337 23851
rect 41337 23817 41371 23851
rect 41371 23817 41380 23851
rect 41328 23808 41380 23817
rect 35164 23740 35216 23792
rect 37740 23740 37792 23792
rect 20168 23715 20220 23724
rect 20168 23681 20177 23715
rect 20177 23681 20211 23715
rect 20211 23681 20220 23715
rect 20168 23672 20220 23681
rect 21088 23672 21140 23724
rect 26424 23672 26476 23724
rect 28264 23672 28316 23724
rect 29000 23715 29052 23724
rect 29000 23681 29009 23715
rect 29009 23681 29043 23715
rect 29043 23681 29052 23715
rect 29000 23672 29052 23681
rect 16580 23604 16632 23656
rect 20536 23604 20588 23656
rect 21364 23647 21416 23656
rect 21364 23613 21373 23647
rect 21373 23613 21407 23647
rect 21407 23613 21416 23647
rect 21364 23604 21416 23613
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 16672 23536 16724 23588
rect 17960 23536 18012 23588
rect 21916 23536 21968 23588
rect 25780 23604 25832 23656
rect 25872 23647 25924 23656
rect 25872 23613 25881 23647
rect 25881 23613 25915 23647
rect 25915 23613 25924 23647
rect 25872 23604 25924 23613
rect 23572 23536 23624 23588
rect 28816 23604 28868 23656
rect 19708 23468 19760 23520
rect 20076 23468 20128 23520
rect 21088 23468 21140 23520
rect 22008 23511 22060 23520
rect 22008 23477 22017 23511
rect 22017 23477 22051 23511
rect 22051 23477 22060 23511
rect 22008 23468 22060 23477
rect 24860 23468 24912 23520
rect 26700 23468 26752 23520
rect 27436 23468 27488 23520
rect 29000 23536 29052 23588
rect 30932 23647 30984 23656
rect 30932 23613 30941 23647
rect 30941 23613 30975 23647
rect 30975 23613 30984 23647
rect 30932 23604 30984 23613
rect 32312 23715 32364 23724
rect 32312 23681 32321 23715
rect 32321 23681 32355 23715
rect 32355 23681 32364 23715
rect 32312 23672 32364 23681
rect 32404 23715 32456 23724
rect 32404 23681 32413 23715
rect 32413 23681 32447 23715
rect 32447 23681 32456 23715
rect 32404 23672 32456 23681
rect 32496 23715 32548 23724
rect 32496 23681 32505 23715
rect 32505 23681 32539 23715
rect 32539 23681 32548 23715
rect 32496 23672 32548 23681
rect 35348 23672 35400 23724
rect 38292 23672 38344 23724
rect 39396 23715 39448 23724
rect 39396 23681 39405 23715
rect 39405 23681 39439 23715
rect 39439 23681 39448 23715
rect 39396 23672 39448 23681
rect 39672 23715 39724 23724
rect 39672 23681 39706 23715
rect 39706 23681 39724 23715
rect 39672 23672 39724 23681
rect 34520 23604 34572 23656
rect 38568 23647 38620 23656
rect 38568 23613 38577 23647
rect 38577 23613 38611 23647
rect 38611 23613 38620 23647
rect 38568 23604 38620 23613
rect 41420 23647 41472 23656
rect 41420 23613 41429 23647
rect 41429 23613 41463 23647
rect 41463 23613 41472 23647
rect 41420 23604 41472 23613
rect 41512 23647 41564 23656
rect 41512 23613 41521 23647
rect 41521 23613 41555 23647
rect 41555 23613 41564 23647
rect 41512 23604 41564 23613
rect 29920 23536 29972 23588
rect 32404 23536 32456 23588
rect 38384 23536 38436 23588
rect 28908 23468 28960 23520
rect 30012 23511 30064 23520
rect 30012 23477 30021 23511
rect 30021 23477 30055 23511
rect 30055 23477 30064 23511
rect 30012 23468 30064 23477
rect 33324 23468 33376 23520
rect 34704 23511 34756 23520
rect 34704 23477 34713 23511
rect 34713 23477 34747 23511
rect 34747 23477 34756 23511
rect 34704 23468 34756 23477
rect 37924 23468 37976 23520
rect 40776 23511 40828 23520
rect 40776 23477 40785 23511
rect 40785 23477 40819 23511
rect 40819 23477 40828 23511
rect 40776 23468 40828 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3240 23264 3292 23316
rect 6460 23264 6512 23316
rect 7196 23264 7248 23316
rect 7748 23264 7800 23316
rect 8208 23264 8260 23316
rect 9864 23264 9916 23316
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 13728 23264 13780 23316
rect 3700 23196 3752 23248
rect 8300 23196 8352 23248
rect 12716 23196 12768 23248
rect 15660 23264 15712 23316
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2780 23128 2832 23180
rect 3240 23060 3292 23112
rect 3148 22992 3200 23044
rect 4620 23128 4672 23180
rect 4988 23128 5040 23180
rect 10508 23171 10560 23180
rect 3608 23103 3660 23112
rect 3608 23069 3617 23103
rect 3617 23069 3651 23103
rect 3651 23069 3660 23103
rect 3608 23060 3660 23069
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 5080 22992 5132 23044
rect 5908 22992 5960 23044
rect 6460 23103 6512 23112
rect 6460 23069 6469 23103
rect 6469 23069 6503 23103
rect 6503 23069 6512 23103
rect 6460 23060 6512 23069
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 7012 23060 7064 23112
rect 6736 22992 6788 23044
rect 7104 23035 7156 23044
rect 7104 23001 7113 23035
rect 7113 23001 7147 23035
rect 7147 23001 7156 23035
rect 7104 22992 7156 23001
rect 7196 22992 7248 23044
rect 7656 23103 7708 23112
rect 7656 23069 7665 23103
rect 7665 23069 7699 23103
rect 7699 23069 7708 23103
rect 7656 23060 7708 23069
rect 7932 23103 7984 23112
rect 7932 23069 7941 23103
rect 7941 23069 7975 23103
rect 7975 23069 7984 23103
rect 7932 23060 7984 23069
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 12440 23128 12492 23180
rect 12992 23128 13044 23180
rect 15936 23196 15988 23248
rect 848 22924 900 22976
rect 5632 22924 5684 22976
rect 6920 22924 6972 22976
rect 7380 22924 7432 22976
rect 8392 23035 8444 23044
rect 8392 23001 8401 23035
rect 8401 23001 8435 23035
rect 8435 23001 8444 23035
rect 8392 22992 8444 23001
rect 8668 22924 8720 22976
rect 9312 23060 9364 23112
rect 11060 23060 11112 23112
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 15200 23103 15252 23112
rect 15200 23069 15218 23103
rect 15218 23069 15252 23103
rect 15200 23060 15252 23069
rect 9128 22992 9180 23044
rect 11428 22924 11480 22976
rect 18604 23264 18656 23316
rect 23112 23264 23164 23316
rect 23296 23264 23348 23316
rect 28264 23264 28316 23316
rect 17224 23196 17276 23248
rect 17592 23128 17644 23180
rect 11888 22967 11940 22976
rect 11888 22933 11897 22967
rect 11897 22933 11931 22967
rect 11931 22933 11940 22967
rect 11888 22924 11940 22933
rect 13268 22924 13320 22976
rect 14832 22924 14884 22976
rect 17500 23103 17552 23112
rect 17500 23069 17509 23103
rect 17509 23069 17543 23103
rect 17543 23069 17552 23103
rect 17500 23060 17552 23069
rect 19800 23103 19852 23112
rect 19800 23069 19809 23103
rect 19809 23069 19843 23103
rect 19843 23069 19852 23103
rect 19800 23060 19852 23069
rect 19892 23060 19944 23112
rect 27436 23171 27488 23180
rect 27436 23137 27445 23171
rect 27445 23137 27479 23171
rect 27479 23137 27488 23171
rect 27436 23128 27488 23137
rect 26424 23060 26476 23112
rect 26976 23103 27028 23112
rect 26976 23069 26994 23103
rect 26994 23069 27028 23103
rect 26976 23060 27028 23069
rect 22008 22992 22060 23044
rect 24492 22992 24544 23044
rect 25964 22992 26016 23044
rect 28264 23035 28316 23044
rect 28264 23001 28273 23035
rect 28273 23001 28307 23035
rect 28307 23001 28316 23035
rect 28264 22992 28316 23001
rect 28908 23103 28960 23112
rect 28908 23069 28917 23103
rect 28917 23069 28951 23103
rect 28951 23069 28960 23103
rect 28908 23060 28960 23069
rect 29000 23060 29052 23112
rect 30104 23060 30156 23112
rect 17684 22924 17736 22976
rect 22836 22924 22888 22976
rect 25780 22967 25832 22976
rect 25780 22933 25789 22967
rect 25789 22933 25823 22967
rect 25823 22933 25832 22967
rect 25780 22924 25832 22933
rect 25872 22967 25924 22976
rect 25872 22933 25881 22967
rect 25881 22933 25915 22967
rect 25915 22933 25924 22967
rect 25872 22924 25924 22933
rect 29184 22992 29236 23044
rect 30012 22992 30064 23044
rect 30932 23307 30984 23316
rect 30932 23273 30941 23307
rect 30941 23273 30975 23307
rect 30975 23273 30984 23307
rect 30932 23264 30984 23273
rect 32036 23264 32088 23316
rect 31668 23171 31720 23180
rect 31668 23137 31677 23171
rect 31677 23137 31711 23171
rect 31711 23137 31720 23171
rect 31668 23128 31720 23137
rect 34796 23264 34848 23316
rect 36084 23264 36136 23316
rect 36452 23264 36504 23316
rect 38292 23264 38344 23316
rect 39672 23264 39724 23316
rect 41420 23264 41472 23316
rect 38660 23128 38712 23180
rect 40776 23171 40828 23180
rect 40776 23137 40785 23171
rect 40785 23137 40819 23171
rect 40819 23137 40828 23171
rect 40776 23128 40828 23137
rect 42064 23171 42116 23180
rect 42064 23137 42073 23171
rect 42073 23137 42107 23171
rect 42107 23137 42116 23171
rect 42064 23128 42116 23137
rect 32496 23060 32548 23112
rect 31208 23035 31260 23044
rect 31208 23001 31217 23035
rect 31217 23001 31251 23035
rect 31251 23001 31260 23035
rect 31208 22992 31260 23001
rect 28816 22924 28868 22976
rect 31392 22924 31444 22976
rect 33324 22992 33376 23044
rect 34888 23060 34940 23112
rect 37924 23103 37976 23112
rect 37924 23069 37958 23103
rect 37958 23069 37976 23103
rect 37924 23060 37976 23069
rect 40040 23060 40092 23112
rect 35440 22992 35492 23044
rect 37004 22992 37056 23044
rect 41972 22992 42024 23044
rect 32772 22924 32824 22976
rect 34520 22967 34572 22976
rect 34520 22933 34529 22967
rect 34529 22933 34563 22967
rect 34563 22933 34572 22967
rect 34520 22924 34572 22933
rect 35348 22967 35400 22976
rect 35348 22933 35357 22967
rect 35357 22933 35391 22967
rect 35391 22933 35400 22967
rect 35348 22924 35400 22933
rect 39028 22967 39080 22976
rect 39028 22933 39037 22967
rect 39037 22933 39071 22967
rect 39071 22933 39080 22967
rect 39028 22924 39080 22933
rect 41052 22924 41104 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 1400 22763 1452 22772
rect 1400 22729 1409 22763
rect 1409 22729 1443 22763
rect 1443 22729 1452 22763
rect 1400 22720 1452 22729
rect 5264 22720 5316 22772
rect 6920 22720 6972 22772
rect 7380 22720 7432 22772
rect 8484 22720 8536 22772
rect 9128 22720 9180 22772
rect 3148 22652 3200 22704
rect 3976 22652 4028 22704
rect 1768 22584 1820 22636
rect 4620 22584 4672 22636
rect 4712 22627 4764 22636
rect 4712 22593 4721 22627
rect 4721 22593 4755 22627
rect 4755 22593 4764 22627
rect 4712 22584 4764 22593
rect 5908 22652 5960 22704
rect 3148 22559 3200 22568
rect 3148 22525 3157 22559
rect 3157 22525 3191 22559
rect 3191 22525 3200 22559
rect 3148 22516 3200 22525
rect 5540 22584 5592 22636
rect 5724 22584 5776 22636
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 7288 22584 7340 22636
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 7472 22584 7524 22636
rect 8392 22652 8444 22704
rect 9312 22695 9364 22704
rect 9312 22661 9321 22695
rect 9321 22661 9355 22695
rect 9355 22661 9364 22695
rect 9312 22652 9364 22661
rect 9772 22720 9824 22772
rect 13268 22763 13320 22772
rect 13268 22729 13277 22763
rect 13277 22729 13311 22763
rect 13311 22729 13320 22763
rect 13268 22720 13320 22729
rect 11888 22652 11940 22704
rect 16672 22652 16724 22704
rect 17500 22652 17552 22704
rect 18144 22652 18196 22704
rect 7012 22516 7064 22568
rect 7656 22559 7708 22568
rect 7656 22525 7665 22559
rect 7665 22525 7699 22559
rect 7699 22525 7708 22559
rect 7656 22516 7708 22525
rect 7748 22559 7800 22568
rect 7748 22525 7757 22559
rect 7757 22525 7791 22559
rect 7791 22525 7800 22559
rect 7748 22516 7800 22525
rect 7932 22448 7984 22500
rect 4804 22380 4856 22432
rect 4988 22423 5040 22432
rect 4988 22389 4997 22423
rect 4997 22389 5031 22423
rect 5031 22389 5040 22423
rect 4988 22380 5040 22389
rect 5080 22380 5132 22432
rect 5356 22423 5408 22432
rect 5356 22389 5365 22423
rect 5365 22389 5399 22423
rect 5399 22389 5408 22423
rect 5356 22380 5408 22389
rect 7012 22380 7064 22432
rect 7196 22380 7248 22432
rect 7748 22380 7800 22432
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 11428 22584 11480 22636
rect 11520 22627 11572 22636
rect 11520 22593 11529 22627
rect 11529 22593 11563 22627
rect 11563 22593 11572 22627
rect 11520 22584 11572 22593
rect 12900 22584 12952 22636
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 17408 22584 17460 22636
rect 17684 22627 17736 22636
rect 17684 22593 17693 22627
rect 17693 22593 17727 22627
rect 17727 22593 17736 22627
rect 17684 22584 17736 22593
rect 18236 22584 18288 22636
rect 19616 22720 19668 22772
rect 19800 22720 19852 22772
rect 20720 22720 20772 22772
rect 21364 22720 21416 22772
rect 32036 22720 32088 22772
rect 34888 22720 34940 22772
rect 35440 22720 35492 22772
rect 41052 22763 41104 22772
rect 41052 22729 41061 22763
rect 41061 22729 41095 22763
rect 41095 22729 41104 22763
rect 41052 22720 41104 22729
rect 41972 22720 42024 22772
rect 26332 22652 26384 22704
rect 20076 22627 20128 22636
rect 20076 22593 20110 22627
rect 20110 22593 20128 22627
rect 20076 22584 20128 22593
rect 26424 22584 26476 22636
rect 27436 22652 27488 22704
rect 30840 22652 30892 22704
rect 34704 22652 34756 22704
rect 27252 22627 27304 22636
rect 27252 22593 27286 22627
rect 27286 22593 27304 22627
rect 27252 22584 27304 22593
rect 30932 22584 30984 22636
rect 35532 22652 35584 22704
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 14832 22559 14884 22568
rect 14832 22525 14841 22559
rect 14841 22525 14875 22559
rect 14875 22525 14884 22559
rect 14832 22516 14884 22525
rect 17592 22516 17644 22568
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 15108 22423 15160 22432
rect 15108 22389 15117 22423
rect 15117 22389 15151 22423
rect 15151 22389 15160 22423
rect 15108 22380 15160 22389
rect 16672 22423 16724 22432
rect 16672 22389 16681 22423
rect 16681 22389 16715 22423
rect 16715 22389 16724 22423
rect 16672 22380 16724 22389
rect 22100 22516 22152 22568
rect 19800 22380 19852 22432
rect 22560 22380 22612 22432
rect 22928 22380 22980 22432
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 26516 22516 26568 22568
rect 26792 22516 26844 22568
rect 25964 22380 26016 22432
rect 28356 22423 28408 22432
rect 28356 22389 28365 22423
rect 28365 22389 28399 22423
rect 28399 22389 28408 22423
rect 28356 22380 28408 22389
rect 29460 22516 29512 22568
rect 30104 22516 30156 22568
rect 32772 22559 32824 22568
rect 32772 22525 32781 22559
rect 32781 22525 32815 22559
rect 32815 22525 32824 22559
rect 32772 22516 32824 22525
rect 37280 22627 37332 22636
rect 37280 22593 37289 22627
rect 37289 22593 37323 22627
rect 37323 22593 37332 22627
rect 37280 22584 37332 22593
rect 37556 22627 37608 22636
rect 37556 22593 37590 22627
rect 37590 22593 37608 22627
rect 37556 22584 37608 22593
rect 39856 22652 39908 22704
rect 41604 22652 41656 22704
rect 39580 22627 39632 22636
rect 39580 22593 39614 22627
rect 39614 22593 39632 22627
rect 39580 22584 39632 22593
rect 41696 22584 41748 22636
rect 36912 22559 36964 22568
rect 36912 22525 36921 22559
rect 36921 22525 36955 22559
rect 36955 22525 36964 22559
rect 36912 22516 36964 22525
rect 40776 22516 40828 22568
rect 30104 22380 30156 22432
rect 30656 22380 30708 22432
rect 32036 22380 32088 22432
rect 34796 22380 34848 22432
rect 38660 22423 38712 22432
rect 38660 22389 38669 22423
rect 38669 22389 38703 22423
rect 38703 22389 38712 22423
rect 38660 22380 38712 22389
rect 40684 22423 40736 22432
rect 40684 22389 40693 22423
rect 40693 22389 40727 22423
rect 40727 22389 40736 22423
rect 40684 22380 40736 22389
rect 41512 22423 41564 22432
rect 41512 22389 41521 22423
rect 41521 22389 41555 22423
rect 41555 22389 41564 22423
rect 41512 22380 41564 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3056 22176 3108 22228
rect 4712 22176 4764 22228
rect 5356 22176 5408 22228
rect 7012 22108 7064 22160
rect 4344 22040 4396 22092
rect 4620 22040 4672 22092
rect 7104 22083 7156 22092
rect 7104 22049 7113 22083
rect 7113 22049 7147 22083
rect 7147 22049 7156 22083
rect 7104 22040 7156 22049
rect 7288 22083 7340 22092
rect 7288 22049 7297 22083
rect 7297 22049 7331 22083
rect 7331 22049 7340 22083
rect 7288 22040 7340 22049
rect 8024 22083 8076 22092
rect 8024 22049 8033 22083
rect 8033 22049 8067 22083
rect 8067 22049 8076 22083
rect 8024 22040 8076 22049
rect 1768 21972 1820 22024
rect 3148 22015 3200 22024
rect 3148 21981 3157 22015
rect 3157 21981 3191 22015
rect 3191 21981 3200 22015
rect 3148 21972 3200 21981
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 7196 21972 7248 22024
rect 4252 21947 4304 21956
rect 4252 21913 4261 21947
rect 4261 21913 4295 21947
rect 4295 21913 4304 21947
rect 4252 21904 4304 21913
rect 1400 21879 1452 21888
rect 1400 21845 1409 21879
rect 1409 21845 1443 21879
rect 1443 21845 1452 21879
rect 1400 21836 1452 21845
rect 3700 21836 3752 21888
rect 7472 21972 7524 22024
rect 7840 22015 7892 22024
rect 7840 21981 7849 22015
rect 7849 21981 7883 22015
rect 7883 21981 7892 22015
rect 7840 21972 7892 21981
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 9312 22176 9364 22228
rect 4620 21836 4672 21888
rect 4988 21836 5040 21888
rect 6552 21836 6604 21888
rect 8576 22015 8628 22024
rect 8576 21981 8585 22015
rect 8585 21981 8619 22015
rect 8619 21981 8628 22015
rect 8576 21972 8628 21981
rect 9772 21972 9824 22024
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 18328 22176 18380 22228
rect 15108 22108 15160 22160
rect 17776 22108 17828 22160
rect 20168 22176 20220 22228
rect 27252 22176 27304 22228
rect 29460 22176 29512 22228
rect 30932 22219 30984 22228
rect 30932 22185 30941 22219
rect 30941 22185 30975 22219
rect 30975 22185 30984 22219
rect 30932 22176 30984 22185
rect 34796 22176 34848 22228
rect 35348 22176 35400 22228
rect 37556 22176 37608 22228
rect 15476 22083 15528 22092
rect 15476 22049 15485 22083
rect 15485 22049 15519 22083
rect 15519 22049 15528 22083
rect 15476 22040 15528 22049
rect 16672 21972 16724 22024
rect 16764 22015 16816 22024
rect 16764 21981 16773 22015
rect 16773 21981 16807 22015
rect 16807 21981 16816 22015
rect 16764 21972 16816 21981
rect 19800 22083 19852 22092
rect 19800 22049 19809 22083
rect 19809 22049 19843 22083
rect 19843 22049 19852 22083
rect 19800 22040 19852 22049
rect 21916 22083 21968 22092
rect 21916 22049 21925 22083
rect 21925 22049 21959 22083
rect 21959 22049 21968 22083
rect 21916 22040 21968 22049
rect 24676 22108 24728 22160
rect 22836 22040 22888 22092
rect 26332 22040 26384 22092
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 28816 22108 28868 22160
rect 31208 22108 31260 22160
rect 28356 22040 28408 22092
rect 30012 22083 30064 22092
rect 30012 22049 30021 22083
rect 30021 22049 30055 22083
rect 30055 22049 30064 22083
rect 30012 22040 30064 22049
rect 31392 22040 31444 22092
rect 17500 21972 17552 22024
rect 18604 22015 18656 22024
rect 18604 21981 18613 22015
rect 18613 21981 18647 22015
rect 18647 21981 18656 22015
rect 18604 21972 18656 21981
rect 21640 22015 21692 22024
rect 21640 21981 21649 22015
rect 21649 21981 21683 22015
rect 21683 21981 21692 22015
rect 21640 21972 21692 21981
rect 22468 22015 22520 22024
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22468 21972 22520 21981
rect 25780 21972 25832 22024
rect 25964 21972 26016 22024
rect 8484 21947 8536 21956
rect 8484 21913 8493 21947
rect 8493 21913 8527 21947
rect 8527 21913 8536 21947
rect 8484 21904 8536 21913
rect 12164 21947 12216 21956
rect 12164 21913 12173 21947
rect 12173 21913 12207 21947
rect 12207 21913 12216 21947
rect 12164 21904 12216 21913
rect 12900 21904 12952 21956
rect 13912 21947 13964 21956
rect 13912 21913 13921 21947
rect 13921 21913 13955 21947
rect 13955 21913 13964 21947
rect 13912 21904 13964 21913
rect 10508 21879 10560 21888
rect 10508 21845 10517 21879
rect 10517 21845 10551 21879
rect 10551 21845 10560 21879
rect 10508 21836 10560 21845
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15292 21836 15344 21888
rect 16580 21836 16632 21888
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 21180 21879 21232 21888
rect 21180 21845 21189 21879
rect 21189 21845 21223 21879
rect 21223 21845 21232 21879
rect 21180 21836 21232 21845
rect 22560 21947 22612 21956
rect 22560 21913 22569 21947
rect 22569 21913 22603 21947
rect 22603 21913 22612 21947
rect 22560 21904 22612 21913
rect 24308 21904 24360 21956
rect 27712 22015 27764 22024
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 31300 22015 31352 22024
rect 31300 21981 31309 22015
rect 31309 21981 31343 22015
rect 31343 21981 31352 22015
rect 31300 21972 31352 21981
rect 32036 22040 32088 22092
rect 33140 22108 33192 22160
rect 32312 21904 32364 21956
rect 33876 22040 33928 22092
rect 33508 21972 33560 22024
rect 35532 21972 35584 22024
rect 35256 21947 35308 21956
rect 35256 21913 35290 21947
rect 35290 21913 35308 21947
rect 35256 21904 35308 21913
rect 21732 21879 21784 21888
rect 21732 21845 21741 21879
rect 21741 21845 21775 21879
rect 21775 21845 21784 21879
rect 21732 21836 21784 21845
rect 24216 21836 24268 21888
rect 24952 21879 25004 21888
rect 24952 21845 24961 21879
rect 24961 21845 24995 21879
rect 24995 21845 25004 21879
rect 24952 21836 25004 21845
rect 25688 21879 25740 21888
rect 25688 21845 25697 21879
rect 25697 21845 25731 21879
rect 25731 21845 25740 21879
rect 25688 21836 25740 21845
rect 28172 21879 28224 21888
rect 28172 21845 28181 21879
rect 28181 21845 28215 21879
rect 28215 21845 28224 21879
rect 28172 21836 28224 21845
rect 29920 21879 29972 21888
rect 29920 21845 29929 21879
rect 29929 21845 29963 21879
rect 29963 21845 29972 21879
rect 29920 21836 29972 21845
rect 31300 21836 31352 21888
rect 32588 21879 32640 21888
rect 32588 21845 32597 21879
rect 32597 21845 32631 21879
rect 32631 21845 32640 21879
rect 32588 21836 32640 21845
rect 33232 21836 33284 21888
rect 33600 21836 33652 21888
rect 36084 21836 36136 21888
rect 38292 22083 38344 22092
rect 38292 22049 38301 22083
rect 38301 22049 38335 22083
rect 38335 22049 38344 22083
rect 38292 22040 38344 22049
rect 38568 22040 38620 22092
rect 38660 22040 38712 22092
rect 41144 22040 41196 22092
rect 41696 22040 41748 22092
rect 41880 22040 41932 22092
rect 38016 21972 38068 22024
rect 39856 21972 39908 22024
rect 40224 22015 40276 22024
rect 40224 21981 40233 22015
rect 40233 21981 40267 22015
rect 40267 21981 40276 22015
rect 40224 21972 40276 21981
rect 36452 21879 36504 21888
rect 36452 21845 36461 21879
rect 36461 21845 36495 21879
rect 36495 21845 36504 21879
rect 36452 21836 36504 21845
rect 37648 21836 37700 21888
rect 40592 21904 40644 21956
rect 40776 21836 40828 21888
rect 41420 21836 41472 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 1308 21632 1360 21684
rect 4344 21675 4396 21684
rect 4344 21641 4353 21675
rect 4353 21641 4387 21675
rect 4387 21641 4396 21675
rect 4344 21632 4396 21641
rect 7840 21632 7892 21684
rect 12164 21632 12216 21684
rect 13912 21632 13964 21684
rect 3608 21564 3660 21616
rect 4620 21564 4672 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 3976 21496 4028 21548
rect 6000 21564 6052 21616
rect 8576 21564 8628 21616
rect 12900 21564 12952 21616
rect 14924 21632 14976 21684
rect 14188 21564 14240 21616
rect 15292 21564 15344 21616
rect 17408 21632 17460 21684
rect 20168 21632 20220 21684
rect 21456 21564 21508 21616
rect 24308 21675 24360 21684
rect 24308 21641 24317 21675
rect 24317 21641 24351 21675
rect 24351 21641 24360 21675
rect 24308 21632 24360 21641
rect 24492 21632 24544 21684
rect 28172 21675 28224 21684
rect 28172 21641 28181 21675
rect 28181 21641 28215 21675
rect 28215 21641 28224 21675
rect 28172 21632 28224 21641
rect 29920 21632 29972 21684
rect 31300 21675 31352 21684
rect 31300 21641 31309 21675
rect 31309 21641 31343 21675
rect 31343 21641 31352 21675
rect 31300 21632 31352 21641
rect 33508 21675 33560 21684
rect 33508 21641 33517 21675
rect 33517 21641 33551 21675
rect 33551 21641 33560 21675
rect 33508 21632 33560 21641
rect 33876 21632 33928 21684
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 7012 21496 7064 21548
rect 8116 21496 8168 21548
rect 10508 21496 10560 21548
rect 14556 21539 14608 21548
rect 14556 21505 14565 21539
rect 14565 21505 14599 21539
rect 14599 21505 14608 21539
rect 14556 21496 14608 21505
rect 21180 21496 21232 21548
rect 6552 21428 6604 21480
rect 8024 21428 8076 21480
rect 12992 21471 13044 21480
rect 12992 21437 13001 21471
rect 13001 21437 13035 21471
rect 13035 21437 13044 21471
rect 12992 21428 13044 21437
rect 13820 21428 13872 21480
rect 16764 21428 16816 21480
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 18144 21428 18196 21480
rect 1032 21360 1084 21412
rect 4252 21360 4304 21412
rect 19892 21360 19944 21412
rect 21640 21471 21692 21480
rect 21640 21437 21649 21471
rect 21649 21437 21683 21471
rect 21683 21437 21692 21471
rect 21640 21428 21692 21437
rect 22192 21496 22244 21548
rect 22928 21539 22980 21548
rect 22928 21505 22937 21539
rect 22937 21505 22971 21539
rect 22971 21505 22980 21539
rect 22928 21496 22980 21505
rect 23480 21496 23532 21548
rect 24400 21496 24452 21548
rect 24584 21539 24636 21548
rect 24584 21505 24593 21539
rect 24593 21505 24627 21539
rect 24627 21505 24636 21539
rect 24584 21496 24636 21505
rect 25044 21564 25096 21616
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 26424 21564 26476 21616
rect 32588 21564 32640 21616
rect 33784 21564 33836 21616
rect 35256 21675 35308 21684
rect 35256 21641 35265 21675
rect 35265 21641 35299 21675
rect 35299 21641 35308 21675
rect 35256 21632 35308 21641
rect 39580 21632 39632 21684
rect 39764 21632 39816 21684
rect 25596 21496 25648 21548
rect 30656 21539 30708 21548
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 31944 21496 31996 21548
rect 34336 21564 34388 21616
rect 35992 21564 36044 21616
rect 40592 21564 40644 21616
rect 41328 21564 41380 21616
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 27252 21428 27304 21480
rect 28908 21428 28960 21480
rect 31392 21471 31444 21480
rect 31392 21437 31401 21471
rect 31401 21437 31435 21471
rect 31435 21437 31444 21471
rect 31392 21428 31444 21437
rect 32128 21471 32180 21480
rect 32128 21437 32137 21471
rect 32137 21437 32171 21471
rect 32171 21437 32180 21471
rect 32128 21428 32180 21437
rect 4528 21335 4580 21344
rect 4528 21301 4537 21335
rect 4537 21301 4571 21335
rect 4571 21301 4580 21335
rect 4528 21292 4580 21301
rect 6920 21292 6972 21344
rect 7564 21335 7616 21344
rect 7564 21301 7573 21335
rect 7573 21301 7607 21335
rect 7607 21301 7616 21335
rect 7564 21292 7616 21301
rect 14096 21292 14148 21344
rect 18144 21292 18196 21344
rect 18696 21292 18748 21344
rect 19708 21335 19760 21344
rect 19708 21301 19717 21335
rect 19717 21301 19751 21335
rect 19751 21301 19760 21335
rect 19708 21292 19760 21301
rect 20812 21292 20864 21344
rect 21180 21292 21232 21344
rect 21732 21292 21784 21344
rect 22100 21292 22152 21344
rect 23204 21292 23256 21344
rect 24676 21292 24728 21344
rect 25228 21292 25280 21344
rect 27252 21292 27304 21344
rect 27528 21292 27580 21344
rect 27712 21335 27764 21344
rect 27712 21301 27721 21335
rect 27721 21301 27755 21335
rect 27755 21301 27764 21335
rect 27712 21292 27764 21301
rect 30380 21292 30432 21344
rect 35348 21496 35400 21548
rect 35624 21539 35676 21548
rect 35624 21505 35633 21539
rect 35633 21505 35667 21539
rect 35667 21505 35676 21539
rect 35624 21496 35676 21505
rect 36452 21496 36504 21548
rect 40132 21496 40184 21548
rect 34704 21428 34756 21480
rect 37280 21471 37332 21480
rect 37280 21437 37289 21471
rect 37289 21437 37323 21471
rect 37323 21437 37332 21471
rect 37280 21428 37332 21437
rect 37556 21471 37608 21480
rect 37556 21437 37565 21471
rect 37565 21437 37599 21471
rect 37599 21437 37608 21471
rect 37556 21428 37608 21437
rect 37924 21428 37976 21480
rect 38292 21428 38344 21480
rect 40224 21428 40276 21480
rect 36912 21360 36964 21412
rect 39212 21360 39264 21412
rect 40592 21471 40644 21480
rect 40592 21437 40601 21471
rect 40601 21437 40635 21471
rect 40635 21437 40644 21471
rect 40592 21428 40644 21437
rect 34336 21292 34388 21344
rect 35624 21292 35676 21344
rect 37924 21292 37976 21344
rect 38568 21292 38620 21344
rect 42064 21335 42116 21344
rect 42064 21301 42073 21335
rect 42073 21301 42107 21335
rect 42107 21301 42116 21335
rect 42064 21292 42116 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1768 21088 1820 21140
rect 4896 21088 4948 21140
rect 2872 20995 2924 21004
rect 2872 20961 2881 20995
rect 2881 20961 2915 20995
rect 2915 20961 2924 20995
rect 2872 20952 2924 20961
rect 3148 20927 3200 20936
rect 3148 20893 3157 20927
rect 3157 20893 3191 20927
rect 3191 20893 3200 20927
rect 3148 20884 3200 20893
rect 3884 20884 3936 20936
rect 4712 20952 4764 21004
rect 4160 20884 4212 20936
rect 1860 20816 1912 20868
rect 4804 20884 4856 20936
rect 4896 20927 4948 20936
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 11152 21131 11204 21140
rect 11152 21097 11161 21131
rect 11161 21097 11195 21131
rect 11195 21097 11204 21131
rect 11152 21088 11204 21097
rect 16580 21131 16632 21140
rect 16580 21097 16589 21131
rect 16589 21097 16623 21131
rect 16623 21097 16632 21131
rect 16580 21088 16632 21097
rect 17408 21088 17460 21140
rect 15476 21020 15528 21072
rect 17868 21020 17920 21072
rect 6368 20952 6420 21004
rect 11888 20952 11940 21004
rect 13820 20952 13872 21004
rect 14832 20952 14884 21004
rect 18144 20995 18196 21004
rect 18144 20961 18153 20995
rect 18153 20961 18187 20995
rect 18187 20961 18196 20995
rect 18144 20952 18196 20961
rect 18236 20995 18288 21004
rect 18236 20961 18245 20995
rect 18245 20961 18279 20995
rect 18279 20961 18288 20995
rect 18236 20952 18288 20961
rect 3332 20748 3384 20800
rect 5356 20884 5408 20936
rect 16580 20884 16632 20936
rect 20996 21088 21048 21140
rect 22284 21088 22336 21140
rect 23480 21131 23532 21140
rect 23480 21097 23489 21131
rect 23489 21097 23523 21131
rect 23523 21097 23532 21131
rect 23480 21088 23532 21097
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 19156 20952 19208 21004
rect 21180 21020 21232 21072
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 20812 20927 20864 20936
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 6644 20816 6696 20868
rect 7564 20816 7616 20868
rect 10968 20859 11020 20868
rect 10968 20825 10977 20859
rect 10977 20825 11011 20859
rect 11011 20825 11020 20859
rect 10968 20816 11020 20825
rect 12164 20816 12216 20868
rect 14924 20816 14976 20868
rect 19708 20816 19760 20868
rect 22192 20952 22244 21004
rect 25688 21020 25740 21072
rect 23756 20884 23808 20936
rect 25228 20952 25280 21004
rect 28908 21131 28960 21140
rect 28908 21097 28917 21131
rect 28917 21097 28951 21131
rect 28951 21097 28960 21131
rect 28908 21088 28960 21097
rect 28724 21020 28776 21072
rect 27436 20952 27488 21004
rect 30104 20995 30156 21004
rect 30104 20961 30113 20995
rect 30113 20961 30147 20995
rect 30147 20961 30156 20995
rect 30104 20952 30156 20961
rect 30380 20995 30432 21004
rect 30380 20961 30389 20995
rect 30389 20961 30423 20995
rect 30423 20961 30432 20995
rect 30380 20952 30432 20961
rect 31944 21131 31996 21140
rect 31944 21097 31953 21131
rect 31953 21097 31987 21131
rect 31987 21097 31996 21131
rect 31944 21088 31996 21097
rect 35624 21088 35676 21140
rect 37556 21088 37608 21140
rect 40592 21088 40644 21140
rect 41144 21088 41196 21140
rect 31484 21020 31536 21072
rect 33600 21020 33652 21072
rect 11336 20791 11388 20800
rect 11336 20757 11345 20791
rect 11345 20757 11379 20791
rect 11379 20757 11388 20791
rect 11336 20748 11388 20757
rect 17132 20748 17184 20800
rect 18236 20748 18288 20800
rect 21548 20859 21600 20868
rect 21548 20825 21557 20859
rect 21557 20825 21591 20859
rect 21591 20825 21600 20859
rect 21548 20816 21600 20825
rect 22100 20816 22152 20868
rect 19984 20791 20036 20800
rect 19984 20757 19993 20791
rect 19993 20757 20027 20791
rect 20027 20757 20036 20791
rect 19984 20748 20036 20757
rect 20444 20791 20496 20800
rect 20444 20757 20453 20791
rect 20453 20757 20487 20791
rect 20487 20757 20496 20791
rect 20444 20748 20496 20757
rect 21916 20748 21968 20800
rect 26792 20884 26844 20936
rect 26976 20927 27028 20936
rect 26976 20893 26985 20927
rect 26985 20893 27019 20927
rect 27019 20893 27028 20927
rect 26976 20884 27028 20893
rect 34888 21020 34940 21072
rect 36728 21020 36780 21072
rect 37280 21020 37332 21072
rect 37648 20995 37700 21004
rect 37648 20961 37657 20995
rect 37657 20961 37691 20995
rect 37691 20961 37700 20995
rect 37648 20952 37700 20961
rect 38568 20952 38620 21004
rect 41512 20952 41564 21004
rect 24216 20816 24268 20868
rect 24032 20748 24084 20800
rect 27712 20816 27764 20868
rect 29460 20816 29512 20868
rect 30380 20816 30432 20868
rect 30840 20816 30892 20868
rect 24952 20748 25004 20800
rect 25596 20791 25648 20800
rect 25596 20757 25605 20791
rect 25605 20757 25639 20791
rect 25639 20757 25648 20791
rect 25596 20748 25648 20757
rect 27528 20748 27580 20800
rect 31760 20748 31812 20800
rect 33784 20884 33836 20936
rect 34060 20884 34112 20936
rect 33600 20748 33652 20800
rect 34980 20927 35032 20936
rect 34980 20893 34989 20927
rect 34989 20893 35023 20927
rect 35023 20893 35032 20927
rect 34980 20884 35032 20893
rect 35256 20884 35308 20936
rect 35348 20927 35400 20936
rect 35348 20893 35357 20927
rect 35357 20893 35391 20927
rect 35391 20893 35400 20927
rect 35348 20884 35400 20893
rect 34888 20859 34940 20868
rect 34888 20825 34897 20859
rect 34897 20825 34931 20859
rect 34931 20825 34940 20859
rect 34888 20816 34940 20825
rect 38016 20859 38068 20868
rect 38016 20825 38025 20859
rect 38025 20825 38059 20859
rect 38059 20825 38068 20859
rect 38016 20816 38068 20825
rect 39212 20816 39264 20868
rect 41512 20816 41564 20868
rect 36268 20748 36320 20800
rect 40132 20748 40184 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 1860 20544 1912 20596
rect 4620 20544 4672 20596
rect 5172 20544 5224 20596
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 5356 20544 5408 20596
rect 5816 20587 5868 20596
rect 5816 20553 5825 20587
rect 5825 20553 5859 20587
rect 5859 20553 5868 20587
rect 5816 20544 5868 20553
rect 8760 20544 8812 20596
rect 3700 20476 3752 20528
rect 2228 20408 2280 20460
rect 3148 20340 3200 20392
rect 3332 20451 3384 20460
rect 3332 20417 3341 20451
rect 3341 20417 3375 20451
rect 3375 20417 3384 20451
rect 3332 20408 3384 20417
rect 4712 20408 4764 20460
rect 5356 20451 5408 20460
rect 5356 20417 5365 20451
rect 5365 20417 5399 20451
rect 5399 20417 5408 20451
rect 5356 20408 5408 20417
rect 6092 20476 6144 20528
rect 5632 20451 5684 20460
rect 5632 20417 5641 20451
rect 5641 20417 5675 20451
rect 5675 20417 5684 20451
rect 5632 20408 5684 20417
rect 5724 20408 5776 20460
rect 14096 20544 14148 20596
rect 14556 20544 14608 20596
rect 16856 20544 16908 20596
rect 11336 20476 11388 20528
rect 13820 20476 13872 20528
rect 15200 20476 15252 20528
rect 10600 20408 10652 20460
rect 11520 20451 11572 20460
rect 11520 20417 11529 20451
rect 11529 20417 11563 20451
rect 11563 20417 11572 20451
rect 11520 20408 11572 20417
rect 11612 20408 11664 20460
rect 12992 20408 13044 20460
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 9956 20383 10008 20392
rect 9956 20349 9965 20383
rect 9965 20349 9999 20383
rect 9999 20349 10008 20383
rect 9956 20340 10008 20349
rect 10324 20383 10376 20392
rect 10324 20349 10333 20383
rect 10333 20349 10367 20383
rect 10367 20349 10376 20383
rect 10324 20340 10376 20349
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 15016 20408 15068 20460
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 4160 20272 4212 20324
rect 5448 20272 5500 20324
rect 8208 20272 8260 20324
rect 16028 20340 16080 20392
rect 17132 20383 17184 20392
rect 17132 20349 17141 20383
rect 17141 20349 17175 20383
rect 17175 20349 17184 20383
rect 17132 20340 17184 20349
rect 17776 20408 17828 20460
rect 17592 20340 17644 20392
rect 17684 20383 17736 20392
rect 17684 20349 17693 20383
rect 17693 20349 17727 20383
rect 17727 20349 17736 20383
rect 17684 20340 17736 20349
rect 5724 20204 5776 20256
rect 8484 20204 8536 20256
rect 9588 20204 9640 20256
rect 10692 20204 10744 20256
rect 10784 20204 10836 20256
rect 12900 20247 12952 20256
rect 12900 20213 12909 20247
rect 12909 20213 12943 20247
rect 12943 20213 12952 20247
rect 12900 20204 12952 20213
rect 14372 20204 14424 20256
rect 16304 20247 16356 20256
rect 16304 20213 16313 20247
rect 16313 20213 16347 20247
rect 16347 20213 16356 20247
rect 16304 20204 16356 20213
rect 16488 20204 16540 20256
rect 18604 20204 18656 20256
rect 18972 20204 19024 20256
rect 19156 20247 19208 20256
rect 19156 20213 19165 20247
rect 19165 20213 19199 20247
rect 19199 20213 19208 20247
rect 19156 20204 19208 20213
rect 22100 20544 22152 20596
rect 22284 20587 22336 20596
rect 22284 20553 22293 20587
rect 22293 20553 22327 20587
rect 22327 20553 22336 20587
rect 22284 20544 22336 20553
rect 23940 20544 23992 20596
rect 26976 20544 27028 20596
rect 27528 20544 27580 20596
rect 29368 20544 29420 20596
rect 31944 20587 31996 20596
rect 31944 20553 31953 20587
rect 31953 20553 31987 20587
rect 31987 20553 31996 20587
rect 31944 20544 31996 20553
rect 32680 20544 32732 20596
rect 33416 20544 33468 20596
rect 34060 20587 34112 20596
rect 34060 20553 34069 20587
rect 34069 20553 34103 20587
rect 34103 20553 34112 20587
rect 34060 20544 34112 20553
rect 20444 20476 20496 20528
rect 21456 20476 21508 20528
rect 21732 20476 21784 20528
rect 23204 20476 23256 20528
rect 23756 20476 23808 20528
rect 25412 20476 25464 20528
rect 29460 20476 29512 20528
rect 36728 20519 36780 20528
rect 36728 20485 36746 20519
rect 36746 20485 36780 20519
rect 36728 20476 36780 20485
rect 37464 20476 37516 20528
rect 37832 20476 37884 20528
rect 40132 20476 40184 20528
rect 41512 20587 41564 20596
rect 41512 20553 41521 20587
rect 41521 20553 41555 20587
rect 41555 20553 41564 20587
rect 41512 20544 41564 20553
rect 41696 20476 41748 20528
rect 22284 20408 22336 20460
rect 20904 20340 20956 20392
rect 21640 20383 21692 20392
rect 21640 20349 21649 20383
rect 21649 20349 21683 20383
rect 21683 20349 21692 20383
rect 21640 20340 21692 20349
rect 22376 20383 22428 20392
rect 22376 20349 22385 20383
rect 22385 20349 22419 20383
rect 22419 20349 22428 20383
rect 22376 20340 22428 20349
rect 26792 20408 26844 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27436 20408 27488 20460
rect 33876 20408 33928 20460
rect 34060 20408 34112 20460
rect 34428 20451 34480 20460
rect 34428 20417 34462 20451
rect 34462 20417 34480 20451
rect 34428 20408 34480 20417
rect 40684 20408 40736 20460
rect 21548 20272 21600 20324
rect 22100 20272 22152 20324
rect 24032 20340 24084 20392
rect 25044 20383 25096 20392
rect 25044 20349 25053 20383
rect 25053 20349 25087 20383
rect 25087 20349 25096 20383
rect 25044 20340 25096 20349
rect 27252 20340 27304 20392
rect 28448 20340 28500 20392
rect 21272 20204 21324 20256
rect 21824 20204 21876 20256
rect 23020 20204 23072 20256
rect 27160 20204 27212 20256
rect 31208 20340 31260 20392
rect 32128 20204 32180 20256
rect 32588 20383 32640 20392
rect 32588 20349 32597 20383
rect 32597 20349 32631 20383
rect 32631 20349 32640 20383
rect 32588 20340 32640 20349
rect 32772 20204 32824 20256
rect 37372 20340 37424 20392
rect 37740 20383 37792 20392
rect 37740 20349 37749 20383
rect 37749 20349 37783 20383
rect 37783 20349 37792 20383
rect 37740 20340 37792 20349
rect 35348 20272 35400 20324
rect 35532 20247 35584 20256
rect 35532 20213 35541 20247
rect 35541 20213 35575 20247
rect 35575 20213 35584 20247
rect 35532 20204 35584 20213
rect 36360 20204 36412 20256
rect 38108 20383 38160 20392
rect 38108 20349 38117 20383
rect 38117 20349 38151 20383
rect 38151 20349 38160 20383
rect 38108 20340 38160 20349
rect 39580 20383 39632 20392
rect 39580 20349 39589 20383
rect 39589 20349 39623 20383
rect 39623 20349 39632 20383
rect 39580 20340 39632 20349
rect 38476 20204 38528 20256
rect 39120 20204 39172 20256
rect 39212 20204 39264 20256
rect 40316 20340 40368 20392
rect 41788 20408 41840 20460
rect 42064 20451 42116 20460
rect 42064 20417 42073 20451
rect 42073 20417 42107 20451
rect 42107 20417 42116 20451
rect 42064 20408 42116 20417
rect 40040 20272 40092 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 5816 20000 5868 20052
rect 5724 19932 5776 19984
rect 9956 20000 10008 20052
rect 12164 20043 12216 20052
rect 12164 20009 12173 20043
rect 12173 20009 12207 20043
rect 12207 20009 12216 20043
rect 12164 20000 12216 20009
rect 16580 20000 16632 20052
rect 17776 20043 17828 20052
rect 17776 20009 17785 20043
rect 17785 20009 17819 20043
rect 17819 20009 17828 20043
rect 17776 20000 17828 20009
rect 18604 20000 18656 20052
rect 19156 20000 19208 20052
rect 22468 20000 22520 20052
rect 27068 20043 27120 20052
rect 27068 20009 27077 20043
rect 27077 20009 27111 20043
rect 27111 20009 27120 20043
rect 27068 20000 27120 20009
rect 27344 20000 27396 20052
rect 28448 20043 28500 20052
rect 28448 20009 28457 20043
rect 28457 20009 28491 20043
rect 28491 20009 28500 20043
rect 28448 20000 28500 20009
rect 31208 20043 31260 20052
rect 31208 20009 31217 20043
rect 31217 20009 31251 20043
rect 31251 20009 31260 20043
rect 31208 20000 31260 20009
rect 32588 20000 32640 20052
rect 34428 20000 34480 20052
rect 37464 20000 37516 20052
rect 39580 20000 39632 20052
rect 10508 19932 10560 19984
rect 6000 19907 6052 19916
rect 6000 19873 6009 19907
rect 6009 19873 6043 19907
rect 6043 19873 6052 19907
rect 6000 19864 6052 19873
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 8300 19864 8352 19916
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 5724 19796 5776 19848
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 2412 19728 2464 19780
rect 3148 19728 3200 19780
rect 4620 19728 4672 19780
rect 6368 19728 6420 19780
rect 6276 19703 6328 19712
rect 6276 19669 6285 19703
rect 6285 19669 6319 19703
rect 6319 19669 6328 19703
rect 6276 19660 6328 19669
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 10692 19796 10744 19848
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 16304 19864 16356 19916
rect 16672 19796 16724 19848
rect 17684 19796 17736 19848
rect 18880 19864 18932 19916
rect 25044 19864 25096 19916
rect 27436 19864 27488 19916
rect 28080 19864 28132 19916
rect 33232 19907 33284 19916
rect 33232 19873 33241 19907
rect 33241 19873 33275 19907
rect 33275 19873 33284 19907
rect 33232 19864 33284 19873
rect 33508 19864 33560 19916
rect 33784 19864 33836 19916
rect 35532 19907 35584 19916
rect 35532 19873 35541 19907
rect 35541 19873 35575 19907
rect 35575 19873 35584 19907
rect 35532 19864 35584 19873
rect 37372 19864 37424 19916
rect 13912 19728 13964 19780
rect 16488 19728 16540 19780
rect 11612 19660 11664 19712
rect 12348 19660 12400 19712
rect 14096 19660 14148 19712
rect 15752 19660 15804 19712
rect 18420 19796 18472 19848
rect 18972 19796 19024 19848
rect 19156 19796 19208 19848
rect 19248 19839 19300 19848
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 19984 19796 20036 19848
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 29276 19796 29328 19848
rect 31944 19796 31996 19848
rect 33600 19796 33652 19848
rect 34152 19839 34204 19848
rect 34152 19805 34161 19839
rect 34161 19805 34195 19839
rect 34195 19805 34204 19839
rect 34152 19796 34204 19805
rect 38108 19839 38160 19848
rect 38108 19805 38117 19839
rect 38117 19805 38151 19839
rect 38151 19805 38160 19839
rect 38108 19796 38160 19805
rect 41328 19932 41380 19984
rect 38292 19864 38344 19916
rect 38936 19796 38988 19848
rect 39120 19864 39172 19916
rect 25596 19771 25648 19780
rect 25596 19737 25605 19771
rect 25605 19737 25639 19771
rect 25639 19737 25648 19771
rect 25596 19728 25648 19737
rect 18512 19660 18564 19712
rect 20904 19660 20956 19712
rect 23756 19660 23808 19712
rect 28724 19728 28776 19780
rect 36360 19771 36412 19780
rect 36360 19737 36369 19771
rect 36369 19737 36403 19771
rect 36403 19737 36412 19771
rect 36360 19728 36412 19737
rect 37832 19728 37884 19780
rect 38292 19771 38344 19780
rect 38292 19737 38301 19771
rect 38301 19737 38335 19771
rect 38335 19737 38344 19771
rect 38292 19728 38344 19737
rect 39396 19796 39448 19848
rect 28172 19660 28224 19712
rect 30380 19660 30432 19712
rect 31668 19703 31720 19712
rect 31668 19669 31677 19703
rect 31677 19669 31711 19703
rect 31711 19669 31720 19703
rect 31668 19660 31720 19669
rect 34796 19660 34848 19712
rect 37924 19703 37976 19712
rect 37924 19669 37933 19703
rect 37933 19669 37967 19703
rect 37967 19669 37976 19703
rect 37924 19660 37976 19669
rect 38016 19660 38068 19712
rect 39396 19660 39448 19712
rect 39488 19660 39540 19712
rect 40592 19796 40644 19848
rect 41144 19839 41196 19848
rect 41144 19805 41153 19839
rect 41153 19805 41187 19839
rect 41187 19805 41196 19839
rect 41144 19796 41196 19805
rect 42156 19839 42208 19848
rect 42156 19805 42165 19839
rect 42165 19805 42199 19839
rect 42199 19805 42208 19839
rect 42156 19796 42208 19805
rect 40224 19771 40276 19780
rect 40224 19737 40233 19771
rect 40233 19737 40267 19771
rect 40267 19737 40276 19771
rect 40224 19728 40276 19737
rect 41512 19703 41564 19712
rect 41512 19669 41521 19703
rect 41521 19669 41555 19703
rect 41555 19669 41564 19703
rect 41512 19660 41564 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 5816 19499 5868 19508
rect 3792 19388 3844 19440
rect 5816 19465 5825 19499
rect 5825 19465 5859 19499
rect 5859 19465 5868 19499
rect 5816 19456 5868 19465
rect 6092 19456 6144 19508
rect 8300 19456 8352 19508
rect 12440 19456 12492 19508
rect 12900 19456 12952 19508
rect 15108 19456 15160 19508
rect 16396 19456 16448 19508
rect 16580 19456 16632 19508
rect 18420 19499 18472 19508
rect 18420 19465 18429 19499
rect 18429 19465 18463 19499
rect 18463 19465 18472 19499
rect 18420 19456 18472 19465
rect 19064 19456 19116 19508
rect 9680 19388 9732 19440
rect 10140 19431 10192 19440
rect 10140 19397 10149 19431
rect 10149 19397 10183 19431
rect 10183 19397 10192 19431
rect 10140 19388 10192 19397
rect 10784 19388 10836 19440
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 4712 19320 4764 19372
rect 6000 19320 6052 19372
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 6644 19363 6696 19372
rect 6644 19329 6678 19363
rect 6678 19329 6696 19363
rect 6644 19320 6696 19329
rect 8024 19363 8076 19372
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 3608 19252 3660 19304
rect 5080 19184 5132 19236
rect 5448 19184 5500 19236
rect 5724 19184 5776 19236
rect 10324 19320 10376 19372
rect 17684 19388 17736 19440
rect 10692 19252 10744 19304
rect 11428 19252 11480 19304
rect 12348 19252 12400 19304
rect 13820 19295 13872 19304
rect 13820 19261 13829 19295
rect 13829 19261 13863 19295
rect 13863 19261 13872 19295
rect 13820 19252 13872 19261
rect 4988 19116 5040 19168
rect 5816 19116 5868 19168
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 8668 19184 8720 19236
rect 11612 19184 11664 19236
rect 11888 19184 11940 19236
rect 12256 19184 12308 19236
rect 13912 19227 13964 19236
rect 13912 19193 13921 19227
rect 13921 19193 13955 19227
rect 13955 19193 13964 19227
rect 13912 19184 13964 19193
rect 7748 19159 7800 19168
rect 7748 19125 7757 19159
rect 7757 19125 7791 19159
rect 7791 19125 7800 19159
rect 7748 19116 7800 19125
rect 12072 19116 12124 19168
rect 13084 19116 13136 19168
rect 15200 19320 15252 19372
rect 15384 19363 15436 19372
rect 15384 19329 15418 19363
rect 15418 19329 15436 19363
rect 15384 19320 15436 19329
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 19248 19320 19300 19372
rect 21180 19388 21232 19440
rect 22376 19456 22428 19508
rect 25596 19499 25648 19508
rect 25596 19465 25605 19499
rect 25605 19465 25639 19499
rect 25639 19465 25648 19499
rect 25596 19456 25648 19465
rect 27068 19456 27120 19508
rect 28724 19456 28776 19508
rect 22100 19388 22152 19440
rect 25044 19388 25096 19440
rect 25412 19388 25464 19440
rect 28172 19388 28224 19440
rect 33048 19456 33100 19508
rect 33692 19456 33744 19508
rect 34336 19456 34388 19508
rect 38292 19456 38344 19508
rect 38936 19456 38988 19508
rect 40776 19456 40828 19508
rect 41144 19456 41196 19508
rect 27436 19363 27488 19372
rect 27436 19329 27445 19363
rect 27445 19329 27479 19363
rect 27479 19329 27488 19363
rect 27436 19320 27488 19329
rect 29920 19320 29972 19372
rect 32128 19320 32180 19372
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 20260 19252 20312 19304
rect 21364 19252 21416 19304
rect 21824 19184 21876 19236
rect 23480 19252 23532 19304
rect 26056 19295 26108 19304
rect 26056 19261 26065 19295
rect 26065 19261 26099 19295
rect 26099 19261 26108 19295
rect 26056 19252 26108 19261
rect 28172 19252 28224 19304
rect 29736 19252 29788 19304
rect 30656 19252 30708 19304
rect 15108 19116 15160 19168
rect 22284 19116 22336 19168
rect 23204 19116 23256 19168
rect 32680 19184 32732 19236
rect 32864 19363 32916 19372
rect 32864 19329 32873 19363
rect 32873 19329 32907 19363
rect 32907 19329 32916 19363
rect 32864 19320 32916 19329
rect 33416 19363 33468 19372
rect 33416 19329 33425 19363
rect 33425 19329 33459 19363
rect 33459 19329 33468 19363
rect 33416 19320 33468 19329
rect 33692 19252 33744 19304
rect 34060 19320 34112 19372
rect 34244 19363 34296 19372
rect 34244 19329 34253 19363
rect 34253 19329 34287 19363
rect 34287 19329 34296 19363
rect 34244 19320 34296 19329
rect 34336 19363 34388 19372
rect 34336 19329 34345 19363
rect 34345 19329 34379 19363
rect 34379 19329 34388 19363
rect 34336 19320 34388 19329
rect 35624 19320 35676 19372
rect 36728 19363 36780 19372
rect 36728 19329 36737 19363
rect 36737 19329 36771 19363
rect 36771 19329 36780 19363
rect 36728 19320 36780 19329
rect 38568 19388 38620 19440
rect 39488 19431 39540 19440
rect 39488 19397 39497 19431
rect 39497 19397 39531 19431
rect 39531 19397 39540 19431
rect 39488 19388 39540 19397
rect 40132 19388 40184 19440
rect 37924 19320 37976 19372
rect 41696 19320 41748 19372
rect 33508 19184 33560 19236
rect 31484 19116 31536 19168
rect 34520 19159 34572 19168
rect 34520 19125 34529 19159
rect 34529 19125 34563 19159
rect 34563 19125 34572 19159
rect 34520 19116 34572 19125
rect 37556 19252 37608 19304
rect 39212 19295 39264 19304
rect 39212 19261 39221 19295
rect 39221 19261 39255 19295
rect 39255 19261 39264 19295
rect 39212 19252 39264 19261
rect 40132 19252 40184 19304
rect 41604 19295 41656 19304
rect 41604 19261 41613 19295
rect 41613 19261 41647 19295
rect 41647 19261 41656 19295
rect 41604 19252 41656 19261
rect 41420 19184 41472 19236
rect 34888 19116 34940 19168
rect 36084 19116 36136 19168
rect 37188 19116 37240 19168
rect 37280 19116 37332 19168
rect 37924 19116 37976 19168
rect 38200 19159 38252 19168
rect 38200 19125 38209 19159
rect 38209 19125 38243 19159
rect 38243 19125 38252 19159
rect 38200 19116 38252 19125
rect 41052 19159 41104 19168
rect 41052 19125 41061 19159
rect 41061 19125 41095 19159
rect 41095 19125 41104 19159
rect 41052 19116 41104 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3608 18912 3660 18964
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2320 18776 2372 18828
rect 4620 18776 4672 18828
rect 1768 18751 1820 18760
rect 1768 18717 1777 18751
rect 1777 18717 1811 18751
rect 1811 18717 1820 18751
rect 1768 18708 1820 18717
rect 5080 18887 5132 18896
rect 5080 18853 5089 18887
rect 5089 18853 5123 18887
rect 5123 18853 5132 18887
rect 5080 18844 5132 18853
rect 5264 18844 5316 18896
rect 4988 18751 5040 18760
rect 4988 18717 4997 18751
rect 4997 18717 5031 18751
rect 5031 18717 5040 18751
rect 4988 18708 5040 18717
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 5264 18751 5316 18760
rect 5264 18717 5273 18751
rect 5273 18717 5307 18751
rect 5307 18717 5316 18751
rect 5264 18708 5316 18717
rect 6276 18912 6328 18964
rect 6644 18912 6696 18964
rect 6184 18887 6236 18896
rect 6184 18853 6193 18887
rect 6193 18853 6227 18887
rect 6227 18853 6236 18887
rect 6184 18844 6236 18853
rect 9772 18912 9824 18964
rect 10140 18912 10192 18964
rect 10324 18955 10376 18964
rect 10324 18921 10333 18955
rect 10333 18921 10367 18955
rect 10367 18921 10376 18955
rect 10324 18912 10376 18921
rect 11152 18912 11204 18964
rect 11704 18955 11756 18964
rect 11704 18921 11713 18955
rect 11713 18921 11747 18955
rect 11747 18921 11756 18955
rect 11704 18912 11756 18921
rect 11888 18955 11940 18964
rect 11888 18921 11897 18955
rect 11897 18921 11931 18955
rect 11931 18921 11940 18955
rect 11888 18912 11940 18921
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 3700 18640 3752 18692
rect 4252 18640 4304 18692
rect 5724 18708 5776 18760
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 11244 18844 11296 18896
rect 12440 18844 12492 18896
rect 8668 18776 8720 18828
rect 8300 18640 8352 18692
rect 4712 18572 4764 18624
rect 5172 18572 5224 18624
rect 5632 18572 5684 18624
rect 8024 18572 8076 18624
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 10324 18776 10376 18828
rect 9588 18708 9640 18760
rect 9680 18640 9732 18692
rect 9956 18708 10008 18760
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 10968 18776 11020 18828
rect 13820 18912 13872 18964
rect 15384 18955 15436 18964
rect 15384 18921 15393 18955
rect 15393 18921 15427 18955
rect 15427 18921 15436 18955
rect 15384 18912 15436 18921
rect 16948 18912 17000 18964
rect 20260 18955 20312 18964
rect 20260 18921 20269 18955
rect 20269 18921 20303 18955
rect 20303 18921 20312 18955
rect 20260 18912 20312 18921
rect 23112 18912 23164 18964
rect 23756 18912 23808 18964
rect 28172 18955 28224 18964
rect 28172 18921 28181 18955
rect 28181 18921 28215 18955
rect 28215 18921 28224 18955
rect 28172 18912 28224 18921
rect 35624 18912 35676 18964
rect 11244 18708 11296 18760
rect 9588 18572 9640 18624
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 10140 18615 10192 18624
rect 10140 18581 10149 18615
rect 10149 18581 10183 18615
rect 10183 18581 10192 18615
rect 10140 18572 10192 18581
rect 10968 18615 11020 18624
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 11612 18640 11664 18692
rect 12072 18640 12124 18692
rect 12532 18708 12584 18760
rect 14556 18708 14608 18760
rect 16304 18776 16356 18828
rect 16948 18776 17000 18828
rect 17500 18776 17552 18828
rect 22284 18844 22336 18896
rect 24124 18819 24176 18828
rect 24124 18785 24133 18819
rect 24133 18785 24167 18819
rect 24167 18785 24176 18819
rect 24124 18776 24176 18785
rect 25136 18776 25188 18828
rect 29276 18776 29328 18828
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 18420 18708 18472 18760
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 12256 18572 12308 18624
rect 17868 18640 17920 18692
rect 20536 18640 20588 18692
rect 22100 18683 22152 18692
rect 22100 18649 22109 18683
rect 22109 18649 22143 18683
rect 22143 18649 22152 18683
rect 28356 18751 28408 18760
rect 28356 18717 28365 18751
rect 28365 18717 28399 18751
rect 28399 18717 28408 18751
rect 28356 18708 28408 18717
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 28724 18708 28776 18760
rect 30564 18844 30616 18896
rect 30380 18776 30432 18828
rect 32772 18776 32824 18828
rect 37648 18844 37700 18896
rect 39764 18844 39816 18896
rect 34520 18776 34572 18828
rect 36176 18819 36228 18828
rect 36176 18785 36185 18819
rect 36185 18785 36219 18819
rect 36219 18785 36228 18819
rect 36176 18776 36228 18785
rect 22100 18640 22152 18649
rect 22560 18640 22612 18692
rect 23112 18640 23164 18692
rect 13176 18572 13228 18624
rect 18880 18572 18932 18624
rect 21364 18572 21416 18624
rect 23664 18572 23716 18624
rect 28448 18683 28500 18692
rect 28448 18649 28457 18683
rect 28457 18649 28491 18683
rect 28491 18649 28500 18683
rect 28448 18640 28500 18649
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 33692 18708 33744 18760
rect 37280 18776 37332 18828
rect 37556 18776 37608 18828
rect 38200 18776 38252 18828
rect 41788 18912 41840 18964
rect 42156 18955 42208 18964
rect 42156 18921 42165 18955
rect 42165 18921 42199 18955
rect 42199 18921 42208 18955
rect 42156 18912 42208 18921
rect 28632 18572 28684 18624
rect 30656 18640 30708 18692
rect 31208 18640 31260 18692
rect 37188 18751 37240 18760
rect 37188 18717 37197 18751
rect 37197 18717 37231 18751
rect 37231 18717 37240 18751
rect 37188 18708 37240 18717
rect 39212 18751 39264 18760
rect 39212 18717 39221 18751
rect 39221 18717 39255 18751
rect 39255 18717 39264 18751
rect 39212 18708 39264 18717
rect 40316 18819 40368 18828
rect 40316 18785 40325 18819
rect 40325 18785 40359 18819
rect 40359 18785 40368 18819
rect 40316 18776 40368 18785
rect 41052 18776 41104 18828
rect 29184 18615 29236 18624
rect 29184 18581 29193 18615
rect 29193 18581 29227 18615
rect 29227 18581 29236 18615
rect 29184 18572 29236 18581
rect 30104 18572 30156 18624
rect 30472 18572 30524 18624
rect 31024 18572 31076 18624
rect 37556 18640 37608 18692
rect 31668 18572 31720 18624
rect 32496 18615 32548 18624
rect 32496 18581 32505 18615
rect 32505 18581 32539 18615
rect 32539 18581 32548 18615
rect 32496 18572 32548 18581
rect 32588 18572 32640 18624
rect 34060 18572 34112 18624
rect 35532 18572 35584 18624
rect 37464 18572 37516 18624
rect 41420 18640 41472 18692
rect 40132 18572 40184 18624
rect 40316 18615 40368 18624
rect 40316 18581 40325 18615
rect 40325 18581 40359 18615
rect 40359 18581 40368 18615
rect 40316 18572 40368 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 1768 18368 1820 18420
rect 4252 18411 4304 18420
rect 4252 18377 4261 18411
rect 4261 18377 4295 18411
rect 4295 18377 4304 18411
rect 4252 18368 4304 18377
rect 3608 18300 3660 18352
rect 4620 18368 4672 18420
rect 5264 18411 5316 18420
rect 5264 18377 5273 18411
rect 5273 18377 5307 18411
rect 5307 18377 5316 18411
rect 5264 18368 5316 18377
rect 4804 18343 4856 18352
rect 4804 18309 4813 18343
rect 4813 18309 4847 18343
rect 4847 18309 4856 18343
rect 4804 18300 4856 18309
rect 5724 18300 5776 18352
rect 5908 18300 5960 18352
rect 1492 18232 1544 18284
rect 4620 18232 4672 18284
rect 2412 18164 2464 18216
rect 3792 18164 3844 18216
rect 4804 18164 4856 18216
rect 6184 18232 6236 18284
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8300 18232 8352 18284
rect 8760 18232 8812 18284
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 5264 18164 5316 18216
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 5724 18207 5776 18216
rect 5724 18173 5733 18207
rect 5733 18173 5767 18207
rect 5767 18173 5776 18207
rect 5724 18164 5776 18173
rect 9588 18232 9640 18284
rect 9864 18232 9916 18284
rect 10048 18368 10100 18420
rect 12348 18368 12400 18420
rect 14096 18368 14148 18420
rect 15108 18368 15160 18420
rect 11980 18300 12032 18352
rect 10508 18232 10560 18284
rect 12256 18232 12308 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 15200 18300 15252 18352
rect 9404 18164 9456 18216
rect 9956 18164 10008 18216
rect 11428 18164 11480 18216
rect 7656 18096 7708 18148
rect 7288 18028 7340 18080
rect 8024 18028 8076 18080
rect 10140 18096 10192 18148
rect 9128 18071 9180 18080
rect 9128 18037 9137 18071
rect 9137 18037 9171 18071
rect 9171 18037 9180 18071
rect 9128 18028 9180 18037
rect 11060 18028 11112 18080
rect 11612 18164 11664 18216
rect 11704 18164 11756 18216
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 19156 18368 19208 18420
rect 21364 18368 21416 18420
rect 21824 18411 21876 18420
rect 21824 18377 21833 18411
rect 21833 18377 21867 18411
rect 21867 18377 21876 18411
rect 21824 18368 21876 18377
rect 22100 18368 22152 18420
rect 22560 18411 22612 18420
rect 22560 18377 22569 18411
rect 22569 18377 22603 18411
rect 22603 18377 22612 18411
rect 22560 18368 22612 18377
rect 27160 18368 27212 18420
rect 28448 18411 28500 18420
rect 28448 18377 28457 18411
rect 28457 18377 28491 18411
rect 28491 18377 28500 18411
rect 28448 18368 28500 18377
rect 28632 18411 28684 18420
rect 28632 18377 28641 18411
rect 28641 18377 28675 18411
rect 28675 18377 28684 18411
rect 28632 18368 28684 18377
rect 19340 18300 19392 18352
rect 18880 18275 18932 18284
rect 18880 18241 18889 18275
rect 18889 18241 18923 18275
rect 18923 18241 18932 18275
rect 18880 18232 18932 18241
rect 18972 18275 19024 18284
rect 18972 18241 18981 18275
rect 18981 18241 19015 18275
rect 19015 18241 19024 18275
rect 18972 18232 19024 18241
rect 19432 18232 19484 18284
rect 19616 18275 19668 18284
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 19892 18275 19944 18284
rect 19892 18241 19901 18275
rect 19901 18241 19935 18275
rect 19935 18241 19944 18275
rect 19892 18232 19944 18241
rect 20720 18232 20772 18284
rect 12900 18028 12952 18080
rect 14556 18028 14608 18080
rect 16580 18164 16632 18216
rect 17960 18164 18012 18216
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 20352 18164 20404 18216
rect 20076 18096 20128 18148
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 22560 18232 22612 18284
rect 22652 18232 22704 18284
rect 23480 18275 23532 18284
rect 23480 18241 23489 18275
rect 23489 18241 23523 18275
rect 23523 18241 23532 18275
rect 23480 18232 23532 18241
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 23664 18275 23716 18284
rect 23664 18241 23673 18275
rect 23673 18241 23707 18275
rect 23707 18241 23716 18275
rect 23664 18232 23716 18241
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 22284 18164 22336 18216
rect 23388 18164 23440 18216
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24124 18232 24176 18241
rect 24860 18300 24912 18352
rect 25044 18300 25096 18352
rect 29184 18368 29236 18420
rect 31208 18411 31260 18420
rect 31208 18377 31217 18411
rect 31217 18377 31251 18411
rect 31251 18377 31260 18411
rect 31208 18368 31260 18377
rect 25320 18164 25372 18216
rect 27068 18232 27120 18284
rect 27252 18275 27304 18284
rect 27252 18241 27261 18275
rect 27261 18241 27295 18275
rect 27295 18241 27304 18275
rect 27252 18232 27304 18241
rect 29460 18300 29512 18352
rect 30104 18343 30156 18352
rect 30104 18309 30113 18343
rect 30113 18309 30147 18343
rect 30147 18309 30156 18343
rect 30104 18300 30156 18309
rect 30564 18300 30616 18352
rect 30656 18343 30708 18352
rect 30656 18309 30665 18343
rect 30665 18309 30699 18343
rect 30699 18309 30708 18343
rect 30656 18300 30708 18309
rect 31484 18343 31536 18352
rect 31484 18309 31493 18343
rect 31493 18309 31527 18343
rect 31527 18309 31536 18343
rect 31484 18300 31536 18309
rect 31668 18343 31720 18352
rect 31668 18309 31703 18343
rect 31703 18309 31720 18343
rect 31668 18300 31720 18309
rect 32588 18300 32640 18352
rect 35440 18368 35492 18420
rect 37740 18368 37792 18420
rect 38384 18368 38436 18420
rect 41604 18368 41656 18420
rect 41788 18411 41840 18420
rect 41788 18377 41797 18411
rect 41797 18377 41831 18411
rect 41831 18377 41840 18411
rect 41788 18368 41840 18377
rect 37464 18300 37516 18352
rect 40500 18300 40552 18352
rect 41328 18343 41380 18352
rect 41328 18309 41337 18343
rect 41337 18309 41371 18343
rect 41371 18309 41380 18343
rect 41328 18300 41380 18309
rect 41512 18300 41564 18352
rect 15292 18028 15344 18080
rect 16580 18028 16632 18080
rect 18788 18028 18840 18080
rect 19340 18028 19392 18080
rect 21916 18028 21968 18080
rect 23664 18096 23716 18148
rect 23848 18096 23900 18148
rect 24124 18096 24176 18148
rect 26148 18139 26200 18148
rect 26148 18105 26157 18139
rect 26157 18105 26191 18139
rect 26191 18105 26200 18139
rect 26148 18096 26200 18105
rect 25596 18028 25648 18080
rect 25688 18028 25740 18080
rect 30380 18275 30432 18284
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 29092 18164 29144 18216
rect 31484 18164 31536 18216
rect 32220 18232 32272 18284
rect 32496 18275 32548 18284
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 31944 18096 31996 18148
rect 32312 18096 32364 18148
rect 28908 18028 28960 18080
rect 30288 18028 30340 18080
rect 32772 18207 32824 18216
rect 32772 18173 32781 18207
rect 32781 18173 32815 18207
rect 32815 18173 32824 18207
rect 32772 18164 32824 18173
rect 34612 18164 34664 18216
rect 37280 18164 37332 18216
rect 38108 18232 38160 18284
rect 39028 18275 39080 18284
rect 39028 18241 39037 18275
rect 39037 18241 39071 18275
rect 39071 18241 39080 18275
rect 39028 18232 39080 18241
rect 40040 18232 40092 18284
rect 41144 18232 41196 18284
rect 39764 18207 39816 18216
rect 39764 18173 39773 18207
rect 39773 18173 39807 18207
rect 39807 18173 39816 18207
rect 39764 18164 39816 18173
rect 40224 18207 40276 18216
rect 40224 18173 40233 18207
rect 40233 18173 40267 18207
rect 40267 18173 40276 18207
rect 40224 18164 40276 18173
rect 40132 18096 40184 18148
rect 40776 18164 40828 18216
rect 42064 18232 42116 18284
rect 42156 18275 42208 18284
rect 42156 18241 42165 18275
rect 42165 18241 42199 18275
rect 42199 18241 42208 18275
rect 42156 18232 42208 18241
rect 40408 18096 40460 18148
rect 33140 18028 33192 18080
rect 33692 18028 33744 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3792 17867 3844 17876
rect 3792 17833 3801 17867
rect 3801 17833 3835 17867
rect 3835 17833 3844 17867
rect 3792 17824 3844 17833
rect 5356 17867 5408 17876
rect 5356 17833 5365 17867
rect 5365 17833 5399 17867
rect 5399 17833 5408 17867
rect 5356 17824 5408 17833
rect 5724 17824 5776 17876
rect 5448 17756 5500 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 5632 17688 5684 17740
rect 5724 17731 5776 17740
rect 5724 17697 5733 17731
rect 5733 17697 5767 17731
rect 5767 17697 5776 17731
rect 5724 17688 5776 17697
rect 7564 17824 7616 17876
rect 8024 17824 8076 17876
rect 9680 17824 9732 17876
rect 10048 17824 10100 17876
rect 10508 17824 10560 17876
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 14004 17824 14056 17876
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 18052 17824 18104 17876
rect 19248 17824 19300 17876
rect 20812 17824 20864 17876
rect 22192 17824 22244 17876
rect 24860 17867 24912 17876
rect 24860 17833 24869 17867
rect 24869 17833 24903 17867
rect 24903 17833 24912 17867
rect 24860 17824 24912 17833
rect 28356 17824 28408 17876
rect 29552 17867 29604 17876
rect 29552 17833 29561 17867
rect 29561 17833 29595 17867
rect 29595 17833 29604 17867
rect 29552 17824 29604 17833
rect 36176 17824 36228 17876
rect 37280 17867 37332 17876
rect 37280 17833 37289 17867
rect 37289 17833 37323 17867
rect 37323 17833 37332 17867
rect 37280 17824 37332 17833
rect 37556 17824 37608 17876
rect 7196 17799 7248 17808
rect 7196 17765 7205 17799
rect 7205 17765 7239 17799
rect 7239 17765 7248 17799
rect 7196 17756 7248 17765
rect 8760 17799 8812 17808
rect 8760 17765 8769 17799
rect 8769 17765 8803 17799
rect 8803 17765 8812 17799
rect 8760 17756 8812 17765
rect 9496 17756 9548 17808
rect 10232 17756 10284 17808
rect 12164 17756 12216 17808
rect 7288 17688 7340 17740
rect 1768 17663 1820 17672
rect 1768 17629 1777 17663
rect 1777 17629 1811 17663
rect 1811 17629 1820 17663
rect 1768 17620 1820 17629
rect 4620 17620 4672 17672
rect 5172 17620 5224 17672
rect 2596 17552 2648 17604
rect 5356 17552 5408 17604
rect 5632 17552 5684 17604
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 11520 17688 11572 17740
rect 21456 17756 21508 17808
rect 15108 17688 15160 17740
rect 15200 17688 15252 17740
rect 18696 17688 18748 17740
rect 18788 17731 18840 17740
rect 18788 17697 18797 17731
rect 18797 17697 18831 17731
rect 18831 17697 18840 17731
rect 18788 17688 18840 17697
rect 20720 17688 20772 17740
rect 9404 17663 9456 17672
rect 9404 17629 9413 17663
rect 9413 17629 9447 17663
rect 9447 17629 9456 17663
rect 9404 17620 9456 17629
rect 9496 17663 9548 17672
rect 9496 17629 9505 17663
rect 9505 17629 9539 17663
rect 9539 17629 9548 17663
rect 9496 17620 9548 17629
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 5724 17484 5776 17536
rect 6460 17484 6512 17536
rect 9588 17552 9640 17604
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 10232 17620 10284 17672
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 13452 17620 13504 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14556 17620 14608 17672
rect 15292 17620 15344 17672
rect 17684 17620 17736 17672
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 19892 17620 19944 17672
rect 20352 17620 20404 17672
rect 20996 17620 21048 17672
rect 21272 17620 21324 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 21732 17731 21784 17740
rect 21732 17697 21741 17731
rect 21741 17697 21775 17731
rect 21775 17697 21784 17731
rect 21732 17688 21784 17697
rect 22560 17756 22612 17808
rect 24952 17756 25004 17808
rect 25688 17756 25740 17808
rect 28540 17756 28592 17808
rect 29368 17756 29420 17808
rect 25136 17688 25188 17740
rect 7748 17484 7800 17536
rect 9404 17484 9456 17536
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 11704 17552 11756 17604
rect 23388 17663 23440 17672
rect 23388 17629 23397 17663
rect 23397 17629 23431 17663
rect 23431 17629 23440 17663
rect 23388 17620 23440 17629
rect 24032 17620 24084 17672
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 24952 17620 25004 17672
rect 26056 17688 26108 17740
rect 28356 17688 28408 17740
rect 28632 17688 28684 17740
rect 15384 17527 15436 17536
rect 15384 17493 15393 17527
rect 15393 17493 15427 17527
rect 15427 17493 15436 17527
rect 15384 17484 15436 17493
rect 17224 17527 17276 17536
rect 17224 17493 17233 17527
rect 17233 17493 17267 17527
rect 17267 17493 17276 17527
rect 17224 17484 17276 17493
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 20168 17484 20220 17536
rect 21272 17484 21324 17536
rect 21732 17484 21784 17536
rect 24124 17552 24176 17604
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 25136 17595 25188 17604
rect 25136 17561 25145 17595
rect 25145 17561 25179 17595
rect 25179 17561 25188 17595
rect 25136 17552 25188 17561
rect 26516 17552 26568 17604
rect 27068 17595 27120 17604
rect 27068 17561 27077 17595
rect 27077 17561 27111 17595
rect 27111 17561 27120 17595
rect 27068 17552 27120 17561
rect 23480 17484 23532 17536
rect 24400 17484 24452 17536
rect 25320 17484 25372 17536
rect 26424 17484 26476 17536
rect 26976 17484 27028 17536
rect 27344 17484 27396 17536
rect 27712 17620 27764 17672
rect 27896 17552 27948 17604
rect 28816 17620 28868 17672
rect 28908 17663 28960 17672
rect 28908 17629 28917 17663
rect 28917 17629 28951 17663
rect 28951 17629 28960 17663
rect 28908 17620 28960 17629
rect 29184 17663 29236 17672
rect 29184 17629 29193 17663
rect 29193 17629 29227 17663
rect 29227 17629 29236 17663
rect 29184 17620 29236 17629
rect 29736 17663 29788 17672
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 29920 17663 29972 17672
rect 29920 17629 29929 17663
rect 29929 17629 29963 17663
rect 29963 17629 29972 17663
rect 29920 17620 29972 17629
rect 30104 17663 30156 17672
rect 30104 17629 30113 17663
rect 30113 17629 30147 17663
rect 30147 17629 30156 17663
rect 30104 17620 30156 17629
rect 29828 17595 29880 17604
rect 29828 17561 29837 17595
rect 29837 17561 29871 17595
rect 29871 17561 29880 17595
rect 29828 17552 29880 17561
rect 27528 17527 27580 17536
rect 27528 17493 27537 17527
rect 27537 17493 27571 17527
rect 27571 17493 27580 17527
rect 27528 17484 27580 17493
rect 29000 17484 29052 17536
rect 29092 17527 29144 17536
rect 29092 17493 29101 17527
rect 29101 17493 29135 17527
rect 29135 17493 29144 17527
rect 30288 17620 30340 17672
rect 30840 17799 30892 17808
rect 30840 17765 30849 17799
rect 30849 17765 30883 17799
rect 30883 17765 30892 17799
rect 30840 17756 30892 17765
rect 32128 17756 32180 17808
rect 32220 17756 32272 17808
rect 32496 17756 32548 17808
rect 37188 17756 37240 17808
rect 32588 17688 32640 17740
rect 37924 17688 37976 17740
rect 31668 17663 31720 17672
rect 31668 17629 31677 17663
rect 31677 17629 31711 17663
rect 31711 17629 31720 17663
rect 31668 17620 31720 17629
rect 33416 17620 33468 17672
rect 33692 17663 33744 17672
rect 33692 17629 33701 17663
rect 33701 17629 33735 17663
rect 33735 17629 33744 17663
rect 33692 17620 33744 17629
rect 32220 17552 32272 17604
rect 32772 17595 32824 17604
rect 32772 17561 32781 17595
rect 32781 17561 32815 17595
rect 32815 17561 32824 17595
rect 32772 17552 32824 17561
rect 34612 17552 34664 17604
rect 34980 17595 35032 17604
rect 34980 17561 34989 17595
rect 34989 17561 35023 17595
rect 35023 17561 35032 17595
rect 34980 17552 35032 17561
rect 35440 17552 35492 17604
rect 37648 17663 37700 17672
rect 37648 17629 37657 17663
rect 37657 17629 37691 17663
rect 37691 17629 37700 17663
rect 37648 17620 37700 17629
rect 38108 17620 38160 17672
rect 40592 17620 40644 17672
rect 41788 17620 41840 17672
rect 37740 17552 37792 17604
rect 41880 17552 41932 17604
rect 29092 17484 29144 17493
rect 33048 17484 33100 17536
rect 36452 17527 36504 17536
rect 36452 17493 36461 17527
rect 36461 17493 36495 17527
rect 36495 17493 36504 17527
rect 36452 17484 36504 17493
rect 36544 17527 36596 17536
rect 36544 17493 36553 17527
rect 36553 17493 36587 17527
rect 36587 17493 36596 17527
rect 36544 17484 36596 17493
rect 37464 17484 37516 17536
rect 38016 17484 38068 17536
rect 40776 17484 40828 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 1768 17280 1820 17332
rect 2596 17280 2648 17332
rect 5264 17280 5316 17332
rect 5540 17280 5592 17332
rect 6552 17280 6604 17332
rect 7196 17280 7248 17332
rect 10692 17280 10744 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 4712 17212 4764 17264
rect 6184 17255 6236 17264
rect 6184 17221 6193 17255
rect 6193 17221 6227 17255
rect 6227 17221 6236 17255
rect 6184 17212 6236 17221
rect 848 17144 900 17196
rect 2412 17144 2464 17196
rect 2964 17119 3016 17128
rect 2964 17085 2973 17119
rect 2973 17085 3007 17119
rect 3007 17085 3016 17119
rect 2964 17076 3016 17085
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 5264 17144 5316 17196
rect 5448 17076 5500 17128
rect 5908 17144 5960 17196
rect 6460 17144 6512 17196
rect 7656 17144 7708 17196
rect 6368 17119 6420 17128
rect 6368 17085 6377 17119
rect 6377 17085 6411 17119
rect 6411 17085 6420 17119
rect 6368 17076 6420 17085
rect 7840 17144 7892 17196
rect 9128 17212 9180 17264
rect 9864 17212 9916 17264
rect 14096 17212 14148 17264
rect 4712 16940 4764 16992
rect 5632 16940 5684 16992
rect 6184 16940 6236 16992
rect 7656 17008 7708 17060
rect 8300 17119 8352 17128
rect 8300 17085 8309 17119
rect 8309 17085 8343 17119
rect 8343 17085 8352 17119
rect 8300 17076 8352 17085
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 9496 17187 9548 17196
rect 8668 17144 8720 17153
rect 9496 17153 9505 17187
rect 9505 17153 9539 17187
rect 9539 17153 9548 17187
rect 9496 17144 9548 17153
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 8760 17076 8812 17128
rect 9680 17076 9732 17128
rect 10600 17076 10652 17128
rect 14004 17144 14056 17196
rect 17132 17323 17184 17332
rect 17132 17289 17141 17323
rect 17141 17289 17175 17323
rect 17175 17289 17184 17323
rect 17132 17280 17184 17289
rect 18696 17323 18748 17332
rect 18696 17289 18705 17323
rect 18705 17289 18739 17323
rect 18739 17289 18748 17323
rect 18696 17280 18748 17289
rect 15016 17212 15068 17264
rect 17224 17212 17276 17264
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 15200 17076 15252 17128
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 18880 17280 18932 17332
rect 19156 17280 19208 17332
rect 19248 17280 19300 17332
rect 19340 17212 19392 17264
rect 20812 17323 20864 17332
rect 20812 17289 20821 17323
rect 20821 17289 20855 17323
rect 20855 17289 20864 17323
rect 20812 17280 20864 17289
rect 19892 17255 19944 17264
rect 19892 17221 19901 17255
rect 19901 17221 19935 17255
rect 19935 17221 19944 17255
rect 19892 17212 19944 17221
rect 21456 17280 21508 17332
rect 24492 17280 24544 17332
rect 24584 17280 24636 17332
rect 8668 17008 8720 17060
rect 7564 16940 7616 16992
rect 9404 16983 9456 16992
rect 9404 16949 9413 16983
rect 9413 16949 9447 16983
rect 9447 16949 9456 16983
rect 9404 16940 9456 16949
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 13820 17008 13872 17060
rect 17776 17076 17828 17128
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 19156 17187 19208 17196
rect 19156 17153 19191 17187
rect 19191 17153 19208 17187
rect 19156 17144 19208 17153
rect 19432 17144 19484 17196
rect 19616 17187 19668 17196
rect 19616 17153 19625 17187
rect 19625 17153 19659 17187
rect 19659 17153 19668 17187
rect 19616 17144 19668 17153
rect 20076 17144 20128 17196
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 13912 16940 13964 16992
rect 14188 16940 14240 16992
rect 14556 16940 14608 16992
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 15568 16940 15620 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20352 17008 20404 17060
rect 20628 17008 20680 17060
rect 20996 17144 21048 17196
rect 21548 17144 21600 17196
rect 23480 17255 23532 17264
rect 23480 17221 23489 17255
rect 23489 17221 23523 17255
rect 23523 17221 23532 17255
rect 23480 17212 23532 17221
rect 25136 17280 25188 17332
rect 27344 17323 27396 17332
rect 27344 17289 27353 17323
rect 27353 17289 27387 17323
rect 27387 17289 27396 17323
rect 27344 17280 27396 17289
rect 22008 17187 22060 17196
rect 22008 17153 22017 17187
rect 22017 17153 22051 17187
rect 22051 17153 22060 17187
rect 22008 17144 22060 17153
rect 24124 17187 24176 17196
rect 24124 17153 24133 17187
rect 24133 17153 24167 17187
rect 24167 17153 24176 17187
rect 24124 17144 24176 17153
rect 24400 17187 24452 17196
rect 24400 17153 24409 17187
rect 24409 17153 24443 17187
rect 24443 17153 24452 17187
rect 24400 17144 24452 17153
rect 21272 17008 21324 17060
rect 24032 17008 24084 17060
rect 24768 17187 24820 17196
rect 24768 17153 24777 17187
rect 24777 17153 24811 17187
rect 24811 17153 24820 17187
rect 24768 17144 24820 17153
rect 24952 17187 25004 17196
rect 24952 17153 24961 17187
rect 24961 17153 24995 17187
rect 24995 17153 25004 17187
rect 24952 17144 25004 17153
rect 25688 17212 25740 17264
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 27252 17212 27304 17264
rect 26424 17144 26476 17153
rect 24676 17119 24728 17128
rect 24676 17085 24685 17119
rect 24685 17085 24719 17119
rect 24719 17085 24728 17119
rect 24676 17076 24728 17085
rect 24860 17076 24912 17128
rect 27712 17187 27764 17196
rect 27712 17153 27721 17187
rect 27721 17153 27755 17187
rect 27755 17153 27764 17187
rect 27712 17144 27764 17153
rect 27896 17187 27948 17196
rect 27896 17153 27905 17187
rect 27905 17153 27939 17187
rect 27939 17153 27948 17187
rect 27896 17144 27948 17153
rect 29184 17280 29236 17332
rect 31944 17280 31996 17332
rect 32680 17280 32732 17332
rect 34980 17280 35032 17332
rect 36544 17280 36596 17332
rect 36636 17280 36688 17332
rect 33692 17212 33744 17264
rect 34796 17212 34848 17264
rect 38108 17212 38160 17264
rect 39856 17212 39908 17264
rect 40316 17255 40368 17264
rect 40316 17221 40325 17255
rect 40325 17221 40359 17255
rect 40359 17221 40368 17255
rect 40316 17212 40368 17221
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 24952 17008 25004 17060
rect 27160 17076 27212 17128
rect 28448 17187 28500 17196
rect 28448 17153 28457 17187
rect 28457 17153 28491 17187
rect 28491 17153 28500 17187
rect 28448 17144 28500 17153
rect 28540 17144 28592 17196
rect 29000 17144 29052 17196
rect 29460 17187 29512 17196
rect 29460 17153 29469 17187
rect 29469 17153 29503 17187
rect 29503 17153 29512 17187
rect 29460 17144 29512 17153
rect 29184 17119 29236 17128
rect 29184 17085 29193 17119
rect 29193 17085 29227 17119
rect 29227 17085 29236 17119
rect 29184 17076 29236 17085
rect 30840 17119 30892 17128
rect 30840 17085 30849 17119
rect 30849 17085 30883 17119
rect 30883 17085 30892 17119
rect 30840 17076 30892 17085
rect 32128 17144 32180 17196
rect 33048 17144 33100 17196
rect 33416 17144 33468 17196
rect 31668 17076 31720 17128
rect 33232 17076 33284 17128
rect 37096 17076 37148 17128
rect 38476 17144 38528 17196
rect 38752 17076 38804 17128
rect 40224 17144 40276 17196
rect 40776 17255 40828 17264
rect 40776 17221 40785 17255
rect 40785 17221 40819 17255
rect 40819 17221 40828 17255
rect 40776 17212 40828 17221
rect 41788 17187 41840 17196
rect 41788 17153 41797 17187
rect 41797 17153 41831 17187
rect 41831 17153 41840 17187
rect 41788 17144 41840 17153
rect 41880 17144 41932 17196
rect 42156 17187 42208 17196
rect 42156 17153 42165 17187
rect 42165 17153 42199 17187
rect 42199 17153 42208 17187
rect 42156 17144 42208 17153
rect 24676 16940 24728 16992
rect 25964 16940 26016 16992
rect 29000 17008 29052 17060
rect 29092 17051 29144 17060
rect 29092 17017 29101 17051
rect 29101 17017 29135 17051
rect 29135 17017 29144 17051
rect 29092 17008 29144 17017
rect 31484 17008 31536 17060
rect 31760 17008 31812 17060
rect 32312 17008 32364 17060
rect 38844 17008 38896 17060
rect 28540 16940 28592 16992
rect 28632 16983 28684 16992
rect 28632 16949 28641 16983
rect 28641 16949 28675 16983
rect 28675 16949 28684 16983
rect 28632 16940 28684 16949
rect 28908 16940 28960 16992
rect 32588 16940 32640 16992
rect 38384 16940 38436 16992
rect 38660 16940 38712 16992
rect 41236 16983 41288 16992
rect 41236 16949 41245 16983
rect 41245 16949 41279 16983
rect 41279 16949 41288 16983
rect 41236 16940 41288 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2964 16736 3016 16788
rect 5356 16779 5408 16788
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 7564 16736 7616 16788
rect 8760 16779 8812 16788
rect 8760 16745 8769 16779
rect 8769 16745 8803 16779
rect 8803 16745 8812 16779
rect 8760 16736 8812 16745
rect 9404 16736 9456 16788
rect 12716 16736 12768 16788
rect 13820 16736 13872 16788
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 17040 16736 17092 16788
rect 19340 16736 19392 16788
rect 20168 16736 20220 16788
rect 3240 16600 3292 16652
rect 12808 16600 12860 16652
rect 17960 16668 18012 16720
rect 24952 16736 25004 16788
rect 27068 16736 27120 16788
rect 28908 16736 28960 16788
rect 29092 16736 29144 16788
rect 31760 16736 31812 16788
rect 32128 16736 32180 16788
rect 32312 16736 32364 16788
rect 33232 16779 33284 16788
rect 33232 16745 33241 16779
rect 33241 16745 33275 16779
rect 33275 16745 33284 16779
rect 33232 16736 33284 16745
rect 36636 16736 36688 16788
rect 38752 16779 38804 16788
rect 38752 16745 38761 16779
rect 38761 16745 38795 16779
rect 38795 16745 38804 16779
rect 38752 16736 38804 16745
rect 42156 16779 42208 16788
rect 42156 16745 42165 16779
rect 42165 16745 42199 16779
rect 42199 16745 42208 16779
rect 42156 16736 42208 16745
rect 4804 16532 4856 16584
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 7380 16575 7432 16584
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 9496 16575 9548 16584
rect 9496 16541 9505 16575
rect 9505 16541 9539 16575
rect 9539 16541 9548 16575
rect 9496 16532 9548 16541
rect 11336 16532 11388 16584
rect 4620 16464 4672 16516
rect 5356 16507 5408 16516
rect 5356 16473 5365 16507
rect 5365 16473 5399 16507
rect 5399 16473 5408 16507
rect 5356 16464 5408 16473
rect 5724 16464 5776 16516
rect 11980 16464 12032 16516
rect 13820 16532 13872 16584
rect 14096 16532 14148 16584
rect 15200 16600 15252 16652
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 9864 16396 9916 16448
rect 13912 16464 13964 16516
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 13820 16396 13872 16448
rect 14740 16464 14792 16516
rect 16304 16464 16356 16516
rect 17868 16575 17920 16584
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 17868 16532 17920 16541
rect 19432 16600 19484 16652
rect 19616 16600 19668 16652
rect 20812 16643 20864 16652
rect 20812 16609 20821 16643
rect 20821 16609 20855 16643
rect 20855 16609 20864 16643
rect 20812 16600 20864 16609
rect 19156 16532 19208 16584
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 28632 16711 28684 16720
rect 28632 16677 28641 16711
rect 28641 16677 28675 16711
rect 28675 16677 28684 16711
rect 28632 16668 28684 16677
rect 28724 16711 28776 16720
rect 28724 16677 28733 16711
rect 28733 16677 28767 16711
rect 28767 16677 28776 16711
rect 28724 16668 28776 16677
rect 28816 16668 28868 16720
rect 24768 16600 24820 16652
rect 24860 16600 24912 16652
rect 26332 16600 26384 16652
rect 28448 16600 28500 16652
rect 29184 16668 29236 16720
rect 24032 16464 24084 16516
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 20076 16396 20128 16448
rect 20444 16396 20496 16448
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 25596 16532 25648 16584
rect 25964 16575 26016 16584
rect 25964 16541 25973 16575
rect 25973 16541 26007 16575
rect 26007 16541 26016 16575
rect 25964 16532 26016 16541
rect 26148 16575 26200 16584
rect 26148 16541 26157 16575
rect 26157 16541 26191 16575
rect 26191 16541 26200 16575
rect 26148 16532 26200 16541
rect 28908 16575 28960 16586
rect 24860 16396 24912 16448
rect 25964 16396 26016 16448
rect 28908 16541 28927 16575
rect 28927 16541 28960 16575
rect 28908 16534 28960 16541
rect 29460 16600 29512 16652
rect 31852 16600 31904 16652
rect 32312 16600 32364 16652
rect 33140 16643 33192 16652
rect 33140 16609 33149 16643
rect 33149 16609 33183 16643
rect 33183 16609 33192 16643
rect 33140 16600 33192 16609
rect 29368 16532 29420 16584
rect 29736 16532 29788 16584
rect 30932 16532 30984 16584
rect 29184 16464 29236 16516
rect 29460 16464 29512 16516
rect 29828 16464 29880 16516
rect 31484 16507 31536 16516
rect 31484 16473 31493 16507
rect 31493 16473 31527 16507
rect 31527 16473 31536 16507
rect 31484 16464 31536 16473
rect 31668 16575 31720 16584
rect 31668 16541 31677 16575
rect 31677 16541 31711 16575
rect 31711 16541 31720 16575
rect 31668 16532 31720 16541
rect 34336 16668 34388 16720
rect 35348 16668 35400 16720
rect 36452 16668 36504 16720
rect 36084 16600 36136 16652
rect 38384 16643 38436 16652
rect 38384 16609 38393 16643
rect 38393 16609 38427 16643
rect 38427 16609 38436 16643
rect 38384 16600 38436 16609
rect 39212 16600 39264 16652
rect 40040 16668 40092 16720
rect 31116 16439 31168 16448
rect 31116 16405 31125 16439
rect 31125 16405 31159 16439
rect 31159 16405 31168 16439
rect 31116 16396 31168 16405
rect 32680 16464 32732 16516
rect 32956 16507 33008 16516
rect 32956 16473 32965 16507
rect 32965 16473 32999 16507
rect 32999 16473 33008 16507
rect 32956 16464 33008 16473
rect 36360 16532 36412 16584
rect 37832 16464 37884 16516
rect 38292 16464 38344 16516
rect 39856 16575 39908 16584
rect 39856 16541 39865 16575
rect 39865 16541 39899 16575
rect 39899 16541 39908 16575
rect 39856 16532 39908 16541
rect 40224 16575 40276 16584
rect 40224 16541 40233 16575
rect 40233 16541 40267 16575
rect 40267 16541 40276 16575
rect 40224 16532 40276 16541
rect 40316 16575 40368 16584
rect 40316 16541 40325 16575
rect 40325 16541 40359 16575
rect 40359 16541 40368 16575
rect 40316 16532 40368 16541
rect 40684 16507 40736 16516
rect 40684 16473 40693 16507
rect 40693 16473 40727 16507
rect 40727 16473 40736 16507
rect 40684 16464 40736 16473
rect 42064 16464 42116 16516
rect 33232 16396 33284 16448
rect 33324 16396 33376 16448
rect 37740 16396 37792 16448
rect 38108 16396 38160 16448
rect 40592 16396 40644 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 2596 16192 2648 16244
rect 4804 16192 4856 16244
rect 6920 16192 6972 16244
rect 10876 16124 10928 16176
rect 17316 16192 17368 16244
rect 19524 16192 19576 16244
rect 24032 16192 24084 16244
rect 848 16056 900 16108
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2412 16056 2464 16108
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 8760 16056 8812 16108
rect 12164 16124 12216 16176
rect 12900 16056 12952 16108
rect 3792 15988 3844 16040
rect 3884 15988 3936 16040
rect 5356 15988 5408 16040
rect 11520 16031 11572 16040
rect 11520 15997 11529 16031
rect 11529 15997 11563 16031
rect 11563 15997 11572 16031
rect 11520 15988 11572 15997
rect 13176 16099 13228 16108
rect 13176 16065 13185 16099
rect 13185 16065 13219 16099
rect 13219 16065 13228 16099
rect 13176 16056 13228 16065
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 11336 15920 11388 15972
rect 1768 15852 1820 15904
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 1860 15852 1912 15861
rect 5264 15852 5316 15904
rect 11428 15852 11480 15904
rect 12716 15920 12768 15972
rect 13268 15963 13320 15972
rect 13268 15929 13277 15963
rect 13277 15929 13311 15963
rect 13311 15929 13320 15963
rect 13268 15920 13320 15929
rect 12256 15852 12308 15904
rect 15200 15988 15252 16040
rect 17040 15988 17092 16040
rect 17316 15988 17368 16040
rect 19064 16056 19116 16108
rect 18788 15988 18840 16040
rect 19524 16099 19576 16108
rect 19524 16065 19533 16099
rect 19533 16065 19567 16099
rect 19567 16065 19576 16099
rect 19524 16056 19576 16065
rect 19616 16099 19668 16108
rect 19616 16065 19625 16099
rect 19625 16065 19659 16099
rect 19659 16065 19668 16099
rect 19616 16056 19668 16065
rect 19984 16124 20036 16176
rect 20168 16124 20220 16176
rect 19892 16099 19944 16108
rect 19892 16065 19901 16099
rect 19901 16065 19935 16099
rect 19935 16065 19944 16099
rect 19892 16056 19944 16065
rect 20444 16167 20496 16176
rect 20444 16133 20453 16167
rect 20453 16133 20487 16167
rect 20487 16133 20496 16167
rect 20444 16124 20496 16133
rect 20536 16167 20588 16176
rect 20536 16133 20545 16167
rect 20545 16133 20579 16167
rect 20579 16133 20588 16167
rect 20536 16124 20588 16133
rect 23940 16124 23992 16176
rect 25228 16192 25280 16244
rect 26240 16192 26292 16244
rect 27344 16235 27396 16244
rect 27344 16201 27353 16235
rect 27353 16201 27387 16235
rect 27387 16201 27396 16235
rect 27344 16192 27396 16201
rect 28908 16192 28960 16244
rect 21916 16056 21968 16108
rect 24676 16167 24728 16176
rect 24676 16133 24685 16167
rect 24685 16133 24719 16167
rect 24719 16133 24728 16167
rect 24676 16124 24728 16133
rect 24860 16124 24912 16176
rect 29920 16192 29972 16244
rect 31392 16192 31444 16244
rect 31668 16192 31720 16244
rect 33968 16192 34020 16244
rect 36360 16235 36412 16244
rect 36360 16201 36369 16235
rect 36369 16201 36403 16235
rect 36403 16201 36412 16235
rect 36360 16192 36412 16201
rect 37832 16192 37884 16244
rect 29644 16124 29696 16176
rect 32588 16124 32640 16176
rect 33324 16124 33376 16176
rect 20444 15988 20496 16040
rect 21456 16031 21508 16040
rect 21456 15997 21465 16031
rect 21465 15997 21499 16031
rect 21499 15997 21508 16031
rect 21456 15988 21508 15997
rect 24768 15988 24820 16040
rect 25504 16056 25556 16108
rect 25688 15988 25740 16040
rect 28080 16056 28132 16108
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 30288 16099 30340 16108
rect 29092 15988 29144 16040
rect 29368 15988 29420 16040
rect 19340 15920 19392 15972
rect 19984 15920 20036 15972
rect 23664 15920 23716 15972
rect 26424 15920 26476 15972
rect 15200 15852 15252 15904
rect 15752 15852 15804 15904
rect 18788 15852 18840 15904
rect 19524 15852 19576 15904
rect 20812 15895 20864 15904
rect 20812 15861 20821 15895
rect 20821 15861 20855 15895
rect 20855 15861 20864 15895
rect 20812 15852 20864 15861
rect 26056 15852 26108 15904
rect 28724 15852 28776 15904
rect 29184 15852 29236 15904
rect 30288 16065 30297 16099
rect 30297 16065 30331 16099
rect 30331 16065 30340 16099
rect 30288 16056 30340 16065
rect 30564 16099 30616 16108
rect 30564 16065 30573 16099
rect 30573 16065 30607 16099
rect 30607 16065 30616 16099
rect 30564 16056 30616 16065
rect 30472 15852 30524 15904
rect 32220 16099 32272 16108
rect 32220 16065 32229 16099
rect 32229 16065 32263 16099
rect 32263 16065 32272 16099
rect 32220 16056 32272 16065
rect 31208 15988 31260 16040
rect 32772 16031 32824 16040
rect 32772 15997 32781 16031
rect 32781 15997 32815 16031
rect 32815 15997 32824 16031
rect 32772 15988 32824 15997
rect 33600 15988 33652 16040
rect 32312 15920 32364 15972
rect 31484 15852 31536 15904
rect 33416 15852 33468 15904
rect 35348 16124 35400 16176
rect 34612 16099 34664 16108
rect 34612 16065 34621 16099
rect 34621 16065 34655 16099
rect 34655 16065 34664 16099
rect 34612 16056 34664 16065
rect 35440 15988 35492 16040
rect 35532 15988 35584 16040
rect 38660 16124 38712 16176
rect 40040 16235 40092 16244
rect 40040 16201 40049 16235
rect 40049 16201 40083 16235
rect 40083 16201 40092 16235
rect 40040 16192 40092 16201
rect 40684 16192 40736 16244
rect 41236 16124 41288 16176
rect 37464 16099 37516 16108
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 37740 16056 37792 16108
rect 40132 16099 40184 16108
rect 40132 16065 40141 16099
rect 40141 16065 40175 16099
rect 40175 16065 40184 16099
rect 40132 16056 40184 16065
rect 40408 16099 40460 16108
rect 40408 16065 40417 16099
rect 40417 16065 40451 16099
rect 40451 16065 40460 16099
rect 40408 16056 40460 16065
rect 38292 16031 38344 16040
rect 38292 15997 38301 16031
rect 38301 15997 38335 16031
rect 38335 15997 38344 16031
rect 38292 15988 38344 15997
rect 40040 15988 40092 16040
rect 40592 16056 40644 16108
rect 37464 15920 37516 15972
rect 41604 16031 41656 16040
rect 41604 15997 41613 16031
rect 41613 15997 41647 16031
rect 41647 15997 41656 16031
rect 41604 15988 41656 15997
rect 35348 15852 35400 15904
rect 37188 15852 37240 15904
rect 38108 15852 38160 15904
rect 39764 15852 39816 15904
rect 40224 15852 40276 15904
rect 41696 15852 41748 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3792 15691 3844 15700
rect 3792 15657 3801 15691
rect 3801 15657 3835 15691
rect 3835 15657 3844 15691
rect 3792 15648 3844 15657
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 11428 15648 11480 15700
rect 11704 15648 11756 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 2320 15512 2372 15564
rect 5724 15555 5776 15564
rect 5724 15521 5733 15555
rect 5733 15521 5767 15555
rect 5767 15521 5776 15555
rect 5724 15512 5776 15521
rect 6460 15512 6512 15564
rect 10876 15512 10928 15564
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 5816 15487 5868 15496
rect 5816 15453 5825 15487
rect 5825 15453 5859 15487
rect 5859 15453 5868 15487
rect 5816 15444 5868 15453
rect 6736 15444 6788 15496
rect 8484 15444 8536 15496
rect 9220 15444 9272 15496
rect 2596 15376 2648 15428
rect 6644 15308 6696 15360
rect 10048 15444 10100 15496
rect 12164 15512 12216 15564
rect 12900 15648 12952 15700
rect 17224 15691 17276 15700
rect 17224 15657 17233 15691
rect 17233 15657 17267 15691
rect 17267 15657 17276 15691
rect 17224 15648 17276 15657
rect 17316 15691 17368 15700
rect 17316 15657 17325 15691
rect 17325 15657 17359 15691
rect 17359 15657 17368 15691
rect 17316 15648 17368 15657
rect 18420 15648 18472 15700
rect 19616 15648 19668 15700
rect 23664 15648 23716 15700
rect 25596 15648 25648 15700
rect 14924 15580 14976 15632
rect 13912 15512 13964 15564
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 21456 15512 21508 15564
rect 23204 15512 23256 15564
rect 25688 15580 25740 15632
rect 24860 15512 24912 15564
rect 26148 15512 26200 15564
rect 11704 15444 11756 15496
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12256 15444 12308 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 9864 15308 9916 15360
rect 11060 15308 11112 15360
rect 11152 15351 11204 15360
rect 11152 15317 11161 15351
rect 11161 15317 11195 15351
rect 11195 15317 11204 15351
rect 11152 15308 11204 15317
rect 12716 15376 12768 15428
rect 11980 15308 12032 15360
rect 12072 15308 12124 15360
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 13268 15376 13320 15428
rect 15200 15444 15252 15496
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 17684 15444 17736 15496
rect 19156 15444 19208 15496
rect 15752 15419 15804 15428
rect 15752 15385 15761 15419
rect 15761 15385 15795 15419
rect 15795 15385 15804 15419
rect 15752 15376 15804 15385
rect 16304 15376 16356 15428
rect 18788 15419 18840 15428
rect 18788 15385 18797 15419
rect 18797 15385 18831 15419
rect 18831 15385 18840 15419
rect 18788 15376 18840 15385
rect 19432 15419 19484 15428
rect 19432 15385 19441 15419
rect 19441 15385 19475 15419
rect 19475 15385 19484 15419
rect 24308 15444 24360 15496
rect 24952 15444 25004 15496
rect 27344 15648 27396 15700
rect 29000 15648 29052 15700
rect 29092 15648 29144 15700
rect 30196 15648 30248 15700
rect 30656 15580 30708 15632
rect 27712 15555 27764 15564
rect 27712 15521 27721 15555
rect 27721 15521 27755 15555
rect 27755 15521 27764 15555
rect 27712 15512 27764 15521
rect 28356 15512 28408 15564
rect 29092 15444 29144 15496
rect 29920 15444 29972 15496
rect 19432 15376 19484 15385
rect 20812 15376 20864 15428
rect 20996 15376 21048 15428
rect 19892 15308 19944 15360
rect 22652 15308 22704 15360
rect 24676 15376 24728 15428
rect 26056 15419 26108 15428
rect 26056 15385 26065 15419
rect 26065 15385 26099 15419
rect 26099 15385 26108 15419
rect 26056 15376 26108 15385
rect 27528 15376 27580 15428
rect 29460 15376 29512 15428
rect 30472 15487 30524 15496
rect 30472 15453 30481 15487
rect 30481 15453 30515 15487
rect 30515 15453 30524 15487
rect 30472 15444 30524 15453
rect 30656 15487 30708 15496
rect 30656 15453 30665 15487
rect 30665 15453 30699 15487
rect 30699 15453 30708 15487
rect 30656 15444 30708 15453
rect 28448 15308 28500 15360
rect 29184 15308 29236 15360
rect 29552 15351 29604 15360
rect 29552 15317 29561 15351
rect 29561 15317 29595 15351
rect 29595 15317 29604 15351
rect 29552 15308 29604 15317
rect 30196 15308 30248 15360
rect 32588 15648 32640 15700
rect 33600 15691 33652 15700
rect 33600 15657 33609 15691
rect 33609 15657 33643 15691
rect 33643 15657 33652 15691
rect 33600 15648 33652 15657
rect 35440 15691 35492 15700
rect 35440 15657 35449 15691
rect 35449 15657 35483 15691
rect 35483 15657 35492 15691
rect 35440 15648 35492 15657
rect 32680 15623 32732 15632
rect 32680 15589 32689 15623
rect 32689 15589 32723 15623
rect 32723 15589 32732 15623
rect 32680 15580 32732 15589
rect 31208 15512 31260 15564
rect 34244 15580 34296 15632
rect 33416 15512 33468 15564
rect 33968 15487 34020 15496
rect 33968 15453 33977 15487
rect 33977 15453 34011 15487
rect 34011 15453 34020 15487
rect 33968 15444 34020 15453
rect 34704 15444 34756 15496
rect 34888 15444 34940 15496
rect 35532 15444 35584 15496
rect 30380 15308 30432 15360
rect 31484 15376 31536 15428
rect 32496 15376 32548 15428
rect 33324 15376 33376 15428
rect 31852 15308 31904 15360
rect 32956 15308 33008 15360
rect 35440 15308 35492 15360
rect 37188 15555 37240 15564
rect 37188 15521 37197 15555
rect 37197 15521 37231 15555
rect 37231 15521 37240 15555
rect 37188 15512 37240 15521
rect 40224 15691 40276 15700
rect 40224 15657 40233 15691
rect 40233 15657 40267 15691
rect 40267 15657 40276 15691
rect 40224 15648 40276 15657
rect 41972 15580 42024 15632
rect 37464 15487 37516 15496
rect 37464 15453 37473 15487
rect 37473 15453 37507 15487
rect 37507 15453 37516 15487
rect 37464 15444 37516 15453
rect 38568 15444 38620 15496
rect 40408 15487 40460 15496
rect 40408 15453 40417 15487
rect 40417 15453 40451 15487
rect 40451 15453 40460 15487
rect 40408 15444 40460 15453
rect 37832 15376 37884 15428
rect 38292 15419 38344 15428
rect 38292 15385 38301 15419
rect 38301 15385 38335 15419
rect 38335 15385 38344 15419
rect 38292 15376 38344 15385
rect 40500 15376 40552 15428
rect 40868 15376 40920 15428
rect 41512 15376 41564 15428
rect 38476 15308 38528 15360
rect 41420 15308 41472 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 3240 15104 3292 15156
rect 5816 15104 5868 15156
rect 6184 15104 6236 15156
rect 6828 15104 6880 15156
rect 2596 15036 2648 15088
rect 10232 15104 10284 15156
rect 11152 15104 11204 15156
rect 12072 15104 12124 15156
rect 14740 15104 14792 15156
rect 19432 15104 19484 15156
rect 20720 15104 20772 15156
rect 20812 15104 20864 15156
rect 21364 15104 21416 15156
rect 23296 15104 23348 15156
rect 17684 15036 17736 15088
rect 19524 15079 19576 15088
rect 19524 15045 19533 15079
rect 19533 15045 19567 15079
rect 19567 15045 19576 15079
rect 19524 15036 19576 15045
rect 23112 15036 23164 15088
rect 1400 15011 1452 15020
rect 1400 14977 1409 15011
rect 1409 14977 1443 15011
rect 1443 14977 1452 15011
rect 1400 14968 1452 14977
rect 1860 14968 1912 15020
rect 11060 14968 11112 15020
rect 11336 15011 11388 15020
rect 11336 14977 11345 15011
rect 11345 14977 11379 15011
rect 11379 14977 11388 15011
rect 11336 14968 11388 14977
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 13912 15011 13964 15020
rect 13912 14977 13946 15011
rect 13946 14977 13964 15011
rect 13912 14968 13964 14977
rect 19984 14968 20036 15020
rect 20168 14968 20220 15020
rect 5816 14900 5868 14952
rect 6368 14943 6420 14952
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 10324 14832 10376 14884
rect 8116 14807 8168 14816
rect 8116 14773 8125 14807
rect 8125 14773 8159 14807
rect 8159 14773 8168 14807
rect 8116 14764 8168 14773
rect 9680 14764 9732 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13912 14764 13964 14816
rect 15476 14832 15528 14884
rect 19432 14764 19484 14816
rect 21456 14968 21508 15020
rect 22008 14968 22060 15020
rect 20720 14900 20772 14952
rect 24492 15036 24544 15088
rect 26148 15036 26200 15088
rect 29552 15036 29604 15088
rect 29644 15036 29696 15088
rect 31208 15036 31260 15088
rect 32220 15104 32272 15156
rect 36544 15104 36596 15156
rect 38292 15104 38344 15156
rect 38568 15104 38620 15156
rect 27528 14968 27580 15020
rect 24492 14900 24544 14952
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24860 14943 24912 14952
rect 24860 14909 24869 14943
rect 24869 14909 24903 14943
rect 24903 14909 24912 14943
rect 24860 14900 24912 14909
rect 24952 14943 25004 14952
rect 24952 14909 24961 14943
rect 24961 14909 24995 14943
rect 24995 14909 25004 14943
rect 24952 14900 25004 14909
rect 26424 14943 26476 14952
rect 26424 14909 26433 14943
rect 26433 14909 26467 14943
rect 26467 14909 26476 14943
rect 26424 14900 26476 14909
rect 27620 14900 27672 14952
rect 29184 15011 29236 15020
rect 29184 14977 29193 15011
rect 29193 14977 29227 15011
rect 29227 14977 29236 15011
rect 29184 14968 29236 14977
rect 23572 14832 23624 14884
rect 29092 14943 29144 14952
rect 29092 14909 29101 14943
rect 29101 14909 29135 14943
rect 29135 14909 29144 14943
rect 29092 14900 29144 14909
rect 29552 14900 29604 14952
rect 35348 15036 35400 15088
rect 37832 15036 37884 15088
rect 31576 15011 31628 15020
rect 31576 14977 31585 15011
rect 31585 14977 31619 15011
rect 31619 14977 31628 15011
rect 31576 14968 31628 14977
rect 34244 15011 34296 15020
rect 34244 14977 34253 15011
rect 34253 14977 34287 15011
rect 34287 14977 34296 15011
rect 34244 14968 34296 14977
rect 35440 15011 35492 15020
rect 32772 14900 32824 14952
rect 33140 14900 33192 14952
rect 35440 14977 35449 15011
rect 35449 14977 35483 15011
rect 35483 14977 35492 15011
rect 35440 14968 35492 14977
rect 36084 14968 36136 15020
rect 40040 15104 40092 15156
rect 40408 15104 40460 15156
rect 40224 14968 40276 15020
rect 40592 14968 40644 15020
rect 34888 14943 34940 14952
rect 34888 14909 34897 14943
rect 34897 14909 34931 14943
rect 34931 14909 34940 14943
rect 34888 14900 34940 14909
rect 20720 14807 20772 14816
rect 20720 14773 20729 14807
rect 20729 14773 20763 14807
rect 20763 14773 20772 14807
rect 20720 14764 20772 14773
rect 24768 14764 24820 14816
rect 28080 14764 28132 14816
rect 29460 14764 29512 14816
rect 29920 14832 29972 14884
rect 33416 14832 33468 14884
rect 34704 14832 34756 14884
rect 36452 14943 36504 14952
rect 36452 14909 36461 14943
rect 36461 14909 36495 14943
rect 36495 14909 36504 14943
rect 36452 14900 36504 14909
rect 37280 14900 37332 14952
rect 37832 14900 37884 14952
rect 40132 14943 40184 14952
rect 40132 14909 40141 14943
rect 40141 14909 40175 14943
rect 40175 14909 40184 14943
rect 40132 14900 40184 14909
rect 37648 14764 37700 14816
rect 39856 14832 39908 14884
rect 41420 14968 41472 15020
rect 41972 15011 42024 15020
rect 41972 14977 41981 15011
rect 41981 14977 42015 15011
rect 42015 14977 42024 15011
rect 41972 14968 42024 14977
rect 41604 14832 41656 14884
rect 40684 14764 40736 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 5816 14560 5868 14612
rect 6644 14560 6696 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 10324 14603 10376 14612
rect 10324 14569 10333 14603
rect 10333 14569 10367 14603
rect 10367 14569 10376 14603
rect 10324 14560 10376 14569
rect 11336 14560 11388 14612
rect 11980 14560 12032 14612
rect 14648 14560 14700 14612
rect 10416 14492 10468 14544
rect 8116 14424 8168 14476
rect 2504 14356 2556 14408
rect 3976 14356 4028 14408
rect 4620 14288 4672 14340
rect 6460 14331 6512 14340
rect 6460 14297 6469 14331
rect 6469 14297 6503 14331
rect 6503 14297 6512 14331
rect 6460 14288 6512 14297
rect 6552 14288 6604 14340
rect 7380 14356 7432 14408
rect 8484 14356 8536 14408
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 2688 14220 2740 14272
rect 5448 14220 5500 14272
rect 9705 14331 9757 14340
rect 9705 14297 9715 14331
rect 9715 14297 9749 14331
rect 9749 14297 9757 14331
rect 9956 14356 10008 14408
rect 12900 14424 12952 14476
rect 22008 14560 22060 14612
rect 24308 14560 24360 14612
rect 24584 14560 24636 14612
rect 25688 14560 25740 14612
rect 26884 14560 26936 14612
rect 27712 14560 27764 14612
rect 28264 14560 28316 14612
rect 32220 14560 32272 14612
rect 32312 14560 32364 14612
rect 32772 14603 32824 14612
rect 32772 14569 32781 14603
rect 32781 14569 32815 14603
rect 32815 14569 32824 14603
rect 32772 14560 32824 14569
rect 24492 14492 24544 14544
rect 26516 14492 26568 14544
rect 27252 14492 27304 14544
rect 29368 14492 29420 14544
rect 17408 14467 17460 14476
rect 17408 14433 17417 14467
rect 17417 14433 17451 14467
rect 17451 14433 17460 14467
rect 17408 14424 17460 14433
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 24860 14424 24912 14476
rect 25136 14424 25188 14476
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 12072 14356 12124 14408
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 18604 14356 18656 14408
rect 19892 14356 19944 14408
rect 9705 14288 9757 14297
rect 11428 14288 11480 14340
rect 7748 14220 7800 14272
rect 9220 14220 9272 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 10324 14220 10376 14272
rect 13728 14220 13780 14272
rect 16304 14220 16356 14272
rect 17960 14288 18012 14340
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 24768 14356 24820 14408
rect 26148 14424 26200 14476
rect 26332 14356 26384 14408
rect 27068 14356 27120 14408
rect 31208 14424 31260 14476
rect 33232 14467 33284 14476
rect 33232 14433 33241 14467
rect 33241 14433 33275 14467
rect 33275 14433 33284 14467
rect 33232 14424 33284 14433
rect 33416 14467 33468 14476
rect 33416 14433 33425 14467
rect 33425 14433 33459 14467
rect 33459 14433 33468 14467
rect 33416 14424 33468 14433
rect 34704 14424 34756 14476
rect 36268 14560 36320 14612
rect 40132 14560 40184 14612
rect 40500 14560 40552 14612
rect 41972 14560 42024 14612
rect 40224 14492 40276 14544
rect 36360 14467 36412 14476
rect 36360 14433 36369 14467
rect 36369 14433 36403 14467
rect 36403 14433 36412 14467
rect 36360 14424 36412 14433
rect 37188 14424 37240 14476
rect 38200 14424 38252 14476
rect 40684 14467 40736 14476
rect 40684 14433 40693 14467
rect 40693 14433 40727 14467
rect 40727 14433 40736 14467
rect 40684 14424 40736 14433
rect 28264 14399 28316 14408
rect 28264 14365 28273 14399
rect 28273 14365 28307 14399
rect 28307 14365 28316 14399
rect 28264 14356 28316 14365
rect 28356 14356 28408 14408
rect 29460 14356 29512 14408
rect 32496 14356 32548 14408
rect 33968 14356 34020 14408
rect 34336 14356 34388 14408
rect 36452 14356 36504 14408
rect 36728 14356 36780 14408
rect 37464 14356 37516 14408
rect 38384 14399 38436 14408
rect 38384 14365 38393 14399
rect 38393 14365 38427 14399
rect 38427 14365 38436 14399
rect 38384 14356 38436 14365
rect 39856 14399 39908 14408
rect 39856 14365 39865 14399
rect 39865 14365 39899 14399
rect 39899 14365 39908 14399
rect 39856 14356 39908 14365
rect 17040 14220 17092 14272
rect 18788 14263 18840 14272
rect 18788 14229 18797 14263
rect 18797 14229 18831 14263
rect 18831 14229 18840 14263
rect 18788 14220 18840 14229
rect 20628 14288 20680 14340
rect 20996 14288 21048 14340
rect 21180 14288 21232 14340
rect 22652 14331 22704 14340
rect 22652 14297 22661 14331
rect 22661 14297 22695 14331
rect 22695 14297 22704 14331
rect 22652 14288 22704 14297
rect 23112 14288 23164 14340
rect 29000 14331 29052 14340
rect 29000 14297 29009 14331
rect 29009 14297 29043 14331
rect 29043 14297 29052 14331
rect 29000 14288 29052 14297
rect 29736 14331 29788 14340
rect 29736 14297 29745 14331
rect 29745 14297 29779 14331
rect 29779 14297 29788 14331
rect 29736 14288 29788 14297
rect 30932 14288 30984 14340
rect 31116 14288 31168 14340
rect 20536 14220 20588 14272
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 26516 14263 26568 14272
rect 26516 14229 26525 14263
rect 26525 14229 26559 14263
rect 26559 14229 26568 14263
rect 26516 14220 26568 14229
rect 29920 14220 29972 14272
rect 33416 14288 33468 14340
rect 41972 14288 42024 14340
rect 34244 14220 34296 14272
rect 35440 14220 35492 14272
rect 36268 14220 36320 14272
rect 36912 14263 36964 14272
rect 36912 14229 36921 14263
rect 36921 14229 36955 14263
rect 36955 14229 36964 14263
rect 36912 14220 36964 14229
rect 37832 14263 37884 14272
rect 37832 14229 37841 14263
rect 37841 14229 37875 14263
rect 37875 14229 37884 14263
rect 37832 14220 37884 14229
rect 39948 14220 40000 14272
rect 40040 14220 40092 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 2688 13991 2740 14000
rect 2688 13957 2697 13991
rect 2697 13957 2731 13991
rect 2731 13957 2740 13991
rect 2688 13948 2740 13957
rect 3976 13948 4028 14000
rect 5724 14016 5776 14068
rect 6736 14059 6788 14068
rect 6736 14025 6738 14059
rect 6738 14025 6772 14059
rect 6772 14025 6788 14059
rect 6736 14016 6788 14025
rect 7104 14016 7156 14068
rect 12992 14016 13044 14068
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 2412 13812 2464 13821
rect 2688 13812 2740 13864
rect 6184 13880 6236 13932
rect 6368 13812 6420 13864
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 7748 13948 7800 14000
rect 10232 13948 10284 14000
rect 4620 13744 4672 13796
rect 7380 13744 7432 13796
rect 4712 13676 4764 13728
rect 6920 13676 6972 13728
rect 11888 13880 11940 13932
rect 11980 13880 12032 13932
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 12992 13880 13044 13932
rect 13728 13923 13780 13932
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 16580 14016 16632 14068
rect 18604 14059 18656 14068
rect 18604 14025 18613 14059
rect 18613 14025 18647 14059
rect 18647 14025 18656 14059
rect 18604 14016 18656 14025
rect 19800 14016 19852 14068
rect 17040 13948 17092 14000
rect 17684 13948 17736 14000
rect 19892 13948 19944 14000
rect 20352 13948 20404 14000
rect 21272 13991 21324 14000
rect 21272 13957 21281 13991
rect 21281 13957 21315 13991
rect 21315 13957 21324 13991
rect 21272 13948 21324 13957
rect 22468 14016 22520 14068
rect 24400 14059 24452 14068
rect 24400 14025 24409 14059
rect 24409 14025 24443 14059
rect 24443 14025 24452 14059
rect 24400 14016 24452 14025
rect 10692 13812 10744 13864
rect 12716 13744 12768 13796
rect 15384 13812 15436 13864
rect 20812 13923 20864 13932
rect 20812 13889 20821 13923
rect 20821 13889 20855 13923
rect 20855 13889 20864 13923
rect 20812 13880 20864 13889
rect 20996 13880 21048 13932
rect 21640 13923 21692 13932
rect 21640 13889 21649 13923
rect 21649 13889 21683 13923
rect 21683 13889 21692 13923
rect 21640 13880 21692 13889
rect 16580 13812 16632 13864
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 16948 13855 17000 13864
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17684 13812 17736 13864
rect 18972 13812 19024 13864
rect 19524 13812 19576 13864
rect 20168 13812 20220 13864
rect 20260 13812 20312 13864
rect 20904 13812 20956 13864
rect 19708 13744 19760 13796
rect 8392 13676 8444 13728
rect 13636 13676 13688 13728
rect 16764 13676 16816 13728
rect 18052 13676 18104 13728
rect 21272 13744 21324 13796
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 24952 14016 25004 14068
rect 25872 14016 25924 14068
rect 26148 14016 26200 14068
rect 25136 13948 25188 14000
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 25504 13880 25556 13932
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 25872 13923 25924 13932
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 26332 13923 26384 13932
rect 26332 13889 26341 13923
rect 26341 13889 26375 13923
rect 26375 13889 26384 13923
rect 26332 13880 26384 13889
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 27252 13991 27304 14000
rect 27252 13957 27261 13991
rect 27261 13957 27295 13991
rect 27295 13957 27304 13991
rect 27252 13948 27304 13957
rect 25872 13744 25924 13796
rect 21548 13676 21600 13728
rect 25688 13719 25740 13728
rect 25688 13685 25697 13719
rect 25697 13685 25731 13719
rect 25731 13685 25740 13719
rect 25688 13676 25740 13685
rect 26056 13719 26108 13728
rect 26056 13685 26065 13719
rect 26065 13685 26099 13719
rect 26099 13685 26108 13719
rect 26056 13676 26108 13685
rect 26792 13812 26844 13864
rect 29460 14016 29512 14068
rect 31576 14016 31628 14068
rect 33416 14059 33468 14068
rect 33416 14025 33425 14059
rect 33425 14025 33459 14059
rect 33459 14025 33468 14059
rect 33416 14016 33468 14025
rect 33508 14059 33560 14068
rect 33508 14025 33517 14059
rect 33517 14025 33551 14059
rect 33551 14025 33560 14059
rect 33508 14016 33560 14025
rect 34244 14059 34296 14068
rect 34244 14025 34253 14059
rect 34253 14025 34287 14059
rect 34287 14025 34296 14059
rect 34244 14016 34296 14025
rect 34428 14016 34480 14068
rect 35440 14016 35492 14068
rect 37280 14016 37332 14068
rect 37556 14016 37608 14068
rect 29000 13948 29052 14000
rect 29552 13948 29604 14000
rect 31024 13948 31076 14000
rect 31484 13991 31536 14000
rect 31484 13957 31493 13991
rect 31493 13957 31527 13991
rect 31527 13957 31536 13991
rect 31484 13948 31536 13957
rect 34520 13948 34572 14000
rect 27988 13812 28040 13864
rect 29552 13812 29604 13864
rect 31944 13880 31996 13932
rect 34060 13880 34112 13932
rect 37924 13948 37976 14000
rect 39304 14059 39356 14068
rect 39304 14025 39313 14059
rect 39313 14025 39347 14059
rect 39347 14025 39356 14059
rect 39304 14016 39356 14025
rect 41512 14016 41564 14068
rect 41972 13948 42024 14000
rect 36636 13880 36688 13932
rect 32312 13812 32364 13864
rect 32404 13855 32456 13864
rect 32404 13821 32413 13855
rect 32413 13821 32447 13855
rect 32447 13821 32456 13855
rect 32404 13812 32456 13821
rect 32864 13744 32916 13796
rect 33140 13744 33192 13796
rect 34428 13744 34480 13796
rect 34612 13812 34664 13864
rect 35256 13855 35308 13864
rect 35256 13821 35265 13855
rect 35265 13821 35299 13855
rect 35299 13821 35308 13855
rect 35256 13812 35308 13821
rect 37464 13812 37516 13864
rect 37832 13855 37884 13864
rect 37832 13821 37841 13855
rect 37841 13821 37875 13855
rect 37875 13821 37884 13855
rect 37832 13812 37884 13821
rect 38384 13812 38436 13864
rect 39948 13855 40000 13864
rect 39948 13821 39957 13855
rect 39957 13821 39991 13855
rect 39991 13821 40000 13855
rect 39948 13812 40000 13821
rect 40408 13812 40460 13864
rect 26240 13676 26292 13728
rect 28816 13676 28868 13728
rect 28908 13676 28960 13728
rect 32956 13719 33008 13728
rect 32956 13685 32965 13719
rect 32965 13685 32999 13719
rect 32999 13685 33008 13719
rect 32956 13676 33008 13685
rect 33416 13676 33468 13728
rect 34888 13719 34940 13728
rect 34888 13685 34897 13719
rect 34897 13685 34931 13719
rect 34931 13685 34940 13719
rect 34888 13676 34940 13685
rect 35532 13676 35584 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4068 13472 4120 13524
rect 5632 13472 5684 13524
rect 6000 13472 6052 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 2412 13336 2464 13388
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 2688 13200 2740 13252
rect 2964 13243 3016 13252
rect 2964 13209 2973 13243
rect 2973 13209 3007 13243
rect 3007 13209 3016 13243
rect 2964 13200 3016 13209
rect 2228 13132 2280 13184
rect 6552 13404 6604 13456
rect 6736 13336 6788 13388
rect 8116 13472 8168 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 16580 13472 16632 13524
rect 17684 13404 17736 13456
rect 19524 13472 19576 13524
rect 19708 13472 19760 13524
rect 21640 13472 21692 13524
rect 23204 13472 23256 13524
rect 26332 13515 26384 13524
rect 26332 13481 26341 13515
rect 26341 13481 26375 13515
rect 26375 13481 26384 13515
rect 26332 13472 26384 13481
rect 26516 13515 26568 13524
rect 26516 13481 26525 13515
rect 26525 13481 26559 13515
rect 26559 13481 26568 13515
rect 26516 13472 26568 13481
rect 28908 13472 28960 13524
rect 6828 13268 6880 13320
rect 7288 13268 7340 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 4620 13200 4672 13252
rect 6644 13200 6696 13252
rect 8392 13311 8444 13320
rect 8392 13277 8401 13311
rect 8401 13277 8435 13311
rect 8435 13277 8444 13311
rect 8392 13268 8444 13277
rect 4344 13132 4396 13184
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 7656 13175 7708 13184
rect 7656 13141 7665 13175
rect 7665 13141 7699 13175
rect 7699 13141 7708 13175
rect 7656 13132 7708 13141
rect 8668 13268 8720 13320
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 16672 13336 16724 13388
rect 17868 13336 17920 13388
rect 13636 13311 13688 13320
rect 13636 13277 13654 13311
rect 13654 13277 13688 13311
rect 13636 13268 13688 13277
rect 10232 13200 10284 13252
rect 11520 13200 11572 13252
rect 13176 13200 13228 13252
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15384 13268 15436 13320
rect 16488 13268 16540 13320
rect 18512 13336 18564 13388
rect 26240 13447 26292 13456
rect 26240 13413 26249 13447
rect 26249 13413 26283 13447
rect 26283 13413 26292 13447
rect 26240 13404 26292 13413
rect 34980 13515 35032 13524
rect 34980 13481 34989 13515
rect 34989 13481 35023 13515
rect 35023 13481 35032 13515
rect 34980 13472 35032 13481
rect 20720 13336 20772 13388
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 26056 13379 26108 13388
rect 26056 13345 26065 13379
rect 26065 13345 26099 13379
rect 26099 13345 26108 13379
rect 26056 13336 26108 13345
rect 19432 13311 19484 13320
rect 17224 13243 17276 13252
rect 17224 13209 17233 13243
rect 17233 13209 17267 13243
rect 17267 13209 17276 13243
rect 17224 13200 17276 13209
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 21180 13268 21232 13320
rect 24768 13268 24820 13320
rect 29552 13404 29604 13456
rect 34336 13447 34388 13456
rect 34336 13413 34345 13447
rect 34345 13413 34379 13447
rect 34379 13413 34388 13447
rect 34336 13404 34388 13413
rect 28356 13336 28408 13388
rect 29000 13336 29052 13388
rect 32404 13336 32456 13388
rect 32864 13379 32916 13388
rect 32864 13345 32873 13379
rect 32873 13345 32907 13379
rect 32907 13345 32916 13379
rect 32864 13336 32916 13345
rect 36176 13472 36228 13524
rect 36912 13472 36964 13524
rect 37832 13472 37884 13524
rect 39948 13472 40000 13524
rect 38660 13404 38712 13456
rect 35348 13379 35400 13388
rect 35348 13345 35357 13379
rect 35357 13345 35391 13379
rect 35391 13345 35400 13379
rect 35348 13336 35400 13345
rect 36268 13336 36320 13388
rect 36636 13336 36688 13388
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 28172 13311 28224 13320
rect 28172 13277 28181 13311
rect 28181 13277 28215 13311
rect 28215 13277 28224 13311
rect 28172 13268 28224 13277
rect 28816 13311 28868 13320
rect 28816 13277 28825 13311
rect 28825 13277 28859 13311
rect 28859 13277 28868 13311
rect 28816 13268 28868 13277
rect 19616 13200 19668 13252
rect 19984 13200 20036 13252
rect 10048 13132 10100 13184
rect 11152 13132 11204 13184
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 12716 13132 12768 13184
rect 14372 13132 14424 13184
rect 18236 13175 18288 13184
rect 18236 13141 18245 13175
rect 18245 13141 18279 13175
rect 18279 13141 18288 13175
rect 18236 13132 18288 13141
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 18972 13132 19024 13184
rect 23112 13200 23164 13252
rect 29460 13268 29512 13320
rect 29828 13268 29880 13320
rect 32128 13268 32180 13320
rect 22468 13132 22520 13184
rect 24032 13132 24084 13184
rect 24676 13132 24728 13184
rect 25964 13132 26016 13184
rect 26424 13132 26476 13184
rect 27436 13132 27488 13184
rect 29644 13132 29696 13184
rect 30932 13200 30984 13252
rect 31024 13243 31076 13252
rect 31024 13209 31033 13243
rect 31033 13209 31067 13243
rect 31067 13209 31076 13243
rect 31024 13200 31076 13209
rect 34152 13268 34204 13320
rect 37924 13336 37976 13388
rect 32864 13200 32916 13252
rect 34428 13200 34480 13252
rect 35532 13200 35584 13252
rect 30564 13132 30616 13184
rect 36268 13132 36320 13184
rect 37004 13132 37056 13184
rect 39304 13268 39356 13320
rect 39488 13336 39540 13388
rect 39764 13336 39816 13388
rect 40040 13311 40092 13320
rect 40040 13277 40049 13311
rect 40049 13277 40083 13311
rect 40083 13277 40092 13311
rect 40040 13268 40092 13277
rect 40408 13404 40460 13456
rect 41972 13447 42024 13456
rect 41972 13413 41981 13447
rect 41981 13413 42015 13447
rect 42015 13413 42024 13447
rect 41972 13404 42024 13413
rect 40500 13311 40552 13320
rect 40500 13277 40509 13311
rect 40509 13277 40543 13311
rect 40543 13277 40552 13311
rect 40500 13268 40552 13277
rect 41788 13311 41840 13320
rect 41788 13277 41797 13311
rect 41797 13277 41831 13311
rect 41831 13277 41840 13311
rect 41788 13268 41840 13277
rect 41696 13132 41748 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 2504 12971 2556 12980
rect 2504 12937 2513 12971
rect 2513 12937 2547 12971
rect 2547 12937 2556 12971
rect 2504 12928 2556 12937
rect 2964 12928 3016 12980
rect 3424 12928 3476 12980
rect 4620 12928 4672 12980
rect 2228 12860 2280 12912
rect 4068 12860 4120 12912
rect 4712 12903 4764 12912
rect 4712 12869 4721 12903
rect 4721 12869 4755 12903
rect 4755 12869 4764 12903
rect 4712 12860 4764 12869
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 11152 12971 11204 12980
rect 11152 12937 11179 12971
rect 11179 12937 11204 12971
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 2596 12835 2648 12844
rect 2596 12801 2605 12835
rect 2605 12801 2639 12835
rect 2639 12801 2648 12835
rect 2596 12792 2648 12801
rect 3516 12792 3568 12844
rect 3976 12792 4028 12844
rect 7380 12860 7432 12912
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 4712 12724 4764 12776
rect 6920 12792 6972 12844
rect 7288 12792 7340 12844
rect 8668 12860 8720 12912
rect 9864 12860 9916 12912
rect 9772 12792 9824 12844
rect 10600 12860 10652 12912
rect 11152 12928 11204 12937
rect 13176 12971 13228 12980
rect 13176 12937 13185 12971
rect 13185 12937 13219 12971
rect 13219 12937 13228 12971
rect 13176 12928 13228 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 16948 12928 17000 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 17684 12928 17736 12980
rect 17960 12928 18012 12980
rect 19248 12928 19300 12980
rect 19984 12928 20036 12980
rect 21088 12971 21140 12980
rect 21088 12937 21097 12971
rect 21097 12937 21131 12971
rect 21131 12937 21140 12971
rect 21088 12928 21140 12937
rect 21180 12928 21232 12980
rect 24032 12971 24084 12980
rect 24032 12937 24041 12971
rect 24041 12937 24075 12971
rect 24075 12937 24084 12971
rect 24032 12928 24084 12937
rect 24124 12971 24176 12980
rect 24124 12937 24133 12971
rect 24133 12937 24167 12971
rect 24167 12937 24176 12971
rect 24124 12928 24176 12937
rect 25044 12971 25096 12980
rect 25044 12937 25053 12971
rect 25053 12937 25087 12971
rect 25087 12937 25096 12971
rect 25044 12928 25096 12937
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 10140 12792 10192 12801
rect 10692 12792 10744 12844
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13912 12860 13964 12912
rect 7104 12724 7156 12776
rect 6368 12699 6420 12708
rect 6368 12665 6377 12699
rect 6377 12665 6411 12699
rect 6411 12665 6420 12699
rect 6368 12656 6420 12665
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12440 12724 12492 12776
rect 4712 12588 4764 12640
rect 7104 12588 7156 12640
rect 9680 12588 9732 12640
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 10232 12588 10284 12597
rect 12716 12656 12768 12708
rect 16764 12792 16816 12844
rect 18144 12860 18196 12912
rect 18788 12860 18840 12912
rect 18972 12860 19024 12912
rect 17960 12792 18012 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 20168 12860 20220 12912
rect 21272 12860 21324 12912
rect 21640 12860 21692 12912
rect 14096 12724 14148 12776
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 17776 12724 17828 12776
rect 17868 12724 17920 12776
rect 19248 12724 19300 12776
rect 20168 12724 20220 12776
rect 23572 12835 23624 12844
rect 23572 12801 23581 12835
rect 23581 12801 23615 12835
rect 23615 12801 23624 12835
rect 23572 12792 23624 12801
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 22468 12724 22520 12733
rect 22744 12724 22796 12776
rect 26424 12860 26476 12912
rect 26792 12860 26844 12912
rect 27436 12903 27488 12912
rect 27436 12869 27445 12903
rect 27445 12869 27479 12903
rect 27479 12869 27488 12903
rect 27436 12860 27488 12869
rect 28908 12860 28960 12912
rect 31024 12928 31076 12980
rect 32956 12928 33008 12980
rect 31944 12860 31996 12912
rect 33416 12860 33468 12912
rect 25780 12792 25832 12844
rect 29828 12792 29880 12844
rect 30564 12835 30616 12844
rect 30564 12801 30579 12835
rect 30579 12801 30613 12835
rect 30613 12801 30616 12835
rect 30564 12792 30616 12801
rect 26240 12767 26292 12776
rect 26240 12733 26249 12767
rect 26249 12733 26283 12767
rect 26283 12733 26292 12767
rect 26240 12724 26292 12733
rect 31024 12792 31076 12844
rect 32496 12792 32548 12844
rect 30840 12767 30892 12776
rect 30840 12733 30849 12767
rect 30849 12733 30883 12767
rect 30883 12733 30892 12767
rect 30840 12724 30892 12733
rect 31484 12724 31536 12776
rect 32956 12792 33008 12844
rect 34428 12792 34480 12844
rect 35164 12971 35216 12980
rect 35164 12937 35173 12971
rect 35173 12937 35207 12971
rect 35207 12937 35216 12971
rect 35164 12928 35216 12937
rect 37188 12928 37240 12980
rect 36084 12860 36136 12912
rect 36544 12860 36596 12912
rect 37004 12860 37056 12912
rect 35532 12835 35584 12844
rect 35532 12801 35541 12835
rect 35541 12801 35575 12835
rect 35575 12801 35584 12835
rect 35532 12792 35584 12801
rect 35900 12792 35952 12844
rect 32864 12724 32916 12776
rect 33968 12724 34020 12776
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 18052 12588 18104 12640
rect 19708 12588 19760 12640
rect 19892 12588 19944 12640
rect 20260 12588 20312 12640
rect 20536 12588 20588 12640
rect 34704 12656 34756 12708
rect 36544 12767 36596 12776
rect 36544 12733 36553 12767
rect 36553 12733 36587 12767
rect 36587 12733 36596 12767
rect 36544 12724 36596 12733
rect 37372 12724 37424 12776
rect 37556 12835 37608 12844
rect 37556 12801 37565 12835
rect 37565 12801 37599 12835
rect 37599 12801 37608 12835
rect 37556 12792 37608 12801
rect 37924 12903 37976 12912
rect 37924 12869 37933 12903
rect 37933 12869 37967 12903
rect 37967 12869 37976 12903
rect 37924 12860 37976 12869
rect 38660 12860 38712 12912
rect 41788 12860 41840 12912
rect 38844 12792 38896 12844
rect 37648 12724 37700 12776
rect 36636 12656 36688 12708
rect 37924 12656 37976 12708
rect 40500 12656 40552 12708
rect 23572 12588 23624 12640
rect 24676 12588 24728 12640
rect 28816 12588 28868 12640
rect 29184 12588 29236 12640
rect 29644 12588 29696 12640
rect 30564 12631 30616 12640
rect 30564 12597 30573 12631
rect 30573 12597 30607 12631
rect 30607 12597 30616 12631
rect 30564 12588 30616 12597
rect 31760 12588 31812 12640
rect 37372 12588 37424 12640
rect 37832 12588 37884 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1676 12384 1728 12436
rect 1952 12427 2004 12436
rect 1952 12393 1961 12427
rect 1961 12393 1995 12427
rect 1995 12393 2004 12427
rect 1952 12384 2004 12393
rect 4620 12384 4672 12436
rect 2780 12316 2832 12368
rect 7104 12384 7156 12436
rect 10140 12384 10192 12436
rect 11520 12384 11572 12436
rect 17224 12384 17276 12436
rect 20720 12384 20772 12436
rect 24676 12427 24728 12436
rect 14096 12359 14148 12368
rect 2228 12248 2280 12300
rect 3792 12248 3844 12300
rect 4344 12248 4396 12300
rect 4620 12248 4672 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 2044 12180 2096 12232
rect 5540 12180 5592 12232
rect 9772 12180 9824 12232
rect 10048 12248 10100 12300
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 11888 12248 11940 12300
rect 14096 12325 14105 12359
rect 14105 12325 14139 12359
rect 14139 12325 14148 12359
rect 14096 12316 14148 12325
rect 24676 12393 24706 12427
rect 24706 12393 24728 12427
rect 24676 12384 24728 12393
rect 26240 12384 26292 12436
rect 28172 12384 28224 12436
rect 31852 12384 31904 12436
rect 35440 12384 35492 12436
rect 35900 12384 35952 12436
rect 23296 12316 23348 12368
rect 26424 12316 26476 12368
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 20536 12291 20588 12300
rect 20536 12257 20545 12291
rect 20545 12257 20579 12291
rect 20579 12257 20588 12291
rect 20536 12248 20588 12257
rect 16856 12180 16908 12232
rect 20444 12180 20496 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 22744 12248 22796 12300
rect 24768 12248 24820 12300
rect 25872 12248 25924 12300
rect 26700 12291 26752 12300
rect 26700 12257 26709 12291
rect 26709 12257 26743 12291
rect 26743 12257 26752 12291
rect 26700 12248 26752 12257
rect 26884 12316 26936 12368
rect 29184 12316 29236 12368
rect 38844 12316 38896 12368
rect 2504 12112 2556 12164
rect 4804 12112 4856 12164
rect 5264 12112 5316 12164
rect 7288 12112 7340 12164
rect 4160 12044 4212 12096
rect 5356 12044 5408 12096
rect 5724 12044 5776 12096
rect 9220 12044 9272 12096
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 9588 12087 9640 12096
rect 9588 12053 9597 12087
rect 9597 12053 9631 12087
rect 9631 12053 9640 12087
rect 9588 12044 9640 12053
rect 9680 12087 9732 12096
rect 9680 12053 9689 12087
rect 9689 12053 9723 12087
rect 9723 12053 9732 12087
rect 9680 12044 9732 12053
rect 15200 12155 15252 12164
rect 15200 12121 15218 12155
rect 15218 12121 15252 12155
rect 15200 12112 15252 12121
rect 9956 12044 10008 12096
rect 10692 12044 10744 12096
rect 13544 12044 13596 12096
rect 17960 12112 18012 12164
rect 18236 12044 18288 12096
rect 19524 12044 19576 12096
rect 20536 12112 20588 12164
rect 21272 12155 21324 12164
rect 21272 12121 21281 12155
rect 21281 12121 21315 12155
rect 21315 12121 21324 12155
rect 21272 12112 21324 12121
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 22100 12180 22152 12189
rect 22284 12180 22336 12232
rect 22468 12180 22520 12232
rect 23020 12112 23072 12164
rect 20076 12044 20128 12096
rect 21640 12087 21692 12096
rect 21640 12053 21649 12087
rect 21649 12053 21683 12087
rect 21683 12053 21692 12087
rect 21640 12044 21692 12053
rect 21824 12044 21876 12096
rect 23480 12223 23532 12232
rect 23480 12189 23489 12223
rect 23489 12189 23523 12223
rect 23523 12189 23532 12223
rect 23480 12180 23532 12189
rect 29000 12248 29052 12300
rect 30564 12248 30616 12300
rect 31484 12248 31536 12300
rect 37096 12248 37148 12300
rect 23388 12112 23440 12164
rect 23664 12044 23716 12096
rect 24308 12044 24360 12096
rect 27712 12180 27764 12232
rect 28816 12180 28868 12232
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 32036 12180 32088 12232
rect 34704 12180 34756 12232
rect 24584 12112 24636 12164
rect 29920 12112 29972 12164
rect 34520 12112 34572 12164
rect 35348 12112 35400 12164
rect 36544 12180 36596 12232
rect 37280 12223 37332 12232
rect 37280 12189 37289 12223
rect 37289 12189 37323 12223
rect 37323 12189 37332 12223
rect 37280 12180 37332 12189
rect 39488 12223 39540 12232
rect 39488 12189 39497 12223
rect 39497 12189 39531 12223
rect 39531 12189 39540 12223
rect 39488 12180 39540 12189
rect 37556 12155 37608 12164
rect 37556 12121 37565 12155
rect 37565 12121 37599 12155
rect 37599 12121 37608 12155
rect 37556 12112 37608 12121
rect 38844 12112 38896 12164
rect 24860 12044 24912 12096
rect 26240 12087 26292 12096
rect 26240 12053 26249 12087
rect 26249 12053 26283 12087
rect 26283 12053 26292 12087
rect 26240 12044 26292 12053
rect 27160 12044 27212 12096
rect 31392 12087 31444 12096
rect 31392 12053 31401 12087
rect 31401 12053 31435 12087
rect 31435 12053 31444 12087
rect 31392 12044 31444 12053
rect 34796 12044 34848 12096
rect 35532 12044 35584 12096
rect 36176 12044 36228 12096
rect 39488 12044 39540 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 3516 11883 3568 11892
rect 3516 11849 3525 11883
rect 3525 11849 3559 11883
rect 3559 11849 3568 11883
rect 3516 11840 3568 11849
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2228 11704 2280 11756
rect 2504 11704 2556 11756
rect 2780 11704 2832 11756
rect 4160 11840 4212 11892
rect 2136 11568 2188 11620
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 4160 11704 4212 11756
rect 10508 11883 10560 11892
rect 10508 11849 10517 11883
rect 10517 11849 10551 11883
rect 10551 11849 10560 11883
rect 10508 11840 10560 11849
rect 11980 11840 12032 11892
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 13912 11840 13964 11892
rect 18604 11840 18656 11892
rect 22284 11840 22336 11892
rect 22468 11883 22520 11892
rect 22468 11849 22477 11883
rect 22477 11849 22511 11883
rect 22511 11849 22520 11883
rect 22468 11840 22520 11849
rect 7012 11772 7064 11824
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 3424 11636 3476 11688
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 9772 11772 9824 11824
rect 11520 11815 11572 11824
rect 11520 11781 11529 11815
rect 11529 11781 11563 11815
rect 11563 11781 11572 11815
rect 11520 11772 11572 11781
rect 12716 11815 12768 11824
rect 12716 11781 12725 11815
rect 12725 11781 12759 11815
rect 12759 11781 12768 11815
rect 12716 11772 12768 11781
rect 14372 11815 14424 11824
rect 14372 11781 14390 11815
rect 14390 11781 14424 11815
rect 14372 11772 14424 11781
rect 18512 11772 18564 11824
rect 20168 11772 20220 11824
rect 20536 11815 20588 11824
rect 20536 11781 20545 11815
rect 20545 11781 20579 11815
rect 20579 11781 20588 11815
rect 20536 11772 20588 11781
rect 21364 11772 21416 11824
rect 23388 11840 23440 11892
rect 24308 11840 24360 11892
rect 23572 11772 23624 11824
rect 7564 11704 7616 11756
rect 9956 11704 10008 11756
rect 19524 11747 19576 11756
rect 19524 11713 19533 11747
rect 19533 11713 19567 11747
rect 19567 11713 19576 11747
rect 19524 11704 19576 11713
rect 848 11500 900 11552
rect 2044 11543 2096 11552
rect 2044 11509 2053 11543
rect 2053 11509 2087 11543
rect 2087 11509 2096 11543
rect 2044 11500 2096 11509
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 9588 11636 9640 11688
rect 16856 11636 16908 11688
rect 20076 11747 20128 11756
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 21824 11747 21876 11756
rect 21824 11713 21833 11747
rect 21833 11713 21867 11747
rect 21867 11713 21876 11747
rect 21824 11704 21876 11713
rect 4344 11568 4396 11620
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 4436 11543 4488 11552
rect 4436 11509 4445 11543
rect 4445 11509 4479 11543
rect 4479 11509 4488 11543
rect 4436 11500 4488 11509
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 7748 11568 7800 11620
rect 19524 11568 19576 11620
rect 7104 11543 7156 11552
rect 7104 11509 7113 11543
rect 7113 11509 7147 11543
rect 7147 11509 7156 11543
rect 7104 11500 7156 11509
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 10416 11500 10468 11552
rect 12440 11500 12492 11552
rect 21456 11636 21508 11688
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 22836 11704 22888 11756
rect 24400 11704 24452 11756
rect 26332 11840 26384 11892
rect 27160 11815 27212 11824
rect 27160 11781 27169 11815
rect 27169 11781 27203 11815
rect 27203 11781 27212 11815
rect 27160 11772 27212 11781
rect 21088 11500 21140 11552
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 23388 11500 23440 11552
rect 23664 11500 23716 11552
rect 25504 11704 25556 11756
rect 27436 11704 27488 11756
rect 27896 11747 27948 11756
rect 27896 11713 27905 11747
rect 27905 11713 27939 11747
rect 27939 11713 27948 11747
rect 27896 11704 27948 11713
rect 30380 11840 30432 11892
rect 29000 11772 29052 11824
rect 29920 11772 29972 11824
rect 31392 11772 31444 11824
rect 32404 11815 32456 11824
rect 32404 11781 32413 11815
rect 32413 11781 32447 11815
rect 32447 11781 32456 11815
rect 32404 11772 32456 11781
rect 28724 11747 28776 11756
rect 28724 11713 28733 11747
rect 28733 11713 28767 11747
rect 28767 11713 28776 11747
rect 28724 11704 28776 11713
rect 28816 11747 28868 11756
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 27528 11636 27580 11688
rect 27988 11636 28040 11688
rect 28356 11543 28408 11552
rect 28356 11509 28365 11543
rect 28365 11509 28399 11543
rect 28399 11509 28408 11543
rect 28356 11500 28408 11509
rect 31852 11704 31904 11756
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 34336 11772 34388 11824
rect 33968 11747 34020 11756
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 33968 11704 34020 11713
rect 34612 11840 34664 11892
rect 36176 11840 36228 11892
rect 34796 11815 34848 11824
rect 34796 11781 34805 11815
rect 34805 11781 34839 11815
rect 34839 11781 34848 11815
rect 34796 11772 34848 11781
rect 37280 11840 37332 11892
rect 38844 11772 38896 11824
rect 31576 11679 31628 11688
rect 31576 11645 31585 11679
rect 31585 11645 31619 11679
rect 31619 11645 31628 11679
rect 31576 11636 31628 11645
rect 32588 11636 32640 11688
rect 34520 11679 34572 11688
rect 34520 11645 34529 11679
rect 34529 11645 34563 11679
rect 34563 11645 34572 11679
rect 34520 11636 34572 11645
rect 35256 11636 35308 11688
rect 35532 11636 35584 11688
rect 37832 11747 37884 11756
rect 37832 11713 37841 11747
rect 37841 11713 37875 11747
rect 37875 11713 37884 11747
rect 37832 11704 37884 11713
rect 37924 11704 37976 11756
rect 36452 11636 36504 11688
rect 37740 11679 37792 11688
rect 37740 11645 37749 11679
rect 37749 11645 37783 11679
rect 37783 11645 37792 11679
rect 37740 11636 37792 11645
rect 32864 11568 32916 11620
rect 37556 11611 37608 11620
rect 37556 11577 37565 11611
rect 37565 11577 37599 11611
rect 37599 11577 37608 11611
rect 37556 11568 37608 11577
rect 38200 11679 38252 11688
rect 38200 11645 38209 11679
rect 38209 11645 38243 11679
rect 38243 11645 38252 11679
rect 38200 11636 38252 11645
rect 40776 11679 40828 11688
rect 40776 11645 40785 11679
rect 40785 11645 40819 11679
rect 40819 11645 40828 11679
rect 40776 11636 40828 11645
rect 38844 11568 38896 11620
rect 30840 11500 30892 11552
rect 31300 11500 31352 11552
rect 32220 11500 32272 11552
rect 34428 11543 34480 11552
rect 34428 11509 34437 11543
rect 34437 11509 34471 11543
rect 34471 11509 34480 11543
rect 34428 11500 34480 11509
rect 36360 11543 36412 11552
rect 36360 11509 36369 11543
rect 36369 11509 36403 11543
rect 36403 11509 36412 11543
rect 36360 11500 36412 11509
rect 38384 11543 38436 11552
rect 38384 11509 38393 11543
rect 38393 11509 38427 11543
rect 38427 11509 38436 11543
rect 38384 11500 38436 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1952 11296 2004 11348
rect 2504 11271 2556 11280
rect 2504 11237 2513 11271
rect 2513 11237 2547 11271
rect 2547 11237 2556 11271
rect 2504 11228 2556 11237
rect 2044 11203 2096 11212
rect 2044 11169 2053 11203
rect 2053 11169 2087 11203
rect 2087 11169 2096 11203
rect 2044 11160 2096 11169
rect 6644 11296 6696 11348
rect 4068 11271 4120 11280
rect 4068 11237 4077 11271
rect 4077 11237 4111 11271
rect 4111 11237 4120 11271
rect 4068 11228 4120 11237
rect 5724 11228 5776 11280
rect 2136 11092 2188 11144
rect 2228 11092 2280 11144
rect 3148 11203 3200 11212
rect 3148 11169 3157 11203
rect 3157 11169 3191 11203
rect 3191 11169 3200 11203
rect 3148 11160 3200 11169
rect 3516 11160 3568 11212
rect 5632 11160 5684 11212
rect 7196 11160 7248 11212
rect 7564 11228 7616 11280
rect 9956 11296 10008 11348
rect 9588 11271 9640 11280
rect 9588 11237 9597 11271
rect 9597 11237 9631 11271
rect 9631 11237 9640 11271
rect 9588 11228 9640 11237
rect 10508 11296 10560 11348
rect 14280 11296 14332 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 21456 11339 21508 11348
rect 21456 11305 21465 11339
rect 21465 11305 21499 11339
rect 21499 11305 21508 11339
rect 21456 11296 21508 11305
rect 27528 11339 27580 11348
rect 27528 11305 27537 11339
rect 27537 11305 27571 11339
rect 27571 11305 27580 11339
rect 27528 11296 27580 11305
rect 27896 11296 27948 11348
rect 32588 11296 32640 11348
rect 33968 11296 34020 11348
rect 34704 11296 34756 11348
rect 3884 11135 3936 11144
rect 3884 11101 3893 11135
rect 3893 11101 3927 11135
rect 3927 11101 3936 11135
rect 3884 11092 3936 11101
rect 3424 11024 3476 11076
rect 6092 11092 6144 11144
rect 4804 11024 4856 11076
rect 6920 11092 6972 11144
rect 7104 11092 7156 11144
rect 7380 11024 7432 11076
rect 7748 11092 7800 11144
rect 9404 11092 9456 11144
rect 9496 11135 9548 11154
rect 9496 11102 9505 11135
rect 9505 11102 9539 11135
rect 9539 11102 9548 11135
rect 8116 11024 8168 11076
rect 14556 11228 14608 11280
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 11428 11160 11480 11212
rect 13176 11160 13228 11212
rect 13084 11092 13136 11144
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 18788 11135 18840 11144
rect 18788 11101 18797 11135
rect 18797 11101 18831 11135
rect 18831 11101 18840 11135
rect 18788 11092 18840 11101
rect 19432 11160 19484 11212
rect 20444 11160 20496 11212
rect 21640 11160 21692 11212
rect 26148 11160 26200 11212
rect 19524 11092 19576 11144
rect 23388 11092 23440 11144
rect 24860 11092 24912 11144
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 25780 11092 25832 11101
rect 33600 11228 33652 11280
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 3148 10956 3200 11008
rect 5264 10956 5316 11008
rect 5816 10956 5868 11008
rect 7564 10956 7616 11008
rect 7932 10999 7984 11008
rect 7932 10965 7941 10999
rect 7941 10965 7975 10999
rect 7975 10965 7984 10999
rect 7932 10956 7984 10965
rect 9634 10956 9686 11008
rect 9772 10956 9824 11008
rect 10232 10956 10284 11008
rect 11888 11024 11940 11076
rect 13912 11024 13964 11076
rect 19340 11024 19392 11076
rect 19616 11024 19668 11076
rect 20168 11024 20220 11076
rect 18880 10956 18932 11008
rect 24400 11024 24452 11076
rect 20812 10956 20864 11008
rect 27436 11024 27488 11076
rect 30380 11160 30432 11212
rect 27988 11135 28040 11144
rect 27988 11101 27997 11135
rect 27997 11101 28031 11135
rect 28031 11101 28040 11135
rect 27988 11092 28040 11101
rect 28080 11135 28132 11144
rect 28080 11101 28089 11135
rect 28089 11101 28123 11135
rect 28123 11101 28132 11135
rect 28080 11092 28132 11101
rect 28724 11092 28776 11144
rect 31300 11135 31352 11144
rect 31300 11101 31309 11135
rect 31309 11101 31343 11135
rect 31343 11101 31352 11135
rect 31300 11092 31352 11101
rect 32404 11160 32456 11212
rect 32496 11160 32548 11212
rect 31760 11092 31812 11144
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 34336 11160 34388 11212
rect 35992 11296 36044 11348
rect 36268 11339 36320 11348
rect 36268 11305 36277 11339
rect 36277 11305 36311 11339
rect 36311 11305 36320 11339
rect 36268 11296 36320 11305
rect 35532 11203 35584 11212
rect 35532 11169 35541 11203
rect 35541 11169 35575 11203
rect 35575 11169 35584 11203
rect 35532 11160 35584 11169
rect 27896 11024 27948 11076
rect 28356 11024 28408 11076
rect 29276 10956 29328 11008
rect 34244 11135 34296 11144
rect 34244 11101 34253 11135
rect 34253 11101 34287 11135
rect 34287 11101 34296 11135
rect 34244 11092 34296 11101
rect 34520 11092 34572 11144
rect 34796 11092 34848 11144
rect 36360 11160 36412 11212
rect 37372 11296 37424 11348
rect 37832 11339 37884 11348
rect 37832 11305 37841 11339
rect 37841 11305 37875 11339
rect 37875 11305 37884 11339
rect 37832 11296 37884 11305
rect 38844 11296 38896 11348
rect 37004 11160 37056 11212
rect 38108 11203 38160 11212
rect 38108 11169 38117 11203
rect 38117 11169 38151 11203
rect 38151 11169 38160 11203
rect 38108 11160 38160 11169
rect 39488 11203 39540 11212
rect 39488 11169 39497 11203
rect 39497 11169 39531 11203
rect 39531 11169 39540 11203
rect 39488 11160 39540 11169
rect 37188 11135 37240 11144
rect 37188 11101 37197 11135
rect 37197 11101 37231 11135
rect 37231 11101 37240 11135
rect 37188 11092 37240 11101
rect 37464 11135 37516 11144
rect 37464 11101 37473 11135
rect 37473 11101 37507 11135
rect 37507 11101 37516 11135
rect 37464 11092 37516 11101
rect 37648 11092 37700 11144
rect 38384 11092 38436 11144
rect 34428 11024 34480 11076
rect 34244 10956 34296 11008
rect 35992 10956 36044 11008
rect 37464 10956 37516 11008
rect 37740 10956 37792 11008
rect 37924 10956 37976 11008
rect 38568 10956 38620 11008
rect 40868 10956 40920 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 2504 10752 2556 10804
rect 3884 10752 3936 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 6092 10795 6144 10804
rect 6092 10761 6101 10795
rect 6101 10761 6135 10795
rect 6135 10761 6144 10795
rect 6092 10752 6144 10761
rect 2964 10684 3016 10736
rect 7656 10752 7708 10804
rect 7748 10752 7800 10804
rect 8116 10752 8168 10804
rect 6736 10727 6788 10736
rect 6736 10693 6745 10727
rect 6745 10693 6779 10727
rect 6779 10693 6788 10727
rect 6736 10684 6788 10693
rect 7012 10684 7064 10736
rect 10048 10752 10100 10804
rect 17960 10752 18012 10804
rect 9956 10727 10008 10736
rect 9956 10693 9965 10727
rect 9965 10693 9999 10727
rect 9999 10693 10008 10727
rect 9956 10684 10008 10693
rect 10692 10727 10744 10736
rect 10692 10693 10701 10727
rect 10701 10693 10735 10727
rect 10735 10693 10744 10727
rect 10692 10684 10744 10693
rect 17868 10684 17920 10736
rect 18788 10752 18840 10804
rect 20536 10752 20588 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 22100 10752 22152 10804
rect 23020 10752 23072 10804
rect 18880 10684 18932 10736
rect 20260 10684 20312 10736
rect 4620 10616 4672 10668
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 10600 10616 10652 10668
rect 1400 10591 1452 10600
rect 1400 10557 1409 10591
rect 1409 10557 1443 10591
rect 1443 10557 1452 10591
rect 1400 10548 1452 10557
rect 6828 10548 6880 10600
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 6276 10412 6328 10464
rect 7380 10480 7432 10532
rect 9864 10548 9916 10600
rect 11428 10548 11480 10600
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 16856 10591 16908 10600
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 18328 10548 18380 10600
rect 20168 10591 20220 10600
rect 20168 10557 20177 10591
rect 20177 10557 20211 10591
rect 20211 10557 20220 10591
rect 20168 10548 20220 10557
rect 11704 10480 11756 10532
rect 7840 10412 7892 10464
rect 9588 10412 9640 10464
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 10508 10412 10560 10421
rect 11152 10412 11204 10464
rect 19156 10412 19208 10464
rect 19524 10412 19576 10464
rect 21364 10684 21416 10736
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 25504 10752 25556 10804
rect 28080 10795 28132 10804
rect 28080 10761 28089 10795
rect 28089 10761 28123 10795
rect 28123 10761 28132 10795
rect 28080 10752 28132 10761
rect 28172 10752 28224 10804
rect 29092 10752 29144 10804
rect 29552 10752 29604 10804
rect 32128 10752 32180 10804
rect 24860 10727 24912 10736
rect 24860 10693 24869 10727
rect 24869 10693 24903 10727
rect 24903 10693 24912 10727
rect 24860 10684 24912 10693
rect 25596 10727 25648 10736
rect 25596 10693 25605 10727
rect 25605 10693 25639 10727
rect 25639 10693 25648 10727
rect 25596 10684 25648 10693
rect 34520 10752 34572 10804
rect 21180 10480 21232 10532
rect 22744 10659 22796 10668
rect 22744 10625 22753 10659
rect 22753 10625 22787 10659
rect 22787 10625 22796 10659
rect 22744 10616 22796 10625
rect 22192 10548 22244 10600
rect 22192 10412 22244 10464
rect 22284 10412 22336 10464
rect 22928 10480 22980 10532
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 23848 10548 23900 10600
rect 24676 10548 24728 10600
rect 25688 10591 25740 10600
rect 25688 10557 25697 10591
rect 25697 10557 25731 10591
rect 25731 10557 25740 10591
rect 25688 10548 25740 10557
rect 26516 10548 26568 10600
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 27528 10659 27580 10668
rect 27528 10625 27537 10659
rect 27537 10625 27571 10659
rect 27571 10625 27580 10659
rect 27528 10616 27580 10625
rect 28816 10616 28868 10668
rect 27620 10548 27672 10600
rect 28724 10548 28776 10600
rect 29092 10659 29144 10668
rect 29092 10625 29101 10659
rect 29101 10625 29135 10659
rect 29135 10625 29144 10659
rect 29092 10616 29144 10625
rect 29736 10616 29788 10668
rect 34152 10684 34204 10736
rect 34980 10684 35032 10736
rect 35348 10684 35400 10736
rect 30656 10616 30708 10668
rect 36176 10752 36228 10804
rect 38108 10752 38160 10804
rect 40776 10752 40828 10804
rect 35992 10727 36044 10736
rect 35992 10693 36001 10727
rect 36001 10693 36035 10727
rect 36035 10693 36044 10727
rect 35992 10684 36044 10693
rect 36176 10659 36228 10668
rect 36176 10625 36185 10659
rect 36185 10625 36219 10659
rect 36219 10625 36228 10659
rect 36176 10616 36228 10625
rect 36912 10616 36964 10668
rect 37372 10616 37424 10668
rect 40684 10684 40736 10736
rect 37740 10616 37792 10668
rect 29092 10480 29144 10532
rect 23940 10455 23992 10464
rect 23940 10421 23949 10455
rect 23949 10421 23983 10455
rect 23983 10421 23992 10455
rect 23940 10412 23992 10421
rect 26976 10455 27028 10464
rect 26976 10421 26985 10455
rect 26985 10421 27019 10455
rect 27019 10421 27028 10455
rect 26976 10412 27028 10421
rect 27344 10412 27396 10464
rect 28172 10412 28224 10464
rect 28908 10412 28960 10464
rect 32404 10591 32456 10600
rect 32404 10557 32413 10591
rect 32413 10557 32447 10591
rect 32447 10557 32456 10591
rect 32404 10548 32456 10557
rect 34796 10548 34848 10600
rect 37924 10659 37976 10668
rect 37924 10625 37933 10659
rect 37933 10625 37967 10659
rect 37967 10625 37976 10659
rect 37924 10616 37976 10625
rect 38016 10659 38068 10668
rect 38016 10625 38025 10659
rect 38025 10625 38059 10659
rect 38059 10625 38068 10659
rect 38016 10616 38068 10625
rect 38384 10616 38436 10668
rect 38476 10659 38528 10668
rect 38476 10625 38485 10659
rect 38485 10625 38519 10659
rect 38519 10625 38528 10659
rect 38476 10616 38528 10625
rect 38568 10659 38620 10668
rect 38568 10625 38577 10659
rect 38577 10625 38611 10659
rect 38611 10625 38620 10659
rect 38568 10616 38620 10625
rect 38844 10616 38896 10668
rect 32588 10412 32640 10464
rect 33876 10455 33928 10464
rect 33876 10421 33885 10455
rect 33885 10421 33919 10455
rect 33919 10421 33928 10455
rect 33876 10412 33928 10421
rect 34152 10412 34204 10464
rect 34704 10412 34756 10464
rect 38108 10548 38160 10600
rect 41880 10616 41932 10668
rect 39396 10480 39448 10532
rect 38476 10412 38528 10464
rect 38936 10412 38988 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 3424 10208 3476 10260
rect 5540 10208 5592 10260
rect 6184 10251 6236 10260
rect 6184 10217 6193 10251
rect 6193 10217 6227 10251
rect 6227 10217 6236 10251
rect 6184 10208 6236 10217
rect 2688 10072 2740 10124
rect 7012 10208 7064 10260
rect 7104 10208 7156 10260
rect 9864 10251 9916 10260
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10600 10208 10652 10260
rect 6644 10140 6696 10192
rect 7196 10072 7248 10124
rect 7472 10140 7524 10192
rect 5448 10004 5500 10056
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 6276 10004 6328 10056
rect 7472 10004 7524 10056
rect 4620 9936 4672 9988
rect 6644 9979 6696 9988
rect 6644 9945 6653 9979
rect 6653 9945 6687 9979
rect 6687 9945 6696 9979
rect 6644 9936 6696 9945
rect 6920 9936 6972 9988
rect 8024 10072 8076 10124
rect 9312 10072 9364 10124
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 12900 10208 12952 10260
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 5264 9868 5316 9920
rect 6552 9868 6604 9920
rect 6828 9868 6880 9920
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 7840 9979 7892 9988
rect 7840 9945 7849 9979
rect 7849 9945 7883 9979
rect 7883 9945 7892 9979
rect 7840 9936 7892 9945
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 10508 9979 10560 9988
rect 10508 9945 10517 9979
rect 10517 9945 10551 9979
rect 10551 9945 10560 9979
rect 10508 9936 10560 9945
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 9772 9868 9824 9920
rect 11336 10072 11388 10124
rect 11980 10072 12032 10124
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11428 10004 11480 10056
rect 17960 9936 18012 9988
rect 18144 10072 18196 10124
rect 19708 10208 19760 10260
rect 20168 10208 20220 10260
rect 22008 10251 22060 10260
rect 22008 10217 22017 10251
rect 22017 10217 22051 10251
rect 22051 10217 22060 10251
rect 22008 10208 22060 10217
rect 23112 10208 23164 10260
rect 24216 10251 24268 10260
rect 24216 10217 24225 10251
rect 24225 10217 24259 10251
rect 24259 10217 24268 10251
rect 24216 10208 24268 10217
rect 25872 10208 25924 10260
rect 26976 10208 27028 10260
rect 27896 10208 27948 10260
rect 29000 10208 29052 10260
rect 29368 10208 29420 10260
rect 30656 10251 30708 10260
rect 30656 10217 30665 10251
rect 30665 10217 30699 10251
rect 30699 10217 30708 10251
rect 30656 10208 30708 10217
rect 31024 10208 31076 10260
rect 32404 10208 32456 10260
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 19248 10072 19300 10124
rect 20260 10047 20312 10056
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 20536 10047 20588 10056
rect 20536 10013 20545 10047
rect 20545 10013 20579 10047
rect 20579 10013 20588 10047
rect 20536 10004 20588 10013
rect 23756 10072 23808 10124
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 22928 10047 22980 10056
rect 22928 10013 22937 10047
rect 22937 10013 22971 10047
rect 22971 10013 22980 10047
rect 22928 10004 22980 10013
rect 28816 10140 28868 10192
rect 31484 10140 31536 10192
rect 24124 10072 24176 10124
rect 24216 10072 24268 10124
rect 24400 10072 24452 10124
rect 25780 10072 25832 10124
rect 34704 10140 34756 10192
rect 13544 9868 13596 9920
rect 18236 9868 18288 9920
rect 19616 9936 19668 9988
rect 21180 9936 21232 9988
rect 19800 9868 19852 9920
rect 21272 9868 21324 9920
rect 28724 10004 28776 10056
rect 29184 10004 29236 10056
rect 29276 10047 29328 10056
rect 29276 10013 29285 10047
rect 29285 10013 29319 10047
rect 29319 10013 29328 10047
rect 29276 10004 29328 10013
rect 26424 9936 26476 9988
rect 27344 9936 27396 9988
rect 27712 9936 27764 9988
rect 27896 9936 27948 9988
rect 30472 9979 30524 9988
rect 30472 9945 30481 9979
rect 30481 9945 30515 9979
rect 30515 9945 30524 9979
rect 30472 9936 30524 9945
rect 29092 9911 29144 9920
rect 29092 9877 29101 9911
rect 29101 9877 29135 9911
rect 29135 9877 29144 9911
rect 29092 9868 29144 9877
rect 29184 9868 29236 9920
rect 31024 10047 31076 10056
rect 31024 10013 31033 10047
rect 31033 10013 31067 10047
rect 31067 10013 31076 10047
rect 31024 10004 31076 10013
rect 31668 10004 31720 10056
rect 31760 10047 31812 10056
rect 31760 10013 31769 10047
rect 31769 10013 31803 10047
rect 31803 10013 31812 10047
rect 31760 10004 31812 10013
rect 31208 9979 31260 9988
rect 31208 9945 31217 9979
rect 31217 9945 31251 9979
rect 31251 9945 31260 9979
rect 31208 9936 31260 9945
rect 33784 10072 33836 10124
rect 33876 10115 33928 10124
rect 33876 10081 33885 10115
rect 33885 10081 33919 10115
rect 33919 10081 33928 10115
rect 33876 10072 33928 10081
rect 32496 10004 32548 10056
rect 33324 10047 33376 10056
rect 33324 10013 33333 10047
rect 33333 10013 33367 10047
rect 33367 10013 33376 10047
rect 33324 10004 33376 10013
rect 31116 9868 31168 9920
rect 32772 9979 32824 9988
rect 32772 9945 32781 9979
rect 32781 9945 32815 9979
rect 32815 9945 32824 9979
rect 32772 9936 32824 9945
rect 33876 9936 33928 9988
rect 36912 10115 36964 10124
rect 36912 10081 36921 10115
rect 36921 10081 36955 10115
rect 36955 10081 36964 10115
rect 36912 10072 36964 10081
rect 37556 10140 37608 10192
rect 37740 10208 37792 10260
rect 38108 10140 38160 10192
rect 38568 10140 38620 10192
rect 40316 10140 40368 10192
rect 37372 10004 37424 10056
rect 37464 10047 37516 10056
rect 37464 10013 37473 10047
rect 37473 10013 37507 10047
rect 37507 10013 37516 10047
rect 37464 10004 37516 10013
rect 37648 10004 37700 10056
rect 38016 10072 38068 10124
rect 38936 10004 38988 10056
rect 39028 10047 39080 10056
rect 39028 10013 39037 10047
rect 39037 10013 39071 10047
rect 39071 10013 39080 10047
rect 39028 10004 39080 10013
rect 40684 10072 40736 10124
rect 40592 10047 40644 10056
rect 40592 10013 40601 10047
rect 40601 10013 40635 10047
rect 40635 10013 40644 10047
rect 40592 10004 40644 10013
rect 31944 9868 31996 9920
rect 32312 9868 32364 9920
rect 34336 9979 34388 9988
rect 34336 9945 34345 9979
rect 34345 9945 34379 9979
rect 34379 9945 34388 9979
rect 34336 9936 34388 9945
rect 34152 9911 34204 9920
rect 34152 9877 34161 9911
rect 34161 9877 34195 9911
rect 34195 9877 34204 9911
rect 34152 9868 34204 9877
rect 37556 9868 37608 9920
rect 37648 9868 37700 9920
rect 38200 9936 38252 9988
rect 39304 9979 39356 9988
rect 39304 9945 39313 9979
rect 39313 9945 39347 9979
rect 39347 9945 39356 9979
rect 41788 10208 41840 10260
rect 39304 9936 39356 9945
rect 38936 9868 38988 9920
rect 39856 9868 39908 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 3424 9664 3476 9716
rect 3240 9596 3292 9648
rect 1400 9528 1452 9580
rect 2688 9528 2740 9580
rect 6644 9664 6696 9716
rect 7104 9707 7156 9716
rect 7104 9673 7113 9707
rect 7113 9673 7147 9707
rect 7147 9673 7156 9707
rect 7104 9664 7156 9673
rect 5448 9596 5500 9648
rect 6000 9639 6052 9648
rect 6000 9605 6009 9639
rect 6009 9605 6043 9639
rect 6043 9605 6052 9639
rect 7840 9664 7892 9716
rect 13544 9664 13596 9716
rect 25688 9664 25740 9716
rect 25872 9664 25924 9716
rect 6000 9596 6052 9605
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 8024 9596 8076 9648
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 5632 9571 5684 9580
rect 5632 9537 5641 9571
rect 5641 9537 5675 9571
rect 5675 9537 5684 9571
rect 5632 9528 5684 9537
rect 5632 9392 5684 9444
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 7932 9528 7984 9580
rect 11704 9596 11756 9648
rect 12440 9596 12492 9648
rect 23940 9596 23992 9648
rect 24216 9596 24268 9648
rect 27528 9664 27580 9716
rect 27712 9664 27764 9716
rect 28264 9664 28316 9716
rect 6644 9460 6696 9469
rect 9772 9460 9824 9512
rect 20904 9528 20956 9580
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 10508 9460 10560 9512
rect 10968 9460 11020 9512
rect 11428 9460 11480 9512
rect 11152 9392 11204 9444
rect 5540 9324 5592 9376
rect 8300 9324 8352 9376
rect 9680 9367 9732 9376
rect 9680 9333 9689 9367
rect 9689 9333 9723 9367
rect 9723 9333 9732 9367
rect 9680 9324 9732 9333
rect 10692 9324 10744 9376
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 21824 9503 21876 9512
rect 21824 9469 21833 9503
rect 21833 9469 21867 9503
rect 21867 9469 21876 9503
rect 21824 9460 21876 9469
rect 22928 9460 22980 9512
rect 23388 9503 23440 9512
rect 23388 9469 23397 9503
rect 23397 9469 23431 9503
rect 23431 9469 23440 9503
rect 23388 9460 23440 9469
rect 26608 9528 26660 9580
rect 27344 9639 27396 9648
rect 27344 9605 27353 9639
rect 27353 9605 27387 9639
rect 27387 9605 27396 9639
rect 27344 9596 27396 9605
rect 28080 9596 28132 9648
rect 27160 9528 27212 9580
rect 28816 9596 28868 9648
rect 28908 9639 28960 9648
rect 28908 9605 28917 9639
rect 28917 9605 28951 9639
rect 28951 9605 28960 9639
rect 28908 9596 28960 9605
rect 29368 9596 29420 9648
rect 30564 9664 30616 9716
rect 30748 9596 30800 9648
rect 31576 9596 31628 9648
rect 31668 9639 31720 9648
rect 31668 9605 31677 9639
rect 31677 9605 31711 9639
rect 31711 9605 31720 9639
rect 31668 9596 31720 9605
rect 31944 9596 31996 9648
rect 33876 9664 33928 9716
rect 36084 9664 36136 9716
rect 36912 9664 36964 9716
rect 37004 9664 37056 9716
rect 38936 9664 38988 9716
rect 39028 9707 39080 9716
rect 39028 9673 39037 9707
rect 39037 9673 39071 9707
rect 39071 9673 39080 9707
rect 39028 9664 39080 9673
rect 40684 9664 40736 9716
rect 31484 9571 31536 9580
rect 31484 9537 31493 9571
rect 31493 9537 31527 9571
rect 31527 9537 31536 9571
rect 31484 9528 31536 9537
rect 33140 9571 33192 9580
rect 33140 9537 33149 9571
rect 33149 9537 33183 9571
rect 33183 9537 33192 9571
rect 33140 9528 33192 9537
rect 33232 9571 33284 9580
rect 33232 9537 33241 9571
rect 33241 9537 33275 9571
rect 33275 9537 33284 9571
rect 33232 9528 33284 9537
rect 33324 9571 33376 9580
rect 33324 9537 33333 9571
rect 33333 9537 33367 9571
rect 33367 9537 33376 9571
rect 33324 9528 33376 9537
rect 34152 9596 34204 9648
rect 34060 9528 34112 9580
rect 34336 9596 34388 9648
rect 34704 9639 34756 9648
rect 34704 9605 34713 9639
rect 34713 9605 34747 9639
rect 34747 9605 34756 9639
rect 34704 9596 34756 9605
rect 37556 9639 37608 9648
rect 37556 9605 37565 9639
rect 37565 9605 37599 9639
rect 37599 9605 37608 9639
rect 37556 9596 37608 9605
rect 39304 9596 39356 9648
rect 39396 9639 39448 9648
rect 39396 9605 39405 9639
rect 39405 9605 39439 9639
rect 39439 9605 39448 9639
rect 39396 9596 39448 9605
rect 39856 9596 39908 9648
rect 26240 9503 26292 9512
rect 26240 9469 26249 9503
rect 26249 9469 26283 9503
rect 26283 9469 26292 9503
rect 26240 9460 26292 9469
rect 26884 9460 26936 9512
rect 27068 9460 27120 9512
rect 28080 9503 28132 9512
rect 28080 9469 28089 9503
rect 28089 9469 28123 9503
rect 28123 9469 28132 9503
rect 28080 9460 28132 9469
rect 28540 9503 28592 9512
rect 28540 9469 28549 9503
rect 28549 9469 28583 9503
rect 28583 9469 28592 9503
rect 28540 9460 28592 9469
rect 28632 9503 28684 9512
rect 28632 9469 28641 9503
rect 28641 9469 28675 9503
rect 28675 9469 28684 9503
rect 28632 9460 28684 9469
rect 29276 9460 29328 9512
rect 29552 9460 29604 9512
rect 30472 9460 30524 9512
rect 31208 9460 31260 9512
rect 31300 9460 31352 9512
rect 32496 9460 32548 9512
rect 22376 9324 22428 9376
rect 22836 9324 22888 9376
rect 24032 9324 24084 9376
rect 24676 9324 24728 9376
rect 26700 9367 26752 9376
rect 26700 9333 26709 9367
rect 26709 9333 26743 9367
rect 26743 9333 26752 9367
rect 26700 9324 26752 9333
rect 27620 9324 27672 9376
rect 29000 9324 29052 9376
rect 33140 9392 33192 9444
rect 30380 9324 30432 9376
rect 31300 9324 31352 9376
rect 31852 9324 31904 9376
rect 33876 9503 33928 9512
rect 33876 9469 33885 9503
rect 33885 9469 33919 9503
rect 33919 9469 33928 9503
rect 33876 9460 33928 9469
rect 34796 9528 34848 9580
rect 35532 9571 35584 9580
rect 35532 9537 35541 9571
rect 35541 9537 35575 9571
rect 35575 9537 35584 9571
rect 35532 9528 35584 9537
rect 37280 9571 37332 9580
rect 37280 9537 37289 9571
rect 37289 9537 37323 9571
rect 37323 9537 37332 9571
rect 37280 9528 37332 9537
rect 35716 9460 35768 9512
rect 35348 9392 35400 9444
rect 34152 9324 34204 9376
rect 34520 9324 34572 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3884 9120 3936 9172
rect 5448 9163 5500 9172
rect 5448 9129 5457 9163
rect 5457 9129 5491 9163
rect 5491 9129 5500 9163
rect 5448 9120 5500 9129
rect 6000 9120 6052 9172
rect 6184 9120 6236 9172
rect 10968 9120 11020 9172
rect 11796 9120 11848 9172
rect 20904 9163 20956 9172
rect 20904 9129 20913 9163
rect 20913 9129 20947 9163
rect 20947 9129 20956 9163
rect 20904 9120 20956 9129
rect 3240 8984 3292 9036
rect 7472 8984 7524 9036
rect 10692 8984 10744 9036
rect 4068 8916 4120 8968
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5540 8916 5592 8968
rect 6000 8959 6052 8968
rect 6000 8925 6009 8959
rect 6009 8925 6043 8959
rect 6043 8925 6052 8959
rect 6000 8916 6052 8925
rect 7104 8916 7156 8968
rect 11152 8916 11204 8968
rect 11336 8916 11388 8968
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 10232 8848 10284 8900
rect 20260 9052 20312 9104
rect 20996 9052 21048 9104
rect 19524 8984 19576 9036
rect 20812 8984 20864 9036
rect 23664 9120 23716 9172
rect 24124 9120 24176 9172
rect 24676 9120 24728 9172
rect 28540 9120 28592 9172
rect 31760 9120 31812 9172
rect 24400 9052 24452 9104
rect 26884 9052 26936 9104
rect 22376 9027 22428 9036
rect 22376 8993 22385 9027
rect 22385 8993 22419 9027
rect 22419 8993 22428 9027
rect 22376 8984 22428 8993
rect 23756 8984 23808 9036
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 19616 8891 19668 8900
rect 19616 8857 19625 8891
rect 19625 8857 19659 8891
rect 19659 8857 19668 8891
rect 19616 8848 19668 8857
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 26608 8916 26660 8968
rect 26700 8959 26752 8968
rect 27620 8984 27672 9036
rect 26700 8925 26739 8959
rect 26739 8925 26752 8959
rect 26700 8916 26752 8925
rect 27528 8959 27580 8968
rect 27528 8925 27537 8959
rect 27537 8925 27571 8959
rect 27571 8925 27580 8959
rect 27528 8916 27580 8925
rect 28448 8916 28500 8968
rect 30472 9052 30524 9104
rect 33140 9120 33192 9172
rect 33324 9120 33376 9172
rect 32956 9052 33008 9104
rect 30748 9027 30800 9036
rect 29000 8959 29052 8968
rect 29000 8925 29009 8959
rect 29009 8925 29043 8959
rect 29043 8925 29052 8959
rect 29000 8916 29052 8925
rect 29092 8959 29144 8968
rect 29092 8925 29101 8959
rect 29101 8925 29135 8959
rect 29135 8925 29144 8959
rect 29092 8916 29144 8925
rect 29184 8959 29236 8968
rect 29184 8925 29193 8959
rect 29193 8925 29227 8959
rect 29227 8925 29236 8959
rect 29184 8916 29236 8925
rect 30748 8993 30757 9027
rect 30757 8993 30791 9027
rect 30791 8993 30800 9027
rect 30748 8984 30800 8993
rect 32128 8916 32180 8968
rect 33048 8984 33100 9036
rect 33876 9120 33928 9172
rect 33968 9120 34020 9172
rect 34612 9120 34664 9172
rect 35256 9120 35308 9172
rect 35532 9120 35584 9172
rect 37372 9120 37424 9172
rect 38476 9120 38528 9172
rect 33600 9052 33652 9104
rect 32864 8916 32916 8968
rect 3608 8780 3660 8832
rect 4804 8780 4856 8832
rect 5724 8780 5776 8832
rect 6460 8780 6512 8832
rect 20352 8780 20404 8832
rect 22100 8780 22152 8832
rect 24124 8848 24176 8900
rect 23848 8780 23900 8832
rect 28080 8848 28132 8900
rect 27160 8780 27212 8832
rect 27436 8780 27488 8832
rect 28172 8823 28224 8832
rect 28172 8789 28181 8823
rect 28181 8789 28215 8823
rect 28215 8789 28224 8823
rect 28172 8780 28224 8789
rect 28356 8780 28408 8832
rect 29276 8780 29328 8832
rect 29460 8780 29512 8832
rect 31668 8780 31720 8832
rect 34336 8959 34388 8968
rect 34336 8925 34345 8959
rect 34345 8925 34379 8959
rect 34379 8925 34388 8959
rect 34336 8916 34388 8925
rect 35348 8916 35400 8968
rect 35716 8984 35768 9036
rect 37372 8984 37424 9036
rect 34612 8848 34664 8900
rect 37280 8848 37332 8900
rect 37832 8916 37884 8968
rect 37924 8848 37976 8900
rect 34428 8780 34480 8832
rect 34704 8780 34756 8832
rect 35164 8780 35216 8832
rect 37648 8780 37700 8832
rect 37740 8823 37792 8832
rect 37740 8789 37749 8823
rect 37749 8789 37783 8823
rect 37783 8789 37792 8823
rect 37740 8780 37792 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 3240 8508 3292 8560
rect 3976 8508 4028 8560
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 3792 8440 3844 8492
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 6644 8576 6696 8628
rect 6920 8576 6972 8628
rect 19524 8576 19576 8628
rect 21364 8576 21416 8628
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2688 8372 2740 8424
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 6828 8508 6880 8560
rect 7012 8508 7064 8560
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 3792 8304 3844 8356
rect 4068 8304 4120 8356
rect 4896 8372 4948 8424
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 7196 8440 7248 8492
rect 8668 8508 8720 8560
rect 20352 8551 20404 8560
rect 20352 8517 20361 8551
rect 20361 8517 20395 8551
rect 20395 8517 20404 8551
rect 20352 8508 20404 8517
rect 20720 8551 20772 8560
rect 20720 8517 20729 8551
rect 20729 8517 20763 8551
rect 20763 8517 20772 8551
rect 20720 8508 20772 8517
rect 23664 8508 23716 8560
rect 6920 8372 6972 8424
rect 5540 8304 5592 8356
rect 5632 8304 5684 8356
rect 7012 8304 7064 8356
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 16856 8440 16908 8492
rect 18328 8440 18380 8492
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 8760 8372 8812 8424
rect 19156 8372 19208 8424
rect 22376 8440 22428 8492
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 26424 8576 26476 8628
rect 28908 8576 28960 8628
rect 26516 8551 26568 8560
rect 23848 8372 23900 8424
rect 24032 8372 24084 8424
rect 24400 8483 24452 8492
rect 24400 8449 24409 8483
rect 24409 8449 24443 8483
rect 24443 8449 24452 8483
rect 24400 8440 24452 8449
rect 25228 8440 25280 8492
rect 26516 8517 26525 8551
rect 26525 8517 26559 8551
rect 26559 8517 26568 8551
rect 26516 8508 26568 8517
rect 26424 8483 26476 8492
rect 26424 8449 26433 8483
rect 26433 8449 26467 8483
rect 26467 8449 26476 8483
rect 26424 8440 26476 8449
rect 28172 8508 28224 8560
rect 28356 8551 28408 8560
rect 28356 8517 28365 8551
rect 28365 8517 28399 8551
rect 28399 8517 28408 8551
rect 28356 8508 28408 8517
rect 27068 8440 27120 8492
rect 27436 8440 27488 8492
rect 5448 8279 5500 8288
rect 5448 8245 5457 8279
rect 5457 8245 5491 8279
rect 5491 8245 5500 8279
rect 5448 8236 5500 8245
rect 6644 8236 6696 8288
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 8208 8236 8260 8245
rect 10324 8304 10376 8356
rect 11152 8304 11204 8356
rect 19340 8304 19392 8356
rect 20996 8304 21048 8356
rect 21364 8304 21416 8356
rect 27160 8372 27212 8424
rect 30380 8576 30432 8628
rect 32864 8619 32916 8628
rect 32864 8585 32873 8619
rect 32873 8585 32907 8619
rect 32907 8585 32916 8619
rect 32864 8576 32916 8585
rect 29460 8483 29512 8492
rect 29460 8449 29469 8483
rect 29469 8449 29503 8483
rect 29503 8449 29512 8483
rect 29460 8440 29512 8449
rect 29552 8440 29604 8492
rect 30748 8508 30800 8560
rect 32956 8508 33008 8560
rect 31576 8440 31628 8492
rect 26332 8304 26384 8356
rect 28080 8304 28132 8356
rect 29184 8415 29236 8424
rect 29184 8381 29193 8415
rect 29193 8381 29227 8415
rect 29227 8381 29236 8415
rect 29184 8372 29236 8381
rect 29276 8415 29328 8424
rect 29276 8381 29285 8415
rect 29285 8381 29319 8415
rect 29319 8381 29328 8415
rect 29276 8372 29328 8381
rect 30472 8415 30524 8424
rect 30472 8381 30481 8415
rect 30481 8381 30515 8415
rect 30515 8381 30524 8415
rect 30472 8372 30524 8381
rect 23480 8279 23532 8288
rect 23480 8245 23489 8279
rect 23489 8245 23523 8279
rect 23523 8245 23532 8279
rect 23480 8236 23532 8245
rect 25412 8236 25464 8288
rect 28264 8236 28316 8288
rect 29828 8236 29880 8288
rect 30564 8236 30616 8288
rect 31944 8236 31996 8288
rect 33140 8483 33192 8492
rect 33140 8449 33149 8483
rect 33149 8449 33183 8483
rect 33183 8449 33192 8483
rect 33140 8440 33192 8449
rect 33324 8440 33376 8492
rect 33968 8508 34020 8560
rect 34336 8576 34388 8628
rect 34428 8576 34480 8628
rect 35440 8508 35492 8560
rect 37832 8551 37884 8560
rect 37832 8517 37841 8551
rect 37841 8517 37875 8551
rect 37875 8517 37884 8551
rect 37832 8508 37884 8517
rect 34244 8440 34296 8492
rect 32956 8372 33008 8424
rect 35164 8440 35216 8492
rect 36268 8440 36320 8492
rect 37648 8440 37700 8492
rect 34796 8415 34848 8424
rect 34796 8381 34805 8415
rect 34805 8381 34839 8415
rect 34839 8381 34848 8415
rect 34796 8372 34848 8381
rect 35440 8415 35492 8424
rect 35440 8381 35449 8415
rect 35449 8381 35483 8415
rect 35483 8381 35492 8415
rect 35440 8372 35492 8381
rect 34060 8304 34112 8356
rect 37464 8415 37516 8424
rect 37464 8381 37473 8415
rect 37473 8381 37507 8415
rect 37507 8381 37516 8415
rect 37464 8372 37516 8381
rect 35900 8304 35952 8356
rect 33232 8236 33284 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2320 8032 2372 8084
rect 4436 8032 4488 8084
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 4620 7896 4672 7948
rect 4804 7896 4856 7948
rect 2964 7760 3016 7812
rect 3608 7803 3660 7812
rect 3608 7769 3617 7803
rect 3617 7769 3651 7803
rect 3651 7769 3660 7803
rect 3608 7760 3660 7769
rect 4068 7828 4120 7880
rect 4528 7828 4580 7880
rect 6092 8032 6144 8084
rect 6828 8032 6880 8084
rect 7380 7964 7432 8016
rect 8024 8032 8076 8084
rect 7840 8007 7892 8016
rect 7840 7973 7849 8007
rect 7849 7973 7883 8007
rect 7883 7973 7892 8007
rect 7840 7964 7892 7973
rect 8668 8032 8720 8084
rect 9036 8032 9088 8084
rect 19432 8032 19484 8084
rect 19892 8032 19944 8084
rect 25228 8075 25280 8084
rect 25228 8041 25237 8075
rect 25237 8041 25271 8075
rect 25271 8041 25280 8075
rect 25228 8032 25280 8041
rect 27528 8032 27580 8084
rect 28632 8032 28684 8084
rect 5632 7828 5684 7880
rect 6092 7828 6144 7880
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7380 7828 7432 7880
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 23388 7896 23440 7948
rect 25688 7939 25740 7948
rect 25688 7905 25697 7939
rect 25697 7905 25731 7939
rect 25731 7905 25740 7939
rect 25688 7896 25740 7905
rect 26332 7896 26384 7948
rect 27436 7896 27488 7948
rect 28908 7896 28960 7948
rect 30472 8032 30524 8084
rect 31208 7964 31260 8016
rect 29552 7939 29604 7948
rect 29552 7905 29561 7939
rect 29561 7905 29595 7939
rect 29595 7905 29604 7939
rect 29552 7896 29604 7905
rect 29828 7939 29880 7948
rect 29828 7905 29837 7939
rect 29837 7905 29871 7939
rect 29871 7905 29880 7939
rect 29828 7896 29880 7905
rect 30564 7896 30616 7948
rect 3976 7760 4028 7812
rect 6920 7760 6972 7812
rect 7196 7760 7248 7812
rect 3792 7692 3844 7744
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 4620 7692 4672 7744
rect 4896 7692 4948 7744
rect 5264 7692 5316 7744
rect 6552 7692 6604 7744
rect 7656 7692 7708 7744
rect 8116 7692 8168 7744
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9312 7871 9364 7880
rect 9312 7837 9321 7871
rect 9321 7837 9355 7871
rect 9355 7837 9364 7871
rect 9312 7828 9364 7837
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 9588 7692 9640 7744
rect 11612 7692 11664 7744
rect 20812 7760 20864 7812
rect 22100 7803 22152 7812
rect 22100 7769 22109 7803
rect 22109 7769 22143 7803
rect 22143 7769 22152 7803
rect 22100 7760 22152 7769
rect 20628 7735 20680 7744
rect 20628 7701 20637 7735
rect 20637 7701 20671 7735
rect 20671 7701 20680 7735
rect 20628 7692 20680 7701
rect 24124 7760 24176 7812
rect 23480 7692 23532 7744
rect 31852 7896 31904 7948
rect 31944 7939 31996 7948
rect 31944 7905 31953 7939
rect 31953 7905 31987 7939
rect 31987 7905 31996 7939
rect 31944 7896 31996 7905
rect 32956 8032 33008 8084
rect 34796 8032 34848 8084
rect 35900 8032 35952 8084
rect 37832 8032 37884 8084
rect 32588 7896 32640 7948
rect 34980 7896 35032 7948
rect 35440 7896 35492 7948
rect 27344 7760 27396 7812
rect 29368 7760 29420 7812
rect 31576 7692 31628 7744
rect 32496 7803 32548 7812
rect 32496 7769 32505 7803
rect 32505 7769 32539 7803
rect 32539 7769 32548 7803
rect 32496 7760 32548 7769
rect 33232 7760 33284 7812
rect 33140 7692 33192 7744
rect 35900 7760 35952 7812
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 2320 7395 2372 7404
rect 2320 7361 2329 7395
rect 2329 7361 2363 7395
rect 2363 7361 2372 7395
rect 2320 7352 2372 7361
rect 2688 7352 2740 7404
rect 4160 7420 4212 7472
rect 3792 7395 3844 7404
rect 3792 7361 3801 7395
rect 3801 7361 3835 7395
rect 3835 7361 3844 7395
rect 3792 7352 3844 7361
rect 3976 7352 4028 7404
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 4528 7488 4580 7540
rect 4620 7463 4672 7472
rect 4620 7429 4629 7463
rect 4629 7429 4663 7463
rect 4663 7429 4672 7463
rect 4620 7420 4672 7429
rect 4528 7395 4580 7404
rect 4528 7361 4537 7395
rect 4537 7361 4571 7395
rect 4571 7361 4580 7395
rect 4528 7352 4580 7361
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 8208 7488 8260 7540
rect 19156 7488 19208 7540
rect 21824 7488 21876 7540
rect 22100 7488 22152 7540
rect 24400 7488 24452 7540
rect 24492 7488 24544 7540
rect 27344 7531 27396 7540
rect 7196 7420 7248 7472
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 3608 7284 3660 7293
rect 5632 7284 5684 7336
rect 4712 7216 4764 7268
rect 4528 7148 4580 7200
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 5264 7148 5316 7200
rect 8024 7352 8076 7404
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 7196 7284 7248 7336
rect 7380 7284 7432 7336
rect 8852 7420 8904 7472
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 11152 7463 11204 7472
rect 11152 7429 11161 7463
rect 11161 7429 11195 7463
rect 11195 7429 11204 7463
rect 11152 7420 11204 7429
rect 19800 7463 19852 7472
rect 19800 7429 19809 7463
rect 19809 7429 19843 7463
rect 19843 7429 19852 7463
rect 19800 7420 19852 7429
rect 19892 7463 19944 7472
rect 19892 7429 19901 7463
rect 19901 7429 19935 7463
rect 19935 7429 19944 7463
rect 19892 7420 19944 7429
rect 21272 7463 21324 7472
rect 21272 7429 21281 7463
rect 21281 7429 21315 7463
rect 21315 7429 21324 7463
rect 21272 7420 21324 7429
rect 21364 7463 21416 7472
rect 21364 7429 21373 7463
rect 21373 7429 21407 7463
rect 21407 7429 21416 7463
rect 21364 7420 21416 7429
rect 11612 7352 11664 7404
rect 12072 7352 12124 7404
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19708 7352 19760 7404
rect 20904 7352 20956 7404
rect 23204 7463 23256 7472
rect 23204 7429 23213 7463
rect 23213 7429 23247 7463
rect 23247 7429 23256 7463
rect 23204 7420 23256 7429
rect 24032 7420 24084 7472
rect 27344 7497 27353 7531
rect 27353 7497 27387 7531
rect 27387 7497 27396 7531
rect 27344 7488 27396 7497
rect 28632 7488 28684 7540
rect 29184 7488 29236 7540
rect 34060 7488 34112 7540
rect 35348 7531 35400 7540
rect 35348 7497 35357 7531
rect 35357 7497 35391 7531
rect 35391 7497 35400 7531
rect 35348 7488 35400 7497
rect 35440 7488 35492 7540
rect 25412 7463 25464 7472
rect 25412 7429 25421 7463
rect 25421 7429 25455 7463
rect 25455 7429 25464 7463
rect 25412 7420 25464 7429
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 12348 7284 12400 7336
rect 20628 7284 20680 7336
rect 23848 7352 23900 7404
rect 25688 7395 25740 7404
rect 25688 7361 25697 7395
rect 25697 7361 25731 7395
rect 25731 7361 25740 7395
rect 25688 7352 25740 7361
rect 33140 7420 33192 7472
rect 34704 7463 34756 7472
rect 34704 7429 34713 7463
rect 34713 7429 34747 7463
rect 34747 7429 34756 7463
rect 34704 7420 34756 7429
rect 36084 7420 36136 7472
rect 11060 7216 11112 7268
rect 11704 7216 11756 7268
rect 8668 7148 8720 7200
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 9220 7148 9272 7200
rect 11244 7191 11296 7200
rect 11244 7157 11253 7191
rect 11253 7157 11287 7191
rect 11287 7157 11296 7191
rect 11244 7148 11296 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 19708 7148 19760 7200
rect 29368 7352 29420 7404
rect 34980 7395 35032 7404
rect 34980 7361 34989 7395
rect 34989 7361 35023 7395
rect 35023 7361 35032 7395
rect 34980 7352 35032 7361
rect 28264 7327 28316 7336
rect 28264 7293 28273 7327
rect 28273 7293 28307 7327
rect 28307 7293 28316 7327
rect 28264 7284 28316 7293
rect 37740 7284 37792 7336
rect 32496 7148 32548 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4620 6944 4672 6996
rect 4896 6944 4948 6996
rect 9312 6944 9364 6996
rect 9864 6944 9916 6996
rect 12072 6944 12124 6996
rect 6092 6876 6144 6928
rect 7288 6876 7340 6928
rect 6000 6808 6052 6860
rect 9588 6808 9640 6860
rect 11704 6808 11756 6860
rect 6368 6740 6420 6792
rect 6828 6740 6880 6792
rect 2964 6604 3016 6656
rect 3516 6604 3568 6656
rect 6092 6672 6144 6724
rect 6552 6715 6604 6724
rect 6552 6681 6561 6715
rect 6561 6681 6595 6715
rect 6595 6681 6604 6715
rect 6552 6672 6604 6681
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 7104 6672 7156 6724
rect 9588 6715 9640 6724
rect 9588 6681 9597 6715
rect 9597 6681 9631 6715
rect 9631 6681 9640 6715
rect 9588 6672 9640 6681
rect 10232 6672 10284 6724
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 9680 6604 9732 6656
rect 9772 6604 9824 6656
rect 10600 6672 10652 6724
rect 11428 6672 11480 6724
rect 11612 6604 11664 6656
rect 12348 6604 12400 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 8300 6400 8352 6452
rect 9680 6400 9732 6452
rect 11888 6400 11940 6452
rect 12348 6400 12400 6452
rect 6828 6196 6880 6248
rect 9496 6196 9548 6248
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 10232 6332 10284 6384
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 12164 6332 12216 6384
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 11060 6264 11112 6316
rect 11244 6307 11296 6316
rect 11244 6273 11253 6307
rect 11253 6273 11287 6307
rect 11287 6273 11296 6307
rect 11244 6264 11296 6273
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12072 6264 12124 6316
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 9036 6128 9088 6180
rect 10048 6128 10100 6180
rect 9588 6060 9640 6112
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 10324 6171 10376 6180
rect 10324 6137 10333 6171
rect 10333 6137 10367 6171
rect 10367 6137 10376 6171
rect 10324 6128 10376 6137
rect 11612 6128 11664 6180
rect 12992 6128 13044 6180
rect 10876 6060 10928 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4436 5856 4488 5908
rect 5724 5856 5776 5908
rect 8944 5856 8996 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 9588 5856 9640 5908
rect 9864 5856 9916 5908
rect 10324 5856 10376 5908
rect 11244 5856 11296 5908
rect 12348 5899 12400 5908
rect 12348 5865 12357 5899
rect 12357 5865 12391 5899
rect 12391 5865 12400 5899
rect 12348 5856 12400 5865
rect 2320 5788 2372 5840
rect 5264 5788 5316 5840
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 2780 5652 2832 5704
rect 4344 5652 4396 5704
rect 4436 5627 4488 5636
rect 4436 5593 4445 5627
rect 4445 5593 4479 5627
rect 4479 5593 4488 5627
rect 4436 5584 4488 5593
rect 4896 5652 4948 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 4988 5627 5040 5636
rect 4988 5593 4997 5627
rect 4997 5593 5031 5627
rect 5031 5593 5040 5627
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 8852 5652 8904 5704
rect 9220 5720 9272 5772
rect 9496 5652 9548 5704
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 4988 5584 5040 5593
rect 9404 5584 9456 5636
rect 2964 5516 3016 5568
rect 4160 5516 4212 5568
rect 4252 5516 4304 5568
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 8668 5516 8720 5568
rect 10876 5627 10928 5636
rect 10876 5593 10885 5627
rect 10885 5593 10919 5627
rect 10919 5593 10928 5627
rect 10876 5584 10928 5593
rect 11428 5584 11480 5636
rect 11520 5516 11572 5568
rect 11796 5516 11848 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 4344 5312 4396 5364
rect 9404 5312 9456 5364
rect 9864 5312 9916 5364
rect 9956 5312 10008 5364
rect 3516 5244 3568 5296
rect 3884 5244 3936 5296
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 6000 5287 6052 5296
rect 6000 5253 6009 5287
rect 6009 5253 6043 5287
rect 6043 5253 6052 5287
rect 6000 5244 6052 5253
rect 6552 5244 6604 5296
rect 7288 5244 7340 5296
rect 8852 5244 8904 5296
rect 1400 5108 1452 5160
rect 2136 5108 2188 5160
rect 2780 5108 2832 5160
rect 4344 5151 4396 5160
rect 4344 5117 4353 5151
rect 4353 5117 4387 5151
rect 4387 5117 4396 5151
rect 4344 5108 4396 5117
rect 4712 5108 4764 5160
rect 9128 5176 9180 5228
rect 9588 5176 9640 5228
rect 9772 5176 9824 5228
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 5540 5108 5592 5160
rect 10048 5176 10100 5228
rect 11980 5244 12032 5296
rect 4620 5040 4672 5092
rect 3792 4972 3844 5024
rect 4252 4972 4304 5024
rect 4436 4972 4488 5024
rect 4896 4972 4948 5024
rect 5356 4972 5408 5024
rect 6828 4972 6880 5024
rect 7380 4972 7432 5024
rect 9220 4972 9272 5024
rect 9312 4972 9364 5024
rect 9864 5015 9916 5024
rect 9864 4981 9873 5015
rect 9873 4981 9907 5015
rect 9907 4981 9916 5015
rect 9864 4972 9916 4981
rect 10232 5015 10284 5024
rect 10232 4981 10241 5015
rect 10241 4981 10275 5015
rect 10275 4981 10284 5015
rect 10232 4972 10284 4981
rect 10784 4972 10836 5024
rect 12440 4972 12492 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 2412 4768 2464 4820
rect 3516 4768 3568 4820
rect 4068 4768 4120 4820
rect 5448 4768 5500 4820
rect 7012 4811 7064 4820
rect 7012 4777 7021 4811
rect 7021 4777 7055 4811
rect 7055 4777 7064 4811
rect 7012 4768 7064 4777
rect 7472 4768 7524 4820
rect 4712 4700 4764 4752
rect 5908 4700 5960 4752
rect 7288 4743 7340 4752
rect 7288 4709 7297 4743
rect 7297 4709 7331 4743
rect 7331 4709 7340 4743
rect 7288 4700 7340 4709
rect 8300 4700 8352 4752
rect 9404 4768 9456 4820
rect 10048 4768 10100 4820
rect 10784 4700 10836 4752
rect 3884 4632 3936 4684
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4252 4564 4304 4616
rect 4896 4632 4948 4684
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 5264 4564 5316 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 7380 4564 7432 4616
rect 8852 4632 8904 4684
rect 2412 4496 2464 4548
rect 2964 4496 3016 4548
rect 2688 4428 2740 4480
rect 4436 4496 4488 4548
rect 7472 4539 7524 4548
rect 7472 4505 7481 4539
rect 7481 4505 7515 4539
rect 7515 4505 7524 4539
rect 7472 4496 7524 4505
rect 9404 4564 9456 4616
rect 9680 4564 9732 4616
rect 10416 4632 10468 4684
rect 10600 4632 10652 4684
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 8852 4496 8904 4548
rect 9220 4496 9272 4548
rect 9588 4496 9640 4548
rect 10508 4564 10560 4616
rect 12440 4564 12492 4616
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 4804 4428 4856 4480
rect 8576 4428 8628 4480
rect 11336 4496 11388 4548
rect 11152 4428 11204 4480
rect 11796 4539 11848 4548
rect 11796 4505 11805 4539
rect 11805 4505 11839 4539
rect 11839 4505 11848 4539
rect 11796 4496 11848 4505
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4620 4224 4672 4276
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 9128 4224 9180 4276
rect 9864 4224 9916 4276
rect 4712 4156 4764 4208
rect 5264 4156 5316 4208
rect 9588 4156 9640 4208
rect 10324 4224 10376 4276
rect 11336 4224 11388 4276
rect 4344 4088 4396 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 3516 3952 3568 4004
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 4712 4063 4764 4072
rect 4712 4029 4721 4063
rect 4721 4029 4755 4063
rect 4755 4029 4764 4063
rect 4712 4020 4764 4029
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 4896 4020 4948 4072
rect 3240 3884 3292 3936
rect 4528 3884 4580 3936
rect 5448 3952 5500 4004
rect 8300 4088 8352 4140
rect 8576 4088 8628 4140
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 10508 4156 10560 4208
rect 7932 3952 7984 4004
rect 5356 3884 5408 3936
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 9404 4020 9456 4072
rect 9956 3952 10008 4004
rect 11244 3952 11296 4004
rect 10508 3884 10560 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2228 3680 2280 3732
rect 4712 3680 4764 3732
rect 4896 3680 4948 3732
rect 5264 3680 5316 3732
rect 3148 3544 3200 3596
rect 3884 3587 3936 3596
rect 3884 3553 3893 3587
rect 3893 3553 3927 3587
rect 3927 3553 3936 3587
rect 3884 3544 3936 3553
rect 5540 3544 5592 3596
rect 3240 3519 3292 3528
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 5448 3476 5500 3528
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 11796 3612 11848 3664
rect 9496 3544 9548 3596
rect 4160 3451 4212 3460
rect 4160 3417 4169 3451
rect 4169 3417 4203 3451
rect 4203 3417 4212 3451
rect 4160 3408 4212 3417
rect 5908 3408 5960 3460
rect 8668 3476 8720 3528
rect 10140 3476 10192 3528
rect 10232 3519 10284 3528
rect 10232 3485 10241 3519
rect 10241 3485 10275 3519
rect 10275 3485 10284 3519
rect 10232 3476 10284 3485
rect 10508 3519 10560 3528
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 11520 3476 11572 3528
rect 42156 3519 42208 3528
rect 42156 3485 42165 3519
rect 42165 3485 42199 3519
rect 42199 3485 42208 3519
rect 42156 3476 42208 3485
rect 3424 3340 3476 3392
rect 4528 3340 4580 3392
rect 6920 3408 6972 3460
rect 8852 3408 8904 3460
rect 9772 3340 9824 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4160 3136 4212 3188
rect 3424 3111 3476 3120
rect 3424 3077 3433 3111
rect 3433 3077 3467 3111
rect 3467 3077 3476 3111
rect 3424 3068 3476 3077
rect 5908 3136 5960 3188
rect 9404 3179 9456 3188
rect 9404 3145 9413 3179
rect 9413 3145 9447 3179
rect 9447 3145 9456 3179
rect 9404 3136 9456 3145
rect 5264 3111 5316 3120
rect 5264 3077 5273 3111
rect 5273 3077 5307 3111
rect 5307 3077 5316 3111
rect 5264 3068 5316 3077
rect 5356 3111 5408 3120
rect 5356 3077 5365 3111
rect 5365 3077 5399 3111
rect 5399 3077 5408 3111
rect 5356 3068 5408 3077
rect 7932 3111 7984 3120
rect 7932 3077 7941 3111
rect 7941 3077 7975 3111
rect 7975 3077 7984 3111
rect 7932 3068 7984 3077
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 4712 3000 4764 3052
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 6828 3000 6880 3052
rect 10600 3136 10652 3188
rect 9772 3111 9824 3120
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 10324 3068 10376 3120
rect 4804 2932 4856 2984
rect 10140 2932 10192 2984
rect 10324 2796 10376 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8760 2388 8812 2440
rect 11612 2252 11664 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 17406 45098 17462 45787
rect 19338 45098 19394 45787
rect 19982 45098 20038 45787
rect 20626 45098 20682 45787
rect 17406 45070 17724 45098
rect 17406 44987 17462 45070
rect 4874 43548 5182 43557
rect 4874 43546 4880 43548
rect 4936 43546 4960 43548
rect 5016 43546 5040 43548
rect 5096 43546 5120 43548
rect 5176 43546 5182 43548
rect 4936 43494 4938 43546
rect 5118 43494 5120 43546
rect 4874 43492 4880 43494
rect 4936 43492 4960 43494
rect 5016 43492 5040 43494
rect 5096 43492 5120 43494
rect 5176 43492 5182 43494
rect 4874 43483 5182 43492
rect 17696 43450 17724 45070
rect 19338 45070 19564 45098
rect 19338 44987 19394 45070
rect 19536 43450 19564 45070
rect 19982 45070 20300 45098
rect 19982 44987 20038 45070
rect 20272 43450 20300 45070
rect 20548 45070 20682 45098
rect 20548 43450 20576 45070
rect 20626 44987 20682 45070
rect 22558 45098 22614 45787
rect 23202 45098 23258 45787
rect 25134 45098 25190 45787
rect 28998 45098 29054 45787
rect 22558 45070 22876 45098
rect 22558 44987 22614 45070
rect 22848 43450 22876 45070
rect 23202 45070 23428 45098
rect 23202 44987 23258 45070
rect 23400 43450 23428 45070
rect 25134 45070 25360 45098
rect 25134 44987 25190 45070
rect 25332 43450 25360 45070
rect 28998 45070 29224 45098
rect 28998 44987 29054 45070
rect 29196 43450 29224 45070
rect 35594 43548 35902 43557
rect 35594 43546 35600 43548
rect 35656 43546 35680 43548
rect 35736 43546 35760 43548
rect 35816 43546 35840 43548
rect 35896 43546 35902 43548
rect 35656 43494 35658 43546
rect 35838 43494 35840 43546
rect 35594 43492 35600 43494
rect 35656 43492 35680 43494
rect 35736 43492 35760 43494
rect 35816 43492 35840 43494
rect 35896 43492 35902 43494
rect 35594 43483 35902 43492
rect 17684 43444 17736 43450
rect 17684 43386 17736 43392
rect 19524 43444 19576 43450
rect 19524 43386 19576 43392
rect 20260 43444 20312 43450
rect 20260 43386 20312 43392
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 22836 43444 22888 43450
rect 22836 43386 22888 43392
rect 23388 43444 23440 43450
rect 23388 43386 23440 43392
rect 25320 43444 25372 43450
rect 25320 43386 25372 43392
rect 29184 43444 29236 43450
rect 29184 43386 29236 43392
rect 24400 43376 24452 43382
rect 24400 43318 24452 43324
rect 28448 43376 28500 43382
rect 28448 43318 28500 43324
rect 17500 43308 17552 43314
rect 17500 43250 17552 43256
rect 19800 43308 19852 43314
rect 19800 43250 19852 43256
rect 20996 43308 21048 43314
rect 20996 43250 21048 43256
rect 22744 43308 22796 43314
rect 22744 43250 22796 43256
rect 23020 43308 23072 43314
rect 23020 43250 23072 43256
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 17512 42906 17540 43250
rect 19340 43240 19392 43246
rect 19340 43182 19392 43188
rect 17500 42900 17552 42906
rect 17500 42842 17552 42848
rect 15660 42696 15712 42702
rect 15660 42638 15712 42644
rect 4874 42460 5182 42469
rect 4874 42458 4880 42460
rect 4936 42458 4960 42460
rect 5016 42458 5040 42460
rect 5096 42458 5120 42460
rect 5176 42458 5182 42460
rect 4936 42406 4938 42458
rect 5118 42406 5120 42458
rect 4874 42404 4880 42406
rect 4936 42404 4960 42406
rect 5016 42404 5040 42406
rect 5096 42404 5120 42406
rect 5176 42404 5182 42406
rect 4874 42395 5182 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 15672 41682 15700 42638
rect 16212 42628 16264 42634
rect 16212 42570 16264 42576
rect 16396 42628 16448 42634
rect 16396 42570 16448 42576
rect 16224 42226 16252 42570
rect 15936 42220 15988 42226
rect 15936 42162 15988 42168
rect 16212 42220 16264 42226
rect 16212 42162 16264 42168
rect 15660 41676 15712 41682
rect 15660 41618 15712 41624
rect 1306 41576 1362 41585
rect 1306 41511 1362 41520
rect 15384 41540 15436 41546
rect 1320 40730 1348 41511
rect 15384 41482 15436 41488
rect 4874 41372 5182 41381
rect 4874 41370 4880 41372
rect 4936 41370 4960 41372
rect 5016 41370 5040 41372
rect 5096 41370 5120 41372
rect 5176 41370 5182 41372
rect 4936 41318 4938 41370
rect 5118 41318 5120 41370
rect 4874 41316 4880 41318
rect 4936 41316 4960 41318
rect 5016 41316 5040 41318
rect 5096 41316 5120 41318
rect 5176 41316 5182 41318
rect 4874 41307 5182 41316
rect 15396 41274 15424 41482
rect 15384 41268 15436 41274
rect 15384 41210 15436 41216
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 1308 40724 1360 40730
rect 1308 40666 1360 40672
rect 4874 40284 5182 40293
rect 4874 40282 4880 40284
rect 4936 40282 4960 40284
rect 5016 40282 5040 40284
rect 5096 40282 5120 40284
rect 5176 40282 5182 40284
rect 4936 40230 4938 40282
rect 5118 40230 5120 40282
rect 4874 40228 4880 40230
rect 4936 40228 4960 40230
rect 5016 40228 5040 40230
rect 5096 40228 5120 40230
rect 5176 40228 5182 40230
rect 4874 40219 5182 40228
rect 14556 40044 14608 40050
rect 14556 39986 14608 39992
rect 12900 39976 12952 39982
rect 12900 39918 12952 39924
rect 13544 39976 13596 39982
rect 13544 39918 13596 39924
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 3608 38956 3660 38962
rect 3608 38898 3660 38904
rect 3240 38752 3292 38758
rect 3240 38694 3292 38700
rect 1400 38412 1452 38418
rect 1400 38354 1452 38360
rect 1412 37330 1440 38354
rect 1952 38276 2004 38282
rect 1952 38218 2004 38224
rect 2964 38276 3016 38282
rect 2964 38218 3016 38224
rect 1964 38010 1992 38218
rect 2596 38208 2648 38214
rect 2596 38150 2648 38156
rect 1952 38004 2004 38010
rect 1952 37946 2004 37952
rect 2608 37874 2636 38150
rect 1860 37868 1912 37874
rect 1860 37810 1912 37816
rect 2044 37868 2096 37874
rect 2044 37810 2096 37816
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 1872 37466 1900 37810
rect 1860 37460 1912 37466
rect 1860 37402 1912 37408
rect 2056 37330 2084 37810
rect 2872 37664 2924 37670
rect 2872 37606 2924 37612
rect 1400 37324 1452 37330
rect 1400 37266 1452 37272
rect 2044 37324 2096 37330
rect 2044 37266 2096 37272
rect 1412 35630 1440 37266
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 1676 37188 1728 37194
rect 1676 37130 1728 37136
rect 1688 36922 1716 37130
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 2792 35698 2820 37198
rect 2884 36922 2912 37606
rect 2976 37262 3004 38218
rect 3148 37664 3200 37670
rect 3148 37606 3200 37612
rect 2964 37256 3016 37262
rect 2964 37198 3016 37204
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 3160 36786 3188 37606
rect 2872 36780 2924 36786
rect 2872 36722 2924 36728
rect 3148 36780 3200 36786
rect 3148 36722 3200 36728
rect 2884 36174 2912 36722
rect 3252 36718 3280 38694
rect 3424 38344 3476 38350
rect 3424 38286 3476 38292
rect 3436 38214 3464 38286
rect 3424 38208 3476 38214
rect 3424 38150 3476 38156
rect 3516 38208 3568 38214
rect 3516 38150 3568 38156
rect 3332 37800 3384 37806
rect 3332 37742 3384 37748
rect 3344 36718 3372 37742
rect 3436 37466 3464 38150
rect 3528 37874 3556 38150
rect 3516 37868 3568 37874
rect 3516 37810 3568 37816
rect 3424 37460 3476 37466
rect 3424 37402 3476 37408
rect 3516 36780 3568 36786
rect 3516 36722 3568 36728
rect 3240 36712 3292 36718
rect 3240 36654 3292 36660
rect 3332 36712 3384 36718
rect 3332 36654 3384 36660
rect 2872 36168 2924 36174
rect 2872 36110 2924 36116
rect 2964 36168 3016 36174
rect 2964 36110 3016 36116
rect 2872 36032 2924 36038
rect 2872 35974 2924 35980
rect 2780 35692 2832 35698
rect 2780 35634 2832 35640
rect 1400 35624 1452 35630
rect 1400 35566 1452 35572
rect 1412 35154 1440 35566
rect 2136 35488 2188 35494
rect 2136 35430 2188 35436
rect 2148 35154 2176 35430
rect 1400 35148 1452 35154
rect 1400 35090 1452 35096
rect 2136 35148 2188 35154
rect 2136 35090 2188 35096
rect 2688 35148 2740 35154
rect 2688 35090 2740 35096
rect 2700 33658 2728 35090
rect 1676 33652 1728 33658
rect 1676 33594 1728 33600
rect 2688 33652 2740 33658
rect 2688 33594 2740 33600
rect 1688 32978 1716 33594
rect 2792 33522 2820 35634
rect 2884 35630 2912 35974
rect 2872 35624 2924 35630
rect 2872 35566 2924 35572
rect 2976 34746 3004 36110
rect 3528 36106 3556 36722
rect 3516 36100 3568 36106
rect 3516 36042 3568 36048
rect 3528 35630 3556 36042
rect 3620 35834 3648 38898
rect 12912 38894 12940 39918
rect 13556 39642 13584 39918
rect 13544 39636 13596 39642
rect 13544 39578 13596 39584
rect 14004 39296 14056 39302
rect 14004 39238 14056 39244
rect 12900 38888 12952 38894
rect 12900 38830 12952 38836
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 7288 38548 7340 38554
rect 7340 38508 7420 38536
rect 7288 38490 7340 38496
rect 3792 38412 3844 38418
rect 3792 38354 3844 38360
rect 5264 38412 5316 38418
rect 5264 38354 5316 38360
rect 7104 38412 7156 38418
rect 7104 38354 7156 38360
rect 3804 37806 3832 38354
rect 4712 38208 4764 38214
rect 4712 38150 4764 38156
rect 4804 38208 4856 38214
rect 4804 38150 4856 38156
rect 3700 37800 3752 37806
rect 3700 37742 3752 37748
rect 3792 37800 3844 37806
rect 3792 37742 3844 37748
rect 4620 37800 4672 37806
rect 4620 37742 4672 37748
rect 3712 37398 3740 37742
rect 3700 37392 3752 37398
rect 3700 37334 3752 37340
rect 3804 37330 3832 37742
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4068 37392 4120 37398
rect 4068 37334 4120 37340
rect 4160 37392 4212 37398
rect 4160 37334 4212 37340
rect 3792 37324 3844 37330
rect 3792 37266 3844 37272
rect 3804 36854 3832 37266
rect 3792 36848 3844 36854
rect 3792 36790 3844 36796
rect 4080 36582 4108 37334
rect 4172 37126 4200 37334
rect 4160 37120 4212 37126
rect 4160 37062 4212 37068
rect 4436 37120 4488 37126
rect 4436 37062 4488 37068
rect 4448 36786 4476 37062
rect 4632 36922 4660 37742
rect 4620 36916 4672 36922
rect 4620 36858 4672 36864
rect 4436 36780 4488 36786
rect 4436 36722 4488 36728
rect 4528 36780 4580 36786
rect 4724 36768 4752 38150
rect 4816 37670 4844 38150
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 5172 37732 5224 37738
rect 5172 37674 5224 37680
rect 4804 37664 4856 37670
rect 4804 37606 4856 37612
rect 4816 37194 4844 37606
rect 5184 37398 5212 37674
rect 5172 37392 5224 37398
rect 5172 37334 5224 37340
rect 5184 37262 5212 37334
rect 5172 37256 5224 37262
rect 5172 37198 5224 37204
rect 4804 37188 4856 37194
rect 4804 37130 4856 37136
rect 4580 36740 4752 36768
rect 4528 36722 4580 36728
rect 4344 36712 4396 36718
rect 4342 36680 4344 36689
rect 4396 36680 4398 36689
rect 4342 36615 4398 36624
rect 4710 36680 4766 36689
rect 4816 36650 4844 37130
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 5172 36916 5224 36922
rect 5276 36904 5304 38354
rect 6092 38344 6144 38350
rect 6092 38286 6144 38292
rect 6828 38344 6880 38350
rect 6828 38286 6880 38292
rect 5448 38276 5500 38282
rect 5448 38218 5500 38224
rect 5460 37738 5488 38218
rect 5908 38208 5960 38214
rect 5908 38150 5960 38156
rect 5816 38004 5868 38010
rect 5816 37946 5868 37952
rect 5540 37868 5592 37874
rect 5540 37810 5592 37816
rect 5448 37732 5500 37738
rect 5448 37674 5500 37680
rect 5552 37126 5580 37810
rect 5356 37120 5408 37126
rect 5356 37062 5408 37068
rect 5540 37120 5592 37126
rect 5540 37062 5592 37068
rect 5368 36922 5396 37062
rect 5224 36876 5304 36904
rect 5356 36916 5408 36922
rect 5172 36858 5224 36864
rect 5356 36858 5408 36864
rect 4988 36780 5040 36786
rect 4988 36722 5040 36728
rect 4710 36615 4766 36624
rect 4804 36644 4856 36650
rect 4068 36576 4120 36582
rect 4068 36518 4120 36524
rect 3976 36304 4028 36310
rect 3804 36252 3976 36258
rect 3804 36246 4028 36252
rect 3804 36242 4016 36246
rect 3792 36236 4016 36242
rect 3844 36230 4016 36236
rect 3792 36178 3844 36184
rect 3884 36168 3936 36174
rect 3884 36110 3936 36116
rect 3700 36100 3752 36106
rect 3700 36042 3752 36048
rect 3608 35828 3660 35834
rect 3608 35770 3660 35776
rect 3424 35624 3476 35630
rect 3424 35566 3476 35572
rect 3516 35624 3568 35630
rect 3516 35566 3568 35572
rect 2964 34740 3016 34746
rect 2964 34682 3016 34688
rect 2780 33516 2832 33522
rect 2780 33458 2832 33464
rect 2136 33448 2188 33454
rect 2136 33390 2188 33396
rect 1676 32972 1728 32978
rect 1676 32914 1728 32920
rect 2148 32570 2176 33390
rect 2792 32858 2820 33458
rect 3148 33312 3200 33318
rect 3148 33254 3200 33260
rect 3240 33312 3292 33318
rect 3240 33254 3292 33260
rect 2792 32842 3004 32858
rect 2792 32836 3016 32842
rect 2792 32830 2964 32836
rect 2964 32778 3016 32784
rect 2136 32564 2188 32570
rect 2136 32506 2188 32512
rect 2596 32496 2648 32502
rect 2596 32438 2648 32444
rect 2608 31482 2636 32438
rect 3056 32360 3108 32366
rect 3056 32302 3108 32308
rect 3160 32314 3188 33254
rect 3252 32434 3280 33254
rect 3332 32768 3384 32774
rect 3332 32710 3384 32716
rect 3344 32570 3372 32710
rect 3332 32564 3384 32570
rect 3332 32506 3384 32512
rect 3240 32428 3292 32434
rect 3240 32370 3292 32376
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 3344 32314 3372 32370
rect 3068 32026 3096 32302
rect 3160 32286 3372 32314
rect 3056 32020 3108 32026
rect 3056 31962 3108 31968
rect 2596 31476 2648 31482
rect 2596 31418 2648 31424
rect 2872 31408 2924 31414
rect 2872 31350 2924 31356
rect 1676 31136 1728 31142
rect 1676 31078 1728 31084
rect 1688 30666 1716 31078
rect 1676 30660 1728 30666
rect 1676 30602 1728 30608
rect 2884 30326 2912 31350
rect 3240 31340 3292 31346
rect 3240 31282 3292 31288
rect 3148 31272 3200 31278
rect 3148 31214 3200 31220
rect 3056 31204 3108 31210
rect 3056 31146 3108 31152
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 2872 30320 2924 30326
rect 2872 30262 2924 30268
rect 2976 30258 3004 31078
rect 3068 30666 3096 31146
rect 3160 30938 3188 31214
rect 3252 30938 3280 31282
rect 3344 31142 3372 32286
rect 3436 31822 3464 35566
rect 3620 35086 3648 35770
rect 3712 35698 3740 36042
rect 3896 35698 3924 36110
rect 3700 35692 3752 35698
rect 3700 35634 3752 35640
rect 3884 35692 3936 35698
rect 3884 35634 3936 35640
rect 3608 35080 3660 35086
rect 3608 35022 3660 35028
rect 3620 34610 3648 35022
rect 3712 35018 3740 35634
rect 3896 35290 3924 35634
rect 3988 35494 4016 36230
rect 4080 36174 4108 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 36168 4120 36174
rect 4068 36110 4120 36116
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 4080 35494 4108 35974
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 3976 35488 4028 35494
rect 3976 35430 4028 35436
rect 4068 35488 4120 35494
rect 4068 35430 4120 35436
rect 3884 35284 3936 35290
rect 3884 35226 3936 35232
rect 3896 35086 3924 35226
rect 3884 35080 3936 35086
rect 3884 35022 3936 35028
rect 3988 35018 4016 35430
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4342 35048 4398 35057
rect 3700 35012 3752 35018
rect 3700 34954 3752 34960
rect 3976 35012 4028 35018
rect 4342 34983 4344 34992
rect 3976 34954 4028 34960
rect 4396 34983 4398 34992
rect 4344 34954 4396 34960
rect 3988 34678 4016 34954
rect 4068 34944 4120 34950
rect 4068 34886 4120 34892
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 4080 34610 4108 34886
rect 4632 34746 4660 35634
rect 4724 35034 4752 36615
rect 4804 36586 4856 36592
rect 5000 36378 5028 36722
rect 4988 36372 5040 36378
rect 4988 36314 5040 36320
rect 5184 36174 5212 36858
rect 5632 36576 5684 36582
rect 5632 36518 5684 36524
rect 5448 36372 5500 36378
rect 5448 36314 5500 36320
rect 5172 36168 5224 36174
rect 5172 36110 5224 36116
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5264 35692 5316 35698
rect 5264 35634 5316 35640
rect 4896 35624 4948 35630
rect 4894 35592 4896 35601
rect 4948 35592 4950 35601
rect 4894 35527 4950 35536
rect 5276 35290 5304 35634
rect 5264 35284 5316 35290
rect 5264 35226 5316 35232
rect 4724 35006 4844 35034
rect 4712 34944 4764 34950
rect 4712 34886 4764 34892
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 4724 34610 4752 34886
rect 3608 34604 3660 34610
rect 3608 34546 3660 34552
rect 4068 34604 4120 34610
rect 4068 34546 4120 34552
rect 4712 34604 4764 34610
rect 4712 34546 4764 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4816 33658 4844 35006
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 5172 34604 5224 34610
rect 5172 34546 5224 34552
rect 5184 34513 5212 34546
rect 5170 34504 5226 34513
rect 5170 34439 5226 34448
rect 5276 34202 5304 34886
rect 5264 34196 5316 34202
rect 5264 34138 5316 34144
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 3516 33652 3568 33658
rect 3516 33594 3568 33600
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 3528 33454 3556 33594
rect 3608 33584 3660 33590
rect 3608 33526 3660 33532
rect 3620 33454 3648 33526
rect 4068 33516 4120 33522
rect 4068 33458 4120 33464
rect 4804 33516 4856 33522
rect 4804 33458 4856 33464
rect 3516 33448 3568 33454
rect 3516 33390 3568 33396
rect 3608 33448 3660 33454
rect 3608 33390 3660 33396
rect 3528 32978 3556 33390
rect 3516 32972 3568 32978
rect 3516 32914 3568 32920
rect 3620 32910 3648 33390
rect 3792 33312 3844 33318
rect 3792 33254 3844 33260
rect 3608 32904 3660 32910
rect 3608 32846 3660 32852
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3608 32768 3660 32774
rect 3608 32710 3660 32716
rect 3424 31816 3476 31822
rect 3424 31758 3476 31764
rect 3332 31136 3384 31142
rect 3332 31078 3384 31084
rect 3148 30932 3200 30938
rect 3148 30874 3200 30880
rect 3240 30932 3292 30938
rect 3240 30874 3292 30880
rect 3056 30660 3108 30666
rect 3056 30602 3108 30608
rect 2964 30252 3016 30258
rect 2964 30194 3016 30200
rect 2686 30152 2742 30161
rect 2686 30087 2742 30096
rect 2700 29646 2728 30087
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 2688 29640 2740 29646
rect 2872 29640 2924 29646
rect 2688 29582 2740 29588
rect 2870 29608 2872 29617
rect 2924 29608 2926 29617
rect 1676 29096 1728 29102
rect 1676 29038 1728 29044
rect 1688 28762 1716 29038
rect 1676 28756 1728 28762
rect 1676 28698 1728 28704
rect 1780 26994 1808 29582
rect 2870 29543 2926 29552
rect 2964 29504 3016 29510
rect 2964 29446 3016 29452
rect 2976 28558 3004 29446
rect 3068 29238 3096 30602
rect 3160 30598 3188 30874
rect 3148 30592 3200 30598
rect 3148 30534 3200 30540
rect 3160 30394 3188 30534
rect 3148 30388 3200 30394
rect 3148 30330 3200 30336
rect 3240 30388 3292 30394
rect 3240 30330 3292 30336
rect 3252 29646 3280 30330
rect 3330 30288 3386 30297
rect 3330 30223 3332 30232
rect 3384 30223 3386 30232
rect 3332 30194 3384 30200
rect 3436 29850 3464 31758
rect 3528 31414 3556 32710
rect 3620 32434 3648 32710
rect 3804 32434 3832 33254
rect 4080 32910 4108 33458
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 3608 32428 3660 32434
rect 3608 32370 3660 32376
rect 3792 32428 3844 32434
rect 3792 32370 3844 32376
rect 3804 32230 3832 32370
rect 3792 32224 3844 32230
rect 3792 32166 3844 32172
rect 3976 31680 4028 31686
rect 3976 31622 4028 31628
rect 3608 31476 3660 31482
rect 3608 31418 3660 31424
rect 3516 31408 3568 31414
rect 3516 31350 3568 31356
rect 3516 30932 3568 30938
rect 3516 30874 3568 30880
rect 3528 30734 3556 30874
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3620 30104 3648 31418
rect 3792 30864 3844 30870
rect 3792 30806 3844 30812
rect 3804 30326 3832 30806
rect 3792 30320 3844 30326
rect 3988 30308 4016 31622
rect 4080 31482 4108 32846
rect 4712 32836 4764 32842
rect 4712 32778 4764 32784
rect 4724 32416 4752 32778
rect 4816 32774 4844 33458
rect 5368 33046 5396 35974
rect 5460 35698 5488 36314
rect 5644 35834 5672 36518
rect 5632 35828 5684 35834
rect 5632 35770 5684 35776
rect 5448 35692 5500 35698
rect 5448 35634 5500 35640
rect 5632 35624 5684 35630
rect 5630 35592 5632 35601
rect 5684 35592 5686 35601
rect 5448 35556 5500 35562
rect 5630 35527 5686 35536
rect 5448 35498 5500 35504
rect 5460 33522 5488 35498
rect 5540 34740 5592 34746
rect 5540 34682 5592 34688
rect 5552 33998 5580 34682
rect 5632 34672 5684 34678
rect 5632 34614 5684 34620
rect 5540 33992 5592 33998
rect 5540 33934 5592 33940
rect 5644 33522 5672 34614
rect 5828 34066 5856 37946
rect 5920 37466 5948 38150
rect 6104 38010 6132 38286
rect 6460 38276 6512 38282
rect 6460 38218 6512 38224
rect 6092 38004 6144 38010
rect 6092 37946 6144 37952
rect 6472 37942 6500 38218
rect 6460 37936 6512 37942
rect 6460 37878 6512 37884
rect 6644 37800 6696 37806
rect 6564 37748 6644 37754
rect 6564 37742 6696 37748
rect 6564 37726 6684 37742
rect 5908 37460 5960 37466
rect 5908 37402 5960 37408
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 6092 36236 6144 36242
rect 6092 36178 6144 36184
rect 6104 35834 6132 36178
rect 6380 36106 6408 37062
rect 6564 36786 6592 37726
rect 6840 37330 6868 38286
rect 7012 38276 7064 38282
rect 7012 38218 7064 38224
rect 7024 38010 7052 38218
rect 7012 38004 7064 38010
rect 7012 37946 7064 37952
rect 6920 37868 6972 37874
rect 6920 37810 6972 37816
rect 6828 37324 6880 37330
rect 6828 37266 6880 37272
rect 6932 37194 6960 37810
rect 7012 37800 7064 37806
rect 7012 37742 7064 37748
rect 7024 37466 7052 37742
rect 7012 37460 7064 37466
rect 7012 37402 7064 37408
rect 7116 37262 7144 38354
rect 7392 37874 7420 38508
rect 8300 38412 8352 38418
rect 8300 38354 8352 38360
rect 7932 38208 7984 38214
rect 7932 38150 7984 38156
rect 7472 38004 7524 38010
rect 7472 37946 7524 37952
rect 7484 37874 7512 37946
rect 7288 37868 7340 37874
rect 7288 37810 7340 37816
rect 7380 37868 7432 37874
rect 7380 37810 7432 37816
rect 7472 37868 7524 37874
rect 7524 37828 7604 37856
rect 7472 37810 7524 37816
rect 7300 37466 7328 37810
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7104 37256 7156 37262
rect 7104 37198 7156 37204
rect 6920 37188 6972 37194
rect 6920 37130 6972 37136
rect 6932 36922 6960 37130
rect 6920 36916 6972 36922
rect 6920 36858 6972 36864
rect 6644 36848 6696 36854
rect 6644 36790 6696 36796
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 6564 36310 6592 36722
rect 6552 36304 6604 36310
rect 6552 36246 6604 36252
rect 6368 36100 6420 36106
rect 6368 36042 6420 36048
rect 6092 35828 6144 35834
rect 6092 35770 6144 35776
rect 5908 35692 5960 35698
rect 5908 35634 5960 35640
rect 5920 35057 5948 35634
rect 6276 35624 6328 35630
rect 6276 35566 6328 35572
rect 5906 35048 5962 35057
rect 5906 34983 5962 34992
rect 6184 34672 6236 34678
rect 6184 34614 6236 34620
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 5908 34400 5960 34406
rect 5908 34342 5960 34348
rect 5920 34066 5948 34342
rect 5724 34060 5776 34066
rect 5724 34002 5776 34008
rect 5816 34060 5868 34066
rect 5816 34002 5868 34008
rect 5908 34060 5960 34066
rect 5908 34002 5960 34008
rect 5736 33658 5764 34002
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 5448 33516 5500 33522
rect 5448 33458 5500 33464
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5356 33040 5408 33046
rect 5356 32982 5408 32988
rect 5356 32904 5408 32910
rect 5356 32846 5408 32852
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 5264 32768 5316 32774
rect 5264 32710 5316 32716
rect 4816 32552 4844 32710
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4816 32524 5120 32552
rect 4724 32388 4844 32416
rect 4620 32360 4672 32366
rect 4672 32308 4752 32314
rect 4620 32302 4752 32308
rect 4632 32286 4752 32302
rect 4620 32224 4672 32230
rect 4620 32166 4672 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 4632 31278 4660 32166
rect 4724 32026 4752 32286
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 4816 31890 4844 32388
rect 5092 32230 5120 32524
rect 5080 32224 5132 32230
rect 5080 32166 5132 32172
rect 4804 31884 4856 31890
rect 4804 31826 4856 31832
rect 4620 31272 4672 31278
rect 4620 31214 4672 31220
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30734 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30802 4660 31214
rect 4816 30938 4844 31826
rect 5276 31822 5304 32710
rect 5368 32026 5396 32846
rect 5356 32020 5408 32026
rect 5356 31962 5408 31968
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5356 31748 5408 31754
rect 5356 31690 5408 31696
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 5368 31482 5396 31690
rect 5172 31476 5224 31482
rect 5172 31418 5224 31424
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 4896 31204 4948 31210
rect 4896 31146 4948 31152
rect 4804 30932 4856 30938
rect 4804 30874 4856 30880
rect 4908 30802 4936 31146
rect 5184 30802 5212 31418
rect 5460 31362 5488 33458
rect 5632 32904 5684 32910
rect 5828 32892 5856 34002
rect 6104 33862 6132 34546
rect 6092 33856 6144 33862
rect 6092 33798 6144 33804
rect 5684 32864 5856 32892
rect 5632 32846 5684 32852
rect 5540 32768 5592 32774
rect 5540 32710 5592 32716
rect 5368 31334 5488 31362
rect 4620 30796 4672 30802
rect 4620 30738 4672 30744
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 5172 30796 5224 30802
rect 5172 30738 5224 30744
rect 4068 30728 4120 30734
rect 4068 30670 4120 30676
rect 4252 30728 4304 30734
rect 4252 30670 4304 30676
rect 4068 30592 4120 30598
rect 4068 30534 4120 30540
rect 4080 30394 4108 30534
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 3792 30262 3844 30268
rect 3896 30280 4016 30308
rect 4264 30297 4292 30670
rect 4620 30592 4672 30598
rect 4908 30580 4936 30738
rect 5264 30660 5316 30666
rect 5264 30602 5316 30608
rect 4620 30534 4672 30540
rect 4816 30552 4936 30580
rect 4250 30288 4306 30297
rect 3700 30116 3752 30122
rect 3620 30076 3700 30104
rect 3700 30058 3752 30064
rect 3792 30048 3844 30054
rect 3792 29990 3844 29996
rect 3424 29844 3476 29850
rect 3424 29786 3476 29792
rect 3516 29776 3568 29782
rect 3516 29718 3568 29724
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 3252 29238 3280 29582
rect 3056 29232 3108 29238
rect 3056 29174 3108 29180
rect 3240 29232 3292 29238
rect 3240 29174 3292 29180
rect 3252 29102 3280 29174
rect 3528 29102 3556 29718
rect 3804 29714 3832 29990
rect 3792 29708 3844 29714
rect 3792 29650 3844 29656
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 3620 29510 3648 29582
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3804 29170 3832 29650
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 3240 29096 3292 29102
rect 3240 29038 3292 29044
rect 3516 29096 3568 29102
rect 3516 29038 3568 29044
rect 3608 29096 3660 29102
rect 3896 29050 3924 30280
rect 4068 30252 4120 30258
rect 4250 30223 4252 30232
rect 4068 30194 4120 30200
rect 4304 30223 4306 30232
rect 4436 30252 4488 30258
rect 4252 30194 4304 30200
rect 4436 30194 4488 30200
rect 4528 30252 4580 30258
rect 4528 30194 4580 30200
rect 4080 30054 4108 30194
rect 4264 30122 4292 30194
rect 4448 30161 4476 30194
rect 4434 30152 4490 30161
rect 4252 30116 4304 30122
rect 4434 30087 4490 30096
rect 4252 30058 4304 30064
rect 4540 30054 4568 30194
rect 3976 30048 4028 30054
rect 3976 29990 4028 29996
rect 4068 30048 4120 30054
rect 4068 29990 4120 29996
rect 4528 30048 4580 30054
rect 4528 29990 4580 29996
rect 3988 29782 4016 29990
rect 3976 29776 4028 29782
rect 3976 29718 4028 29724
rect 3988 29646 4016 29718
rect 4080 29646 4108 29990
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3976 29640 4028 29646
rect 3976 29582 4028 29588
rect 4068 29640 4120 29646
rect 4068 29582 4120 29588
rect 4344 29640 4396 29646
rect 4632 29617 4660 30534
rect 4712 30252 4764 30258
rect 4816 30240 4844 30552
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4764 30212 4844 30240
rect 4896 30252 4948 30258
rect 4712 30194 4764 30200
rect 5276 30240 5304 30602
rect 4896 30194 4948 30200
rect 5092 30212 5304 30240
rect 4344 29582 4396 29588
rect 4618 29608 4674 29617
rect 4080 29510 4108 29582
rect 4252 29572 4304 29578
rect 4252 29514 4304 29520
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 3660 29044 3924 29050
rect 3608 29038 3924 29044
rect 3240 28960 3292 28966
rect 3240 28902 3292 28908
rect 3252 28762 3280 28902
rect 3240 28756 3292 28762
rect 3240 28698 3292 28704
rect 3528 28694 3556 29038
rect 3620 29022 3924 29038
rect 3516 28688 3568 28694
rect 3516 28630 3568 28636
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 3056 28552 3108 28558
rect 3056 28494 3108 28500
rect 3068 28150 3096 28494
rect 3896 28490 3924 29022
rect 3884 28484 3936 28490
rect 3884 28426 3936 28432
rect 3056 28144 3108 28150
rect 3056 28086 3108 28092
rect 3068 27130 3096 28086
rect 3896 28082 3924 28426
rect 3976 28212 4028 28218
rect 3976 28154 4028 28160
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3056 27124 3108 27130
rect 3056 27066 3108 27072
rect 3516 27056 3568 27062
rect 3516 26998 3568 27004
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 848 26784 900 26790
rect 846 26752 848 26761
rect 900 26752 902 26761
rect 846 26687 902 26696
rect 1676 24744 1728 24750
rect 1676 24686 1728 24692
rect 1688 24410 1716 24686
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1780 24342 1808 26930
rect 2596 26852 2648 26858
rect 2596 26794 2648 26800
rect 2044 26240 2096 26246
rect 2044 26182 2096 26188
rect 2056 25906 2084 26182
rect 2608 25906 2636 26794
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2884 26246 2912 26726
rect 3056 26308 3108 26314
rect 3056 26250 3108 26256
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2884 25906 2912 26182
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 2596 25900 2648 25906
rect 2872 25900 2924 25906
rect 2596 25842 2648 25848
rect 2792 25860 2872 25888
rect 2608 24954 2636 25842
rect 2596 24948 2648 24954
rect 2596 24890 2648 24896
rect 1768 24336 1820 24342
rect 1768 24278 1820 24284
rect 2792 24206 2820 25860
rect 2872 25842 2924 25848
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 24274 2912 25094
rect 3068 24818 3096 26250
rect 3344 25906 3372 26930
rect 3528 25906 3556 26998
rect 3896 26994 3924 28018
rect 3988 27674 4016 28154
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 4080 27470 4108 29446
rect 4264 29170 4292 29514
rect 4252 29164 4304 29170
rect 4252 29106 4304 29112
rect 4356 29102 4384 29582
rect 4618 29543 4674 29552
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4632 28966 4660 29543
rect 4908 29492 4936 30194
rect 5092 29714 5120 30212
rect 5368 30172 5396 31334
rect 5552 30870 5580 32710
rect 5828 32570 5856 32864
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5816 32564 5868 32570
rect 5816 32506 5868 32512
rect 5920 32230 5948 32846
rect 5632 32224 5684 32230
rect 5632 32166 5684 32172
rect 5908 32224 5960 32230
rect 5908 32166 5960 32172
rect 5644 31822 5672 32166
rect 5724 32020 5776 32026
rect 5724 31962 5776 31968
rect 5632 31816 5684 31822
rect 5632 31758 5684 31764
rect 5632 31136 5684 31142
rect 5632 31078 5684 31084
rect 5644 30938 5672 31078
rect 5632 30932 5684 30938
rect 5632 30874 5684 30880
rect 5540 30864 5592 30870
rect 5736 30818 5764 31962
rect 5920 31958 5948 32166
rect 5908 31952 5960 31958
rect 5908 31894 5960 31900
rect 5920 31482 5948 31894
rect 6000 31748 6052 31754
rect 6000 31690 6052 31696
rect 5908 31476 5960 31482
rect 5908 31418 5960 31424
rect 5816 31340 5868 31346
rect 5816 31282 5868 31288
rect 5828 31142 5856 31282
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 5540 30806 5592 30812
rect 5644 30790 5764 30818
rect 5644 30734 5672 30790
rect 6012 30734 6040 31690
rect 6092 31408 6144 31414
rect 6092 31350 6144 31356
rect 6104 31210 6132 31350
rect 6092 31204 6144 31210
rect 6092 31146 6144 31152
rect 6104 30734 6132 31146
rect 5632 30728 5684 30734
rect 5446 30696 5502 30705
rect 5632 30670 5684 30676
rect 6000 30728 6052 30734
rect 6000 30670 6052 30676
rect 6092 30728 6144 30734
rect 6092 30670 6144 30676
rect 5446 30631 5502 30640
rect 5460 30598 5488 30631
rect 5448 30592 5500 30598
rect 5448 30534 5500 30540
rect 5276 30144 5396 30172
rect 5080 29708 5132 29714
rect 5080 29650 5132 29656
rect 4816 29464 4936 29492
rect 4816 29102 4844 29464
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5172 29300 5224 29306
rect 5172 29242 5224 29248
rect 4804 29096 4856 29102
rect 4804 29038 4856 29044
rect 4620 28960 4672 28966
rect 4672 28920 4752 28948
rect 4620 28902 4672 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4620 28620 4672 28626
rect 4620 28562 4672 28568
rect 4344 28484 4396 28490
rect 4344 28426 4396 28432
rect 4356 28218 4384 28426
rect 4344 28212 4396 28218
rect 4344 28154 4396 28160
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4344 27668 4396 27674
rect 4344 27610 4396 27616
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 3884 26988 3936 26994
rect 3884 26930 3936 26936
rect 3792 26784 3844 26790
rect 3792 26726 3844 26732
rect 3804 26450 3832 26726
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 3896 26042 3924 26930
rect 3974 26344 4030 26353
rect 3974 26279 4030 26288
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3332 25900 3384 25906
rect 3516 25900 3568 25906
rect 3332 25842 3384 25848
rect 3436 25860 3516 25888
rect 3240 24948 3292 24954
rect 3240 24890 3292 24896
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 2872 24268 2924 24274
rect 2872 24210 2924 24216
rect 3252 24206 3280 24890
rect 3344 24834 3372 25842
rect 3436 25294 3464 25860
rect 3516 25842 3568 25848
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 3516 25288 3568 25294
rect 3516 25230 3568 25236
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3436 24954 3464 25094
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 3344 24806 3464 24834
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2700 23730 2728 24006
rect 2792 23866 2820 24142
rect 2872 24064 2924 24070
rect 2872 24006 2924 24012
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2792 23186 2820 23802
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 848 22976 900 22982
rect 848 22918 900 22924
rect 860 22681 888 22918
rect 1412 22778 1440 23054
rect 1400 22772 1452 22778
rect 1400 22714 1452 22720
rect 846 22672 902 22681
rect 846 22607 902 22616
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1780 22030 1808 22578
rect 1768 22024 1820 22030
rect 1820 21984 1900 22012
rect 1768 21966 1820 21972
rect 1400 21888 1452 21894
rect 1306 21856 1362 21865
rect 1400 21830 1452 21836
rect 1306 21791 1362 21800
rect 1320 21690 1348 21791
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1412 21554 1440 21830
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1032 21412 1084 21418
rect 1032 21354 1084 21360
rect 1044 21185 1072 21354
rect 1030 21176 1086 21185
rect 1780 21146 1808 21490
rect 1030 21111 1086 21120
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1872 20874 1900 21984
rect 2884 21010 2912 24006
rect 2976 23594 3004 24142
rect 3056 24132 3108 24138
rect 3056 24074 3108 24080
rect 3068 23866 3096 24074
rect 3056 23860 3108 23866
rect 3056 23802 3108 23808
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 3068 22234 3096 23802
rect 3252 23730 3280 24142
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3148 23656 3200 23662
rect 3148 23598 3200 23604
rect 3160 23050 3188 23598
rect 3252 23322 3280 23666
rect 3344 23662 3372 24806
rect 3436 24750 3464 24806
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3528 24410 3556 25230
rect 3988 25158 4016 26279
rect 4080 25974 4108 27406
rect 4356 26994 4384 27610
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4540 26994 4568 27270
rect 4344 26988 4396 26994
rect 4344 26930 4396 26936
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26382 4660 28562
rect 4724 27470 4752 28920
rect 4816 27538 4844 29038
rect 4896 28960 4948 28966
rect 4896 28902 4948 28908
rect 4908 28558 4936 28902
rect 5184 28626 5212 29242
rect 5276 28762 5304 30144
rect 5356 30048 5408 30054
rect 5356 29990 5408 29996
rect 5368 29646 5396 29990
rect 5356 29640 5408 29646
rect 5356 29582 5408 29588
rect 5460 29306 5488 30534
rect 5644 30394 5672 30670
rect 6104 30394 6132 30670
rect 6196 30666 6224 34614
rect 6288 34610 6316 35566
rect 6380 35018 6408 36042
rect 6368 35012 6420 35018
rect 6368 34954 6420 34960
rect 6460 34944 6512 34950
rect 6460 34886 6512 34892
rect 6276 34604 6328 34610
rect 6276 34546 6328 34552
rect 6472 34474 6500 34886
rect 6656 34678 6684 36790
rect 6828 36712 6880 36718
rect 6828 36654 6880 36660
rect 7196 36712 7248 36718
rect 7392 36689 7420 37810
rect 7472 37120 7524 37126
rect 7472 37062 7524 37068
rect 7484 36718 7512 37062
rect 7472 36712 7524 36718
rect 7196 36654 7248 36660
rect 7378 36680 7434 36689
rect 6840 35154 6868 36654
rect 7104 36576 7156 36582
rect 7104 36518 7156 36524
rect 7012 36304 7064 36310
rect 7012 36246 7064 36252
rect 6828 35148 6880 35154
rect 6828 35090 6880 35096
rect 6644 34672 6696 34678
rect 6644 34614 6696 34620
rect 6460 34468 6512 34474
rect 6460 34410 6512 34416
rect 6368 34400 6420 34406
rect 6368 34342 6420 34348
rect 6380 33930 6408 34342
rect 6472 33998 6500 34410
rect 6644 34128 6696 34134
rect 6644 34070 6696 34076
rect 6460 33992 6512 33998
rect 6460 33934 6512 33940
rect 6368 33924 6420 33930
rect 6368 33866 6420 33872
rect 6380 33046 6408 33866
rect 6472 33590 6500 33934
rect 6460 33584 6512 33590
rect 6460 33526 6512 33532
rect 6368 33040 6420 33046
rect 6368 32982 6420 32988
rect 6276 32496 6328 32502
rect 6276 32438 6328 32444
rect 6184 30660 6236 30666
rect 6184 30602 6236 30608
rect 5632 30388 5684 30394
rect 5632 30330 5684 30336
rect 6092 30388 6144 30394
rect 6092 30330 6144 30336
rect 5632 30116 5684 30122
rect 5632 30058 5684 30064
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5552 29850 5580 29990
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 5448 29300 5500 29306
rect 5448 29242 5500 29248
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5264 28756 5316 28762
rect 5264 28698 5316 28704
rect 5172 28620 5224 28626
rect 5172 28562 5224 28568
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5368 28218 5396 29106
rect 5540 28484 5592 28490
rect 5540 28426 5592 28432
rect 5552 28218 5580 28426
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5540 28212 5592 28218
rect 5540 28154 5592 28160
rect 4896 28008 4948 28014
rect 4896 27950 4948 27956
rect 5264 28008 5316 28014
rect 5368 27996 5396 28154
rect 5644 28150 5672 30058
rect 5724 29164 5776 29170
rect 5724 29106 5776 29112
rect 5736 28422 5764 29106
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 5448 28144 5500 28150
rect 5448 28086 5500 28092
rect 5632 28144 5684 28150
rect 5632 28086 5684 28092
rect 5316 27968 5396 27996
rect 5264 27950 5316 27956
rect 4908 27674 4936 27950
rect 5172 27940 5224 27946
rect 5172 27882 5224 27888
rect 4896 27668 4948 27674
rect 4896 27610 4948 27616
rect 5184 27606 5212 27882
rect 5264 27872 5316 27878
rect 5264 27814 5316 27820
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 4804 27532 4856 27538
rect 4804 27474 4856 27480
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4724 26858 4752 27406
rect 4816 27130 4844 27474
rect 5276 27470 5304 27814
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4804 27124 4856 27130
rect 4804 27066 4856 27072
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4712 26852 4764 26858
rect 4712 26794 4764 26800
rect 4816 26586 4844 26862
rect 5264 26852 5316 26858
rect 5264 26794 5316 26800
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 5080 26376 5132 26382
rect 5172 26376 5224 26382
rect 5080 26318 5132 26324
rect 5170 26344 5172 26353
rect 5224 26344 5226 26353
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 4632 25906 4660 26318
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4080 25226 4108 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25362 4660 25842
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 4620 25356 4672 25362
rect 4620 25298 4672 25304
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3516 24404 3568 24410
rect 3516 24346 3568 24352
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3436 23798 3464 24142
rect 3424 23792 3476 23798
rect 3424 23734 3476 23740
rect 3712 23662 3740 24754
rect 3332 23656 3384 23662
rect 3332 23598 3384 23604
rect 3700 23656 3752 23662
rect 3700 23598 3752 23604
rect 3240 23316 3292 23322
rect 3240 23258 3292 23264
rect 3252 23118 3280 23258
rect 3712 23254 3740 23598
rect 3792 23588 3844 23594
rect 3792 23530 3844 23536
rect 3700 23248 3752 23254
rect 3700 23190 3752 23196
rect 3804 23118 3832 23530
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 3608 23112 3660 23118
rect 3608 23054 3660 23060
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3148 23044 3200 23050
rect 3148 22986 3200 22992
rect 3160 22710 3188 22986
rect 3148 22704 3200 22710
rect 3148 22646 3200 22652
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3160 22030 3188 22510
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 3160 20942 3188 21966
rect 3620 21622 3648 23054
rect 3988 22710 4016 25094
rect 4172 24682 4200 25298
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23186 4660 25298
rect 4724 24818 4752 26318
rect 5092 26246 5120 26318
rect 5170 26279 5226 26288
rect 5080 26240 5132 26246
rect 5080 26182 5132 26188
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5276 25906 5304 26794
rect 5368 25906 5396 27968
rect 5460 27334 5488 28086
rect 5736 28014 5764 28358
rect 5724 28008 5776 28014
rect 5552 27968 5724 27996
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5460 26994 5488 27270
rect 5448 26988 5500 26994
rect 5448 26930 5500 26936
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 5264 25900 5316 25906
rect 5264 25842 5316 25848
rect 5356 25900 5408 25906
rect 5356 25842 5408 25848
rect 4816 24886 4844 25842
rect 5276 25498 5304 25842
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 5356 25288 5408 25294
rect 5356 25230 5408 25236
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5368 24954 5396 25230
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4816 24206 4844 24822
rect 5356 24744 5408 24750
rect 5356 24686 5408 24692
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 5368 24138 5396 24686
rect 5552 24206 5580 27968
rect 5724 27950 5776 27956
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5736 26858 5764 27270
rect 6000 26920 6052 26926
rect 6000 26862 6052 26868
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5736 26450 5764 26794
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5736 26042 5764 26250
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5724 26036 5776 26042
rect 5724 25978 5776 25984
rect 5632 25968 5684 25974
rect 5632 25910 5684 25916
rect 5644 25158 5672 25910
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5644 24818 5672 25094
rect 5632 24812 5684 24818
rect 5632 24754 5684 24760
rect 5644 24206 5672 24754
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5356 24132 5408 24138
rect 5356 24074 5408 24080
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5172 23656 5224 23662
rect 5092 23604 5172 23610
rect 5092 23598 5224 23604
rect 5092 23582 5212 23598
rect 4988 23520 5040 23526
rect 4988 23462 5040 23468
rect 5000 23186 5028 23462
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 5092 23050 5120 23582
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22778 5304 23666
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 3976 22704 4028 22710
rect 3896 22664 3976 22692
rect 3700 21888 3752 21894
rect 3700 21830 3752 21836
rect 3608 21616 3660 21622
rect 3608 21558 3660 21564
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1872 20602 1900 20810
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17746 1440 18770
rect 1768 18760 1820 18766
rect 1768 18702 1820 18708
rect 1780 18426 1808 18702
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 17785 1532 18226
rect 1490 17776 1546 17785
rect 1400 17740 1452 17746
rect 1490 17711 1546 17720
rect 1400 17682 1452 17688
rect 1768 17672 1820 17678
rect 1768 17614 1820 17620
rect 1780 17338 1808 17614
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 848 17196 900 17202
rect 848 17138 900 17144
rect 860 16969 888 17138
rect 846 16960 902 16969
rect 846 16895 902 16904
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 860 15881 888 16050
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1412 15026 1440 15506
rect 1688 15065 1716 16050
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1780 15502 1808 15846
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1674 15056 1730 15065
rect 1400 15020 1452 15026
rect 1872 15026 1900 15846
rect 1674 14991 1730 15000
rect 1860 15020 1912 15026
rect 1400 14962 1452 14968
rect 1860 14962 1912 14968
rect 2240 13190 2268 20402
rect 3160 20398 3188 20878
rect 3332 20800 3384 20806
rect 3332 20742 3384 20748
rect 3344 20466 3372 20742
rect 3712 20534 3740 21830
rect 3896 20942 3924 22664
rect 3976 22646 4028 22652
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4526 22128 4582 22137
rect 4344 22092 4396 22098
rect 4632 22098 4660 22578
rect 4724 22234 4752 22578
rect 5172 22568 5224 22574
rect 5224 22516 5304 22522
rect 5172 22510 5304 22516
rect 5184 22494 5304 22510
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4526 22063 4582 22072
rect 4620 22092 4672 22098
rect 4344 22034 4396 22040
rect 4252 21956 4304 21962
rect 4252 21898 4304 21904
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 3700 20528 3752 20534
rect 3752 20488 3832 20516
rect 3700 20470 3752 20476
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3160 19786 3188 20334
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 2424 19378 2452 19722
rect 3804 19446 3832 20488
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 2412 19372 2464 19378
rect 3804 19334 3832 19382
rect 2412 19314 2464 19320
rect 2424 18850 2452 19314
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3712 19306 3832 19334
rect 3620 18970 3648 19246
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 2332 18834 2452 18850
rect 2320 18828 2452 18834
rect 2372 18822 2452 18828
rect 2320 18770 2372 18776
rect 2424 18222 2452 18822
rect 3712 18698 3740 19306
rect 3700 18692 3752 18698
rect 3700 18634 3752 18640
rect 3712 18578 3740 18634
rect 3620 18550 3740 18578
rect 3620 18358 3648 18550
rect 3608 18352 3660 18358
rect 3608 18294 3660 18300
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 2424 17202 2452 18158
rect 3804 17882 3832 18158
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 2608 17338 2636 17546
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2424 16114 2452 17138
rect 2608 16250 2636 17274
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16794 3004 17070
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2424 15586 2452 16050
rect 2332 15570 2452 15586
rect 2320 15564 2452 15570
rect 2372 15558 2452 15564
rect 2320 15506 2372 15512
rect 2608 15434 2636 16186
rect 2596 15428 2648 15434
rect 2596 15370 2648 15376
rect 2608 15094 2636 15370
rect 3252 15162 3280 16594
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3804 15706 3832 15982
rect 3792 15700 3844 15706
rect 3792 15642 3844 15648
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2424 13394 2452 13806
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12918 2268 13126
rect 2516 12986 2544 14350
rect 2608 13818 2636 15030
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2700 14006 2728 14214
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2688 13864 2740 13870
rect 2608 13812 2688 13818
rect 2608 13806 2740 13812
rect 2608 13790 2728 13806
rect 2700 13258 2728 13790
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2976 12986 3004 13194
rect 3436 12986 3464 13262
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1688 12442 1716 12786
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1964 11762 1992 12378
rect 2240 12306 2268 12854
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 848 11552 900 11558
rect 846 11520 848 11529
rect 900 11520 902 11529
rect 846 11455 902 11464
rect 1964 11354 1992 11698
rect 2056 11558 2084 12174
rect 2240 11762 2268 12242
rect 2516 12170 2544 12922
rect 2596 12844 2648 12850
rect 3516 12844 3568 12850
rect 2648 12804 2820 12832
rect 2596 12786 2648 12792
rect 2792 12374 2820 12804
rect 3516 12786 3568 12792
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2516 11762 2544 12106
rect 2792 11762 2820 12310
rect 3528 11898 3556 12786
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2056 11218 2084 11494
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2148 11150 2176 11562
rect 2240 11150 2268 11698
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1544 10976 1546 10985
rect 1490 10911 1546 10920
rect 2516 10810 2544 11222
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 3160 11014 3188 11154
rect 3436 11082 3464 11630
rect 3528 11218 3556 11834
rect 3804 11762 3832 12242
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3896 11150 3924 15982
rect 3988 14414 4016 21490
rect 4264 21418 4292 21898
rect 4356 21690 4384 22034
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4252 21412 4304 21418
rect 4252 21354 4304 21360
rect 4540 21350 4568 22063
rect 4620 22034 4672 22040
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4632 21622 4660 21830
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 4528 21344 4580 21350
rect 4528 21286 4580 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4172 20330 4200 20878
rect 4632 20602 4660 21558
rect 4816 21554 4844 22374
rect 5000 21894 5028 22374
rect 5092 22137 5120 22374
rect 5078 22128 5134 22137
rect 5078 22063 5134 22072
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4724 20466 4752 20946
rect 4908 20942 4936 21082
rect 5000 20942 5028 21490
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18834 4660 19722
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4724 18714 4752 19314
rect 4816 18970 4844 20878
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20602 5304 22494
rect 5368 22438 5396 24074
rect 5552 22642 5580 24142
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5356 22432 5408 22438
rect 5356 22374 5408 22380
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5368 21026 5396 22170
rect 5368 20998 5488 21026
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5368 20602 5396 20878
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5184 20482 5212 20538
rect 5184 20454 5304 20482
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 5000 18766 5028 19110
rect 5092 18902 5120 19178
rect 5276 18902 5304 20454
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 4988 18760 5040 18766
rect 4252 18692 4304 18698
rect 4252 18634 4304 18640
rect 4632 18686 4752 18714
rect 4816 18720 4988 18748
rect 4264 18426 4292 18634
rect 4632 18426 4660 18686
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17678 4660 18226
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16522 4660 17614
rect 4724 17270 4752 18566
rect 4816 18358 4844 18720
rect 4988 18702 5040 18708
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 5184 18630 5212 18702
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18426 5304 18702
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 4712 17264 4764 17270
rect 4712 17206 4764 17212
rect 4816 17202 4844 18158
rect 5184 17678 5212 18158
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5276 17338 5304 18158
rect 5368 17882 5396 20402
rect 5460 20330 5488 20998
rect 5644 20466 5672 22918
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5736 20466 5764 22578
rect 5828 20602 5856 26182
rect 6012 24614 6040 26862
rect 6196 26586 6224 30602
rect 6288 30326 6316 32438
rect 6380 32026 6408 32982
rect 6368 32020 6420 32026
rect 6368 31962 6420 31968
rect 6368 31884 6420 31890
rect 6368 31826 6420 31832
rect 6380 31346 6408 31826
rect 6656 31822 6684 34070
rect 6920 33924 6972 33930
rect 6920 33866 6972 33872
rect 6736 33652 6788 33658
rect 6736 33594 6788 33600
rect 6748 32910 6776 33594
rect 6932 33454 6960 33866
rect 6920 33448 6972 33454
rect 6920 33390 6972 33396
rect 6828 33312 6880 33318
rect 6828 33254 6880 33260
rect 6840 33114 6868 33254
rect 6828 33108 6880 33114
rect 6828 33050 6880 33056
rect 6932 32910 6960 33390
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 7024 32722 7052 36246
rect 7116 36174 7144 36518
rect 7208 36378 7236 36654
rect 7472 36654 7524 36660
rect 7378 36615 7434 36624
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7392 36242 7420 36615
rect 7380 36236 7432 36242
rect 7380 36178 7432 36184
rect 7104 36168 7156 36174
rect 7104 36110 7156 36116
rect 7576 36106 7604 37828
rect 7944 37398 7972 38150
rect 8024 37868 8076 37874
rect 8312 37856 8340 38354
rect 11612 38344 11664 38350
rect 11612 38286 11664 38292
rect 9680 38276 9732 38282
rect 9680 38218 9732 38224
rect 8944 38208 8996 38214
rect 8944 38150 8996 38156
rect 8956 37942 8984 38150
rect 8944 37936 8996 37942
rect 8944 37878 8996 37884
rect 8076 37828 8340 37856
rect 8024 37810 8076 37816
rect 8036 37738 8064 37810
rect 8024 37732 8076 37738
rect 8024 37674 8076 37680
rect 8116 37732 8168 37738
rect 8116 37674 8168 37680
rect 8128 37618 8156 37674
rect 8036 37590 8156 37618
rect 7932 37392 7984 37398
rect 7932 37334 7984 37340
rect 8036 37126 8064 37590
rect 8312 37262 8340 37828
rect 8576 37732 8628 37738
rect 8576 37674 8628 37680
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 8404 37126 8432 37606
rect 8588 37262 8616 37674
rect 9692 37330 9720 38218
rect 9680 37324 9732 37330
rect 9680 37266 9732 37272
rect 8576 37256 8628 37262
rect 8576 37198 8628 37204
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 8116 37120 8168 37126
rect 8116 37062 8168 37068
rect 8392 37120 8444 37126
rect 8392 37062 8444 37068
rect 8036 36310 8064 37062
rect 8128 36922 8156 37062
rect 8116 36916 8168 36922
rect 8116 36858 8168 36864
rect 8024 36304 8076 36310
rect 8024 36246 8076 36252
rect 8128 36242 8156 36858
rect 8116 36236 8168 36242
rect 8116 36178 8168 36184
rect 9588 36168 9640 36174
rect 9588 36110 9640 36116
rect 7564 36100 7616 36106
rect 7484 36060 7564 36088
rect 7288 35148 7340 35154
rect 7288 35090 7340 35096
rect 7300 34542 7328 35090
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 7378 34504 7434 34513
rect 7300 33998 7328 34478
rect 7378 34439 7434 34448
rect 7392 33998 7420 34439
rect 7288 33992 7340 33998
rect 7288 33934 7340 33940
rect 7380 33992 7432 33998
rect 7380 33934 7432 33940
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 7116 33318 7144 33594
rect 7196 33516 7248 33522
rect 7196 33458 7248 33464
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 7116 32910 7144 33254
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7024 32694 7144 32722
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 6932 31906 6960 32370
rect 6840 31878 6960 31906
rect 6840 31822 6868 31878
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6920 31816 6972 31822
rect 6972 31764 7052 31770
rect 6920 31758 7052 31764
rect 6932 31726 7052 31758
rect 6368 31340 6420 31346
rect 6368 31282 6420 31288
rect 6932 31278 6960 31726
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6932 30802 6960 31214
rect 6920 30796 6972 30802
rect 6920 30738 6972 30744
rect 6932 30394 6960 30738
rect 6920 30388 6972 30394
rect 6920 30330 6972 30336
rect 6276 30320 6328 30326
rect 6276 30262 6328 30268
rect 6552 30320 6604 30326
rect 6552 30262 6604 30268
rect 6564 28558 6592 30262
rect 6932 29170 6960 30330
rect 6920 29164 6972 29170
rect 6920 29106 6972 29112
rect 7116 28762 7144 32694
rect 7208 32434 7236 33458
rect 7300 33386 7328 33934
rect 7484 33454 7512 36060
rect 7564 36042 7616 36048
rect 7656 35692 7708 35698
rect 7656 35634 7708 35640
rect 8208 35692 8260 35698
rect 8208 35634 8260 35640
rect 7668 35578 7696 35634
rect 7668 35550 7788 35578
rect 7564 35012 7616 35018
rect 7564 34954 7616 34960
rect 7576 34542 7604 34954
rect 7564 34536 7616 34542
rect 7564 34478 7616 34484
rect 7760 34474 7788 35550
rect 7840 35488 7892 35494
rect 7840 35430 7892 35436
rect 7852 34610 7880 35430
rect 8220 34678 8248 35634
rect 9496 35624 9548 35630
rect 9600 35578 9628 36110
rect 9692 36088 9720 37266
rect 10048 36712 10100 36718
rect 10048 36654 10100 36660
rect 11336 36712 11388 36718
rect 11336 36654 11388 36660
rect 9864 36576 9916 36582
rect 9864 36518 9916 36524
rect 9876 36242 9904 36518
rect 9864 36236 9916 36242
rect 9864 36178 9916 36184
rect 9772 36100 9824 36106
rect 9692 36060 9772 36088
rect 9692 35834 9720 36060
rect 9772 36042 9824 36048
rect 9680 35828 9732 35834
rect 9680 35770 9732 35776
rect 9548 35572 9628 35578
rect 9496 35566 9628 35572
rect 9508 35550 9628 35566
rect 9600 35154 9628 35550
rect 9692 35222 9720 35770
rect 9864 35624 9916 35630
rect 9864 35566 9916 35572
rect 9876 35290 9904 35566
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 9680 35216 9732 35222
rect 9680 35158 9732 35164
rect 9588 35148 9640 35154
rect 9588 35090 9640 35096
rect 9692 35018 9720 35158
rect 10060 35086 10088 36654
rect 10508 36576 10560 36582
rect 10508 36518 10560 36524
rect 11060 36576 11112 36582
rect 11060 36518 11112 36524
rect 10520 36242 10548 36518
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 10520 35086 10548 36178
rect 10048 35080 10100 35086
rect 10048 35022 10100 35028
rect 10508 35080 10560 35086
rect 10508 35022 10560 35028
rect 9128 35012 9180 35018
rect 9128 34954 9180 34960
rect 9680 35012 9732 35018
rect 9680 34954 9732 34960
rect 8576 34944 8628 34950
rect 8576 34886 8628 34892
rect 8208 34672 8260 34678
rect 8036 34632 8208 34660
rect 7840 34604 7892 34610
rect 7840 34546 7892 34552
rect 7932 34604 7984 34610
rect 7932 34546 7984 34552
rect 7748 34468 7800 34474
rect 7748 34410 7800 34416
rect 7656 34060 7708 34066
rect 7656 34002 7708 34008
rect 7380 33448 7432 33454
rect 7380 33390 7432 33396
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7288 33380 7340 33386
rect 7288 33322 7340 33328
rect 7392 33114 7420 33390
rect 7380 33108 7432 33114
rect 7380 33050 7432 33056
rect 7668 32910 7696 34002
rect 7760 33998 7788 34410
rect 7944 34202 7972 34546
rect 7932 34196 7984 34202
rect 7932 34138 7984 34144
rect 8036 33998 8064 34632
rect 8208 34614 8260 34620
rect 8588 34406 8616 34886
rect 8116 34400 8168 34406
rect 8116 34342 8168 34348
rect 8392 34400 8444 34406
rect 8392 34342 8444 34348
rect 8576 34400 8628 34406
rect 8576 34342 8628 34348
rect 8128 34202 8156 34342
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 7748 33992 7800 33998
rect 7748 33934 7800 33940
rect 7840 33992 7892 33998
rect 7840 33934 7892 33940
rect 8024 33992 8076 33998
rect 8024 33934 8076 33940
rect 7852 33590 7880 33934
rect 7932 33924 7984 33930
rect 7932 33866 7984 33872
rect 7840 33584 7892 33590
rect 7840 33526 7892 33532
rect 7944 33522 7972 33866
rect 7932 33516 7984 33522
rect 7932 33458 7984 33464
rect 8024 33448 8076 33454
rect 8024 33390 8076 33396
rect 7656 32904 7708 32910
rect 7656 32846 7708 32852
rect 7668 32502 7696 32846
rect 7656 32496 7708 32502
rect 7656 32438 7708 32444
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 7380 32360 7432 32366
rect 7380 32302 7432 32308
rect 7392 32026 7420 32302
rect 7748 32292 7800 32298
rect 7748 32234 7800 32240
rect 7380 32020 7432 32026
rect 7380 31962 7432 31968
rect 7760 31890 7788 32234
rect 7932 32224 7984 32230
rect 7932 32166 7984 32172
rect 7748 31884 7800 31890
rect 7748 31826 7800 31832
rect 7196 31748 7248 31754
rect 7196 31690 7248 31696
rect 7208 31482 7236 31690
rect 7196 31476 7248 31482
rect 7196 31418 7248 31424
rect 7760 31346 7788 31826
rect 7944 31346 7972 32166
rect 8036 31414 8064 33390
rect 8404 32910 8432 34342
rect 8588 33998 8616 34342
rect 8576 33992 8628 33998
rect 8576 33934 8628 33940
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8404 32434 8432 32846
rect 8496 32842 8524 33798
rect 9140 33590 9168 34954
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 9416 33998 9444 34614
rect 10060 34610 10088 35022
rect 10968 35012 11020 35018
rect 10968 34954 11020 34960
rect 10980 34678 11008 34954
rect 11072 34950 11100 36518
rect 11348 36378 11376 36654
rect 11624 36650 11652 38286
rect 12072 38276 12124 38282
rect 12072 38218 12124 38224
rect 12084 37466 12112 38218
rect 12912 37806 12940 38830
rect 13820 38480 13872 38486
rect 13820 38422 13872 38428
rect 12900 37800 12952 37806
rect 12900 37742 12952 37748
rect 12072 37460 12124 37466
rect 12072 37402 12124 37408
rect 12084 36802 12112 37402
rect 12256 37256 12308 37262
rect 12532 37256 12584 37262
rect 12308 37216 12388 37244
rect 12256 37198 12308 37204
rect 12164 37188 12216 37194
rect 12164 37130 12216 37136
rect 11992 36786 12112 36802
rect 11980 36780 12112 36786
rect 12032 36774 12112 36780
rect 11980 36722 12032 36728
rect 12072 36712 12124 36718
rect 12072 36654 12124 36660
rect 11612 36644 11664 36650
rect 11612 36586 11664 36592
rect 11336 36372 11388 36378
rect 11336 36314 11388 36320
rect 11520 35624 11572 35630
rect 11624 35612 11652 36586
rect 11704 36032 11756 36038
rect 11704 35974 11756 35980
rect 11716 35766 11744 35974
rect 12084 35834 12112 36654
rect 12072 35828 12124 35834
rect 12072 35770 12124 35776
rect 11704 35760 11756 35766
rect 11704 35702 11756 35708
rect 11572 35584 11652 35612
rect 11520 35566 11572 35572
rect 11532 35154 11560 35566
rect 11520 35148 11572 35154
rect 11520 35090 11572 35096
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 10968 34672 11020 34678
rect 10968 34614 11020 34620
rect 11072 34610 11100 34886
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 11060 34604 11112 34610
rect 11060 34546 11112 34552
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9416 33658 9444 33934
rect 9404 33652 9456 33658
rect 9404 33594 9456 33600
rect 9128 33584 9180 33590
rect 9128 33526 9180 33532
rect 10232 33516 10284 33522
rect 10232 33458 10284 33464
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9968 33046 9996 33390
rect 10244 33114 10272 33458
rect 10336 33114 10364 34546
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 11060 33312 11112 33318
rect 11060 33254 11112 33260
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 10324 33108 10376 33114
rect 10324 33050 10376 33056
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 9956 33040 10008 33046
rect 9956 32982 10008 32988
rect 10336 32978 10364 33050
rect 10324 32972 10376 32978
rect 10324 32914 10376 32920
rect 10888 32842 10916 33050
rect 11072 32994 11100 33254
rect 10980 32978 11100 32994
rect 10968 32972 11100 32978
rect 11020 32966 11100 32972
rect 10968 32914 11020 32920
rect 11164 32910 11192 33798
rect 11532 33522 11560 35090
rect 11612 34740 11664 34746
rect 11612 34682 11664 34688
rect 11624 34066 11652 34682
rect 12176 34678 12204 37130
rect 12256 36576 12308 36582
rect 12256 36518 12308 36524
rect 12268 36242 12296 36518
rect 12360 36310 12388 37216
rect 12532 37198 12584 37204
rect 12544 36922 12572 37198
rect 12912 37194 12940 37742
rect 12900 37188 12952 37194
rect 12900 37130 12952 37136
rect 12532 36916 12584 36922
rect 12532 36858 12584 36864
rect 12348 36304 12400 36310
rect 12348 36246 12400 36252
rect 12256 36236 12308 36242
rect 12256 36178 12308 36184
rect 12360 36122 12388 36246
rect 12268 36094 12388 36122
rect 12268 35290 12296 36094
rect 12256 35284 12308 35290
rect 12256 35226 12308 35232
rect 12164 34672 12216 34678
rect 12164 34614 12216 34620
rect 11612 34060 11664 34066
rect 11612 34002 11664 34008
rect 11520 33516 11572 33522
rect 11520 33458 11572 33464
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 8484 32836 8536 32842
rect 8484 32778 8536 32784
rect 10876 32836 10928 32842
rect 10876 32778 10928 32784
rect 12164 32836 12216 32842
rect 12164 32778 12216 32784
rect 8392 32428 8444 32434
rect 8392 32370 8444 32376
rect 8208 32360 8260 32366
rect 8208 32302 8260 32308
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 12072 32360 12124 32366
rect 12072 32302 12124 32308
rect 8220 32026 8248 32302
rect 8668 32224 8720 32230
rect 8668 32166 8720 32172
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8208 31680 8260 31686
rect 8208 31622 8260 31628
rect 8024 31408 8076 31414
rect 8024 31350 8076 31356
rect 7748 31340 7800 31346
rect 7748 31282 7800 31288
rect 7932 31340 7984 31346
rect 7932 31282 7984 31288
rect 8220 31142 8248 31622
rect 8680 31482 8708 32166
rect 9324 32026 9352 32302
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 9312 32020 9364 32026
rect 9312 31962 9364 31968
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 8668 31476 8720 31482
rect 8668 31418 8720 31424
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 7840 30184 7892 30190
rect 7840 30126 7892 30132
rect 7852 29850 7880 30126
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 7104 28756 7156 28762
rect 7104 28698 7156 28704
rect 6552 28552 6604 28558
rect 6472 28512 6552 28540
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6472 26330 6500 28512
rect 6552 28494 6604 28500
rect 7116 28082 7144 28698
rect 8036 28490 8064 29446
rect 8024 28484 8076 28490
rect 8024 28426 8076 28432
rect 7104 28076 7156 28082
rect 7104 28018 7156 28024
rect 8116 28008 8168 28014
rect 8116 27950 8168 27956
rect 8128 27130 8156 27950
rect 8116 27124 8168 27130
rect 8116 27066 8168 27072
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 6552 26784 6604 26790
rect 6552 26726 6604 26732
rect 6288 26314 6500 26330
rect 6288 26308 6512 26314
rect 6288 26302 6460 26308
rect 6288 25294 6316 26302
rect 6460 26250 6512 26256
rect 6564 25906 6592 26726
rect 7104 26308 7156 26314
rect 7104 26250 7156 26256
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 7024 25906 7052 26182
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 6012 24274 6040 24550
rect 6288 24274 6316 25230
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6472 24954 6500 25162
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 6564 24886 6592 25842
rect 7116 25838 7144 26250
rect 7104 25832 7156 25838
rect 7104 25774 7156 25780
rect 6644 25764 6696 25770
rect 6644 25706 6696 25712
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 6276 24268 6328 24274
rect 6276 24210 6328 24216
rect 5908 23044 5960 23050
rect 5908 22986 5960 22992
rect 5920 22710 5948 22986
rect 5908 22704 5960 22710
rect 5908 22646 5960 22652
rect 6012 21622 6040 24210
rect 6288 23730 6316 24210
rect 6564 23798 6592 24822
rect 6656 24818 6684 25706
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6644 24676 6696 24682
rect 6644 24618 6696 24624
rect 6656 24206 6684 24618
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6840 23866 6868 24754
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6932 23866 6960 24346
rect 7116 24342 7144 25774
rect 7104 24336 7156 24342
rect 7104 24278 7156 24284
rect 7208 24138 7236 26862
rect 7564 26512 7616 26518
rect 7564 26454 7616 26460
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7484 24800 7512 25638
rect 7576 25498 7604 26454
rect 8128 26382 8156 27066
rect 8220 27062 8248 31078
rect 10152 30326 10180 31214
rect 10140 30320 10192 30326
rect 10140 30262 10192 30268
rect 10428 30258 10456 31826
rect 10520 30802 10548 32166
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 10784 31748 10836 31754
rect 10784 31690 10836 31696
rect 10876 31748 10928 31754
rect 10876 31690 10928 31696
rect 10796 30938 10824 31690
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10888 30802 10916 31690
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 10980 31414 11008 31622
rect 10968 31408 11020 31414
rect 10968 31350 11020 31356
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 10876 30796 10928 30802
rect 10876 30738 10928 30744
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10612 30190 10640 30670
rect 10692 30592 10744 30598
rect 10692 30534 10744 30540
rect 10704 30258 10732 30534
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8404 28558 8432 29106
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 8496 28218 8524 29446
rect 8680 28218 8708 29514
rect 8944 29504 8996 29510
rect 8944 29446 8996 29452
rect 8956 29306 8984 29446
rect 8944 29300 8996 29306
rect 8944 29242 8996 29248
rect 9048 28966 9076 30126
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9324 29646 9352 29990
rect 9588 29708 9640 29714
rect 9588 29650 9640 29656
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9128 29164 9180 29170
rect 9128 29106 9180 29112
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 9140 28762 9168 29106
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 9416 28218 9444 29446
rect 9600 28626 9628 29650
rect 10232 29640 10284 29646
rect 10232 29582 10284 29588
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 10048 29504 10100 29510
rect 10048 29446 10100 29452
rect 9680 28756 9732 28762
rect 9680 28698 9732 28704
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9692 28082 9720 28698
rect 9784 28558 9812 29446
rect 10060 29170 10088 29446
rect 10244 29306 10272 29582
rect 10704 29306 10732 30194
rect 10888 30122 10916 30738
rect 10980 30598 11008 31350
rect 11532 31346 11560 31758
rect 12084 31754 12112 32302
rect 12176 31822 12204 32778
rect 12164 31816 12216 31822
rect 12164 31758 12216 31764
rect 12072 31748 12124 31754
rect 12072 31690 12124 31696
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 12084 31278 12112 31690
rect 12072 31272 12124 31278
rect 12072 31214 12124 31220
rect 12176 31142 12204 31758
rect 11980 31136 12032 31142
rect 11980 31078 12032 31084
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 11152 30660 11204 30666
rect 11152 30602 11204 30608
rect 10968 30592 11020 30598
rect 10968 30534 11020 30540
rect 11164 30394 11192 30602
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 10876 30116 10928 30122
rect 10876 30058 10928 30064
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10692 29300 10744 29306
rect 10692 29242 10744 29248
rect 10244 29170 10272 29242
rect 10784 29232 10836 29238
rect 10888 29220 10916 30058
rect 10980 29306 11008 30194
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 11060 29640 11112 29646
rect 11164 29628 11192 30126
rect 11112 29600 11192 29628
rect 11060 29582 11112 29588
rect 10968 29300 11020 29306
rect 10968 29242 11020 29248
rect 10836 29192 10916 29220
rect 10784 29174 10836 29180
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10692 29164 10744 29170
rect 10692 29106 10744 29112
rect 10060 28558 10088 29106
rect 10508 29096 10560 29102
rect 10508 29038 10560 29044
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 10048 28552 10100 28558
rect 10048 28494 10100 28500
rect 10140 28552 10192 28558
rect 10140 28494 10192 28500
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 10152 28014 10180 28494
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 8208 27056 8260 27062
rect 8208 26998 8260 27004
rect 8220 26926 8248 26998
rect 10060 26994 10088 27882
rect 10152 26994 10180 27950
rect 10244 27130 10272 28970
rect 10324 28960 10376 28966
rect 10324 28902 10376 28908
rect 10336 28694 10364 28902
rect 10324 28688 10376 28694
rect 10324 28630 10376 28636
rect 10520 27878 10548 29038
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10612 28626 10640 28902
rect 10600 28620 10652 28626
rect 10600 28562 10652 28568
rect 10704 27946 10732 29106
rect 10692 27940 10744 27946
rect 10692 27882 10744 27888
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 10428 27130 10456 27338
rect 10232 27124 10284 27130
rect 10232 27066 10284 27072
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10520 26994 10548 27814
rect 10784 27464 10836 27470
rect 10888 27452 10916 29192
rect 10968 28416 11020 28422
rect 10968 28358 11020 28364
rect 10836 27424 10916 27452
rect 10784 27406 10836 27412
rect 10600 27328 10652 27334
rect 10600 27270 10652 27276
rect 10612 27130 10640 27270
rect 10600 27124 10652 27130
rect 10600 27066 10652 27072
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 10048 26988 10100 26994
rect 10048 26930 10100 26936
rect 10140 26988 10192 26994
rect 10140 26930 10192 26936
rect 10508 26988 10560 26994
rect 10508 26930 10560 26936
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8116 26376 8168 26382
rect 8116 26318 8168 26324
rect 8036 26042 8064 26318
rect 8024 26036 8076 26042
rect 8024 25978 8076 25984
rect 8404 25974 8432 26726
rect 8588 26586 8616 26862
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 9692 26382 9720 26930
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8496 26042 8524 26250
rect 8484 26036 8536 26042
rect 8484 25978 8536 25984
rect 8392 25968 8444 25974
rect 8392 25910 8444 25916
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 7564 25492 7616 25498
rect 7564 25434 7616 25440
rect 7576 24954 7604 25434
rect 7668 24954 7696 25842
rect 7564 24948 7616 24954
rect 7564 24890 7616 24896
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7562 24848 7618 24857
rect 7852 24818 7880 25842
rect 8208 25832 8260 25838
rect 8208 25774 8260 25780
rect 8220 24954 8248 25774
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 7484 24792 7562 24800
rect 7484 24772 7564 24792
rect 7392 24698 7420 24754
rect 7300 24670 7420 24698
rect 7300 24274 7328 24670
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 6552 23792 6604 23798
rect 6552 23734 6604 23740
rect 6276 23724 6328 23730
rect 6828 23724 6880 23730
rect 6276 23666 6328 23672
rect 6748 23684 6828 23712
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6472 23118 6500 23258
rect 6460 23112 6512 23118
rect 6460 23054 6512 23060
rect 6564 21894 6592 23598
rect 6748 23050 6776 23684
rect 6828 23666 6880 23672
rect 6826 23216 6882 23225
rect 7024 23202 7052 24074
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7116 23662 7144 24006
rect 7300 23798 7328 24074
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7392 23730 7420 24550
rect 7484 24138 7512 24772
rect 7616 24783 7618 24792
rect 7656 24812 7708 24818
rect 7564 24754 7616 24760
rect 7656 24754 7708 24760
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7668 24274 7696 24754
rect 7656 24268 7708 24274
rect 7656 24210 7708 24216
rect 7668 24138 7696 24210
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7196 23656 7248 23662
rect 7196 23598 7248 23604
rect 7208 23322 7236 23598
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 6826 23151 6882 23160
rect 6932 23174 7052 23202
rect 6840 23118 6868 23151
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6932 22982 6960 23174
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 22024 6880 22030
rect 6932 21978 6960 22714
rect 7024 22574 7052 23054
rect 7208 23050 7236 23258
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7196 23044 7248 23050
rect 7196 22986 7248 22992
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7024 22166 7052 22374
rect 7012 22160 7064 22166
rect 7012 22102 7064 22108
rect 7116 22098 7144 22986
rect 7208 22438 7236 22986
rect 7392 22982 7420 23666
rect 7668 23118 7696 24074
rect 7852 23866 7880 24754
rect 8312 24682 8340 25842
rect 8300 24676 8352 24682
rect 8300 24618 8352 24624
rect 8312 24274 8340 24618
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7852 23526 7880 23802
rect 7932 23724 7984 23730
rect 7932 23666 7984 23672
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7380 22976 7432 22982
rect 7380 22918 7432 22924
rect 7392 22778 7420 22918
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7392 22642 7420 22714
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7104 22092 7156 22098
rect 7104 22034 7156 22040
rect 7208 22030 7236 22374
rect 7300 22098 7328 22578
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 7484 22030 7512 22578
rect 7668 22574 7696 23054
rect 7760 22574 7788 23258
rect 7944 23118 7972 23666
rect 8220 23322 8248 24210
rect 8588 24206 8616 26318
rect 9692 25906 9720 26318
rect 10060 25974 10088 26930
rect 10232 26852 10284 26858
rect 10232 26794 10284 26800
rect 10244 26586 10272 26794
rect 10520 26586 10548 26930
rect 10888 26586 10916 27424
rect 10980 26926 11008 28358
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10232 26580 10284 26586
rect 10232 26522 10284 26528
rect 10508 26580 10560 26586
rect 10508 26522 10560 26528
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 9312 25764 9364 25770
rect 9312 25706 9364 25712
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 8864 25226 8892 25638
rect 8852 25220 8904 25226
rect 8852 25162 8904 25168
rect 9324 24818 9352 25706
rect 9692 25294 9720 25842
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9586 24848 9642 24857
rect 8760 24812 8812 24818
rect 8760 24754 8812 24760
rect 9312 24812 9364 24818
rect 9586 24783 9588 24792
rect 9312 24754 9364 24760
rect 9640 24783 9642 24792
rect 9588 24754 9640 24760
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 23594 8616 24142
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8300 23248 8352 23254
rect 8298 23216 8300 23225
rect 8352 23216 8354 23225
rect 8298 23151 8354 23160
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7760 22438 7788 22510
rect 7944 22506 7972 23054
rect 8392 23044 8444 23050
rect 8392 22986 8444 22992
rect 8404 22710 8432 22986
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8392 22704 8444 22710
rect 8392 22646 8444 22652
rect 7932 22500 7984 22506
rect 7932 22442 7984 22448
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 6880 21972 6960 21978
rect 6828 21966 6960 21972
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7840 22024 7892 22030
rect 7840 21966 7892 21972
rect 6840 21950 6960 21966
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6000 21616 6052 21622
rect 6000 21558 6052 21564
rect 6564 21486 6592 21830
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6932 21350 6960 21950
rect 7024 21554 7052 21966
rect 7852 21690 7880 21966
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 8036 21486 8064 22034
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 21554 8156 21966
rect 8496 21962 8524 22714
rect 8680 22642 8708 22918
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8484 21956 8536 21962
rect 8484 21898 8536 21904
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5448 20324 5500 20330
rect 5448 20266 5500 20272
rect 5736 20262 5764 20402
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5736 19990 5764 20198
rect 5828 20058 5856 20538
rect 6092 20528 6144 20534
rect 6092 20470 6144 20476
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 6104 19922 6132 20470
rect 6000 19916 6052 19922
rect 6000 19858 6052 19864
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 5724 19848 5776 19854
rect 5908 19848 5960 19854
rect 5724 19790 5776 19796
rect 5828 19808 5908 19836
rect 5736 19242 5764 19790
rect 5828 19514 5856 19808
rect 5908 19790 5960 19796
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 6012 19378 6040 19858
rect 6104 19514 6132 19858
rect 6380 19786 6408 20946
rect 7576 20874 7604 21286
rect 6644 20868 6696 20874
rect 6644 20810 6696 20816
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 6656 19854 6684 20810
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 8220 19854 8248 20266
rect 8496 20262 8524 21898
rect 8588 21622 8616 21966
rect 8576 21616 8628 21622
rect 8576 21558 8628 21564
rect 8772 20602 8800 24754
rect 9324 24290 9352 24754
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9600 24290 9628 24618
rect 9692 24410 9720 25230
rect 9784 24614 9812 25842
rect 10060 25498 10088 25910
rect 11072 25702 11100 29582
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11256 26450 11284 26726
rect 11336 26580 11388 26586
rect 11336 26522 11388 26528
rect 11244 26444 11296 26450
rect 11244 26386 11296 26392
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 10048 25492 10100 25498
rect 10048 25434 10100 25440
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 10704 24410 10732 24754
rect 11072 24750 11100 25638
rect 11348 24818 11376 26522
rect 11440 25498 11468 27338
rect 11532 26926 11560 28358
rect 11624 28218 11652 28494
rect 11992 28422 12020 31078
rect 12256 30184 12308 30190
rect 12256 30126 12308 30132
rect 12268 28558 12296 30126
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 12256 28552 12308 28558
rect 12308 28512 12388 28540
rect 12256 28494 12308 28500
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11612 28212 11664 28218
rect 11612 28154 11664 28160
rect 11978 28112 12034 28121
rect 12084 28082 12112 28494
rect 12256 28416 12308 28422
rect 12254 28384 12256 28393
rect 12308 28384 12310 28393
rect 12254 28319 12310 28328
rect 12360 28150 12388 28512
rect 12452 28257 12480 29446
rect 12544 29209 12572 36858
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12636 36106 12664 36722
rect 12912 36718 12940 37130
rect 13176 36848 13228 36854
rect 13176 36790 13228 36796
rect 12900 36712 12952 36718
rect 12900 36654 12952 36660
rect 13188 36378 13216 36790
rect 13176 36372 13228 36378
rect 13176 36314 13228 36320
rect 13832 36174 13860 38422
rect 13268 36168 13320 36174
rect 13268 36110 13320 36116
rect 13820 36168 13872 36174
rect 13820 36110 13872 36116
rect 12624 36100 12676 36106
rect 12624 36042 12676 36048
rect 13084 36032 13136 36038
rect 13084 35974 13136 35980
rect 12624 34672 12676 34678
rect 12624 34614 12676 34620
rect 12636 34066 12664 34614
rect 12900 34604 12952 34610
rect 12900 34546 12952 34552
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 12530 29200 12586 29209
rect 12530 29135 12586 29144
rect 12530 29064 12586 29073
rect 12530 28999 12532 29008
rect 12584 28999 12586 29008
rect 12532 28970 12584 28976
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12544 28558 12572 28630
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12532 28416 12584 28422
rect 12532 28358 12584 28364
rect 12438 28248 12494 28257
rect 12544 28218 12572 28358
rect 12438 28183 12494 28192
rect 12532 28212 12584 28218
rect 12348 28144 12400 28150
rect 12348 28086 12400 28092
rect 11978 28047 11980 28056
rect 12032 28047 12034 28056
rect 12072 28076 12124 28082
rect 11980 28018 12032 28024
rect 12072 28018 12124 28024
rect 12084 27674 12112 28018
rect 12072 27668 12124 27674
rect 12072 27610 12124 27616
rect 12256 27532 12308 27538
rect 12256 27474 12308 27480
rect 11520 26920 11572 26926
rect 11520 26862 11572 26868
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11716 25362 11744 26726
rect 12268 26586 12296 27474
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12360 26994 12388 27270
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12254 26480 12310 26489
rect 12452 26450 12480 28183
rect 12532 28154 12584 28160
rect 12636 27470 12664 34002
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12820 33114 12848 33458
rect 12808 33108 12860 33114
rect 12808 33050 12860 33056
rect 12912 32026 12940 34546
rect 12992 34536 13044 34542
rect 12992 34478 13044 34484
rect 13004 34202 13032 34478
rect 12992 34196 13044 34202
rect 12992 34138 13044 34144
rect 12900 32020 12952 32026
rect 12900 31962 12952 31968
rect 12912 30938 12940 31962
rect 12900 30932 12952 30938
rect 12900 30874 12952 30880
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12728 30326 12756 30534
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12992 30184 13044 30190
rect 12992 30126 13044 30132
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 12716 29572 12768 29578
rect 12716 29514 12768 29520
rect 12728 29238 12756 29514
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12716 29028 12768 29034
rect 12716 28970 12768 28976
rect 12728 28558 12756 28970
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12820 28218 12848 28698
rect 12912 28422 12940 29650
rect 13004 29306 13032 30126
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 13096 29170 13124 35974
rect 13280 35494 13308 36110
rect 13268 35488 13320 35494
rect 13268 35430 13320 35436
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 13188 32978 13216 34478
rect 13176 32972 13228 32978
rect 13176 32914 13228 32920
rect 13174 29744 13230 29753
rect 13174 29679 13176 29688
rect 13228 29679 13230 29688
rect 13176 29650 13228 29656
rect 13176 29232 13228 29238
rect 13176 29174 13228 29180
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 13188 28490 13216 29174
rect 13280 29034 13308 35430
rect 14016 35222 14044 39238
rect 14568 38962 14596 39986
rect 14832 39840 14884 39846
rect 14832 39782 14884 39788
rect 15108 39840 15160 39846
rect 15108 39782 15160 39788
rect 14844 39506 14872 39782
rect 14740 39500 14792 39506
rect 14740 39442 14792 39448
rect 14832 39500 14884 39506
rect 14832 39442 14884 39448
rect 14556 38956 14608 38962
rect 14476 38916 14556 38944
rect 14096 38888 14148 38894
rect 14096 38830 14148 38836
rect 14108 38554 14136 38830
rect 14096 38548 14148 38554
rect 14096 38490 14148 38496
rect 14372 38276 14424 38282
rect 14476 38264 14504 38916
rect 14556 38898 14608 38904
rect 14752 38826 14780 39442
rect 15120 39438 15148 39782
rect 15108 39432 15160 39438
rect 15108 39374 15160 39380
rect 15200 39364 15252 39370
rect 15200 39306 15252 39312
rect 15752 39364 15804 39370
rect 15752 39306 15804 39312
rect 15108 39296 15160 39302
rect 15108 39238 15160 39244
rect 14740 38820 14792 38826
rect 14740 38762 14792 38768
rect 14752 38418 14780 38762
rect 15016 38752 15068 38758
rect 15016 38694 15068 38700
rect 14740 38412 14792 38418
rect 14740 38354 14792 38360
rect 14752 38298 14780 38354
rect 15028 38350 15056 38694
rect 14424 38236 14504 38264
rect 14372 38218 14424 38224
rect 14476 37874 14504 38236
rect 14568 38270 14780 38298
rect 15016 38344 15068 38350
rect 15016 38286 15068 38292
rect 14464 37868 14516 37874
rect 14464 37810 14516 37816
rect 14096 37800 14148 37806
rect 14096 37742 14148 37748
rect 14108 37466 14136 37742
rect 14476 37466 14504 37810
rect 14096 37460 14148 37466
rect 14096 37402 14148 37408
rect 14464 37460 14516 37466
rect 14464 37402 14516 37408
rect 14568 37398 14596 38270
rect 14648 38208 14700 38214
rect 14648 38150 14700 38156
rect 14556 37392 14608 37398
rect 14556 37334 14608 37340
rect 14568 37262 14596 37334
rect 14372 37256 14424 37262
rect 14556 37256 14608 37262
rect 14372 37198 14424 37204
rect 14476 37216 14556 37244
rect 14188 36916 14240 36922
rect 14188 36858 14240 36864
rect 14200 35766 14228 36858
rect 14384 36666 14412 37198
rect 14292 36638 14412 36666
rect 14292 36174 14320 36638
rect 14280 36168 14332 36174
rect 14476 36122 14504 37216
rect 14556 37198 14608 37204
rect 14556 37120 14608 37126
rect 14556 37062 14608 37068
rect 14568 36242 14596 37062
rect 14556 36236 14608 36242
rect 14556 36178 14608 36184
rect 14280 36110 14332 36116
rect 14292 35834 14320 36110
rect 14384 36094 14504 36122
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14188 35760 14240 35766
rect 14188 35702 14240 35708
rect 14280 35692 14332 35698
rect 14280 35634 14332 35640
rect 14004 35216 14056 35222
rect 14004 35158 14056 35164
rect 14292 35086 14320 35634
rect 14384 35630 14412 36094
rect 14464 36032 14516 36038
rect 14464 35974 14516 35980
rect 14372 35624 14424 35630
rect 14372 35566 14424 35572
rect 13544 35080 13596 35086
rect 13544 35022 13596 35028
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 13556 33658 13584 35022
rect 13912 34944 13964 34950
rect 13912 34886 13964 34892
rect 13924 34066 13952 34886
rect 14016 34542 14044 35022
rect 14004 34536 14056 34542
rect 14004 34478 14056 34484
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 13544 33652 13596 33658
rect 13544 33594 13596 33600
rect 13452 33312 13504 33318
rect 13452 33254 13504 33260
rect 13464 32910 13492 33254
rect 13832 33046 13860 33934
rect 13912 33108 13964 33114
rect 13912 33050 13964 33056
rect 13820 33040 13872 33046
rect 13820 32982 13872 32988
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13452 32904 13504 32910
rect 13452 32846 13504 32852
rect 13556 32502 13584 32914
rect 13924 32858 13952 33050
rect 14016 32910 14044 34478
rect 14292 34202 14320 35022
rect 14476 34746 14504 35974
rect 14660 35834 14688 38150
rect 15120 38010 15148 39238
rect 15212 38962 15240 39306
rect 15764 39098 15792 39306
rect 15752 39092 15804 39098
rect 15752 39034 15804 39040
rect 15200 38956 15252 38962
rect 15200 38898 15252 38904
rect 15108 38004 15160 38010
rect 15108 37946 15160 37952
rect 15120 37618 15148 37946
rect 15028 37590 15148 37618
rect 14740 37392 14792 37398
rect 14740 37334 14792 37340
rect 14752 36718 14780 37334
rect 15028 37330 15056 37590
rect 15108 37460 15160 37466
rect 15108 37402 15160 37408
rect 15016 37324 15068 37330
rect 15016 37266 15068 37272
rect 15120 36854 15148 37402
rect 15384 37120 15436 37126
rect 15384 37062 15436 37068
rect 15396 36922 15424 37062
rect 15384 36916 15436 36922
rect 15384 36858 15436 36864
rect 15108 36848 15160 36854
rect 15108 36790 15160 36796
rect 14740 36712 14792 36718
rect 14740 36654 14792 36660
rect 15752 36712 15804 36718
rect 15752 36654 15804 36660
rect 15764 36378 15792 36654
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 15660 36100 15712 36106
rect 15660 36042 15712 36048
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 14648 35828 14700 35834
rect 14648 35770 14700 35776
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 15108 35624 15160 35630
rect 15108 35566 15160 35572
rect 15120 35086 15148 35566
rect 15108 35080 15160 35086
rect 15108 35022 15160 35028
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 14936 34202 14964 34546
rect 14280 34196 14332 34202
rect 14280 34138 14332 34144
rect 14924 34196 14976 34202
rect 14924 34138 14976 34144
rect 15120 33998 15148 35022
rect 15212 34950 15240 35634
rect 15304 35630 15332 35974
rect 15476 35692 15528 35698
rect 15476 35634 15528 35640
rect 15292 35624 15344 35630
rect 15292 35566 15344 35572
rect 15304 35154 15332 35566
rect 15488 35290 15516 35634
rect 15672 35494 15700 36042
rect 15660 35488 15712 35494
rect 15660 35430 15712 35436
rect 15476 35284 15528 35290
rect 15476 35226 15528 35232
rect 15292 35148 15344 35154
rect 15292 35090 15344 35096
rect 15672 35086 15700 35430
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 15200 34944 15252 34950
rect 15200 34886 15252 34892
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 15568 34672 15620 34678
rect 15568 34614 15620 34620
rect 15476 34536 15528 34542
rect 15476 34478 15528 34484
rect 15488 34066 15516 34478
rect 15476 34060 15528 34066
rect 15476 34002 15528 34008
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15120 33658 15148 33934
rect 15292 33856 15344 33862
rect 15292 33798 15344 33804
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15304 33318 15332 33798
rect 15488 33522 15516 34002
rect 15476 33516 15528 33522
rect 15476 33458 15528 33464
rect 15292 33312 15344 33318
rect 15292 33254 15344 33260
rect 13832 32830 13952 32858
rect 14004 32904 14056 32910
rect 14004 32846 14056 32852
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 13556 32026 13584 32438
rect 13544 32020 13596 32026
rect 13544 31962 13596 31968
rect 13832 31822 13860 32830
rect 14016 32570 14044 32846
rect 14280 32768 14332 32774
rect 14280 32710 14332 32716
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 13464 30734 13492 31622
rect 13832 31482 13860 31758
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13728 31204 13780 31210
rect 13780 31164 13860 31192
rect 13728 31146 13780 31152
rect 13832 30734 13860 31164
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 13820 30728 13872 30734
rect 13820 30670 13872 30676
rect 14188 30728 14240 30734
rect 14188 30670 14240 30676
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13268 29028 13320 29034
rect 13268 28970 13320 28976
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 12992 28484 13044 28490
rect 12992 28426 13044 28432
rect 13084 28484 13136 28490
rect 13084 28426 13136 28432
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 13004 28218 13032 28426
rect 12808 28212 12860 28218
rect 12808 28154 12860 28160
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 12900 28144 12952 28150
rect 12900 28086 12952 28092
rect 12716 27940 12768 27946
rect 12716 27882 12768 27888
rect 12728 27713 12756 27882
rect 12912 27849 12940 28086
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 13004 27985 13032 28018
rect 12990 27976 13046 27985
rect 12990 27911 13046 27920
rect 12898 27840 12954 27849
rect 12898 27775 12954 27784
rect 12714 27704 12770 27713
rect 12714 27639 12770 27648
rect 12714 27568 12770 27577
rect 12714 27503 12770 27512
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12636 26586 12664 26794
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12254 26415 12310 26424
rect 12440 26444 12492 26450
rect 12268 25702 12296 26415
rect 12440 26386 12492 26392
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 9140 24262 9352 24290
rect 9508 24262 9628 24290
rect 9140 23662 9168 24262
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9324 23798 9352 24006
rect 9312 23792 9364 23798
rect 9312 23734 9364 23740
rect 9508 23730 9536 24262
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9600 23866 9628 24074
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9692 23730 9720 24346
rect 11348 24274 11376 24754
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11440 24070 11468 25162
rect 11796 25152 11848 25158
rect 11796 25094 11848 25100
rect 11808 24886 11836 25094
rect 11796 24880 11848 24886
rect 11796 24822 11848 24828
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23798 11468 24006
rect 11808 23866 11836 24074
rect 11796 23860 11848 23866
rect 11796 23802 11848 23808
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9140 23050 9168 23598
rect 9324 23118 9352 23598
rect 9876 23322 9904 23666
rect 10508 23520 10560 23526
rect 10508 23462 10560 23468
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 10520 23186 10548 23462
rect 11072 23322 11100 23666
rect 12452 23662 12480 25298
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 11072 23118 11100 23258
rect 12452 23186 12480 23598
rect 12728 23254 12756 27503
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 12820 27130 12848 27270
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12820 26518 12848 27066
rect 13096 26994 13124 28426
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 13188 27130 13216 28018
rect 13280 27470 13308 28494
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13372 28121 13400 28358
rect 13358 28112 13414 28121
rect 13358 28047 13414 28056
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 13372 26994 13400 28047
rect 13464 27849 13492 29106
rect 13740 29050 13768 30534
rect 14200 29170 14228 30670
rect 14292 29306 14320 32710
rect 14384 32434 14412 32846
rect 15200 32836 15252 32842
rect 15200 32778 15252 32784
rect 15292 32836 15344 32842
rect 15292 32778 15344 32784
rect 14556 32768 14608 32774
rect 14556 32710 14608 32716
rect 14568 32570 14596 32710
rect 14556 32564 14608 32570
rect 14556 32506 14608 32512
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14372 31136 14424 31142
rect 14372 31078 14424 31084
rect 14384 30802 14412 31078
rect 14476 30938 14504 32370
rect 15212 32026 15240 32778
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 15304 31482 15332 32778
rect 15488 32366 15516 33458
rect 15580 33454 15608 34614
rect 15672 34406 15700 34886
rect 15660 34400 15712 34406
rect 15660 34342 15712 34348
rect 15568 33448 15620 33454
rect 15568 33390 15620 33396
rect 15580 32978 15608 33390
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15844 31816 15896 31822
rect 15844 31758 15896 31764
rect 15292 31476 15344 31482
rect 15292 31418 15344 31424
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15200 31272 15252 31278
rect 15120 31232 15200 31260
rect 14464 30932 14516 30938
rect 14464 30874 14516 30880
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 14372 30796 14424 30802
rect 14372 30738 14424 30744
rect 15028 30258 15056 30874
rect 15120 30666 15148 31232
rect 15200 31214 15252 31220
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 14844 29306 14872 30194
rect 14924 30184 14976 30190
rect 14924 30126 14976 30132
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 13740 29022 13860 29050
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13728 28960 13780 28966
rect 13728 28902 13780 28908
rect 13648 28762 13676 28902
rect 13636 28756 13688 28762
rect 13636 28698 13688 28704
rect 13544 28552 13596 28558
rect 13648 28540 13676 28698
rect 13740 28694 13768 28902
rect 13728 28688 13780 28694
rect 13728 28630 13780 28636
rect 13596 28512 13676 28540
rect 13544 28494 13596 28500
rect 13542 28248 13598 28257
rect 13542 28183 13598 28192
rect 13556 28082 13584 28183
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13636 28076 13688 28082
rect 13636 28018 13688 28024
rect 13450 27840 13506 27849
rect 13450 27775 13506 27784
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 12808 26512 12860 26518
rect 12808 26454 12860 26460
rect 13096 26450 13124 26930
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 13084 26444 13136 26450
rect 13084 26386 13136 26392
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 13096 24886 13124 26250
rect 13188 25362 13216 26862
rect 13648 26450 13676 28018
rect 13740 26586 13768 28630
rect 13832 28490 13860 29022
rect 13912 28960 13964 28966
rect 13912 28902 13964 28908
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13924 28422 13952 28902
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 13912 28416 13964 28422
rect 13818 28384 13874 28393
rect 13912 28358 13964 28364
rect 13818 28319 13874 28328
rect 13728 26580 13780 26586
rect 13728 26522 13780 26528
rect 13636 26444 13688 26450
rect 13636 26386 13688 26392
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13464 25974 13492 26182
rect 13452 25968 13504 25974
rect 13452 25910 13504 25916
rect 13176 25356 13228 25362
rect 13176 25298 13228 25304
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 13096 24138 13124 24822
rect 13372 24614 13400 25094
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13084 24132 13136 24138
rect 13084 24074 13136 24080
rect 13268 24064 13320 24070
rect 13372 24041 13400 24550
rect 13556 24206 13584 24550
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13268 24006 13320 24012
rect 13358 24032 13414 24041
rect 13280 23866 13308 24006
rect 13358 23967 13414 23976
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 13740 23730 13768 24686
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13740 23322 13768 23666
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 9128 23044 9180 23050
rect 9128 22986 9180 22992
rect 9140 22778 9168 22986
rect 9128 22772 9180 22778
rect 9128 22714 9180 22720
rect 9324 22710 9352 23054
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9312 22704 9364 22710
rect 9312 22646 9364 22652
rect 9324 22234 9352 22646
rect 9784 22574 9812 22714
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9312 22228 9364 22234
rect 9312 22170 9364 22176
rect 9784 22030 9812 22510
rect 11164 22438 11192 23054
rect 11428 22976 11480 22982
rect 11428 22918 11480 22924
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11440 22642 11468 22918
rect 11900 22710 11928 22918
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 11152 22432 11204 22438
rect 11152 22374 11204 22380
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21554 10548 21830
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5460 17814 5488 19178
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 5828 18766 5856 19110
rect 6196 18902 6224 19110
rect 6288 18970 6316 19654
rect 6380 19378 6408 19722
rect 6656 19496 6684 19790
rect 8312 19514 8340 19858
rect 8300 19508 8352 19514
rect 6656 19468 6868 19496
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6656 18970 6684 19314
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4724 16114 4752 16934
rect 4816 16590 4844 17138
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 16250 4844 16526
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 5276 15910 5304 17138
rect 5368 16794 5396 17546
rect 5460 17134 5488 17750
rect 5552 17338 5580 18158
rect 5644 17746 5672 18566
rect 5736 18358 5764 18702
rect 5724 18352 5776 18358
rect 5724 18294 5776 18300
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5736 17882 5764 18158
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5828 17762 5856 18702
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5736 17746 5856 17762
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5724 17740 5856 17746
rect 5776 17734 5856 17740
rect 5724 17682 5776 17688
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5644 16998 5672 17546
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5368 16046 5396 16458
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14006 4016 14350
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 4632 13802 4660 14282
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4080 12918 4108 13466
rect 4632 13258 4660 13738
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3988 11540 4016 12786
rect 4080 11744 4108 12854
rect 4356 12764 4384 13126
rect 4632 12986 4660 13194
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12918 4752 13670
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4712 12776 4764 12782
rect 4356 12736 4712 12764
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12736
rect 4712 12718 4764 12724
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4724 12322 4752 12582
rect 4632 12306 4752 12322
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4620 12300 4752 12306
rect 4672 12294 4752 12300
rect 4620 12242 4672 12248
rect 4160 12096 4212 12102
rect 4160 12038 4212 12044
rect 4172 11898 4200 12038
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4250 11792 4306 11801
rect 4160 11756 4212 11762
rect 4080 11716 4160 11744
rect 4250 11727 4306 11736
rect 4160 11698 4212 11704
rect 4264 11558 4292 11727
rect 4356 11626 4384 12242
rect 4632 11914 4660 12242
rect 5276 12170 5304 15846
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 4540 11886 4660 11914
rect 4434 11656 4490 11665
rect 4344 11620 4396 11626
rect 4434 11591 4490 11600
rect 4344 11562 4396 11568
rect 4448 11558 4476 11591
rect 4252 11552 4304 11558
rect 3988 11512 4252 11540
rect 4080 11286 4108 11512
rect 4252 11494 4304 11500
rect 4436 11552 4488 11558
rect 4540 11540 4568 11886
rect 4710 11792 4766 11801
rect 4710 11727 4712 11736
rect 4764 11727 4766 11736
rect 4712 11698 4764 11704
rect 4540 11512 4660 11540
rect 4436 11494 4488 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9586 1440 10542
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2700 9586 2728 10066
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 1412 8430 1440 9522
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 1412 7954 1440 8366
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 2332 7410 2360 8026
rect 2700 7546 2728 8366
rect 2976 7818 3004 10678
rect 3436 10266 3464 11018
rect 3896 10810 3924 11086
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4632 10674 4660 11512
rect 4816 11082 4844 12106
rect 5356 12096 5408 12102
rect 5276 12044 5356 12050
rect 5276 12038 5408 12044
rect 5276 12022 5396 12038
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 5276 11014 5304 12022
rect 5354 11792 5410 11801
rect 5354 11727 5410 11736
rect 5368 11694 5396 11727
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3436 9722 3464 10202
rect 4632 9994 4660 10610
rect 5368 10538 5396 11630
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5460 10062 5488 14214
rect 5644 13530 5672 16934
rect 5736 16522 5764 17478
rect 5920 17202 5948 18294
rect 6196 18290 6224 18838
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 6196 17270 6224 18226
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6196 16998 6224 17206
rect 6472 17202 6500 17478
rect 6564 17338 6592 17614
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5736 14074 5764 15506
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5828 15162 5856 15438
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5828 14618 5856 14894
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 6196 13938 6224 15098
rect 6380 14958 6408 17070
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6380 14226 6408 14894
rect 6472 14346 6500 15506
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 14958 6684 15302
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6564 14226 6592 14282
rect 6380 14198 6592 14226
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6012 12306 6040 13466
rect 6380 12714 6408 13806
rect 6564 13462 6592 14198
rect 6656 13938 6684 14554
rect 6748 14074 6776 15438
rect 6840 15162 6868 19468
rect 8300 19450 8352 19456
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7208 17338 7236 17750
rect 7300 17746 7328 18022
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7576 16998 7604 17818
rect 7668 17202 7696 18090
rect 7760 17542 7788 19110
rect 8036 18630 8064 19314
rect 8312 18698 8340 19450
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8680 18834 8708 19178
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 9600 18766 9628 20198
rect 9968 20058 9996 20334
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9692 18834 9720 19382
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9588 18760 9640 18766
rect 9586 18728 9588 18737
rect 9640 18728 9642 18737
rect 8300 18692 8352 18698
rect 9586 18663 9642 18672
rect 9680 18692 9732 18698
rect 8300 18634 8352 18640
rect 9680 18634 9732 18640
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7852 17898 7880 18226
rect 8036 18086 8064 18566
rect 9600 18290 9628 18566
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7852 17882 8064 17898
rect 7852 17876 8076 17882
rect 7852 17870 8024 17876
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7852 17202 7880 17870
rect 8024 17818 8076 17824
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7668 17066 7696 17138
rect 8312 17134 8340 18226
rect 8772 17814 8800 18226
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 9140 17270 9168 18022
rect 9416 17678 9444 18158
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9508 17678 9536 17750
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9600 17610 9628 18226
rect 9692 17882 9720 18634
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9680 17536 9732 17542
rect 9784 17524 9812 18906
rect 9968 18766 9996 19994
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10152 18970 10180 19382
rect 10336 19378 10364 20334
rect 10508 19984 10560 19990
rect 10508 19926 10560 19932
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10336 18970 10364 19314
rect 10520 19122 10548 19926
rect 10612 19854 10640 20402
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10704 19854 10732 20198
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10612 19334 10640 19790
rect 10796 19446 10824 20198
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10612 19310 10732 19334
rect 10612 19306 10744 19310
rect 10692 19304 10744 19306
rect 10692 19246 10744 19252
rect 10520 19094 10640 19122
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18834 10364 18906
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9876 17678 9904 18226
rect 9968 18222 9996 18702
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10060 18426 10088 18566
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9968 17678 9996 18158
rect 10152 18154 10180 18566
rect 10508 18284 10560 18290
rect 10508 18226 10560 18232
rect 10140 18148 10192 18154
rect 10140 18090 10192 18096
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9784 17496 9996 17524
rect 9680 17478 9732 17484
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8680 17066 8708 17138
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16794 7604 16934
rect 8772 16794 8800 17070
rect 9416 16998 9444 17478
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16794 9444 16934
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 6932 16250 6960 16526
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 7392 14414 7420 16526
rect 8772 16114 8800 16730
rect 9508 16590 9536 17138
rect 9692 17134 9720 17478
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9876 16454 9904 17206
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14482 8156 14758
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6656 13258 6684 13874
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13410 6960 13670
rect 7116 13530 7144 14010
rect 7760 14006 7788 14214
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 6748 13394 6960 13410
rect 6736 13388 6960 13394
rect 6788 13382 6960 13388
rect 6736 13330 6788 13336
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6840 12986 6868 13262
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6932 12850 6960 13382
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7116 12782 7144 13466
rect 7392 13326 7420 13738
rect 8128 13530 8156 14418
rect 8496 14414 8524 15438
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 9232 14278 9260 15438
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14464 9720 14758
rect 9876 14618 9904 15302
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9646 14436 9720 14464
rect 9496 14408 9548 14414
rect 9646 14396 9674 14436
rect 9968 14414 9996 17496
rect 10060 15502 10088 17818
rect 10152 17678 10180 18090
rect 10520 17882 10548 18226
rect 10612 17882 10640 19094
rect 10704 18766 10732 19246
rect 10980 18834 11008 20810
rect 11164 18970 11192 21082
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11348 20534 11376 20742
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 11532 20466 11560 22578
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 21010 11928 21966
rect 12912 21962 12940 22578
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12900 21956 12952 21962
rect 12900 21898 12952 21904
rect 12176 21690 12204 21898
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12912 21622 12940 21898
rect 12900 21616 12952 21622
rect 12900 21558 12952 21564
rect 13004 21486 13032 23122
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13280 22778 13308 22918
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 13832 22094 13860 28319
rect 13924 28082 13952 28358
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13910 27976 13966 27985
rect 13910 27911 13966 27920
rect 13924 27878 13952 27911
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13910 27704 13966 27713
rect 13910 27639 13966 27648
rect 13924 27062 13952 27639
rect 14016 27606 14044 28018
rect 14004 27600 14056 27606
rect 14004 27542 14056 27548
rect 14108 27538 14136 28494
rect 14200 27606 14228 29106
rect 14464 28484 14516 28490
rect 14464 28426 14516 28432
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 14096 27532 14148 27538
rect 14096 27474 14148 27480
rect 13912 27056 13964 27062
rect 13912 26998 13964 27004
rect 14108 26926 14136 27474
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 14108 25838 14136 26862
rect 14200 26586 14228 26930
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 14384 25430 14412 27950
rect 14476 25838 14504 28426
rect 14936 28150 14964 30126
rect 15120 28994 15148 30602
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15212 30258 15240 30534
rect 15304 30394 15332 31418
rect 15292 30388 15344 30394
rect 15292 30330 15344 30336
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15304 30054 15332 30194
rect 15292 30048 15344 30054
rect 15292 29990 15344 29996
rect 15396 29238 15424 31418
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15488 30190 15516 31146
rect 15660 31136 15712 31142
rect 15752 31136 15804 31142
rect 15660 31078 15712 31084
rect 15750 31104 15752 31113
rect 15804 31104 15806 31113
rect 15672 30802 15700 31078
rect 15750 31039 15806 31048
rect 15856 30938 15884 31758
rect 15948 31482 15976 42162
rect 16408 41614 16436 42570
rect 16580 42288 16632 42294
rect 16580 42230 16632 42236
rect 16396 41608 16448 41614
rect 16396 41550 16448 41556
rect 16408 41414 16436 41550
rect 16592 41478 16620 42230
rect 17512 42226 17540 42842
rect 19064 42696 19116 42702
rect 19064 42638 19116 42644
rect 18144 42560 18196 42566
rect 18144 42502 18196 42508
rect 18156 42294 18184 42502
rect 18788 42356 18840 42362
rect 18788 42298 18840 42304
rect 18144 42288 18196 42294
rect 18144 42230 18196 42236
rect 17500 42220 17552 42226
rect 17500 42162 17552 42168
rect 18800 41682 18828 42298
rect 18788 41676 18840 41682
rect 18788 41618 18840 41624
rect 17408 41540 17460 41546
rect 17408 41482 17460 41488
rect 16580 41472 16632 41478
rect 16580 41414 16632 41420
rect 16316 41386 16436 41414
rect 16316 40050 16344 41386
rect 16592 41070 16620 41414
rect 17040 41200 17092 41206
rect 17040 41142 17092 41148
rect 16580 41064 16632 41070
rect 16580 41006 16632 41012
rect 16028 40044 16080 40050
rect 16028 39986 16080 39992
rect 16304 40044 16356 40050
rect 16304 39986 16356 39992
rect 16040 38962 16068 39986
rect 16316 39370 16344 39986
rect 16304 39364 16356 39370
rect 16304 39306 16356 39312
rect 16028 38956 16080 38962
rect 16028 38898 16080 38904
rect 16212 37188 16264 37194
rect 16212 37130 16264 37136
rect 16224 36650 16252 37130
rect 16304 36712 16356 36718
rect 16304 36654 16356 36660
rect 16212 36644 16264 36650
rect 16212 36586 16264 36592
rect 16316 36242 16344 36654
rect 16304 36236 16356 36242
rect 16304 36178 16356 36184
rect 16592 35986 16620 41006
rect 17052 40526 17080 41142
rect 17420 40730 17448 41482
rect 18328 41472 18380 41478
rect 18328 41414 18380 41420
rect 17592 41200 17644 41206
rect 17592 41142 17644 41148
rect 17604 41041 17632 41142
rect 17960 41132 18012 41138
rect 17960 41074 18012 41080
rect 17590 41032 17646 41041
rect 17590 40967 17646 40976
rect 17500 40928 17552 40934
rect 17500 40870 17552 40876
rect 17512 40730 17540 40870
rect 17132 40724 17184 40730
rect 17132 40666 17184 40672
rect 17408 40724 17460 40730
rect 17408 40666 17460 40672
rect 17500 40724 17552 40730
rect 17500 40666 17552 40672
rect 17144 40610 17172 40666
rect 17512 40610 17540 40666
rect 17144 40582 17264 40610
rect 17420 40594 17540 40610
rect 17040 40520 17092 40526
rect 17040 40462 17092 40468
rect 17052 39982 17080 40462
rect 17132 40044 17184 40050
rect 17132 39986 17184 39992
rect 17040 39976 17092 39982
rect 17040 39918 17092 39924
rect 17144 39506 17172 39986
rect 17132 39500 17184 39506
rect 17132 39442 17184 39448
rect 17144 39302 17172 39442
rect 17132 39296 17184 39302
rect 17132 39238 17184 39244
rect 17132 38888 17184 38894
rect 17132 38830 17184 38836
rect 16856 37868 16908 37874
rect 16856 37810 16908 37816
rect 16868 36922 16896 37810
rect 16856 36916 16908 36922
rect 16856 36858 16908 36864
rect 16672 36576 16724 36582
rect 16672 36518 16724 36524
rect 16684 36174 16712 36518
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16868 36106 16896 36178
rect 16856 36100 16908 36106
rect 16856 36042 16908 36048
rect 16592 35958 16712 35986
rect 16580 35624 16632 35630
rect 16580 35566 16632 35572
rect 16028 35488 16080 35494
rect 16028 35430 16080 35436
rect 16040 34746 16068 35430
rect 16592 35290 16620 35566
rect 16580 35284 16632 35290
rect 16580 35226 16632 35232
rect 16488 35012 16540 35018
rect 16488 34954 16540 34960
rect 16500 34746 16528 34954
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 16488 34740 16540 34746
rect 16488 34682 16540 34688
rect 16028 34400 16080 34406
rect 16028 34342 16080 34348
rect 16040 33998 16068 34342
rect 16028 33992 16080 33998
rect 16028 33934 16080 33940
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 16132 33658 16160 33798
rect 16120 33652 16172 33658
rect 16120 33594 16172 33600
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16500 33114 16528 33458
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16028 32292 16080 32298
rect 16028 32234 16080 32240
rect 16040 32026 16068 32234
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 15936 31476 15988 31482
rect 15936 31418 15988 31424
rect 15844 30932 15896 30938
rect 15844 30874 15896 30880
rect 15660 30796 15712 30802
rect 15660 30738 15712 30744
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15476 30184 15528 30190
rect 15476 30126 15528 30132
rect 15580 30122 15608 30670
rect 15672 30394 15700 30738
rect 15660 30388 15712 30394
rect 15660 30330 15712 30336
rect 15752 30320 15804 30326
rect 15752 30262 15804 30268
rect 15568 30116 15620 30122
rect 15568 30058 15620 30064
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15292 29096 15344 29102
rect 15292 29038 15344 29044
rect 15028 28966 15148 28994
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14568 27849 14596 28018
rect 14648 27872 14700 27878
rect 14554 27840 14610 27849
rect 14648 27814 14700 27820
rect 14554 27775 14610 27784
rect 14568 26382 14596 27775
rect 14660 27062 14688 27814
rect 14936 27674 14964 28086
rect 14924 27668 14976 27674
rect 14924 27610 14976 27616
rect 15028 27554 15056 28966
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15212 28200 15240 28358
rect 15120 28172 15240 28200
rect 15120 27826 15148 28172
rect 15198 28112 15254 28121
rect 15198 28047 15200 28056
rect 15252 28047 15254 28056
rect 15200 28018 15252 28024
rect 15120 27798 15240 27826
rect 14936 27526 15056 27554
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14648 27056 14700 27062
rect 14648 26998 14700 27004
rect 14752 26382 14780 27270
rect 14936 26790 14964 27526
rect 15212 27062 15240 27798
rect 15200 27056 15252 27062
rect 15200 26998 15252 27004
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 15212 26602 15240 26998
rect 15120 26574 15240 26602
rect 14556 26376 14608 26382
rect 14740 26376 14792 26382
rect 14608 26336 14688 26364
rect 14556 26318 14608 26324
rect 14464 25832 14516 25838
rect 14464 25774 14516 25780
rect 14372 25424 14424 25430
rect 14372 25366 14424 25372
rect 14556 25152 14608 25158
rect 14556 25094 14608 25100
rect 14568 24886 14596 25094
rect 14556 24880 14608 24886
rect 14556 24822 14608 24828
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14016 23730 14044 24006
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13832 22066 14228 22094
rect 13912 21956 13964 21962
rect 13912 21898 13964 21904
rect 13924 21690 13952 21898
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 14200 21622 14228 22066
rect 14188 21616 14240 21622
rect 14188 21558 14240 21564
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 12164 20868 12216 20874
rect 12164 20810 12216 20816
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11624 19718 11652 20402
rect 12176 20058 12204 20810
rect 13004 20466 13032 21422
rect 13832 21010 13860 21422
rect 14096 21344 14148 21350
rect 14096 21286 14148 21292
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13832 20534 13860 20946
rect 14108 20602 14136 21286
rect 14568 20602 14596 21490
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11244 18896 11296 18902
rect 11244 18838 11296 18844
rect 10968 18828 11020 18834
rect 10888 18788 10968 18816
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10244 17678 10272 17750
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10612 17134 10640 17818
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10704 17338 10732 17614
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 9548 14368 9674 14396
rect 9496 14350 9548 14356
rect 9646 14328 9674 14368
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 9705 14340 9757 14346
rect 9646 14300 9705 14328
rect 9692 14288 9705 14300
rect 9692 14282 9757 14288
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8404 13326 8432 13670
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 7300 12850 7328 13262
rect 7392 12918 7420 13262
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 7116 12646 7144 12718
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12442 7144 12582
rect 7104 12436 7156 12442
rect 6932 12406 7104 12434
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 10266 5580 12174
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11218 5672 11494
rect 5736 11286 5764 12038
rect 6932 11762 6960 12406
rect 7104 12378 7156 12384
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6736 11688 6788 11694
rect 6734 11656 6736 11665
rect 6788 11656 6790 11665
rect 6734 11591 6790 11600
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3252 9042 3280 9590
rect 5276 9586 5304 9862
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5460 9178 5488 9590
rect 5552 9382 5580 9998
rect 5632 9580 5684 9586
rect 5736 9568 5764 11222
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5828 10810 5856 10950
rect 6104 10810 6132 11086
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 5684 9540 5764 9568
rect 5632 9522 5684 9528
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 3240 9036 3292 9042
rect 3240 8978 3292 8984
rect 3252 8566 3280 8978
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3620 8498 3648 8774
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 7993 3740 8366
rect 3804 8362 3832 8434
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3698 7984 3754 7993
rect 3698 7919 3754 7928
rect 3896 7868 3924 9114
rect 5552 8974 5580 9318
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3804 7840 3924 7868
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2332 5846 2360 7346
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2700 5710 2728 7346
rect 2976 6662 3004 7754
rect 3620 7342 3648 7754
rect 3804 7750 3832 7840
rect 3988 7818 4016 8502
rect 4080 8362 4108 8910
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 7886 4108 8298
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 3988 7528 4016 7754
rect 3804 7500 4016 7528
rect 3804 7410 3832 7500
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3896 7290 3924 7500
rect 3976 7404 4028 7410
rect 4080 7392 4108 7822
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4172 7478 4200 7686
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4028 7364 4108 7392
rect 4252 7404 4304 7410
rect 3976 7346 4028 7352
rect 4448 7392 4476 8026
rect 4526 7984 4582 7993
rect 4632 7954 4660 8910
rect 4526 7919 4582 7928
rect 4620 7948 4672 7954
rect 4540 7886 4568 7919
rect 4620 7890 4672 7896
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7546 4568 7822
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4632 7478 4660 7686
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 4528 7404 4580 7410
rect 4448 7364 4528 7392
rect 4252 7346 4304 7352
rect 4528 7346 4580 7352
rect 4264 7290 4292 7346
rect 3896 7262 4292 7290
rect 4540 7206 4568 7346
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 7002 4660 7414
rect 4724 7274 4752 8910
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 7954 4844 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4908 7750 4936 8366
rect 5552 8362 5580 8910
rect 5644 8634 5672 9386
rect 5736 8838 5764 9540
rect 6012 9178 6040 9590
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6012 8974 6040 9114
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7410 5304 7686
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4908 7002 4936 7142
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2148 5166 2176 5646
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1412 4826 1440 5102
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 2240 3738 2268 5170
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2424 4554 2452 4762
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2700 4486 2728 5646
rect 2792 5166 2820 5646
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2976 4554 3004 5510
rect 3528 5302 3556 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3528 4826 3556 5238
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3804 4622 3832 4966
rect 3896 4690 3924 5238
rect 4172 5012 4200 5510
rect 4264 5030 4292 5510
rect 4356 5370 4384 5646
rect 4448 5642 4476 5850
rect 5276 5846 5304 7142
rect 5264 5840 5316 5846
rect 4724 5766 5028 5794
rect 5264 5782 5316 5788
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4356 5166 4384 5306
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 4448 5030 4476 5578
rect 4724 5166 4752 5766
rect 4896 5704 4948 5710
rect 4816 5664 4896 5692
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4080 4984 4200 5012
rect 4252 5024 4304 5030
rect 4080 4826 4108 4984
rect 4252 4966 4304 4972
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3058 3188 3538
rect 3252 3534 3280 3878
rect 3528 3534 3556 3946
rect 3896 3602 3924 4626
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4264 4026 4292 4558
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4146 4384 4422
rect 4448 4162 4476 4490
rect 4632 4282 4660 5034
rect 4724 4758 4752 5102
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4816 4622 4844 5664
rect 4896 5646 4948 5652
rect 5000 5642 5028 5766
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4690 4936 4966
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 5276 4622 5304 5646
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4804 4616 4856 4622
rect 4724 4576 4804 4604
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4724 4214 4752 4576
rect 4804 4558 4856 4564
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4712 4208 4764 4214
rect 4344 4140 4396 4146
rect 4448 4134 4660 4162
rect 4712 4150 4764 4156
rect 4344 4082 4396 4088
rect 4632 4078 4660 4134
rect 4724 4078 4752 4150
rect 4816 4078 4844 4422
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5368 4282 5396 4966
rect 5460 4826 5488 8230
rect 5644 7886 5672 8298
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7342 5672 7822
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5552 4622 5580 5102
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 4528 4072 4580 4078
rect 4264 4020 4528 4026
rect 4264 4014 4580 4020
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4264 3998 4568 4014
rect 4540 3942 4568 3998
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3618 4660 4014
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 4540 3590 4660 3618
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 3126 3464 3334
rect 4172 3194 4200 3402
rect 4540 3398 4568 3590
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 4724 3058 4752 3674
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4816 2990 4844 4014
rect 4908 3738 4936 4014
rect 5276 3738 5304 4150
rect 5448 4140 5500 4146
rect 5644 4128 5672 7278
rect 5736 5914 5764 8434
rect 6104 8090 6132 10746
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6196 9178 6224 10202
rect 6288 10062 6316 10406
rect 6656 10198 6684 11290
rect 6748 10742 6776 11591
rect 6932 11150 6960 11698
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 7024 10742 7052 11766
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7116 11150 7144 11494
rect 7208 11218 7236 11494
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6656 9994 6684 10134
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9518 6592 9862
rect 6656 9722 6684 9930
rect 6840 9926 6868 10542
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6472 8498 6500 8774
rect 6656 8634 6684 9454
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6840 8566 6868 9862
rect 6932 8634 6960 9930
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7024 8566 7052 10202
rect 7116 9722 7144 10202
rect 7208 10130 7236 11154
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7116 8974 7144 9658
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6104 7886 6132 8026
rect 6656 7954 6684 8230
rect 6840 8090 6868 8502
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6932 7818 6960 8366
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 6012 5302 6040 6802
rect 6104 6730 6132 6870
rect 6380 6798 6408 7278
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6564 6730 6592 7686
rect 7024 6798 7052 8298
rect 7208 7818 7236 8434
rect 7196 7812 7248 7818
rect 7116 7772 7196 7800
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6840 6254 6868 6734
rect 7116 6730 7144 7772
rect 7196 7754 7248 7760
rect 7300 7562 7328 12106
rect 7576 11762 7604 13126
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11286 7604 11698
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7668 11098 7696 13126
rect 8680 12918 8708 13262
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 9232 12102 9260 14214
rect 9692 12730 9720 14282
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13190 10088 14214
rect 10244 14006 10272 15098
rect 10324 14884 10376 14890
rect 10324 14826 10376 14832
rect 10336 14618 10364 14826
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10428 14550 10456 16934
rect 10888 16182 10916 18788
rect 10968 18770 11020 18776
rect 11256 18766 11284 18838
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 10968 18624 11020 18630
rect 11020 18572 11100 18578
rect 10968 18566 11100 18572
rect 10980 18550 11100 18566
rect 11072 18086 11100 18550
rect 11440 18222 11468 19246
rect 11624 19242 11652 19654
rect 12268 19242 12296 19790
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12360 19310 12388 19654
rect 12912 19514 12940 20198
rect 13832 19922 13860 20470
rect 14108 20398 14136 20538
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 11624 18698 11652 19178
rect 11900 18970 11928 19178
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11624 18222 11652 18634
rect 11716 18222 11744 18906
rect 12084 18698 12112 19110
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18358 12020 18566
rect 11980 18352 12032 18358
rect 11980 18294 12032 18300
rect 11428 18216 11480 18222
rect 11612 18216 11664 18222
rect 11480 18176 11560 18204
rect 11428 18158 11480 18164
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11532 17746 11560 18176
rect 11612 18158 11664 18164
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 10888 15570 10916 16118
rect 11348 15978 11376 16526
rect 11532 16046 11560 17682
rect 11716 17610 11744 18158
rect 12176 17814 12204 18906
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 18290 12296 18566
rect 12360 18426 12388 19246
rect 12452 18902 12480 19450
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12532 18760 12584 18766
rect 12530 18728 12532 18737
rect 12584 18728 12586 18737
rect 12530 18663 12586 18672
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 13096 18222 13124 19110
rect 13832 18970 13860 19246
rect 13924 19242 13952 19722
rect 14108 19718 14136 20334
rect 14384 20262 14412 20402
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18290 13216 18566
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12164 17808 12216 17814
rect 12164 17750 12216 17756
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 12912 17202 12940 18022
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13464 17338 13492 17614
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 14016 17202 14044 17818
rect 14108 17678 14136 18362
rect 14568 18086 14596 18702
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16794 13860 17002
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11348 15706 11376 15914
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11440 15706 11468 15846
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11072 15026 11100 15302
rect 11164 15162 11192 15302
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11532 15026 11560 15982
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11716 15502 11744 15642
rect 11992 15502 12020 16458
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12176 15570 12204 16118
rect 12728 15978 12756 16730
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 15972 12768 15978
rect 12716 15914 12768 15920
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12268 15502 12296 15846
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 11992 15366 12020 15438
rect 12728 15434 12756 15914
rect 12820 15586 12848 16594
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13832 16454 13860 16526
rect 13924 16522 13952 16934
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13188 16114 13216 16390
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 12912 15706 12940 16050
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12820 15558 12940 15586
rect 12912 15502 12940 15558
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 15162 12112 15302
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11348 14618 11376 14962
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10336 14278 10364 14350
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10244 13258 10272 13942
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9864 12912 9916 12918
rect 9916 12860 9996 12866
rect 9864 12854 9996 12860
rect 9772 12844 9824 12850
rect 9876 12838 9996 12854
rect 9772 12786 9824 12792
rect 9600 12702 9720 12730
rect 9784 12730 9812 12786
rect 9784 12702 9904 12730
rect 9600 12458 9628 12702
rect 9680 12640 9732 12646
rect 9732 12588 9812 12594
rect 9680 12582 9812 12588
rect 9692 12566 9812 12582
rect 9600 12430 9720 12458
rect 9692 12102 9720 12430
rect 9784 12238 9812 12566
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7760 11150 7788 11562
rect 7392 11082 7696 11098
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7380 11076 7696 11082
rect 7432 11070 7696 11076
rect 7380 11018 7432 11024
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10674 7604 10950
rect 7760 10810 7788 11086
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7392 9926 7420 10474
rect 7484 10198 7512 10542
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 8022 7420 9862
rect 7484 9636 7512 9998
rect 7564 9648 7616 9654
rect 7484 9608 7564 9636
rect 7564 9590 7616 9596
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7208 7534 7328 7562
rect 7208 7478 7236 7534
rect 7196 7472 7248 7478
rect 7248 7420 7328 7426
rect 7196 7414 7328 7420
rect 7208 7398 7328 7414
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7208 6798 7236 7278
rect 7300 6934 7328 7398
rect 7392 7342 7420 7822
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5302 6592 5510
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6840 5030 6868 6190
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5500 4100 5672 4128
rect 5448 4082 5500 4088
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5276 3126 5304 3674
rect 5368 3126 5396 3878
rect 5460 3534 5488 3946
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5552 3058 5580 3538
rect 5920 3466 5948 4694
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 3194 5948 3402
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6840 3058 6868 4966
rect 6932 3466 6960 5510
rect 7024 4826 7052 5646
rect 7300 5302 7328 6870
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7300 4758 7328 5238
rect 7392 5030 7420 5646
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7392 4622 7420 4966
rect 7484 4826 7512 8978
rect 7668 7750 7696 10746
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 9994 7880 10406
rect 7944 10112 7972 10950
rect 8128 10810 8156 11018
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8024 10124 8076 10130
rect 7944 10084 8024 10112
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7852 9722 7880 9930
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7944 9586 7972 10084
rect 8024 10066 8076 10072
rect 8128 10062 8156 10746
rect 9324 10130 9352 12038
rect 9600 11694 9628 12038
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9600 11529 9628 11630
rect 9692 11558 9720 12038
rect 9784 11830 9812 12174
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9680 11552 9732 11558
rect 9586 11520 9642 11529
rect 9680 11494 9732 11500
rect 9586 11455 9642 11464
rect 9588 11280 9640 11286
rect 9416 11240 9588 11268
rect 9416 11150 9444 11240
rect 9588 11222 9640 11228
rect 9496 11154 9548 11160
rect 9404 11144 9456 11150
rect 9876 11150 9904 12702
rect 9968 12186 9996 12838
rect 10060 12306 10088 13126
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10152 12442 10180 12786
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10244 12238 10272 12582
rect 10428 12434 10456 14486
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10704 13530 10732 13806
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10336 12406 10456 12434
rect 10232 12232 10284 12238
rect 9968 12158 10088 12186
rect 10232 12174 10284 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9968 11762 9996 12038
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9772 11144 9824 11150
rect 9600 11121 9772 11132
rect 9496 11096 9548 11102
rect 9586 11112 9772 11121
rect 9404 11086 9456 11092
rect 9508 10996 9536 11096
rect 9642 11104 9772 11112
rect 9772 11086 9824 11092
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9586 11047 9642 11056
rect 9634 11008 9686 11014
rect 9508 10968 9634 10996
rect 9634 10950 9686 10956
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10130 9628 10406
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 9784 9926 9812 10950
rect 9968 10742 9996 11290
rect 10060 10962 10088 12158
rect 10232 11008 10284 11014
rect 10060 10956 10232 10962
rect 10060 10950 10284 10956
rect 10060 10934 10272 10950
rect 10060 10810 10088 10934
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9956 10736 10008 10742
rect 9956 10678 10008 10684
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9876 10266 9904 10542
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 8036 9654 8064 9862
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 9784 9518 9812 9862
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 8312 8498 8340 9318
rect 9692 8906 9720 9318
rect 10244 8906 10272 10934
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8208 8424 8260 8430
rect 8260 8372 8340 8378
rect 8208 8366 8340 8372
rect 8220 8350 8340 8366
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7840 8016 7892 8022
rect 7838 7984 7840 7993
rect 7892 7984 7894 7993
rect 7838 7919 7894 7928
rect 7840 7880 7892 7886
rect 7838 7848 7840 7857
rect 7892 7848 7894 7857
rect 7838 7783 7894 7792
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 8036 7410 8064 8026
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8128 7546 8156 7686
rect 8220 7546 8248 8230
rect 8312 7886 8340 8350
rect 8680 8090 8708 8502
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8300 7880 8352 7886
rect 8298 7848 8300 7857
rect 8352 7848 8354 7857
rect 8298 7783 8354 7792
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8312 6458 8340 7783
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8680 5574 8708 7142
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7484 4554 7512 4762
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 8312 4146 8340 4694
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8588 4146 8616 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 7944 3126 7972 3946
rect 8680 3534 8708 4082
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8772 2446 8800 8366
rect 9048 8090 9076 8434
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9034 7984 9090 7993
rect 9034 7919 9036 7928
rect 9088 7919 9090 7928
rect 9036 7890 9088 7896
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8864 5710 8892 7414
rect 9232 7206 9260 7822
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9140 6798 9168 7142
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8956 5914 8984 6734
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6186 9076 6598
rect 9036 6180 9088 6186
rect 9036 6122 9088 6128
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9232 5778 9260 7142
rect 9324 7002 9352 7822
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9508 6746 9536 7414
rect 9600 6866 9628 7686
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9508 6730 9628 6746
rect 9508 6724 9640 6730
rect 9508 6718 9588 6724
rect 9588 6666 9640 6672
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5914 9536 6190
rect 9600 6118 9628 6666
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5914 9628 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9600 5794 9628 5850
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9416 5766 9628 5794
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8864 5302 8892 5646
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8864 4690 8892 5238
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8864 4554 8892 4626
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 9140 4282 9168 5170
rect 9232 5114 9260 5714
rect 9416 5642 9444 5766
rect 9496 5704 9548 5710
rect 9692 5658 9720 6258
rect 9784 5710 9812 6598
rect 9876 6118 9904 6938
rect 10244 6730 10272 8842
rect 10336 8362 10364 12406
rect 10612 12306 10640 12854
rect 10704 12850 10732 13466
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12986 11192 13126
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11898 10548 12174
rect 10704 12102 10732 12786
rect 11440 12424 11468 14282
rect 11992 13938 12020 14554
rect 12084 14414 12112 15098
rect 12912 14822 12940 15438
rect 13280 15434 13308 15914
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13924 15026 13952 15506
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 12912 14482 12940 14758
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 13740 13938 13768 14214
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12782 11560 13194
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11520 12436 11572 12442
rect 11440 12396 11520 12424
rect 11900 12434 11928 13874
rect 11992 12782 12020 13874
rect 12440 13184 12492 13190
rect 12544 13172 12572 13874
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13190 12756 13738
rect 12492 13144 12572 13172
rect 12716 13184 12768 13190
rect 12440 13126 12492 13132
rect 12716 13126 12768 13132
rect 12452 12782 12480 13126
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 11520 12378 11572 12384
rect 11808 12406 11928 12434
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 11532 11830 11560 12378
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 10062 10456 11494
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10520 10470 10548 11290
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10612 10266 10640 10610
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10416 10056 10468 10062
rect 10704 10010 10732 10678
rect 11440 10606 11468 11154
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10062 11192 10406
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 10416 9998 10468 10004
rect 10520 9994 10732 10010
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 10508 9988 10732 9994
rect 10560 9982 10732 9988
rect 10508 9930 10560 9936
rect 10520 9518 10548 9930
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10704 9042 10732 9318
rect 10980 9178 11008 9454
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10704 7886 10732 8978
rect 11164 8974 11192 9386
rect 11348 8974 11376 10066
rect 11440 10062 11468 10542
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11440 9518 11468 9998
rect 11532 9674 11560 11766
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11532 9646 11652 9674
rect 11716 9654 11744 10474
rect 11808 10112 11836 12406
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11900 11082 11928 12242
rect 11992 11898 12020 12718
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12452 11558 12480 12718
rect 12728 12714 12756 13126
rect 13004 12850 13032 13874
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13326 13676 13670
rect 13924 13394 13952 14758
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13188 12986 13216 13194
rect 14016 12986 14044 17138
rect 14108 16590 14136 17206
rect 14200 16998 14228 17818
rect 14568 17678 14596 18022
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14568 16998 14596 17614
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14568 16794 14596 16934
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14660 14618 14688 26336
rect 15120 26330 15148 26574
rect 15198 26480 15254 26489
rect 15304 26466 15332 29038
rect 15488 27470 15516 29242
rect 15568 29232 15620 29238
rect 15568 29174 15620 29180
rect 15476 27464 15528 27470
rect 15476 27406 15528 27412
rect 15254 26438 15332 26466
rect 15198 26415 15200 26424
rect 15252 26415 15254 26424
rect 15200 26386 15252 26392
rect 14740 26318 14792 26324
rect 14752 25906 14780 26318
rect 15028 26302 15148 26330
rect 15028 25974 15056 26302
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15384 26240 15436 26246
rect 15488 26228 15516 27406
rect 15436 26200 15516 26228
rect 15384 26182 15436 26188
rect 15016 25968 15068 25974
rect 15016 25910 15068 25916
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 15028 24886 15056 25910
rect 15120 25294 15148 26182
rect 15580 25294 15608 29174
rect 15660 29096 15712 29102
rect 15658 29064 15660 29073
rect 15712 29064 15714 29073
rect 15658 28999 15714 29008
rect 15672 26450 15700 28999
rect 15764 28490 15792 30262
rect 15936 30252 15988 30258
rect 15936 30194 15988 30200
rect 15948 30025 15976 30194
rect 15934 30016 15990 30025
rect 15856 29974 15934 30002
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15856 28150 15884 29974
rect 15934 29951 15990 29960
rect 16040 29306 16068 31962
rect 16396 31816 16448 31822
rect 16500 31804 16528 33050
rect 16448 31776 16528 31804
rect 16580 31816 16632 31822
rect 16396 31758 16448 31764
rect 16684 31804 16712 35958
rect 16868 35630 16896 36042
rect 16948 36032 17000 36038
rect 16948 35974 17000 35980
rect 17040 36032 17092 36038
rect 17040 35974 17092 35980
rect 16960 35834 16988 35974
rect 16948 35828 17000 35834
rect 16948 35770 17000 35776
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 16960 35290 16988 35770
rect 17052 35698 17080 35974
rect 17144 35834 17172 38830
rect 17132 35828 17184 35834
rect 17132 35770 17184 35776
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 16948 35284 17000 35290
rect 16948 35226 17000 35232
rect 16948 34604 17000 34610
rect 16948 34546 17000 34552
rect 16960 33658 16988 34546
rect 16948 33652 17000 33658
rect 16948 33594 17000 33600
rect 17040 33312 17092 33318
rect 17040 33254 17092 33260
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16776 31822 16804 31962
rect 16948 31952 17000 31958
rect 16948 31894 17000 31900
rect 16632 31776 16712 31804
rect 16764 31816 16816 31822
rect 16580 31758 16632 31764
rect 16764 31758 16816 31764
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16672 31680 16724 31686
rect 16578 31648 16634 31657
rect 16672 31622 16724 31628
rect 16578 31583 16634 31592
rect 16486 31376 16542 31385
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 16396 31340 16448 31346
rect 16486 31311 16542 31320
rect 16396 31282 16448 31288
rect 16224 30938 16252 31282
rect 16408 31210 16436 31282
rect 16396 31204 16448 31210
rect 16396 31146 16448 31152
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 16396 30932 16448 30938
rect 16396 30874 16448 30880
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 16304 30728 16356 30734
rect 16304 30670 16356 30676
rect 16132 30258 16160 30670
rect 16210 30288 16266 30297
rect 16120 30252 16172 30258
rect 16210 30223 16266 30232
rect 16120 30194 16172 30200
rect 16132 29889 16160 30194
rect 16118 29880 16174 29889
rect 16118 29815 16174 29824
rect 16028 29300 16080 29306
rect 16028 29242 16080 29248
rect 16224 29238 16252 30223
rect 16316 30054 16344 30670
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16212 29232 16264 29238
rect 16212 29174 16264 29180
rect 16224 29050 16252 29174
rect 16408 29050 16436 30874
rect 16500 30598 16528 31311
rect 16592 30802 16620 31583
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16684 30734 16712 31622
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16488 30592 16540 30598
rect 16488 30534 16540 30540
rect 16488 30320 16540 30326
rect 16488 30262 16540 30268
rect 16040 29022 16252 29050
rect 16316 29022 16436 29050
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 15948 28150 15976 28358
rect 15844 28144 15896 28150
rect 15844 28086 15896 28092
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 15844 27872 15896 27878
rect 15844 27814 15896 27820
rect 15764 27470 15792 27814
rect 15856 27674 15884 27814
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15948 27402 15976 28086
rect 16040 27606 16068 29022
rect 16316 28966 16344 29022
rect 16304 28960 16356 28966
rect 16304 28902 16356 28908
rect 16396 28960 16448 28966
rect 16396 28902 16448 28908
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 16224 28558 16252 28630
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 16132 27470 16160 28018
rect 16224 28014 16252 28494
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16316 28082 16344 28426
rect 16408 28121 16436 28902
rect 16500 28694 16528 30262
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16488 28688 16540 28694
rect 16488 28630 16540 28636
rect 16592 28218 16620 28698
rect 16684 28626 16712 29106
rect 16776 28966 16804 31758
rect 16868 31346 16896 31758
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16868 31249 16896 31282
rect 16854 31240 16910 31249
rect 16854 31175 16910 31184
rect 16856 31136 16908 31142
rect 16856 31078 16908 31084
rect 16764 28960 16816 28966
rect 16764 28902 16816 28908
rect 16764 28688 16816 28694
rect 16764 28630 16816 28636
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 16488 28212 16540 28218
rect 16488 28154 16540 28160
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 16394 28112 16450 28121
rect 16304 28076 16356 28082
rect 16394 28047 16450 28056
rect 16304 28018 16356 28024
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16224 27538 16252 27950
rect 16304 27940 16356 27946
rect 16304 27882 16356 27888
rect 16212 27532 16264 27538
rect 16212 27474 16264 27480
rect 16120 27464 16172 27470
rect 16120 27406 16172 27412
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 16316 27062 16344 27882
rect 16408 27470 16436 28047
rect 16500 28014 16528 28154
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16500 27402 16528 27950
rect 16776 27946 16804 28630
rect 16764 27940 16816 27946
rect 16764 27882 16816 27888
rect 16488 27396 16540 27402
rect 16488 27338 16540 27344
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16684 27130 16712 27338
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16304 27056 16356 27062
rect 16304 26998 16356 27004
rect 15660 26444 15712 26450
rect 15660 26386 15712 26392
rect 16684 26042 16712 27066
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 15108 25288 15160 25294
rect 15476 25288 15528 25294
rect 15108 25230 15160 25236
rect 15474 25256 15476 25265
rect 15568 25288 15620 25294
rect 15528 25256 15530 25265
rect 15568 25230 15620 25236
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15474 25191 15530 25200
rect 16040 24954 16068 25230
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 15566 24848 15622 24857
rect 15028 24410 15056 24822
rect 15566 24783 15622 24792
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15028 23866 15056 24142
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14752 22642 14780 23462
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14844 22574 14872 22918
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21010 14872 21830
rect 14924 21684 14976 21690
rect 14924 21626 14976 21632
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14936 20874 14964 21626
rect 14924 20868 14976 20874
rect 14924 20810 14976 20816
rect 14936 20346 14964 20810
rect 15028 20466 15056 23802
rect 15120 23526 15148 24142
rect 15580 23730 15608 24783
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15764 23662 15792 24550
rect 16040 24274 16068 24890
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15936 23656 15988 23662
rect 15936 23598 15988 23604
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23118 15240 23462
rect 15672 23322 15700 23598
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15948 23254 15976 23598
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15120 22166 15148 22374
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15304 21622 15332 21830
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15488 21078 15516 22034
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15016 20460 15068 20466
rect 15016 20402 15068 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15120 20346 15148 20402
rect 14936 20318 15148 20346
rect 15120 19514 15148 20318
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15212 19378 15240 20470
rect 16028 20392 16080 20398
rect 16224 20380 16252 24754
rect 16408 23769 16436 25774
rect 16578 25392 16634 25401
rect 16684 25362 16712 25842
rect 16776 25430 16804 26726
rect 16764 25424 16816 25430
rect 16764 25366 16816 25372
rect 16578 25327 16634 25336
rect 16672 25356 16724 25362
rect 16592 25294 16620 25327
rect 16672 25298 16724 25304
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16776 25226 16804 25366
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16684 24954 16712 25162
rect 16672 24948 16724 24954
rect 16672 24890 16724 24896
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16394 23760 16450 23769
rect 16394 23695 16396 23704
rect 16448 23695 16450 23704
rect 16396 23666 16448 23672
rect 16592 23662 16620 24074
rect 16684 23730 16712 24142
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16672 23588 16724 23594
rect 16672 23530 16724 23536
rect 16684 22710 16712 23530
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16684 22030 16712 22374
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21146 16620 21830
rect 16776 21486 16804 21966
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16080 20352 16252 20380
rect 16028 20334 16080 20340
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16316 19922 16344 20198
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15120 18426 15148 19110
rect 15108 18420 15160 18426
rect 15028 18380 15108 18408
rect 15028 17270 15056 18380
rect 15108 18362 15160 18368
rect 15212 18358 15240 19314
rect 15396 18970 15424 19314
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15764 18766 15792 19654
rect 16316 18834 16344 19858
rect 16500 19786 16528 20198
rect 16592 20058 16620 20878
rect 16868 20602 16896 31078
rect 16960 30054 16988 31894
rect 17052 31482 17080 33254
rect 17132 31816 17184 31822
rect 17132 31758 17184 31764
rect 17040 31476 17092 31482
rect 17040 31418 17092 31424
rect 17052 31142 17080 31418
rect 17040 31136 17092 31142
rect 17040 31078 17092 31084
rect 17144 30841 17172 31758
rect 17130 30832 17186 30841
rect 17130 30767 17186 30776
rect 17040 30660 17092 30666
rect 17040 30602 17092 30608
rect 17132 30660 17184 30666
rect 17132 30602 17184 30608
rect 17052 30326 17080 30602
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 17040 30184 17092 30190
rect 17144 30161 17172 30602
rect 17040 30126 17092 30132
rect 17130 30152 17186 30161
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 17052 29306 17080 30126
rect 17130 30087 17186 30096
rect 17144 29345 17172 30087
rect 17130 29336 17186 29345
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 17040 29300 17092 29306
rect 17130 29271 17186 29280
rect 17040 29242 17092 29248
rect 16960 29073 16988 29242
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 17132 29164 17184 29170
rect 17132 29106 17184 29112
rect 16946 29064 17002 29073
rect 16946 28999 17002 29008
rect 17052 28762 17080 29106
rect 17040 28756 17092 28762
rect 17040 28698 17092 28704
rect 17144 28694 17172 29106
rect 16948 28688 17000 28694
rect 16948 28630 17000 28636
rect 17132 28688 17184 28694
rect 17132 28630 17184 28636
rect 16960 27674 16988 28630
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 16948 27668 17000 27674
rect 16948 27610 17000 27616
rect 17144 27470 17172 28018
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 16948 26512 17000 26518
rect 16948 26454 17000 26460
rect 16960 24274 16988 26454
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17040 25696 17092 25702
rect 17040 25638 17092 25644
rect 17052 25362 17080 25638
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 17052 24954 17080 25298
rect 17040 24948 17092 24954
rect 17040 24890 17092 24896
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17052 24721 17080 24754
rect 17038 24712 17094 24721
rect 17038 24647 17094 24656
rect 16948 24268 17000 24274
rect 16948 24210 17000 24216
rect 17144 24206 17172 25774
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23798 16988 24006
rect 16948 23792 17000 23798
rect 16948 23734 17000 23740
rect 17236 23254 17264 40582
rect 17408 40588 17540 40594
rect 17460 40582 17540 40588
rect 17408 40530 17460 40536
rect 17316 39976 17368 39982
rect 17316 39918 17368 39924
rect 17328 39574 17356 39918
rect 17316 39568 17368 39574
rect 17316 39510 17368 39516
rect 17316 37324 17368 37330
rect 17316 37266 17368 37272
rect 17328 36922 17356 37266
rect 17316 36916 17368 36922
rect 17316 36858 17368 36864
rect 17420 36786 17448 40530
rect 17604 40458 17632 40967
rect 17776 40928 17828 40934
rect 17776 40870 17828 40876
rect 17868 40928 17920 40934
rect 17868 40870 17920 40876
rect 17788 40662 17816 40870
rect 17776 40656 17828 40662
rect 17776 40598 17828 40604
rect 17880 40526 17908 40870
rect 17868 40520 17920 40526
rect 17868 40462 17920 40468
rect 17592 40452 17644 40458
rect 17592 40394 17644 40400
rect 17604 40186 17632 40394
rect 17592 40180 17644 40186
rect 17592 40122 17644 40128
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17500 39364 17552 39370
rect 17500 39306 17552 39312
rect 17512 38962 17540 39306
rect 17500 38956 17552 38962
rect 17604 38944 17632 39442
rect 17684 38956 17736 38962
rect 17604 38916 17684 38944
rect 17500 38898 17552 38904
rect 17684 38898 17736 38904
rect 17500 38820 17552 38826
rect 17500 38762 17552 38768
rect 17408 36780 17460 36786
rect 17408 36722 17460 36728
rect 17512 36242 17540 38762
rect 17696 37806 17724 38898
rect 17684 37800 17736 37806
rect 17684 37742 17736 37748
rect 17684 37324 17736 37330
rect 17684 37266 17736 37272
rect 17592 37256 17644 37262
rect 17592 37198 17644 37204
rect 17604 36922 17632 37198
rect 17592 36916 17644 36922
rect 17592 36858 17644 36864
rect 17696 36786 17724 37266
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17788 37126 17816 37198
rect 17776 37120 17828 37126
rect 17776 37062 17828 37068
rect 17868 37120 17920 37126
rect 17868 37062 17920 37068
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 17316 35624 17368 35630
rect 17316 35566 17368 35572
rect 17328 35086 17356 35566
rect 17788 35306 17816 37062
rect 17880 36718 17908 37062
rect 17868 36712 17920 36718
rect 17868 36654 17920 36660
rect 17696 35278 17816 35306
rect 17868 35284 17920 35290
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17328 34678 17356 35022
rect 17592 34944 17644 34950
rect 17592 34886 17644 34892
rect 17316 34672 17368 34678
rect 17316 34614 17368 34620
rect 17328 33998 17356 34614
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17604 33658 17632 34886
rect 17592 33652 17644 33658
rect 17592 33594 17644 33600
rect 17316 32836 17368 32842
rect 17316 32778 17368 32784
rect 17328 32570 17356 32778
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17500 32224 17552 32230
rect 17500 32166 17552 32172
rect 17316 31816 17368 31822
rect 17316 31758 17368 31764
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17328 31686 17356 31758
rect 17316 31680 17368 31686
rect 17420 31657 17448 31758
rect 17316 31622 17368 31628
rect 17406 31648 17462 31657
rect 17328 31482 17356 31622
rect 17406 31583 17462 31592
rect 17512 31498 17540 32166
rect 17696 31754 17724 35278
rect 17868 35226 17920 35232
rect 17880 34746 17908 35226
rect 17868 34740 17920 34746
rect 17868 34682 17920 34688
rect 17868 34196 17920 34202
rect 17868 34138 17920 34144
rect 17880 33998 17908 34138
rect 17972 34134 18000 41074
rect 18144 41064 18196 41070
rect 18144 41006 18196 41012
rect 18052 40996 18104 41002
rect 18052 40938 18104 40944
rect 18064 36650 18092 40938
rect 18156 40526 18184 41006
rect 18144 40520 18196 40526
rect 18144 40462 18196 40468
rect 18156 39642 18184 40462
rect 18144 39636 18196 39642
rect 18144 39578 18196 39584
rect 18156 36786 18184 39578
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 18052 36644 18104 36650
rect 18052 36586 18104 36592
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 18248 35766 18276 35974
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 18236 34672 18288 34678
rect 18236 34614 18288 34620
rect 17960 34128 18012 34134
rect 17960 34070 18012 34076
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17880 33522 17908 33934
rect 17972 33862 18000 34070
rect 17960 33856 18012 33862
rect 17960 33798 18012 33804
rect 18144 33856 18196 33862
rect 18144 33798 18196 33804
rect 18052 33584 18104 33590
rect 18052 33526 18104 33532
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 18064 32774 18092 33526
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32570 18092 32710
rect 18052 32564 18104 32570
rect 18052 32506 18104 32512
rect 18064 32450 18092 32506
rect 17972 32422 18092 32450
rect 17776 32224 17828 32230
rect 17776 32166 17828 32172
rect 17316 31476 17368 31482
rect 17316 31418 17368 31424
rect 17420 31470 17540 31498
rect 17604 31726 17724 31754
rect 17314 31376 17370 31385
rect 17314 31311 17316 31320
rect 17368 31311 17370 31320
rect 17316 31282 17368 31288
rect 17314 31240 17370 31249
rect 17314 31175 17370 31184
rect 17328 25276 17356 31175
rect 17420 30938 17448 31470
rect 17498 31376 17554 31385
rect 17498 31311 17500 31320
rect 17552 31311 17554 31320
rect 17500 31282 17552 31288
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17498 30832 17554 30841
rect 17498 30767 17554 30776
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17420 30326 17448 30534
rect 17408 30320 17460 30326
rect 17408 30262 17460 30268
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17420 29850 17448 30126
rect 17408 29844 17460 29850
rect 17408 29786 17460 29792
rect 17512 29209 17540 30767
rect 17498 29200 17554 29209
rect 17604 29170 17632 31726
rect 17684 31680 17736 31686
rect 17684 31622 17736 31628
rect 17696 30734 17724 31622
rect 17788 31346 17816 32166
rect 17776 31340 17828 31346
rect 17776 31282 17828 31288
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17684 30728 17736 30734
rect 17684 30670 17736 30676
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 17696 29850 17724 30670
rect 17788 30394 17816 30670
rect 17776 30388 17828 30394
rect 17776 30330 17828 30336
rect 17684 29844 17736 29850
rect 17684 29786 17736 29792
rect 17788 29714 17816 30330
rect 17880 30172 17908 31282
rect 17972 30326 18000 32422
rect 18052 32360 18104 32366
rect 18052 32302 18104 32308
rect 18064 32026 18092 32302
rect 18052 32020 18104 32026
rect 18052 31962 18104 31968
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 17880 30144 18000 30172
rect 17972 30054 18000 30144
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17776 29708 17828 29714
rect 17776 29650 17828 29656
rect 18064 29510 18092 31758
rect 18156 30734 18184 33798
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18142 30288 18198 30297
rect 18248 30258 18276 34614
rect 18340 31822 18368 41414
rect 18800 41070 18828 41618
rect 18788 41064 18840 41070
rect 18788 41006 18840 41012
rect 18788 40452 18840 40458
rect 18788 40394 18840 40400
rect 18604 40044 18656 40050
rect 18604 39986 18656 39992
rect 18616 39574 18644 39986
rect 18696 39976 18748 39982
rect 18696 39918 18748 39924
rect 18708 39574 18736 39918
rect 18604 39568 18656 39574
rect 18604 39510 18656 39516
rect 18696 39568 18748 39574
rect 18696 39510 18748 39516
rect 18420 39432 18472 39438
rect 18420 39374 18472 39380
rect 18432 39098 18460 39374
rect 18420 39092 18472 39098
rect 18420 39034 18472 39040
rect 18800 37262 18828 40394
rect 18972 37664 19024 37670
rect 18972 37606 19024 37612
rect 18984 37262 19012 37606
rect 18788 37256 18840 37262
rect 18972 37256 19024 37262
rect 18788 37198 18840 37204
rect 18970 37224 18972 37233
rect 19024 37224 19026 37233
rect 18970 37159 19026 37168
rect 18512 33992 18564 33998
rect 18512 33934 18564 33940
rect 18524 33658 18552 33934
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 18420 33448 18472 33454
rect 18420 33390 18472 33396
rect 18432 32570 18460 33390
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 18420 32428 18472 32434
rect 18420 32370 18472 32376
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18328 31136 18380 31142
rect 18432 31113 18460 32370
rect 18788 32292 18840 32298
rect 18788 32234 18840 32240
rect 18972 32292 19024 32298
rect 18972 32234 19024 32240
rect 18800 32026 18828 32234
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18604 31816 18656 31822
rect 18604 31758 18656 31764
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18616 31385 18644 31758
rect 18602 31376 18658 31385
rect 18602 31311 18658 31320
rect 18328 31078 18380 31084
rect 18418 31104 18474 31113
rect 18142 30223 18198 30232
rect 18236 30252 18288 30258
rect 18156 30025 18184 30223
rect 18236 30194 18288 30200
rect 18142 30016 18198 30025
rect 18142 29951 18198 29960
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 17682 29336 17738 29345
rect 17682 29271 17738 29280
rect 17498 29135 17554 29144
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 17408 29096 17460 29102
rect 17460 29056 17540 29084
rect 17408 29038 17460 29044
rect 17512 28490 17540 29056
rect 17696 29050 17724 29271
rect 17960 29164 18012 29170
rect 17960 29106 18012 29112
rect 17604 29022 17724 29050
rect 17500 28484 17552 28490
rect 17500 28426 17552 28432
rect 17408 28076 17460 28082
rect 17512 28064 17540 28426
rect 17604 28422 17632 29022
rect 17868 28756 17920 28762
rect 17868 28698 17920 28704
rect 17684 28552 17736 28558
rect 17684 28494 17736 28500
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17696 28082 17724 28494
rect 17684 28076 17736 28082
rect 17460 28036 17540 28064
rect 17408 28018 17460 28024
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17420 27062 17448 27270
rect 17512 27130 17540 28036
rect 17604 28036 17684 28064
rect 17604 27878 17632 28036
rect 17684 28018 17736 28024
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17776 27872 17828 27878
rect 17776 27814 17828 27820
rect 17604 27470 17632 27814
rect 17788 27674 17816 27814
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17604 27334 17632 27406
rect 17880 27402 17908 28698
rect 17776 27396 17828 27402
rect 17776 27338 17828 27344
rect 17868 27396 17920 27402
rect 17868 27338 17920 27344
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17788 27130 17816 27338
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17408 27056 17460 27062
rect 17408 26998 17460 27004
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17788 26518 17816 26862
rect 17776 26512 17828 26518
rect 17776 26454 17828 26460
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17408 26240 17460 26246
rect 17408 26182 17460 26188
rect 17420 25974 17448 26182
rect 17408 25968 17460 25974
rect 17408 25910 17460 25916
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17408 25424 17460 25430
rect 17406 25392 17408 25401
rect 17460 25392 17462 25401
rect 17406 25327 17462 25336
rect 17408 25288 17460 25294
rect 17328 25248 17408 25276
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 17144 20398 17172 20742
rect 17132 20392 17184 20398
rect 17132 20334 17184 20340
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 15752 18760 15804 18766
rect 16408 18714 16436 19450
rect 15752 18702 15804 18708
rect 16316 18686 16436 18714
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15120 17746 15148 18226
rect 15212 17746 15240 18294
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 15212 17134 15240 17682
rect 15304 17678 15332 18022
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15396 17202 15424 17478
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15212 16658 15240 17070
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14752 15502 14780 16458
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 15638 14964 16050
rect 15212 16046 15240 16594
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15200 15904 15252 15910
rect 15304 15858 15332 16934
rect 15580 16658 15608 16934
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 16316 16522 16344 18686
rect 16592 18222 16620 19450
rect 16684 19378 16712 19790
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16960 18970 16988 19246
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 15252 15852 15332 15858
rect 15200 15846 15332 15852
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15212 15830 15332 15846
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 15212 15502 15240 15830
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 14752 15162 14780 15438
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 15488 14890 15516 15438
rect 15764 15434 15792 15846
rect 16316 15434 16344 16458
rect 15752 15428 15804 15434
rect 15752 15370 15804 15376
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 15476 14884 15528 14890
rect 15476 14826 15528 14832
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 16316 14278 16344 15370
rect 16304 14272 16356 14278
rect 16356 14232 16528 14260
rect 16304 14214 16356 14220
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15396 13326 15424 13806
rect 16500 13326 16528 14232
rect 16592 14074 16620 18022
rect 16960 16674 16988 18770
rect 17144 17338 17172 20334
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 17236 17270 17264 17478
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16794 17080 17138
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 16960 16646 17080 16674
rect 17052 16046 17080 16646
rect 17328 16250 17356 25248
rect 17408 25230 17460 25236
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17420 22642 17448 24890
rect 17512 23118 17540 25434
rect 17604 25430 17632 26318
rect 17696 25498 17724 26318
rect 17880 26314 17908 27338
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17972 25702 18000 29106
rect 18064 29084 18092 29446
rect 18248 29345 18276 30194
rect 18234 29336 18290 29345
rect 18234 29271 18290 29280
rect 18236 29164 18288 29170
rect 18236 29106 18288 29112
rect 18144 29096 18196 29102
rect 18064 29056 18144 29084
rect 18144 29038 18196 29044
rect 18248 28558 18276 29106
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18052 28484 18104 28490
rect 18052 28426 18104 28432
rect 18064 28082 18092 28426
rect 18248 28150 18276 28494
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18052 28076 18104 28082
rect 18052 28018 18104 28024
rect 18236 27940 18288 27946
rect 18236 27882 18288 27888
rect 18144 27532 18196 27538
rect 18144 27474 18196 27480
rect 18156 27062 18184 27474
rect 18248 27470 18276 27882
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 18144 27056 18196 27062
rect 18144 26998 18196 27004
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 18064 25974 18092 26930
rect 18144 26512 18196 26518
rect 18144 26454 18196 26460
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 17960 25696 18012 25702
rect 17960 25638 18012 25644
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17592 25424 17644 25430
rect 17592 25366 17644 25372
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 17972 25265 18000 25298
rect 17958 25256 18014 25265
rect 17684 25220 17736 25226
rect 17958 25191 18014 25200
rect 17684 25162 17736 25168
rect 17592 25152 17644 25158
rect 17592 25094 17644 25100
rect 17604 24886 17632 25094
rect 17592 24880 17644 24886
rect 17592 24822 17644 24828
rect 17696 24721 17724 25162
rect 17774 24848 17830 24857
rect 17774 24783 17830 24792
rect 17682 24712 17738 24721
rect 17682 24647 17738 24656
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17604 23186 17632 24142
rect 17788 24138 17816 24783
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17972 23594 18000 24550
rect 18064 23730 18092 25910
rect 18156 25294 18184 26454
rect 18236 26444 18288 26450
rect 18340 26432 18368 31078
rect 18418 31039 18474 31048
rect 18420 30796 18472 30802
rect 18420 30738 18472 30744
rect 18288 26404 18368 26432
rect 18432 26432 18460 30738
rect 18512 30728 18564 30734
rect 18512 30670 18564 30676
rect 18524 30190 18552 30670
rect 18616 30569 18644 31311
rect 18800 30938 18828 31758
rect 18984 31754 19012 32234
rect 18892 31726 19012 31754
rect 18892 31346 18920 31726
rect 19076 31482 19104 42638
rect 19156 42288 19208 42294
rect 19156 42230 19208 42236
rect 19168 36582 19196 42230
rect 19248 41064 19300 41070
rect 19246 41032 19248 41041
rect 19300 41032 19302 41041
rect 19246 40967 19302 40976
rect 19248 39500 19300 39506
rect 19248 39442 19300 39448
rect 19260 38962 19288 39442
rect 19248 38956 19300 38962
rect 19248 38898 19300 38904
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 19260 38214 19288 38286
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 19260 38010 19288 38150
rect 19248 38004 19300 38010
rect 19248 37946 19300 37952
rect 19248 37120 19300 37126
rect 19248 37062 19300 37068
rect 19260 36922 19288 37062
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 19156 36576 19208 36582
rect 19156 36518 19208 36524
rect 19352 35816 19380 43182
rect 19812 42702 19840 43250
rect 21008 42945 21036 43250
rect 20994 42936 21050 42945
rect 20994 42871 21050 42880
rect 19800 42696 19852 42702
rect 19800 42638 19852 42644
rect 19892 42696 19944 42702
rect 19892 42638 19944 42644
rect 19524 42628 19576 42634
rect 19524 42570 19576 42576
rect 19432 42560 19484 42566
rect 19432 42502 19484 42508
rect 19444 42158 19472 42502
rect 19432 42152 19484 42158
rect 19432 42094 19484 42100
rect 19432 41472 19484 41478
rect 19536 41460 19564 42570
rect 19812 42158 19840 42638
rect 19904 42362 19932 42638
rect 20812 42628 20864 42634
rect 20812 42570 20864 42576
rect 21548 42628 21600 42634
rect 21548 42570 21600 42576
rect 19892 42356 19944 42362
rect 19892 42298 19944 42304
rect 19904 42226 19932 42298
rect 20720 42288 20772 42294
rect 20720 42230 20772 42236
rect 19892 42220 19944 42226
rect 19892 42162 19944 42168
rect 19800 42152 19852 42158
rect 19800 42094 19852 42100
rect 20168 42152 20220 42158
rect 20168 42094 20220 42100
rect 20180 41818 20208 42094
rect 20168 41812 20220 41818
rect 20168 41754 20220 41760
rect 20076 41676 20128 41682
rect 20076 41618 20128 41624
rect 19984 41608 20036 41614
rect 19984 41550 20036 41556
rect 19484 41432 19564 41460
rect 19432 41414 19484 41420
rect 19444 41274 19472 41414
rect 19996 41274 20024 41550
rect 19432 41268 19484 41274
rect 19432 41210 19484 41216
rect 19984 41268 20036 41274
rect 19984 41210 20036 41216
rect 19984 41064 20036 41070
rect 19984 41006 20036 41012
rect 19800 40996 19852 41002
rect 19800 40938 19852 40944
rect 19812 40594 19840 40938
rect 19996 40730 20024 41006
rect 20088 40730 20116 41618
rect 20732 41614 20760 42230
rect 20824 42022 20852 42570
rect 20812 42016 20864 42022
rect 20812 41958 20864 41964
rect 20720 41608 20772 41614
rect 20824 41585 20852 41958
rect 21560 41818 21588 42570
rect 22756 42566 22784 43250
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22744 42560 22796 42566
rect 22744 42502 22796 42508
rect 22008 42356 22060 42362
rect 22008 42298 22060 42304
rect 21732 42016 21784 42022
rect 21732 41958 21784 41964
rect 21824 42016 21876 42022
rect 21824 41958 21876 41964
rect 21548 41812 21600 41818
rect 21548 41754 21600 41760
rect 21744 41682 21772 41958
rect 21088 41676 21140 41682
rect 21088 41618 21140 41624
rect 21732 41676 21784 41682
rect 21732 41618 21784 41624
rect 20720 41550 20772 41556
rect 20810 41576 20866 41585
rect 19984 40724 20036 40730
rect 19984 40666 20036 40672
rect 20076 40724 20128 40730
rect 20076 40666 20128 40672
rect 19800 40588 19852 40594
rect 19800 40530 19852 40536
rect 20088 40458 20116 40666
rect 20076 40452 20128 40458
rect 20076 40394 20128 40400
rect 20628 40452 20680 40458
rect 20628 40394 20680 40400
rect 20088 40186 20116 40394
rect 20640 40186 20668 40394
rect 20076 40180 20128 40186
rect 20076 40122 20128 40128
rect 20628 40180 20680 40186
rect 20628 40122 20680 40128
rect 20640 39574 20668 40122
rect 20732 39846 20760 41550
rect 20810 41511 20866 41520
rect 20904 41132 20956 41138
rect 20904 41074 20956 41080
rect 20916 40730 20944 41074
rect 20996 41064 21048 41070
rect 20996 41006 21048 41012
rect 20904 40724 20956 40730
rect 20904 40666 20956 40672
rect 20812 40656 20864 40662
rect 20812 40598 20864 40604
rect 20824 40118 20852 40598
rect 20812 40112 20864 40118
rect 20812 40054 20864 40060
rect 21008 40050 21036 41006
rect 21100 40934 21128 41618
rect 21364 41540 21416 41546
rect 21364 41482 21416 41488
rect 21376 41414 21404 41482
rect 21376 41386 21496 41414
rect 21088 40928 21140 40934
rect 21088 40870 21140 40876
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 20996 40044 21048 40050
rect 20996 39986 21048 39992
rect 20720 39840 20772 39846
rect 20720 39782 20772 39788
rect 20628 39568 20680 39574
rect 20628 39510 20680 39516
rect 21100 39506 21128 40666
rect 21272 40520 21324 40526
rect 21272 40462 21324 40468
rect 21284 40186 21312 40462
rect 21272 40180 21324 40186
rect 21272 40122 21324 40128
rect 20260 39500 20312 39506
rect 20260 39442 20312 39448
rect 21088 39500 21140 39506
rect 21088 39442 21140 39448
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19524 39432 19576 39438
rect 19524 39374 19576 39380
rect 19708 39432 19760 39438
rect 19708 39374 19760 39380
rect 20168 39432 20220 39438
rect 20168 39374 20220 39380
rect 19444 38944 19472 39374
rect 19536 39098 19564 39374
rect 19524 39092 19576 39098
rect 19524 39034 19576 39040
rect 19524 38956 19576 38962
rect 19444 38916 19524 38944
rect 19524 38898 19576 38904
rect 19536 38554 19564 38898
rect 19720 38894 19748 39374
rect 20180 39098 20208 39374
rect 20272 39098 20300 39442
rect 20996 39364 21048 39370
rect 20996 39306 21048 39312
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20260 39092 20312 39098
rect 20260 39034 20312 39040
rect 21008 38962 21036 39306
rect 20996 38956 21048 38962
rect 20996 38898 21048 38904
rect 19708 38888 19760 38894
rect 19708 38830 19760 38836
rect 19720 38554 19748 38830
rect 21008 38554 21036 38898
rect 19524 38548 19576 38554
rect 19524 38490 19576 38496
rect 19708 38548 19760 38554
rect 19708 38490 19760 38496
rect 20996 38548 21048 38554
rect 20996 38490 21048 38496
rect 21272 38548 21324 38554
rect 21272 38490 21324 38496
rect 19616 38480 19668 38486
rect 19616 38422 19668 38428
rect 19524 38412 19576 38418
rect 19524 38354 19576 38360
rect 19432 38344 19484 38350
rect 19432 38286 19484 38292
rect 19444 38010 19472 38286
rect 19536 38282 19564 38354
rect 19524 38276 19576 38282
rect 19524 38218 19576 38224
rect 19628 38010 19656 38422
rect 21284 38350 21312 38490
rect 19892 38344 19944 38350
rect 19892 38286 19944 38292
rect 20996 38344 21048 38350
rect 20996 38286 21048 38292
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 21362 38312 21418 38321
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 19616 38004 19668 38010
rect 19616 37946 19668 37952
rect 19904 37806 19932 38286
rect 20076 37936 20128 37942
rect 20076 37878 20128 37884
rect 19892 37800 19944 37806
rect 19892 37742 19944 37748
rect 19616 37664 19668 37670
rect 19616 37606 19668 37612
rect 19628 37262 19656 37606
rect 19708 37324 19760 37330
rect 19708 37266 19760 37272
rect 19616 37256 19668 37262
rect 19616 37198 19668 37204
rect 19524 36644 19576 36650
rect 19524 36586 19576 36592
rect 19352 35788 19472 35816
rect 19444 33454 19472 35788
rect 19536 35766 19564 36586
rect 19616 36576 19668 36582
rect 19616 36518 19668 36524
rect 19524 35760 19576 35766
rect 19524 35702 19576 35708
rect 19536 33522 19564 35702
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19432 32836 19484 32842
rect 19536 32824 19564 33458
rect 19484 32796 19564 32824
rect 19432 32778 19484 32784
rect 19156 32768 19208 32774
rect 19156 32710 19208 32716
rect 19168 32434 19196 32710
rect 19444 32502 19472 32778
rect 19628 32502 19656 36518
rect 19720 36242 19748 37266
rect 19800 37120 19852 37126
rect 19800 37062 19852 37068
rect 19708 36236 19760 36242
rect 19708 36178 19760 36184
rect 19708 36032 19760 36038
rect 19708 35974 19760 35980
rect 19720 35290 19748 35974
rect 19812 35562 19840 37062
rect 19904 36922 19932 37742
rect 19892 36916 19944 36922
rect 19892 36858 19944 36864
rect 20088 36718 20116 37878
rect 21008 37806 21036 38286
rect 21362 38247 21364 38256
rect 21416 38247 21418 38256
rect 21364 38218 21416 38224
rect 21376 37874 21404 38218
rect 21364 37868 21416 37874
rect 21364 37810 21416 37816
rect 20996 37800 21048 37806
rect 20996 37742 21048 37748
rect 21008 37466 21036 37742
rect 20996 37460 21048 37466
rect 20996 37402 21048 37408
rect 20076 36712 20128 36718
rect 20076 36654 20128 36660
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 19892 36236 19944 36242
rect 19892 36178 19944 36184
rect 19904 35698 19932 36178
rect 19996 36174 20024 36518
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19892 35692 19944 35698
rect 19892 35634 19944 35640
rect 20088 35630 20116 36654
rect 20904 36100 20956 36106
rect 20904 36042 20956 36048
rect 20916 35834 20944 36042
rect 20904 35828 20956 35834
rect 20904 35770 20956 35776
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 20076 35624 20128 35630
rect 20076 35566 20128 35572
rect 19800 35556 19852 35562
rect 19800 35498 19852 35504
rect 19708 35284 19760 35290
rect 19708 35226 19760 35232
rect 20180 35154 20208 35634
rect 20444 35624 20496 35630
rect 20444 35566 20496 35572
rect 20456 35494 20484 35566
rect 20444 35488 20496 35494
rect 20444 35430 20496 35436
rect 20456 35222 20484 35430
rect 20444 35216 20496 35222
rect 20444 35158 20496 35164
rect 20168 35148 20220 35154
rect 20168 35090 20220 35096
rect 20180 34762 20208 35090
rect 20548 34950 20576 35634
rect 20536 34944 20588 34950
rect 20536 34886 20588 34892
rect 20628 34944 20680 34950
rect 20628 34886 20680 34892
rect 20088 34746 20208 34762
rect 20076 34740 20208 34746
rect 20128 34734 20208 34740
rect 20076 34682 20128 34688
rect 20548 34626 20576 34886
rect 20640 34746 20668 34886
rect 20628 34740 20680 34746
rect 20628 34682 20680 34688
rect 20444 34604 20496 34610
rect 20548 34598 20668 34626
rect 20444 34546 20496 34552
rect 20076 33448 20128 33454
rect 20076 33390 20128 33396
rect 20088 32978 20116 33390
rect 20076 32972 20128 32978
rect 20076 32914 20128 32920
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19616 32496 19668 32502
rect 19616 32438 19668 32444
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 18892 30802 18920 31282
rect 18880 30796 18932 30802
rect 18880 30738 18932 30744
rect 18696 30592 18748 30598
rect 18602 30560 18658 30569
rect 18696 30534 18748 30540
rect 18602 30495 18658 30504
rect 18708 30394 18736 30534
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18604 30048 18656 30054
rect 18602 30016 18604 30025
rect 18656 30016 18658 30025
rect 18602 29951 18658 29960
rect 18696 29096 18748 29102
rect 18696 29038 18748 29044
rect 18788 29096 18840 29102
rect 18788 29038 18840 29044
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18524 28422 18552 28902
rect 18708 28762 18736 29038
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18524 27878 18552 28358
rect 18616 28082 18644 28494
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18708 27690 18736 28698
rect 18800 28694 18828 29038
rect 18788 28688 18840 28694
rect 18788 28630 18840 28636
rect 18892 28626 18920 30738
rect 19062 30560 19118 30569
rect 19062 30495 19118 30504
rect 18972 30184 19024 30190
rect 18972 30126 19024 30132
rect 18880 28620 18932 28626
rect 18880 28562 18932 28568
rect 18788 28552 18840 28558
rect 18788 28494 18840 28500
rect 18800 28150 18828 28494
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 18708 27662 18828 27690
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18708 26994 18736 27542
rect 18800 27538 18828 27662
rect 18788 27532 18840 27538
rect 18788 27474 18840 27480
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18604 26852 18656 26858
rect 18604 26794 18656 26800
rect 18512 26444 18564 26450
rect 18432 26404 18512 26432
rect 18236 26386 18288 26392
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18248 25362 18276 26182
rect 18340 25820 18368 26404
rect 18512 26386 18564 26392
rect 18420 25832 18472 25838
rect 18340 25792 18420 25820
rect 18340 25514 18368 25792
rect 18420 25774 18472 25780
rect 18340 25486 18460 25514
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18340 24954 18368 25298
rect 18432 25294 18460 25486
rect 18524 25362 18552 26386
rect 18616 26382 18644 26794
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18432 24954 18460 25230
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18234 24304 18290 24313
rect 18234 24239 18290 24248
rect 18142 24168 18198 24177
rect 18248 24138 18276 24239
rect 18142 24103 18198 24112
rect 18236 24132 18288 24138
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 17500 23112 17552 23118
rect 17500 23054 17552 23060
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17420 21690 17448 22578
rect 17512 22386 17540 22646
rect 17604 22574 17632 23122
rect 17684 22976 17736 22982
rect 17684 22918 17736 22924
rect 17696 22642 17724 22918
rect 18156 22710 18184 24103
rect 18236 24074 18288 24080
rect 18340 23905 18368 24890
rect 18432 24177 18460 24890
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18524 24206 18552 24618
rect 18616 24410 18644 25638
rect 18708 25401 18736 26930
rect 18788 26512 18840 26518
rect 18788 26454 18840 26460
rect 18800 25770 18828 26454
rect 18788 25764 18840 25770
rect 18788 25706 18840 25712
rect 18694 25392 18750 25401
rect 18694 25327 18750 25336
rect 18800 25226 18828 25706
rect 18788 25220 18840 25226
rect 18788 25162 18840 25168
rect 18694 24848 18750 24857
rect 18694 24783 18696 24792
rect 18748 24783 18750 24792
rect 18696 24754 18748 24760
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18512 24200 18564 24206
rect 18418 24168 18474 24177
rect 18512 24142 18564 24148
rect 18418 24103 18474 24112
rect 18326 23896 18382 23905
rect 18708 23866 18736 24754
rect 18800 24138 18828 25162
rect 18880 24948 18932 24954
rect 18984 24936 19012 30126
rect 18932 24908 19012 24936
rect 18880 24890 18932 24896
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18326 23831 18382 23840
rect 18420 23860 18472 23866
rect 18236 23792 18288 23798
rect 18236 23734 18288 23740
rect 18144 22704 18196 22710
rect 18144 22646 18196 22652
rect 18248 22642 18276 23734
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 17592 22568 17644 22574
rect 17592 22510 17644 22516
rect 17512 22358 17632 22386
rect 17604 22114 17632 22358
rect 18340 22234 18368 23831
rect 18420 23802 18472 23808
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18328 22228 18380 22234
rect 18328 22170 18380 22176
rect 17776 22160 17828 22166
rect 17604 22108 17776 22114
rect 17604 22102 17828 22108
rect 17604 22086 17816 22102
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17420 21146 17448 21422
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17512 18834 17540 21966
rect 17604 20398 17632 22086
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18156 21486 18184 21830
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17696 19854 17724 20334
rect 17788 20058 17816 20402
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17684 19440 17736 19446
rect 17684 19382 17736 19388
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17696 17678 17724 19382
rect 17880 18816 17908 21014
rect 18156 21010 18184 21286
rect 18144 21004 18196 21010
rect 18144 20946 18196 20952
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18248 20806 18276 20946
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 18432 19854 18460 23802
rect 18708 23730 18736 23802
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18616 23610 18644 23666
rect 18892 23610 18920 24890
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18984 24342 19012 24686
rect 19076 24410 19104 30495
rect 19260 29306 19288 32370
rect 19628 32348 19656 32438
rect 19352 32320 19656 32348
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19352 28642 19380 32320
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19444 31278 19472 31758
rect 20088 31754 20116 32438
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 20180 31958 20208 32302
rect 20168 31952 20220 31958
rect 20168 31894 20220 31900
rect 19616 31748 19668 31754
rect 19616 31690 19668 31696
rect 19996 31726 20116 31754
rect 19628 31482 19656 31690
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19800 31408 19852 31414
rect 19800 31350 19852 31356
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 19432 31272 19484 31278
rect 19432 31214 19484 31220
rect 19444 30938 19472 31214
rect 19432 30932 19484 30938
rect 19432 30874 19484 30880
rect 19524 30660 19576 30666
rect 19576 30620 19656 30648
rect 19524 30602 19576 30608
rect 19628 30326 19656 30620
rect 19616 30320 19668 30326
rect 19616 30262 19668 30268
rect 19352 28614 19564 28642
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19444 28218 19472 28426
rect 19432 28212 19484 28218
rect 19432 28154 19484 28160
rect 19338 28112 19394 28121
rect 19338 28047 19394 28056
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 19156 26784 19208 26790
rect 19156 26726 19208 26732
rect 19168 26586 19196 26726
rect 19156 26580 19208 26586
rect 19156 26522 19208 26528
rect 19168 25974 19196 26522
rect 19260 26382 19288 27814
rect 19352 27674 19380 28047
rect 19340 27668 19392 27674
rect 19340 27610 19392 27616
rect 19536 27470 19564 28614
rect 19628 27996 19656 30262
rect 19720 28121 19748 31282
rect 19812 30938 19840 31350
rect 19892 31136 19944 31142
rect 19892 31078 19944 31084
rect 19800 30932 19852 30938
rect 19800 30874 19852 30880
rect 19904 30666 19932 31078
rect 19800 30660 19852 30666
rect 19800 30602 19852 30608
rect 19892 30660 19944 30666
rect 19892 30602 19944 30608
rect 19812 30190 19840 30602
rect 19800 30184 19852 30190
rect 19800 30126 19852 30132
rect 19996 28490 20024 31726
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20076 31204 20128 31210
rect 20076 31146 20128 31152
rect 20088 30802 20116 31146
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 20180 30716 20208 31282
rect 20364 30938 20392 31282
rect 20352 30932 20404 30938
rect 20352 30874 20404 30880
rect 20352 30728 20404 30734
rect 20180 30688 20352 30716
rect 20180 30394 20208 30688
rect 20352 30670 20404 30676
rect 20456 30598 20484 34546
rect 20640 33862 20668 34598
rect 21180 34400 21232 34406
rect 21180 34342 21232 34348
rect 21192 33998 21220 34342
rect 21180 33992 21232 33998
rect 21180 33934 21232 33940
rect 20628 33856 20680 33862
rect 20628 33798 20680 33804
rect 20640 33590 20668 33798
rect 20536 33584 20588 33590
rect 20536 33526 20588 33532
rect 20628 33584 20680 33590
rect 20628 33526 20680 33532
rect 20548 32366 20576 33526
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 20640 32978 20668 33390
rect 20628 32972 20680 32978
rect 20628 32914 20680 32920
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20812 31816 20864 31822
rect 20916 31804 20944 32166
rect 21192 32026 21312 32042
rect 21180 32020 21312 32026
rect 21232 32014 21312 32020
rect 21180 31962 21232 31968
rect 20996 31816 21048 31822
rect 20916 31776 20996 31804
rect 20812 31758 20864 31764
rect 21048 31776 21128 31804
rect 20996 31758 21048 31764
rect 20720 31680 20772 31686
rect 20720 31622 20772 31628
rect 20732 31521 20760 31622
rect 20718 31512 20774 31521
rect 20718 31447 20774 31456
rect 20824 31362 20852 31758
rect 20994 31512 21050 31521
rect 20994 31447 21050 31456
rect 21008 31414 21036 31447
rect 20996 31408 21048 31414
rect 20824 31346 20944 31362
rect 20996 31350 21048 31356
rect 20824 31340 20956 31346
rect 20824 31334 20904 31340
rect 20904 31282 20956 31288
rect 20720 31204 20772 31210
rect 20720 31146 20772 31152
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 20444 30592 20496 30598
rect 20444 30534 20496 30540
rect 20168 30388 20220 30394
rect 20168 30330 20220 30336
rect 20260 30116 20312 30122
rect 20260 30058 20312 30064
rect 20272 29850 20300 30058
rect 20260 29844 20312 29850
rect 20260 29786 20312 29792
rect 20272 29170 20300 29786
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19706 28112 19762 28121
rect 19706 28047 19762 28056
rect 19628 27968 19748 27996
rect 19524 27464 19576 27470
rect 19524 27406 19576 27412
rect 19616 27396 19668 27402
rect 19616 27338 19668 27344
rect 19432 26920 19484 26926
rect 19432 26862 19484 26868
rect 19524 26920 19576 26926
rect 19524 26862 19576 26868
rect 19444 26450 19472 26862
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19168 25702 19196 25910
rect 19156 25696 19208 25702
rect 19156 25638 19208 25644
rect 19536 24818 19564 26862
rect 19628 26586 19656 27338
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19720 24834 19748 27968
rect 19996 27130 20024 28426
rect 20352 27328 20404 27334
rect 20352 27270 20404 27276
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 20364 26450 20392 27270
rect 20456 26926 20484 30534
rect 20548 30394 20576 31078
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20536 30388 20588 30394
rect 20536 30330 20588 30336
rect 20640 30258 20668 30874
rect 20732 30734 20760 31146
rect 20812 31136 20864 31142
rect 20812 31078 20864 31084
rect 20824 30802 20852 31078
rect 20812 30796 20864 30802
rect 20812 30738 20864 30744
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20732 30394 20760 30670
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20628 30252 20680 30258
rect 20628 30194 20680 30200
rect 20640 29646 20668 30194
rect 20628 29640 20680 29646
rect 20628 29582 20680 29588
rect 20810 29608 20866 29617
rect 20810 29543 20812 29552
rect 20864 29543 20866 29552
rect 20812 29514 20864 29520
rect 20536 29504 20588 29510
rect 20536 29446 20588 29452
rect 20548 29170 20576 29446
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20824 28150 20852 29514
rect 20812 28144 20864 28150
rect 20812 28086 20864 28092
rect 20536 27464 20588 27470
rect 20536 27406 20588 27412
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20260 25900 20312 25906
rect 20260 25842 20312 25848
rect 20272 25498 20300 25842
rect 20364 25770 20392 26386
rect 20456 26246 20484 26862
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20272 24954 20300 25230
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 19720 24818 19840 24834
rect 20088 24818 20116 24890
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19708 24812 19840 24818
rect 19760 24806 19840 24812
rect 19708 24754 19760 24760
rect 19536 24698 19564 24754
rect 19536 24670 19748 24698
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19064 24404 19116 24410
rect 19064 24346 19116 24352
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 18972 24336 19024 24342
rect 19260 24313 19288 24346
rect 18972 24278 19024 24284
rect 19246 24304 19302 24313
rect 18984 23866 19012 24278
rect 19246 24239 19302 24248
rect 19628 24206 19656 24550
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19156 24200 19208 24206
rect 19616 24200 19668 24206
rect 19156 24142 19208 24148
rect 19292 24168 19348 24177
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18616 23582 18920 23610
rect 18616 23322 18644 23582
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18604 22024 18656 22030
rect 18602 21992 18604 22001
rect 18656 21992 18658 22001
rect 18602 21927 18658 21936
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18708 21350 18736 21830
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18616 20262 18644 20946
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18616 20058 18644 20198
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18892 19922 18920 20878
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18984 19854 19012 20198
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 17788 18788 17908 18816
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17328 16130 17356 16186
rect 17236 16102 17356 16130
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16684 13870 16712 14350
rect 17052 14278 17080 15982
rect 17236 15706 17264 16102
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17328 15706 17356 15982
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17696 15502 17724 17614
rect 17788 17134 17816 18788
rect 18432 18766 18460 19450
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17776 17128 17828 17134
rect 17776 17070 17828 17076
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 15094 17724 15438
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 14006 17080 14214
rect 17040 14000 17092 14006
rect 17040 13942 17092 13948
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16592 13530 16620 13806
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16684 13394 16712 13806
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12728 11830 12756 12650
rect 13004 11880 13032 12786
rect 13084 11892 13136 11898
rect 13004 11852 13084 11880
rect 13084 11834 13136 11840
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 13096 11150 13124 11834
rect 13188 11218 13216 12922
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13556 11150 13584 12038
rect 13924 11898 13952 12854
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14108 12374 14136 12718
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13924 11082 13952 11834
rect 14292 11354 14320 13262
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14384 11830 14412 13126
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14568 11286 14596 12718
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12170 15240 12582
rect 16684 12434 16712 13330
rect 16776 12850 16804 13670
rect 16960 12986 16988 13806
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 17236 12442 17264 13194
rect 17420 12986 17448 14418
rect 17696 14006 17724 15030
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17696 13870 17724 13942
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17788 13682 17816 17070
rect 17880 16590 17908 18634
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17972 16726 18000 18158
rect 18064 17882 18092 18158
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17696 13654 17816 13682
rect 17696 13462 17724 13654
rect 17880 13546 17908 16526
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18432 15706 18460 16050
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17788 13518 17908 13546
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17696 12986 17724 13398
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17788 12782 17816 13518
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12782 17908 13330
rect 17972 12986 18000 14282
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 17972 12850 18000 12922
rect 18064 12850 18092 13670
rect 18524 13394 18552 19654
rect 19076 19514 19104 24142
rect 19168 23905 19196 24142
rect 19348 24138 19564 24154
rect 19616 24142 19668 24148
rect 19720 24138 19748 24670
rect 19348 24132 19576 24138
rect 19348 24126 19524 24132
rect 19292 24103 19348 24112
rect 19524 24074 19576 24080
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19248 24064 19300 24070
rect 19246 24032 19248 24041
rect 19300 24032 19302 24041
rect 19812 24018 19840 24806
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24614 20208 24754
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 24410 20484 24550
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19904 24018 19932 24210
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19246 23967 19302 23976
rect 19720 23990 19932 24018
rect 19154 23896 19210 23905
rect 19154 23831 19210 23840
rect 19720 23526 19748 23990
rect 20088 23798 20116 24142
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19812 22778 19840 23054
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19156 21004 19208 21010
rect 19156 20946 19208 20952
rect 19168 20262 19196 20946
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 20058 19196 20198
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18892 18290 18920 18566
rect 19168 18426 19196 19790
rect 19260 19378 19288 19790
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19628 19334 19656 22714
rect 19904 22658 19932 23054
rect 19812 22630 19932 22658
rect 20088 22642 20116 23462
rect 20076 22636 20128 22642
rect 19812 22438 19840 22630
rect 20076 22578 20128 22584
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 19812 22098 19840 22374
rect 20180 22234 20208 23666
rect 20548 23662 20576 27406
rect 20720 26308 20772 26314
rect 20720 26250 20772 26256
rect 20732 26042 20760 26250
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20916 25974 20944 31282
rect 21008 29866 21036 31350
rect 21100 31210 21128 31776
rect 21178 31784 21234 31793
rect 21178 31719 21234 31728
rect 21088 31204 21140 31210
rect 21088 31146 21140 31152
rect 21088 30796 21140 30802
rect 21088 30738 21140 30744
rect 21100 30258 21128 30738
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 21192 30122 21220 31719
rect 21180 30116 21232 30122
rect 21180 30058 21232 30064
rect 21008 29838 21128 29866
rect 20994 29744 21050 29753
rect 20994 29679 21050 29688
rect 21008 29578 21036 29679
rect 20996 29572 21048 29578
rect 20996 29514 21048 29520
rect 21100 28966 21128 29838
rect 21180 29708 21232 29714
rect 21180 29650 21232 29656
rect 21192 29510 21220 29650
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21180 29028 21232 29034
rect 21180 28970 21232 28976
rect 21088 28960 21140 28966
rect 21088 28902 21140 28908
rect 20994 28792 21050 28801
rect 20994 28727 20996 28736
rect 21048 28727 21050 28736
rect 20996 28698 21048 28704
rect 21008 28082 21036 28698
rect 21192 28558 21220 28970
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 21192 27674 21220 28494
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 21284 27606 21312 32014
rect 21468 31958 21496 41386
rect 21548 39840 21600 39846
rect 21548 39782 21600 39788
rect 21560 39370 21588 39782
rect 21548 39364 21600 39370
rect 21548 39306 21600 39312
rect 21560 37194 21588 39306
rect 21638 38448 21694 38457
rect 21638 38383 21694 38392
rect 21652 38350 21680 38383
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21548 37188 21600 37194
rect 21548 37130 21600 37136
rect 21560 36854 21588 37130
rect 21548 36848 21600 36854
rect 21548 36790 21600 36796
rect 21560 36088 21588 36790
rect 21640 36100 21692 36106
rect 21560 36060 21640 36088
rect 21640 36042 21692 36048
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21548 31816 21600 31822
rect 21546 31784 21548 31793
rect 21640 31816 21692 31822
rect 21600 31784 21602 31793
rect 21456 31748 21508 31754
rect 21640 31758 21692 31764
rect 21546 31719 21602 31728
rect 21456 31690 21508 31696
rect 21468 30598 21496 31690
rect 21652 31482 21680 31758
rect 21640 31476 21692 31482
rect 21640 31418 21692 31424
rect 21744 31414 21772 41618
rect 21836 41614 21864 41958
rect 22020 41614 22048 42298
rect 21824 41608 21876 41614
rect 22008 41608 22060 41614
rect 21824 41550 21876 41556
rect 22006 41576 22008 41585
rect 22060 41576 22062 41585
rect 22204 41546 22232 42502
rect 22652 42152 22704 42158
rect 22652 42094 22704 42100
rect 22006 41511 22062 41520
rect 22192 41540 22244 41546
rect 22192 41482 22244 41488
rect 22558 41168 22614 41177
rect 22558 41103 22560 41112
rect 22612 41103 22614 41112
rect 22560 41074 22612 41080
rect 22100 40588 22152 40594
rect 22100 40530 22152 40536
rect 21824 40452 21876 40458
rect 21824 40394 21876 40400
rect 21836 39506 21864 40394
rect 22112 40050 22140 40530
rect 22100 40044 22152 40050
rect 22100 39986 22152 39992
rect 21824 39500 21876 39506
rect 21824 39442 21876 39448
rect 21836 39409 21864 39442
rect 21822 39400 21878 39409
rect 21822 39335 21878 39344
rect 22100 38956 22152 38962
rect 22100 38898 22152 38904
rect 22112 38554 22140 38898
rect 22100 38548 22152 38554
rect 22100 38490 22152 38496
rect 22284 38480 22336 38486
rect 22282 38448 22284 38457
rect 22336 38448 22338 38457
rect 22282 38383 22338 38392
rect 22296 38350 22324 38383
rect 22284 38344 22336 38350
rect 22376 38344 22428 38350
rect 22284 38286 22336 38292
rect 22374 38312 22376 38321
rect 22428 38312 22430 38321
rect 22374 38247 22430 38256
rect 21824 38208 21876 38214
rect 21822 38176 21824 38185
rect 22560 38208 22612 38214
rect 21876 38176 21878 38185
rect 21822 38111 21878 38120
rect 22558 38176 22560 38185
rect 22612 38176 22614 38185
rect 22558 38111 22614 38120
rect 22376 37936 22428 37942
rect 22376 37878 22428 37884
rect 22100 37664 22152 37670
rect 22100 37606 22152 37612
rect 22112 37330 22140 37606
rect 22100 37324 22152 37330
rect 22100 37266 22152 37272
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 21916 36780 21968 36786
rect 21916 36722 21968 36728
rect 21928 36378 21956 36722
rect 21916 36372 21968 36378
rect 21916 36314 21968 36320
rect 22204 36242 22232 37130
rect 22192 36236 22244 36242
rect 22192 36178 22244 36184
rect 22284 35624 22336 35630
rect 22284 35566 22336 35572
rect 22296 35290 22324 35566
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22388 35222 22416 37878
rect 22468 37800 22520 37806
rect 22468 37742 22520 37748
rect 22480 36786 22508 37742
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22468 36100 22520 36106
rect 22468 36042 22520 36048
rect 22480 35834 22508 36042
rect 22572 36038 22600 38111
rect 22664 37874 22692 42094
rect 22756 41614 22784 42502
rect 22744 41608 22796 41614
rect 22744 41550 22796 41556
rect 22836 41540 22888 41546
rect 22836 41482 22888 41488
rect 22652 37868 22704 37874
rect 22652 37810 22704 37816
rect 22664 37194 22692 37810
rect 22652 37188 22704 37194
rect 22652 37130 22704 37136
rect 22744 37188 22796 37194
rect 22744 37130 22796 37136
rect 22664 36854 22692 37130
rect 22756 36922 22784 37130
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 22652 36848 22704 36854
rect 22652 36790 22704 36796
rect 22560 36032 22612 36038
rect 22560 35974 22612 35980
rect 22848 35850 22876 41482
rect 22928 41132 22980 41138
rect 22928 41074 22980 41080
rect 22940 40594 22968 41074
rect 22928 40588 22980 40594
rect 22928 40530 22980 40536
rect 22928 39432 22980 39438
rect 22928 39374 22980 39380
rect 22940 38962 22968 39374
rect 22928 38956 22980 38962
rect 22928 38898 22980 38904
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22664 35822 22876 35850
rect 22376 35216 22428 35222
rect 22376 35158 22428 35164
rect 22284 35012 22336 35018
rect 22284 34954 22336 34960
rect 22296 34202 22324 34954
rect 22376 34536 22428 34542
rect 22376 34478 22428 34484
rect 22284 34196 22336 34202
rect 22284 34138 22336 34144
rect 22388 33522 22416 34478
rect 22100 33516 22152 33522
rect 22100 33458 22152 33464
rect 22376 33516 22428 33522
rect 22376 33458 22428 33464
rect 22112 33114 22140 33458
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 22388 32978 22416 33458
rect 22376 32972 22428 32978
rect 22376 32914 22428 32920
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21836 32230 21864 32846
rect 22100 32768 22152 32774
rect 22100 32710 22152 32716
rect 21916 32360 21968 32366
rect 21916 32302 21968 32308
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21928 31822 21956 32302
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21652 30870 21680 31282
rect 21640 30864 21692 30870
rect 21640 30806 21692 30812
rect 21456 30592 21508 30598
rect 21454 30560 21456 30569
rect 21508 30560 21510 30569
rect 21454 30495 21510 30504
rect 21548 29572 21600 29578
rect 21548 29514 21600 29520
rect 21364 28008 21416 28014
rect 21364 27950 21416 27956
rect 21272 27600 21324 27606
rect 21178 27568 21234 27577
rect 21272 27542 21324 27548
rect 21178 27503 21234 27512
rect 21192 27402 21220 27503
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 21376 26926 21404 27950
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21468 27062 21496 27406
rect 21456 27056 21508 27062
rect 21456 26998 21508 27004
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 21364 26920 21416 26926
rect 21364 26862 21416 26868
rect 21008 26586 21036 26862
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 21376 26450 21404 26862
rect 21560 26790 21588 29514
rect 21652 29238 21680 30806
rect 21928 30802 21956 31758
rect 21916 30796 21968 30802
rect 21916 30738 21968 30744
rect 22112 30734 22140 32710
rect 22664 32570 22692 35822
rect 22836 35760 22888 35766
rect 22836 35702 22888 35708
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22756 33862 22784 34886
rect 22848 34066 22876 35702
rect 22836 34060 22888 34066
rect 22836 34002 22888 34008
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22848 33590 22876 34002
rect 22836 33584 22888 33590
rect 22836 33526 22888 33532
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22100 30728 22152 30734
rect 22100 30670 22152 30676
rect 21732 30592 21784 30598
rect 21732 30534 21784 30540
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21744 30326 21772 30534
rect 21732 30320 21784 30326
rect 21732 30262 21784 30268
rect 21744 29646 21772 30262
rect 21836 30258 21864 30534
rect 22112 30394 22140 30670
rect 22388 30598 22416 31622
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 22928 31272 22980 31278
rect 22928 31214 22980 31220
rect 22376 30592 22428 30598
rect 22376 30534 22428 30540
rect 22100 30388 22152 30394
rect 22100 30330 22152 30336
rect 22376 30388 22428 30394
rect 22376 30330 22428 30336
rect 22388 30258 22416 30330
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 21836 29714 21864 30194
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21928 29646 21956 30126
rect 22008 30116 22060 30122
rect 22008 30058 22060 30064
rect 22192 30116 22244 30122
rect 22192 30058 22244 30064
rect 22020 29782 22048 30058
rect 22008 29776 22060 29782
rect 22008 29718 22060 29724
rect 21732 29640 21784 29646
rect 21732 29582 21784 29588
rect 21916 29640 21968 29646
rect 21916 29582 21968 29588
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21914 29200 21970 29209
rect 21652 28558 21680 29174
rect 21914 29135 21916 29144
rect 21968 29135 21970 29144
rect 21916 29106 21968 29112
rect 21928 28558 21956 29106
rect 22008 28960 22060 28966
rect 22008 28902 22060 28908
rect 22020 28558 22048 28902
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 21916 28416 21968 28422
rect 21916 28358 21968 28364
rect 21928 27470 21956 28358
rect 22100 28008 22152 28014
rect 22100 27950 22152 27956
rect 22112 27674 22140 27950
rect 22100 27668 22152 27674
rect 22100 27610 22152 27616
rect 22204 27470 22232 30058
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22296 28422 22324 29514
rect 22388 29238 22416 30194
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22480 28762 22508 31214
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22664 30394 22692 30602
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 22664 30054 22692 30330
rect 22836 30320 22888 30326
rect 22836 30262 22888 30268
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22468 28756 22520 28762
rect 22468 28698 22520 28704
rect 22480 28558 22508 28698
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22284 28416 22336 28422
rect 22284 28358 22336 28364
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21548 26784 21600 26790
rect 21548 26726 21600 26732
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21548 26580 21600 26586
rect 21548 26522 21600 26528
rect 21468 26450 21496 26522
rect 21364 26444 21416 26450
rect 21364 26386 21416 26392
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21560 26330 21588 26522
rect 21468 26314 21588 26330
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21456 26308 21588 26314
rect 21508 26302 21588 26308
rect 21456 26250 21508 26256
rect 21376 26042 21404 26250
rect 21364 26036 21416 26042
rect 21364 25978 21416 25984
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 21272 25968 21324 25974
rect 21272 25910 21324 25916
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21008 24886 21036 25230
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20168 22228 20220 22234
rect 20168 22170 20220 22176
rect 19800 22092 19852 22098
rect 19800 22034 19852 22040
rect 20180 21690 20208 22170
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19720 20874 19748 21286
rect 19708 20868 19760 20874
rect 19708 20810 19760 20816
rect 19628 19306 19748 19334
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19340 18352 19392 18358
rect 19260 18312 19340 18340
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18800 17746 18828 18022
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18708 17338 18736 17682
rect 18892 17338 18920 18226
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 16046 18828 16390
rect 18984 16153 19012 18226
rect 19260 17882 19288 18312
rect 19340 18294 19392 18300
rect 19432 18284 19484 18290
rect 19616 18284 19668 18290
rect 19484 18244 19564 18272
rect 19432 18226 19484 18232
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19260 17678 19288 17818
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19260 17338 19288 17614
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19168 17202 19196 17274
rect 19352 17270 19380 18022
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 18970 16144 19026 16153
rect 19076 16114 19104 17138
rect 19340 17128 19392 17134
rect 19154 17096 19210 17105
rect 19444 17105 19472 17138
rect 19340 17070 19392 17076
rect 19430 17096 19486 17105
rect 19154 17031 19210 17040
rect 19168 16590 19196 17031
rect 19352 16794 19380 17070
rect 19430 17031 19486 17040
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 18970 16079 19026 16088
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18800 15434 18828 15846
rect 19168 15502 19196 16526
rect 19352 15978 19380 16730
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 19444 15434 19472 16594
rect 19536 16250 19564 18244
rect 19616 18226 19668 18232
rect 19628 17542 19656 18226
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19628 16658 19656 17138
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19536 16017 19564 16050
rect 19522 16008 19578 16017
rect 19522 15943 19578 15952
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 19432 15428 19484 15434
rect 19432 15370 19484 15376
rect 19444 15162 19472 15370
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19536 15094 19564 15846
rect 19628 15706 19656 16050
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19524 15088 19576 15094
rect 19524 15030 19576 15036
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18616 14074 18644 14350
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 18064 12646 18092 12786
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 17224 12436 17276 12442
rect 16684 12406 16896 12434
rect 16868 12238 16896 12406
rect 17224 12378 17276 12384
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 16868 11694 16896 12174
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 16868 10606 16896 11630
rect 17972 10810 18000 12106
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17868 10736 17920 10742
rect 17972 10690 18000 10746
rect 17920 10684 18000 10690
rect 17868 10678 18000 10684
rect 17880 10662 18000 10678
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 12912 10266 12940 10542
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 11980 10124 12032 10130
rect 11808 10084 11980 10112
rect 11980 10066 12032 10072
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 6798 10732 7822
rect 11164 7478 11192 8298
rect 11624 7750 11652 9646
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11808 9178 11836 9454
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10244 6390 10272 6666
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10612 6322 10640 6666
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9496 5646 9548 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9232 5086 9352 5114
rect 9324 5030 9352 5086
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9232 4554 9260 4966
rect 9416 4826 9444 5306
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9416 4622 9444 4762
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 3466 8892 4082
rect 9416 4078 9444 4558
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 9416 3194 9444 4014
rect 9508 3602 9536 5646
rect 9600 5630 9720 5658
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9600 5234 9628 5630
rect 9876 5522 9904 5850
rect 9784 5494 9904 5522
rect 9784 5234 9812 5494
rect 9968 5370 9996 6258
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10060 5710 10088 6122
rect 10336 5914 10364 6122
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10600 5704 10652 5710
rect 10704 5692 10732 6734
rect 11072 6322 11100 7210
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 6322 11284 7142
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10652 5664 10732 5692
rect 10600 5646 10652 5652
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9876 5234 9904 5306
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9600 5114 9628 5170
rect 9600 5086 9720 5114
rect 9692 4622 9720 5086
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9600 4214 9628 4490
rect 9876 4282 9904 4966
rect 10060 4826 10088 5170
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9968 4010 9996 4558
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 10152 3534 10180 4082
rect 10244 3534 10272 4966
rect 10612 4690 10640 5646
rect 10888 5642 10916 6054
rect 11256 5914 11284 6258
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11440 5642 11468 6666
rect 11624 6662 11652 7346
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11716 6866 11744 7210
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 6186 11652 6598
rect 11716 6322 11744 6802
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 6322 11928 6394
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11440 5522 11468 5578
rect 11808 5574 11836 6190
rect 11348 5494 11468 5522
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4758 10824 4966
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9784 3126 9812 3334
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10152 2990 10180 3470
rect 10336 3126 10364 4218
rect 10428 4146 10456 4626
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10520 4214 10548 4558
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3534 10548 3878
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10612 3194 10640 4626
rect 11348 4554 11376 5494
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 3602 11192 4422
rect 11348 4282 11376 4490
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11256 3738 11284 3946
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11532 3534 11560 5510
rect 11992 5302 12020 10066
rect 13556 9926 13584 10542
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13556 9722 13584 9862
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7002 12112 7346
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6322 12112 6938
rect 12176 6390 12204 7142
rect 12360 6662 12388 7278
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6458 12388 6598
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12360 5914 12388 6394
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 12452 5030 12480 9590
rect 16868 8498 16896 10542
rect 17972 9994 18000 10662
rect 18156 10130 18184 12854
rect 18248 12102 18276 13126
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18616 11898 18644 13126
rect 18800 12918 18828 14214
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 18984 13190 19012 13806
rect 19444 13326 19472 14758
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13530 19564 13806
rect 19720 13802 19748 19306
rect 19904 18290 19932 21354
rect 19984 20800 20036 20806
rect 19984 20742 20036 20748
rect 20444 20800 20496 20806
rect 20444 20742 20496 20748
rect 19996 19854 20024 20742
rect 20456 20534 20484 20742
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20272 18970 20300 19246
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19904 17678 19932 18226
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19904 17270 19932 17614
rect 19892 17264 19944 17270
rect 19892 17206 19944 17212
rect 20088 17202 20116 18090
rect 20364 17678 20392 18158
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20088 16454 20116 17138
rect 20180 16998 20208 17478
rect 20364 17202 20392 17614
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20180 16182 20208 16730
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19904 15366 19932 16050
rect 19996 15978 20024 16118
rect 20166 16008 20222 16017
rect 19984 15972 20036 15978
rect 20166 15943 20222 15952
rect 19984 15914 20036 15920
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 14414 19932 15302
rect 19996 15026 20024 15914
rect 20180 15026 20208 15943
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19432 13320 19484 13326
rect 19720 13274 19748 13466
rect 19432 13262 19484 13268
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12918 19012 13126
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 19260 12866 19288 12922
rect 19260 12838 19380 12866
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19260 12306 19288 12718
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18524 11354 18552 11766
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18340 10266 18368 10542
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18524 10010 18552 11290
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18800 10810 18828 11086
rect 19352 11082 19380 12838
rect 19444 11218 19472 13262
rect 19628 13258 19748 13274
rect 19616 13252 19748 13258
rect 19668 13246 19748 13252
rect 19616 13194 19668 13200
rect 19706 12744 19762 12753
rect 19706 12679 19762 12688
rect 19720 12646 19748 12679
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19812 12306 19840 14010
rect 20364 14006 20392 17002
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20456 16182 20484 16390
rect 20548 16182 20576 18634
rect 20732 18408 20760 22714
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 20942 20852 21286
rect 21008 21146 21036 24142
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21100 23526 21128 23666
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20916 19718 20944 20334
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20640 18380 20760 18408
rect 20640 17066 20668 18380
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20732 17746 20760 18226
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20628 17060 20680 17066
rect 20628 17002 20680 17008
rect 20732 16266 20760 17682
rect 20824 17338 20852 17818
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20824 16658 20852 17274
rect 20916 17082 20944 19654
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17202 21036 17614
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20916 17054 21036 17082
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20916 16590 20944 16934
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 21008 16402 21036 17054
rect 20640 16238 20760 16266
rect 20916 16374 21036 16402
rect 20444 16176 20496 16182
rect 20444 16118 20496 16124
rect 20536 16176 20588 16182
rect 20536 16118 20588 16124
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 19904 12646 19932 13942
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19996 12986 20024 13194
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 20180 12918 20208 13806
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20168 12776 20220 12782
rect 20272 12764 20300 13806
rect 20220 12736 20300 12764
rect 20168 12718 20220 12724
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19536 11762 19564 12038
rect 20088 11762 20116 12038
rect 20180 11830 20208 12718
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19536 11150 19564 11562
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18892 10742 18920 10950
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 19536 10470 19564 11086
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 19156 10464 19208 10470
rect 19524 10464 19576 10470
rect 19208 10424 19288 10452
rect 19156 10406 19208 10412
rect 19260 10130 19288 10424
rect 19524 10406 19576 10412
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 18604 10056 18656 10062
rect 18524 10004 18604 10010
rect 18524 9998 18656 10004
rect 17960 9988 18012 9994
rect 18524 9982 18644 9998
rect 17960 9930 18012 9936
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 16856 8492 16908 8498
rect 18248 8480 18276 9862
rect 19536 9042 19564 10406
rect 19628 9994 19656 11018
rect 20180 10985 20208 11018
rect 20166 10976 20222 10985
rect 20166 10911 20222 10920
rect 20272 10742 20300 12582
rect 20456 12238 20484 15982
rect 20640 15570 20668 16238
rect 20812 15904 20864 15910
rect 20812 15846 20864 15852
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 14346 20668 15506
rect 20824 15434 20852 15846
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20732 14958 20760 15098
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14482 20760 14758
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20548 12646 20576 14214
rect 20640 13410 20668 14282
rect 20824 13938 20852 15098
rect 20812 13932 20864 13938
rect 20812 13874 20864 13880
rect 20916 13870 20944 16374
rect 20996 15428 21048 15434
rect 20996 15370 21048 15376
rect 21008 14346 21036 15370
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20640 13394 20760 13410
rect 20640 13388 20772 13394
rect 20640 13382 20720 13388
rect 20720 13330 20772 13336
rect 20536 12640 20588 12646
rect 20536 12582 20588 12588
rect 20548 12306 20576 12582
rect 20720 12436 20772 12442
rect 21008 12434 21036 13874
rect 21100 12986 21128 23462
rect 21284 22094 21312 25910
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 21560 25498 21588 25774
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21744 24954 21772 25230
rect 21732 24948 21784 24954
rect 21732 24890 21784 24896
rect 21456 24812 21508 24818
rect 21456 24754 21508 24760
rect 21468 24410 21496 24754
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21744 24410 21772 24686
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 21376 22778 21404 23598
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21284 22066 21404 22094
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 21554 21220 21830
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21192 21078 21220 21286
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21192 15178 21220 19382
rect 21284 18766 21312 20198
rect 21376 19310 21404 22066
rect 21640 22024 21692 22030
rect 21638 21992 21640 22001
rect 21692 21992 21694 22001
rect 21638 21927 21694 21936
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21456 21616 21508 21622
rect 21456 21558 21508 21564
rect 21468 20534 21496 21558
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 21560 20330 21588 20810
rect 21652 20398 21680 21422
rect 21744 21350 21772 21830
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21376 18630 21404 19246
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21284 17542 21312 17614
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 17066 21312 17478
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21376 16946 21404 18362
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21468 17678 21496 17750
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17338 21496 17614
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21652 17218 21680 20334
rect 21744 18306 21772 20470
rect 21836 20262 21864 27270
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22112 25498 22140 25638
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22296 25294 22324 28358
rect 22572 28014 22600 28426
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21928 22098 21956 23530
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 22020 23050 22048 23462
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21928 20806 21956 22034
rect 22112 21350 22140 22510
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22112 20874 22140 21286
rect 22204 21010 22232 21490
rect 22296 21146 22324 25230
rect 22388 23866 22416 27406
rect 22664 25362 22692 29990
rect 22756 29850 22784 29990
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 22848 29782 22876 30262
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 22756 27606 22784 29582
rect 22940 29238 22968 31214
rect 23032 29714 23060 43250
rect 24032 43104 24084 43110
rect 24032 43046 24084 43052
rect 24044 42702 24072 43046
rect 24032 42696 24084 42702
rect 24032 42638 24084 42644
rect 23664 42628 23716 42634
rect 23664 42570 23716 42576
rect 23296 42152 23348 42158
rect 23296 42094 23348 42100
rect 23308 41818 23336 42094
rect 23296 41812 23348 41818
rect 23296 41754 23348 41760
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 23400 40186 23428 41074
rect 23388 40180 23440 40186
rect 23388 40122 23440 40128
rect 23112 40044 23164 40050
rect 23112 39986 23164 39992
rect 23124 39642 23152 39986
rect 23204 39976 23256 39982
rect 23204 39918 23256 39924
rect 23112 39636 23164 39642
rect 23112 39578 23164 39584
rect 23216 39574 23244 39918
rect 23204 39568 23256 39574
rect 23204 39510 23256 39516
rect 23572 39296 23624 39302
rect 23572 39238 23624 39244
rect 23584 38826 23612 39238
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 23572 37664 23624 37670
rect 23572 37606 23624 37612
rect 23584 36922 23612 37606
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23204 36848 23256 36854
rect 23204 36790 23256 36796
rect 23112 36712 23164 36718
rect 23112 36654 23164 36660
rect 23124 35630 23152 36654
rect 23216 35766 23244 36790
rect 23480 36644 23532 36650
rect 23480 36586 23532 36592
rect 23204 35760 23256 35766
rect 23204 35702 23256 35708
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 23112 35624 23164 35630
rect 23112 35566 23164 35572
rect 23308 35290 23336 35634
rect 23296 35284 23348 35290
rect 23296 35226 23348 35232
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23204 35012 23256 35018
rect 23204 34954 23256 34960
rect 23216 34610 23244 34954
rect 23296 34672 23348 34678
rect 23296 34614 23348 34620
rect 23204 34604 23256 34610
rect 23204 34546 23256 34552
rect 23112 33924 23164 33930
rect 23112 33866 23164 33872
rect 23204 33924 23256 33930
rect 23204 33866 23256 33872
rect 23124 33658 23152 33866
rect 23112 33652 23164 33658
rect 23112 33594 23164 33600
rect 23216 33130 23244 33866
rect 23124 33102 23244 33130
rect 23020 29708 23072 29714
rect 23020 29650 23072 29656
rect 22928 29232 22980 29238
rect 22848 29192 22928 29220
rect 22848 28626 22876 29192
rect 22928 29174 22980 29180
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22848 28218 22876 28562
rect 23032 28422 23060 29650
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 22836 28212 22888 28218
rect 22836 28154 22888 28160
rect 22836 28008 22888 28014
rect 22888 27968 22968 27996
rect 22836 27950 22888 27956
rect 22744 27600 22796 27606
rect 22744 27542 22796 27548
rect 22940 27062 22968 27968
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22940 26314 22968 26998
rect 22928 26308 22980 26314
rect 22928 26250 22980 26256
rect 22836 26036 22888 26042
rect 22836 25978 22888 25984
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22848 25294 22876 25978
rect 22468 25288 22520 25294
rect 22468 25230 22520 25236
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 22480 24954 22508 25230
rect 22468 24948 22520 24954
rect 22468 24890 22520 24896
rect 22848 24274 22876 25230
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22940 23798 22968 26250
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25702 23060 26182
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 23032 24206 23060 25230
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 22928 23792 22980 23798
rect 22928 23734 22980 23740
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22480 22030 22508 23598
rect 23124 23322 23152 33102
rect 23204 32564 23256 32570
rect 23204 32506 23256 32512
rect 23216 29646 23244 32506
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 23216 29306 23244 29446
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 23308 28642 23336 34614
rect 23400 34474 23428 35090
rect 23492 34746 23520 36586
rect 23480 34740 23532 34746
rect 23480 34682 23532 34688
rect 23388 34468 23440 34474
rect 23388 34410 23440 34416
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23400 33386 23428 33798
rect 23388 33380 23440 33386
rect 23388 33322 23440 33328
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23492 32910 23520 33254
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23388 32836 23440 32842
rect 23388 32778 23440 32784
rect 23400 32570 23428 32778
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23492 31414 23520 31622
rect 23480 31408 23532 31414
rect 23480 31350 23532 31356
rect 23676 30938 23704 42570
rect 24032 42560 24084 42566
rect 24032 42502 24084 42508
rect 24044 42226 24072 42502
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 24412 42022 24440 43318
rect 24584 43308 24636 43314
rect 24584 43250 24636 43256
rect 26148 43308 26200 43314
rect 26148 43250 26200 43256
rect 28356 43308 28408 43314
rect 28356 43250 28408 43256
rect 24596 42362 24624 43250
rect 24676 43240 24728 43246
rect 24676 43182 24728 43188
rect 24688 42362 24716 43182
rect 26160 42906 26188 43250
rect 28080 43104 28132 43110
rect 28080 43046 28132 43052
rect 26148 42900 26200 42906
rect 26148 42842 26200 42848
rect 24768 42764 24820 42770
rect 24768 42706 24820 42712
rect 27620 42764 27672 42770
rect 27620 42706 27672 42712
rect 24584 42356 24636 42362
rect 24584 42298 24636 42304
rect 24676 42356 24728 42362
rect 24676 42298 24728 42304
rect 24400 42016 24452 42022
rect 24400 41958 24452 41964
rect 24032 41676 24084 41682
rect 24032 41618 24084 41624
rect 23756 41472 23808 41478
rect 23756 41414 23808 41420
rect 23768 41274 23796 41414
rect 23756 41268 23808 41274
rect 23756 41210 23808 41216
rect 24044 41206 24072 41618
rect 24412 41614 24440 41958
rect 24400 41608 24452 41614
rect 24400 41550 24452 41556
rect 24688 41546 24716 42298
rect 24676 41540 24728 41546
rect 24676 41482 24728 41488
rect 24032 41200 24084 41206
rect 23754 41168 23810 41177
rect 24032 41142 24084 41148
rect 24780 41138 24808 42706
rect 25688 42696 25740 42702
rect 25608 42656 25688 42684
rect 25608 42226 25636 42656
rect 25688 42638 25740 42644
rect 26608 42628 26660 42634
rect 26608 42570 26660 42576
rect 26620 42362 26648 42570
rect 26608 42356 26660 42362
rect 26608 42298 26660 42304
rect 25596 42220 25648 42226
rect 25596 42162 25648 42168
rect 27436 42220 27488 42226
rect 27436 42162 27488 42168
rect 25320 42016 25372 42022
rect 25320 41958 25372 41964
rect 23754 41103 23756 41112
rect 23808 41103 23810 41112
rect 24768 41132 24820 41138
rect 23756 41074 23808 41080
rect 24768 41074 24820 41080
rect 25044 41064 25096 41070
rect 25044 41006 25096 41012
rect 25056 40730 25084 41006
rect 25044 40724 25096 40730
rect 25044 40666 25096 40672
rect 25044 40044 25096 40050
rect 25044 39986 25096 39992
rect 24320 39630 24716 39658
rect 25056 39642 25084 39986
rect 25136 39976 25188 39982
rect 25136 39918 25188 39924
rect 25148 39642 25176 39918
rect 23848 39568 23900 39574
rect 23900 39528 24164 39556
rect 23848 39510 23900 39516
rect 23756 39432 23808 39438
rect 23756 39374 23808 39380
rect 24032 39432 24084 39438
rect 24032 39374 24084 39380
rect 23768 39098 23796 39374
rect 24044 39302 24072 39374
rect 24136 39370 24164 39528
rect 24320 39506 24348 39630
rect 24688 39574 24716 39630
rect 25044 39636 25096 39642
rect 25044 39578 25096 39584
rect 25136 39636 25188 39642
rect 25136 39578 25188 39584
rect 24676 39568 24728 39574
rect 24676 39510 24728 39516
rect 25228 39568 25280 39574
rect 25228 39510 25280 39516
rect 24308 39500 24360 39506
rect 24308 39442 24360 39448
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 24124 39364 24176 39370
rect 24124 39306 24176 39312
rect 24032 39296 24084 39302
rect 24032 39238 24084 39244
rect 24596 39098 24624 39374
rect 25240 39098 25268 39510
rect 23756 39092 23808 39098
rect 23756 39034 23808 39040
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 25228 39092 25280 39098
rect 25228 39034 25280 39040
rect 23756 38956 23808 38962
rect 23756 38898 23808 38904
rect 23940 38956 23992 38962
rect 23940 38898 23992 38904
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 23768 38554 23796 38898
rect 23952 38554 23980 38898
rect 24124 38888 24176 38894
rect 24124 38830 24176 38836
rect 23756 38548 23808 38554
rect 23756 38490 23808 38496
rect 23940 38548 23992 38554
rect 23940 38490 23992 38496
rect 23940 38276 23992 38282
rect 23940 38218 23992 38224
rect 23952 36242 23980 38218
rect 24136 37874 24164 38830
rect 25148 38214 25176 38898
rect 25240 38554 25268 38898
rect 25228 38548 25280 38554
rect 25228 38490 25280 38496
rect 25136 38208 25188 38214
rect 25136 38150 25188 38156
rect 24124 37868 24176 37874
rect 24124 37810 24176 37816
rect 24136 37466 24164 37810
rect 24124 37460 24176 37466
rect 24124 37402 24176 37408
rect 25044 37324 25096 37330
rect 25044 37266 25096 37272
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24412 37126 24440 37198
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24412 36854 24440 37062
rect 25056 36922 25084 37266
rect 25136 37188 25188 37194
rect 25136 37130 25188 37136
rect 25044 36916 25096 36922
rect 25044 36858 25096 36864
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 23940 36236 23992 36242
rect 23940 36178 23992 36184
rect 24032 36032 24084 36038
rect 24032 35974 24084 35980
rect 24044 35562 24072 35974
rect 24032 35556 24084 35562
rect 24032 35498 24084 35504
rect 24032 35148 24084 35154
rect 24032 35090 24084 35096
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23940 34944 23992 34950
rect 23940 34886 23992 34892
rect 23860 34542 23888 34886
rect 23952 34746 23980 34886
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23860 33114 23888 34478
rect 23952 34202 23980 34682
rect 24044 34542 24072 35090
rect 24032 34536 24084 34542
rect 24032 34478 24084 34484
rect 23940 34196 23992 34202
rect 23940 34138 23992 34144
rect 24044 34105 24072 34478
rect 24308 34400 24360 34406
rect 24308 34342 24360 34348
rect 24030 34096 24086 34105
rect 24030 34031 24086 34040
rect 24320 33658 24348 34342
rect 24308 33652 24360 33658
rect 24308 33594 24360 33600
rect 23940 33584 23992 33590
rect 23940 33526 23992 33532
rect 23848 33108 23900 33114
rect 23848 33050 23900 33056
rect 23756 31816 23808 31822
rect 23756 31758 23808 31764
rect 23848 31816 23900 31822
rect 23848 31758 23900 31764
rect 23768 30938 23796 31758
rect 23860 31482 23888 31758
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23756 30728 23808 30734
rect 23756 30670 23808 30676
rect 23768 30054 23796 30670
rect 23860 30666 23888 31214
rect 23848 30660 23900 30666
rect 23848 30602 23900 30608
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23400 29322 23428 29582
rect 23400 29294 23520 29322
rect 23388 29164 23440 29170
rect 23388 29106 23440 29112
rect 23216 28614 23336 28642
rect 23216 28234 23244 28614
rect 23216 28206 23336 28234
rect 23400 28218 23428 29106
rect 23492 29102 23520 29294
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 23308 27470 23336 28206
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23296 27464 23348 27470
rect 23216 27424 23296 27452
rect 23216 26518 23244 27424
rect 23296 27406 23348 27412
rect 23400 27334 23428 28154
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23296 26852 23348 26858
rect 23296 26794 23348 26800
rect 23204 26512 23256 26518
rect 23204 26454 23256 26460
rect 23216 26042 23244 26454
rect 23308 26042 23336 26794
rect 23204 26036 23256 26042
rect 23204 25978 23256 25984
rect 23296 26036 23348 26042
rect 23296 25978 23348 25984
rect 23308 25294 23336 25978
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23400 24886 23428 25842
rect 23480 25832 23532 25838
rect 23478 25800 23480 25809
rect 23572 25832 23624 25838
rect 23532 25800 23534 25809
rect 23572 25774 23624 25780
rect 23478 25735 23534 25744
rect 23492 25362 23520 25735
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23492 24750 23520 25298
rect 23584 24857 23612 25774
rect 23664 25696 23716 25702
rect 23664 25638 23716 25644
rect 23676 25294 23704 25638
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23570 24848 23626 24857
rect 23570 24783 23572 24792
rect 23624 24783 23626 24792
rect 23572 24754 23624 24760
rect 23480 24744 23532 24750
rect 23202 24712 23258 24721
rect 23480 24686 23532 24692
rect 23202 24647 23258 24656
rect 23216 24274 23244 24647
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23584 23594 23612 24754
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22572 21962 22600 22374
rect 22848 22098 22876 22918
rect 22928 22432 22980 22438
rect 22928 22374 22980 22380
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22560 21956 22612 21962
rect 22560 21898 22612 21904
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 22100 20596 22152 20602
rect 22204 20584 22232 20946
rect 22296 20602 22324 21082
rect 22152 20556 22232 20584
rect 22284 20596 22336 20602
rect 22100 20538 22152 20544
rect 22284 20538 22336 20544
rect 22112 20330 22140 20538
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 22112 19446 22140 20266
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 21836 18426 21864 19178
rect 22112 18698 22140 19382
rect 22296 19174 22324 20402
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22388 19514 22416 20334
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 18902 22324 19110
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22100 18692 22152 18698
rect 22100 18634 22152 18640
rect 22112 18426 22140 18634
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 21744 18278 21864 18306
rect 21732 17740 21784 17746
rect 21732 17682 21784 17688
rect 21744 17542 21772 17682
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21560 17202 21680 17218
rect 21548 17196 21680 17202
rect 21600 17190 21680 17196
rect 21548 17138 21600 17144
rect 21284 16918 21404 16946
rect 21284 15314 21312 16918
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21468 15570 21496 15982
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21284 15286 21404 15314
rect 21192 15150 21312 15178
rect 21376 15162 21404 15286
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21192 13326 21220 14282
rect 21284 14006 21312 15150
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21468 15026 21496 15506
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21272 14000 21324 14006
rect 21272 13942 21324 13948
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21272 13796 21324 13802
rect 21272 13738 21324 13744
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12986 21220 13262
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21284 12918 21312 13738
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21560 13394 21588 13670
rect 21652 13530 21680 13874
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21652 12918 21680 13466
rect 21272 12912 21324 12918
rect 21272 12854 21324 12860
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21284 12782 21312 12854
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 20720 12378 20772 12384
rect 20824 12406 21036 12434
rect 21836 12434 21864 18278
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 16114 21956 18022
rect 22204 17882 22232 18226
rect 22284 18216 22336 18222
rect 22388 18170 22416 19450
rect 22336 18164 22416 18170
rect 22284 18158 22416 18164
rect 22296 18142 22416 18158
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22008 17196 22060 17202
rect 22008 17138 22060 17144
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22020 15026 22048 17138
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 14618 22048 14962
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 22480 14074 22508 19994
rect 22572 18850 22600 21898
rect 22940 21554 22968 22374
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 23216 20534 23244 21286
rect 23204 20528 23256 20534
rect 23204 20470 23256 20476
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 22572 18822 22692 18850
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22572 18426 22600 18634
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22664 18290 22692 18822
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22572 17814 22600 18226
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 14346 22692 15302
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12782 22508 13126
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 21836 12406 22048 12434
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20548 11830 20576 12106
rect 20536 11824 20588 11830
rect 20536 11766 20588 11772
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20180 10266 20208 10542
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19524 9036 19576 9042
rect 19524 8978 19576 8984
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 18328 8492 18380 8498
rect 18248 8452 18328 8480
rect 16856 8434 16908 8440
rect 18328 8434 18380 8440
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19168 7546 19196 8366
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19352 7954 19380 8298
rect 19444 8090 19472 8910
rect 19536 8634 19564 8978
rect 19628 8906 19656 9930
rect 19616 8900 19668 8906
rect 19616 8842 19668 8848
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19432 7404 19484 7410
rect 19536 7392 19564 8570
rect 19720 7410 19748 10202
rect 20272 10062 20300 10678
rect 20456 10674 20484 11154
rect 20548 10810 20576 11766
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 20548 10062 20576 10746
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19812 7478 19840 9862
rect 20272 9110 20300 9998
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20364 8566 20392 8774
rect 20732 8566 20760 12378
rect 20824 11014 20852 12406
rect 21362 12336 21418 12345
rect 21362 12271 21418 12280
rect 21376 12238 21404 12271
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21100 11558 21128 12174
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20902 10976 20958 10985
rect 20824 9042 20852 10950
rect 20902 10911 20958 10920
rect 20916 10810 20944 10911
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21100 10674 21128 11494
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21192 9994 21220 10474
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21192 9674 21220 9930
rect 21284 9926 21312 12106
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21376 11354 21404 11766
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21468 11354 21496 11630
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21376 10742 21404 11290
rect 21652 11218 21680 12038
rect 21836 11762 21864 12038
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21640 11212 21692 11218
rect 21640 11154 21692 11160
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 22020 10266 22048 12406
rect 22756 12306 22784 12718
rect 23032 12434 23060 20198
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23124 18698 23152 18906
rect 23112 18692 23164 18698
rect 23112 18634 23164 18640
rect 23124 15094 23152 18634
rect 23216 15570 23244 19110
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 23308 15162 23336 23258
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23492 21146 23520 21490
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23768 20942 23796 29990
rect 23860 28150 23888 30602
rect 23952 30258 23980 33526
rect 24032 33448 24084 33454
rect 24032 33390 24084 33396
rect 24044 32366 24072 33390
rect 24124 32904 24176 32910
rect 24124 32846 24176 32852
rect 24136 32502 24164 32846
rect 24504 32842 24532 36722
rect 25148 36310 25176 37130
rect 25136 36304 25188 36310
rect 25136 36246 25188 36252
rect 24584 36032 24636 36038
rect 24584 35974 24636 35980
rect 24596 35834 24624 35974
rect 24584 35828 24636 35834
rect 24584 35770 24636 35776
rect 24768 35624 24820 35630
rect 24768 35566 24820 35572
rect 24780 35290 24808 35566
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 25228 34944 25280 34950
rect 25228 34886 25280 34892
rect 25240 34746 25268 34886
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 25044 33924 25096 33930
rect 25044 33866 25096 33872
rect 25056 33658 25084 33866
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 24492 32836 24544 32842
rect 24492 32778 24544 32784
rect 24400 32768 24452 32774
rect 24400 32710 24452 32716
rect 24412 32570 24440 32710
rect 24400 32564 24452 32570
rect 24400 32506 24452 32512
rect 24124 32496 24176 32502
rect 24124 32438 24176 32444
rect 24032 32360 24084 32366
rect 24032 32302 24084 32308
rect 24124 32360 24176 32366
rect 24124 32302 24176 32308
rect 24136 31822 24164 32302
rect 24124 31816 24176 31822
rect 24124 31758 24176 31764
rect 24136 31226 24164 31758
rect 24400 31272 24452 31278
rect 24136 31210 24256 31226
rect 24400 31214 24452 31220
rect 24136 31204 24268 31210
rect 24136 31198 24216 31204
rect 24216 31146 24268 31152
rect 24308 31136 24360 31142
rect 24308 31078 24360 31084
rect 24032 30728 24084 30734
rect 24032 30670 24084 30676
rect 23940 30252 23992 30258
rect 23940 30194 23992 30200
rect 23848 28144 23900 28150
rect 23848 28086 23900 28092
rect 23848 25832 23900 25838
rect 23952 25820 23980 30194
rect 23900 25792 23980 25820
rect 23848 25774 23900 25780
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23860 25498 23888 25638
rect 23848 25492 23900 25498
rect 23848 25434 23900 25440
rect 23860 25362 23888 25434
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23860 24750 23888 25298
rect 23940 25288 23992 25294
rect 24044 25276 24072 30670
rect 24124 30592 24176 30598
rect 24124 30534 24176 30540
rect 24136 29578 24164 30534
rect 24320 30190 24348 31078
rect 24412 30734 24440 31214
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24308 30184 24360 30190
rect 24228 30144 24308 30172
rect 24124 29572 24176 29578
rect 24124 29514 24176 29520
rect 24124 28076 24176 28082
rect 24124 28018 24176 28024
rect 24136 27470 24164 28018
rect 24228 27606 24256 30144
rect 24308 30126 24360 30132
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24308 29164 24360 29170
rect 24308 29106 24360 29112
rect 24320 27985 24348 29106
rect 24412 28150 24440 29446
rect 24504 29238 24532 32778
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 25056 32026 25084 32370
rect 25044 32020 25096 32026
rect 25044 31962 25096 31968
rect 25332 31482 25360 41958
rect 25504 41540 25556 41546
rect 25504 41482 25556 41488
rect 25516 40458 25544 41482
rect 25608 41070 25636 42162
rect 27344 42152 27396 42158
rect 27344 42094 27396 42100
rect 26884 42016 26936 42022
rect 26884 41958 26936 41964
rect 26896 41682 26924 41958
rect 27356 41818 27384 42094
rect 27448 41818 27476 42162
rect 27632 42140 27660 42706
rect 27896 42696 27948 42702
rect 27896 42638 27948 42644
rect 27712 42152 27764 42158
rect 27632 42112 27712 42140
rect 27344 41812 27396 41818
rect 27344 41754 27396 41760
rect 27436 41812 27488 41818
rect 27436 41754 27488 41760
rect 27632 41682 27660 42112
rect 27712 42094 27764 42100
rect 26884 41676 26936 41682
rect 26884 41618 26936 41624
rect 27344 41676 27396 41682
rect 27344 41618 27396 41624
rect 27620 41676 27672 41682
rect 27620 41618 27672 41624
rect 25872 41608 25924 41614
rect 25872 41550 25924 41556
rect 25964 41608 26016 41614
rect 25964 41550 26016 41556
rect 26056 41608 26108 41614
rect 27068 41608 27120 41614
rect 26108 41568 26372 41596
rect 26056 41550 26108 41556
rect 25688 41472 25740 41478
rect 25688 41414 25740 41420
rect 25596 41064 25648 41070
rect 25596 41006 25648 41012
rect 25700 40594 25728 41414
rect 25884 41274 25912 41550
rect 25872 41268 25924 41274
rect 25872 41210 25924 41216
rect 25780 41064 25832 41070
rect 25780 41006 25832 41012
rect 25688 40588 25740 40594
rect 25688 40530 25740 40536
rect 25504 40452 25556 40458
rect 25504 40394 25556 40400
rect 25688 38956 25740 38962
rect 25688 38898 25740 38904
rect 25700 38554 25728 38898
rect 25596 38548 25648 38554
rect 25596 38490 25648 38496
rect 25688 38548 25740 38554
rect 25688 38490 25740 38496
rect 25608 38418 25636 38490
rect 25596 38412 25648 38418
rect 25596 38354 25648 38360
rect 25700 38350 25728 38490
rect 25412 38344 25464 38350
rect 25412 38286 25464 38292
rect 25688 38344 25740 38350
rect 25688 38286 25740 38292
rect 25424 37738 25452 38286
rect 25412 37732 25464 37738
rect 25412 37674 25464 37680
rect 25792 37262 25820 41006
rect 25884 40730 25912 41210
rect 25976 41018 26004 41550
rect 25976 40990 26188 41018
rect 26160 40934 26188 40990
rect 26148 40928 26200 40934
rect 26148 40870 26200 40876
rect 26240 40928 26292 40934
rect 26240 40870 26292 40876
rect 25872 40724 25924 40730
rect 25872 40666 25924 40672
rect 25884 40440 25912 40666
rect 25962 40624 26018 40633
rect 25962 40559 25964 40568
rect 26016 40559 26018 40568
rect 25964 40530 26016 40536
rect 26160 40526 26188 40870
rect 26252 40633 26280 40870
rect 26238 40624 26294 40633
rect 26238 40559 26294 40568
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 26056 40452 26108 40458
rect 25884 40412 26056 40440
rect 26056 40394 26108 40400
rect 26068 40186 26096 40394
rect 26240 40384 26292 40390
rect 26344 40372 26372 41568
rect 27068 41550 27120 41556
rect 27080 41414 27108 41550
rect 27356 41414 27384 41618
rect 27080 41386 27384 41414
rect 27356 41274 27384 41386
rect 27344 41268 27396 41274
rect 27344 41210 27396 41216
rect 27632 41206 27660 41618
rect 27804 41540 27856 41546
rect 27804 41482 27856 41488
rect 27620 41200 27672 41206
rect 27620 41142 27672 41148
rect 27816 40594 27844 41482
rect 27804 40588 27856 40594
rect 27804 40530 27856 40536
rect 26292 40344 26372 40372
rect 26240 40326 26292 40332
rect 26056 40180 26108 40186
rect 26056 40122 26108 40128
rect 26252 40118 26280 40326
rect 26240 40112 26292 40118
rect 26240 40054 26292 40060
rect 26516 40044 26568 40050
rect 26516 39986 26568 39992
rect 26528 39642 26556 39986
rect 26792 39976 26844 39982
rect 26792 39918 26844 39924
rect 26804 39642 26832 39918
rect 27816 39914 27844 40530
rect 27804 39908 27856 39914
rect 27804 39850 27856 39856
rect 26516 39636 26568 39642
rect 26516 39578 26568 39584
rect 26792 39636 26844 39642
rect 26792 39578 26844 39584
rect 27252 39568 27304 39574
rect 27252 39510 27304 39516
rect 27160 39432 27212 39438
rect 27160 39374 27212 39380
rect 25964 39364 26016 39370
rect 25964 39306 26016 39312
rect 25976 38894 26004 39306
rect 27172 39302 27200 39374
rect 27160 39296 27212 39302
rect 27160 39238 27212 39244
rect 27172 39030 27200 39238
rect 27160 39024 27212 39030
rect 27160 38966 27212 38972
rect 25964 38888 26016 38894
rect 25964 38830 26016 38836
rect 25976 38486 26004 38830
rect 27264 38826 27292 39510
rect 27528 39432 27580 39438
rect 27580 39392 27660 39420
rect 27528 39374 27580 39380
rect 27528 38956 27580 38962
rect 27632 38944 27660 39392
rect 27580 38916 27660 38944
rect 27528 38898 27580 38904
rect 27252 38820 27304 38826
rect 27252 38762 27304 38768
rect 25964 38480 26016 38486
rect 25964 38422 26016 38428
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26056 38208 26108 38214
rect 26056 38150 26108 38156
rect 26068 37466 26096 38150
rect 26056 37460 26108 37466
rect 26056 37402 26108 37408
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 25596 36712 25648 36718
rect 25596 36654 25648 36660
rect 25412 35556 25464 35562
rect 25412 35498 25464 35504
rect 25424 35086 25452 35498
rect 25608 35154 25636 36654
rect 25792 36650 25820 37198
rect 26056 36848 26108 36854
rect 26056 36790 26108 36796
rect 25780 36644 25832 36650
rect 25780 36586 25832 36592
rect 25792 35766 25820 36586
rect 25780 35760 25832 35766
rect 25780 35702 25832 35708
rect 25596 35148 25648 35154
rect 25596 35090 25648 35096
rect 25412 35080 25464 35086
rect 25412 35022 25464 35028
rect 26068 34746 26096 36790
rect 26160 35630 26188 38286
rect 27632 38010 27660 38916
rect 27908 38026 27936 42638
rect 28092 42294 28120 43046
rect 28368 42906 28396 43250
rect 28356 42900 28408 42906
rect 28356 42842 28408 42848
rect 28264 42560 28316 42566
rect 28264 42502 28316 42508
rect 28276 42362 28304 42502
rect 28264 42356 28316 42362
rect 28264 42298 28316 42304
rect 28080 42288 28132 42294
rect 28080 42230 28132 42236
rect 28172 41608 28224 41614
rect 28172 41550 28224 41556
rect 28184 41070 28212 41550
rect 28172 41064 28224 41070
rect 28172 41006 28224 41012
rect 28172 40520 28224 40526
rect 28172 40462 28224 40468
rect 28184 39642 28212 40462
rect 28172 39636 28224 39642
rect 28172 39578 28224 39584
rect 27988 38888 28040 38894
rect 27988 38830 28040 38836
rect 27620 38004 27672 38010
rect 27620 37946 27672 37952
rect 27816 37998 27936 38026
rect 28000 38010 28028 38830
rect 28172 38344 28224 38350
rect 28172 38286 28224 38292
rect 27988 38004 28040 38010
rect 27068 37868 27120 37874
rect 27068 37810 27120 37816
rect 26332 37460 26384 37466
rect 26332 37402 26384 37408
rect 26344 36786 26372 37402
rect 26516 37188 26568 37194
rect 26516 37130 26568 37136
rect 26528 36922 26556 37130
rect 26516 36916 26568 36922
rect 26516 36858 26568 36864
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 27080 36106 27108 37810
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27712 36780 27764 36786
rect 27712 36722 27764 36728
rect 27344 36712 27396 36718
rect 27344 36654 27396 36660
rect 27356 36310 27384 36654
rect 27344 36304 27396 36310
rect 27344 36246 27396 36252
rect 27068 36100 27120 36106
rect 27068 36042 27120 36048
rect 26148 35624 26200 35630
rect 26148 35566 26200 35572
rect 26976 35624 27028 35630
rect 26976 35566 27028 35572
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 26160 35018 26188 35430
rect 26148 35012 26200 35018
rect 26148 34954 26200 34960
rect 26056 34740 26108 34746
rect 26056 34682 26108 34688
rect 26148 34672 26200 34678
rect 26148 34614 26200 34620
rect 25688 34536 25740 34542
rect 25688 34478 25740 34484
rect 25700 34134 25728 34478
rect 25688 34128 25740 34134
rect 25688 34070 25740 34076
rect 26056 33856 26108 33862
rect 26056 33798 26108 33804
rect 26068 33658 26096 33798
rect 26056 33652 26108 33658
rect 26056 33594 26108 33600
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 25780 33448 25832 33454
rect 25780 33390 25832 33396
rect 25688 32768 25740 32774
rect 25688 32710 25740 32716
rect 25700 31890 25728 32710
rect 25792 31890 25820 33390
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 25688 31884 25740 31890
rect 25688 31826 25740 31832
rect 25780 31884 25832 31890
rect 25780 31826 25832 31832
rect 25136 31476 25188 31482
rect 25136 31418 25188 31424
rect 25320 31476 25372 31482
rect 25320 31418 25372 31424
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24584 31204 24636 31210
rect 24584 31146 24636 31152
rect 24596 30870 24624 31146
rect 24964 30938 24992 31282
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 24584 30864 24636 30870
rect 24584 30806 24636 30812
rect 24596 30734 24624 30806
rect 24952 30796 25004 30802
rect 24952 30738 25004 30744
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24596 30394 24624 30670
rect 24584 30388 24636 30394
rect 24584 30330 24636 30336
rect 24688 30326 24716 30670
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 24872 29850 24900 30670
rect 24964 30122 24992 30738
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 24492 29232 24544 29238
rect 24492 29174 24544 29180
rect 24688 29034 24716 29514
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24676 29028 24728 29034
rect 24676 28970 24728 28976
rect 24596 28150 24624 28970
rect 24872 28694 24900 29582
rect 24860 28688 24912 28694
rect 24860 28630 24912 28636
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24780 28218 24808 28426
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24584 28144 24636 28150
rect 24584 28086 24636 28092
rect 24964 28082 24992 28494
rect 25148 28218 25176 31418
rect 25228 31340 25280 31346
rect 25228 31282 25280 31288
rect 25240 30666 25268 31282
rect 25228 30660 25280 30666
rect 25228 30602 25280 30608
rect 25240 28966 25268 30602
rect 25228 28960 25280 28966
rect 25228 28902 25280 28908
rect 25320 28960 25372 28966
rect 25320 28902 25372 28908
rect 25240 28626 25268 28902
rect 25228 28620 25280 28626
rect 25228 28562 25280 28568
rect 25332 28558 25360 28902
rect 25516 28762 25544 31826
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25608 30394 25636 31622
rect 25596 30388 25648 30394
rect 25596 30330 25648 30336
rect 25608 29646 25636 30330
rect 25780 30252 25832 30258
rect 25780 30194 25832 30200
rect 25792 29714 25820 30194
rect 25780 29708 25832 29714
rect 25780 29650 25832 29656
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25608 28540 25636 29582
rect 25780 29504 25832 29510
rect 25780 29446 25832 29452
rect 25792 29170 25820 29446
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 25688 28552 25740 28558
rect 25608 28512 25688 28540
rect 25228 28416 25280 28422
rect 25228 28358 25280 28364
rect 25136 28212 25188 28218
rect 25136 28154 25188 28160
rect 25240 28150 25268 28358
rect 25608 28218 25636 28512
rect 25688 28494 25740 28500
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 25228 28144 25280 28150
rect 25228 28086 25280 28092
rect 25688 28144 25740 28150
rect 25688 28086 25740 28092
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 24306 27976 24362 27985
rect 24306 27911 24308 27920
rect 24360 27911 24362 27920
rect 24308 27882 24360 27888
rect 24216 27600 24268 27606
rect 24216 27542 24268 27548
rect 24780 27470 24808 28018
rect 25700 28014 25728 28086
rect 25688 28008 25740 28014
rect 25688 27950 25740 27956
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24136 26382 24164 27406
rect 24584 27328 24636 27334
rect 24584 27270 24636 27276
rect 24596 27062 24624 27270
rect 24584 27056 24636 27062
rect 24584 26998 24636 27004
rect 24308 26920 24360 26926
rect 24308 26862 24360 26868
rect 24320 26586 24348 26862
rect 24688 26586 24716 27406
rect 25700 27334 25728 27950
rect 25884 27334 25912 33458
rect 26160 32978 26188 34614
rect 26988 34134 27016 35566
rect 27356 35562 27384 36246
rect 27436 36168 27488 36174
rect 27436 36110 27488 36116
rect 27344 35556 27396 35562
rect 27344 35498 27396 35504
rect 27448 35154 27476 36110
rect 27528 36032 27580 36038
rect 27528 35974 27580 35980
rect 27540 35834 27568 35974
rect 27528 35828 27580 35834
rect 27528 35770 27580 35776
rect 27436 35148 27488 35154
rect 27436 35090 27488 35096
rect 27448 34542 27476 35090
rect 27436 34536 27488 34542
rect 27436 34478 27488 34484
rect 27448 34202 27476 34478
rect 27632 34202 27660 36722
rect 27724 36038 27752 36722
rect 27712 36032 27764 36038
rect 27712 35974 27764 35980
rect 27724 35290 27752 35974
rect 27712 35284 27764 35290
rect 27712 35226 27764 35232
rect 27712 34944 27764 34950
rect 27712 34886 27764 34892
rect 27724 34678 27752 34886
rect 27712 34672 27764 34678
rect 27712 34614 27764 34620
rect 27436 34196 27488 34202
rect 27436 34138 27488 34144
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 26976 34128 27028 34134
rect 26976 34070 27028 34076
rect 26148 32972 26200 32978
rect 26148 32914 26200 32920
rect 26700 32972 26752 32978
rect 26700 32914 26752 32920
rect 26160 32570 26188 32914
rect 26148 32564 26200 32570
rect 26148 32506 26200 32512
rect 26712 32026 26740 32914
rect 27252 32768 27304 32774
rect 27252 32710 27304 32716
rect 27264 32434 27292 32710
rect 27448 32502 27476 34138
rect 27526 34096 27582 34105
rect 27526 34031 27528 34040
rect 27580 34031 27582 34040
rect 27528 34002 27580 34008
rect 27436 32496 27488 32502
rect 27436 32438 27488 32444
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 27252 32428 27304 32434
rect 27252 32370 27304 32376
rect 26700 32020 26752 32026
rect 26700 31962 26752 31968
rect 26988 31822 27016 32370
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 27540 31822 27568 31962
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 27528 31816 27580 31822
rect 27528 31758 27580 31764
rect 26240 31748 26292 31754
rect 26240 31690 26292 31696
rect 26252 31482 26280 31690
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 25964 30592 26016 30598
rect 25964 30534 26016 30540
rect 25976 30258 26004 30534
rect 25964 30252 26016 30258
rect 25964 30194 26016 30200
rect 25976 29782 26004 30194
rect 25964 29776 26016 29782
rect 25964 29718 26016 29724
rect 26068 28744 26096 30670
rect 26884 30320 26936 30326
rect 26884 30262 26936 30268
rect 26240 30252 26292 30258
rect 26240 30194 26292 30200
rect 26252 29578 26280 30194
rect 26792 30184 26844 30190
rect 26792 30126 26844 30132
rect 26608 30116 26660 30122
rect 26608 30058 26660 30064
rect 26620 29714 26648 30058
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26240 29572 26292 29578
rect 26240 29514 26292 29520
rect 26804 29306 26832 30126
rect 26896 29850 26924 30262
rect 26988 30190 27016 31758
rect 27540 31278 27568 31758
rect 27712 31408 27764 31414
rect 27712 31350 27764 31356
rect 27528 31272 27580 31278
rect 27528 31214 27580 31220
rect 27620 30728 27672 30734
rect 27620 30670 27672 30676
rect 27160 30592 27212 30598
rect 27160 30534 27212 30540
rect 26976 30184 27028 30190
rect 26976 30126 27028 30132
rect 26884 29844 26936 29850
rect 26884 29786 26936 29792
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 25976 28716 26096 28744
rect 25976 28558 26004 28716
rect 26054 28656 26110 28665
rect 26054 28591 26110 28600
rect 26068 28558 26096 28591
rect 25964 28552 26016 28558
rect 25964 28494 26016 28500
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 26056 28212 26108 28218
rect 26056 28154 26108 28160
rect 26068 27538 26096 28154
rect 26344 27946 26372 28494
rect 26332 27940 26384 27946
rect 26332 27882 26384 27888
rect 26056 27532 26108 27538
rect 26056 27474 26108 27480
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25884 27130 25912 27270
rect 24952 27124 25004 27130
rect 24872 27084 24952 27112
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24676 26580 24728 26586
rect 24676 26522 24728 26528
rect 24872 26466 24900 27084
rect 24952 27066 25004 27072
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25884 26926 25912 27066
rect 25872 26920 25924 26926
rect 25872 26862 25924 26868
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25504 26512 25556 26518
rect 24872 26438 25176 26466
rect 25504 26454 25556 26460
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24400 26308 24452 26314
rect 24400 26250 24452 26256
rect 24412 25906 24440 26250
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 24400 25764 24452 25770
rect 24400 25706 24452 25712
rect 24412 25430 24440 25706
rect 24780 25702 24808 26318
rect 24872 25906 24900 26438
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24964 25770 24992 26318
rect 25044 26036 25096 26042
rect 25044 25978 25096 25984
rect 25056 25945 25084 25978
rect 25042 25936 25098 25945
rect 25042 25871 25044 25880
rect 25096 25871 25098 25880
rect 25148 25888 25176 26438
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25240 26042 25268 26318
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25516 25906 25544 26454
rect 25976 26450 26004 26726
rect 25964 26444 26016 26450
rect 25964 26386 26016 26392
rect 26344 26382 26372 27882
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 25686 25936 25742 25945
rect 25412 25900 25464 25906
rect 25148 25860 25268 25888
rect 25044 25842 25096 25848
rect 24860 25764 24912 25770
rect 24860 25706 24912 25712
rect 24952 25764 25004 25770
rect 24952 25706 25004 25712
rect 25136 25764 25188 25770
rect 25136 25706 25188 25712
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24872 25650 24900 25706
rect 25148 25650 25176 25706
rect 24872 25622 25176 25650
rect 24400 25424 24452 25430
rect 24400 25366 24452 25372
rect 23992 25248 24072 25276
rect 23940 25230 23992 25236
rect 23952 24954 23980 25230
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 23940 24948 23992 24954
rect 23940 24890 23992 24896
rect 24044 24818 24072 25094
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24412 24750 24440 25366
rect 24872 25294 24900 25622
rect 24676 25288 24728 25294
rect 24676 25230 24728 25236
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24688 24886 24716 25230
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24676 24880 24728 24886
rect 24490 24848 24546 24857
rect 24676 24822 24728 24828
rect 24490 24783 24492 24792
rect 24544 24783 24546 24792
rect 24492 24754 24544 24760
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 24400 24744 24452 24750
rect 24400 24686 24452 24692
rect 24584 24676 24636 24682
rect 24584 24618 24636 24624
rect 24400 24132 24452 24138
rect 24400 24074 24452 24080
rect 24216 22568 24268 22574
rect 24216 22510 24268 22516
rect 24228 21894 24256 22510
rect 24308 21956 24360 21962
rect 24308 21898 24360 21904
rect 24216 21888 24268 21894
rect 24216 21830 24268 21836
rect 24320 21690 24348 21898
rect 24308 21684 24360 21690
rect 24308 21626 24360 21632
rect 24412 21554 24440 24074
rect 24492 23860 24544 23866
rect 24492 23802 24544 23808
rect 24504 23304 24532 23802
rect 24596 23798 24624 24618
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 24504 23276 24624 23304
rect 24492 23044 24544 23050
rect 24492 22986 24544 22992
rect 24504 21690 24532 22986
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24596 21554 24624 23276
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24584 21548 24636 21554
rect 24584 21490 24636 21496
rect 24688 21350 24716 22102
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 24216 20868 24268 20874
rect 24216 20810 24268 20816
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23768 19718 23796 20470
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18290 23520 19246
rect 23768 18970 23796 19654
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23676 18290 23704 18566
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23664 18284 23716 18290
rect 23664 18226 23716 18232
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23388 18216 23440 18222
rect 23388 18158 23440 18164
rect 23400 17678 23428 18158
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23492 17270 23520 17478
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23584 16425 23612 18226
rect 23860 18154 23888 18226
rect 23664 18148 23716 18154
rect 23664 18090 23716 18096
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23570 16416 23626 16425
rect 23570 16351 23626 16360
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 23124 14346 23152 15030
rect 23112 14340 23164 14346
rect 23112 14282 23164 14288
rect 23124 13258 23152 14282
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23216 13530 23244 13806
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23112 13252 23164 13258
rect 23112 13194 23164 13200
rect 23032 12406 23152 12434
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22100 12232 22152 12238
rect 22284 12232 22336 12238
rect 22152 12192 22232 12220
rect 22100 12174 22152 12180
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22112 10810 22140 11698
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22204 10606 22232 12192
rect 22284 12174 22336 12180
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22296 11898 22324 12174
rect 22480 11898 22508 12174
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22204 10470 22232 10542
rect 22296 10470 22324 11834
rect 22756 10674 22784 12242
rect 22834 12200 22890 12209
rect 22834 12135 22890 12144
rect 23020 12164 23072 12170
rect 22848 11762 22876 12135
rect 23020 12106 23072 12112
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22192 10464 22244 10470
rect 22192 10406 22244 10412
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22008 10260 22060 10266
rect 22060 10220 22140 10248
rect 22008 10202 22060 10208
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21192 9646 21404 9674
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20916 9178 20944 9522
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19904 7478 19932 8026
rect 20824 7818 20852 8978
rect 20812 7812 20864 7818
rect 20812 7754 20864 7760
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 19800 7472 19852 7478
rect 19798 7440 19800 7449
rect 19892 7472 19944 7478
rect 19852 7440 19854 7449
rect 19484 7364 19564 7392
rect 19708 7404 19760 7410
rect 19432 7346 19484 7352
rect 19892 7414 19944 7420
rect 19798 7375 19854 7384
rect 19708 7346 19760 7352
rect 19720 7206 19748 7346
rect 20640 7342 20668 7686
rect 20916 7410 20944 9114
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21008 8362 21036 9046
rect 21376 8634 21404 9646
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21376 8514 21404 8570
rect 21284 8486 21404 8514
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 21284 7478 21312 8486
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21376 7478 21404 8298
rect 21836 7546 21864 9454
rect 22112 8838 22140 10220
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9586 22784 9998
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22848 9382 22876 11698
rect 23032 10810 23060 12106
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22928 10532 22980 10538
rect 22928 10474 22980 10480
rect 22940 10062 22968 10474
rect 23124 10266 23152 12406
rect 23216 12186 23244 13466
rect 23308 12374 23336 15098
rect 23584 14890 23612 16351
rect 23676 15978 23704 18090
rect 23952 16182 23980 20538
rect 24044 20398 24072 20742
rect 24032 20392 24084 20398
rect 24032 20334 24084 20340
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 24136 18290 24164 18770
rect 24124 18284 24176 18290
rect 24044 18244 24124 18272
rect 24044 17678 24072 18244
rect 24124 18226 24176 18232
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 24136 17610 24164 18090
rect 24124 17604 24176 17610
rect 24124 17546 24176 17552
rect 24136 17202 24164 17546
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24228 17082 24256 20810
rect 24780 17762 24808 24890
rect 25056 24857 25084 25230
rect 25240 25226 25268 25860
rect 25412 25842 25464 25848
rect 25504 25900 25556 25906
rect 25686 25871 25688 25880
rect 25504 25842 25556 25848
rect 25740 25871 25742 25880
rect 25688 25842 25740 25848
rect 25424 25809 25452 25842
rect 25792 25838 25820 26318
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26332 25900 26384 25906
rect 26436 25888 26464 29106
rect 26988 28626 27016 30126
rect 27068 30048 27120 30054
rect 27068 29990 27120 29996
rect 27080 29646 27108 29990
rect 27172 29646 27200 30534
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 27160 29640 27212 29646
rect 27160 29582 27212 29588
rect 27528 29164 27580 29170
rect 27632 29152 27660 30670
rect 27724 30054 27752 31350
rect 27712 30048 27764 30054
rect 27712 29990 27764 29996
rect 27724 29646 27752 29990
rect 27816 29782 27844 37998
rect 27988 37946 28040 37952
rect 27896 37868 27948 37874
rect 27896 37810 27948 37816
rect 27908 36922 27936 37810
rect 27988 37800 28040 37806
rect 27988 37742 28040 37748
rect 28000 37466 28028 37742
rect 27988 37460 28040 37466
rect 27988 37402 28040 37408
rect 28184 37194 28212 38286
rect 28172 37188 28224 37194
rect 28172 37130 28224 37136
rect 28080 37120 28132 37126
rect 28080 37062 28132 37068
rect 27896 36916 27948 36922
rect 27896 36858 27948 36864
rect 28092 36854 28120 37062
rect 28080 36848 28132 36854
rect 28080 36790 28132 36796
rect 27896 36100 27948 36106
rect 27896 36042 27948 36048
rect 27908 35834 27936 36042
rect 27896 35828 27948 35834
rect 27896 35770 27948 35776
rect 28172 33856 28224 33862
rect 28172 33798 28224 33804
rect 28184 32978 28212 33798
rect 28172 32972 28224 32978
rect 28172 32914 28224 32920
rect 27896 32904 27948 32910
rect 27896 32846 27948 32852
rect 27804 29776 27856 29782
rect 27804 29718 27856 29724
rect 27712 29640 27764 29646
rect 27816 29617 27844 29718
rect 27712 29582 27764 29588
rect 27802 29608 27858 29617
rect 27802 29543 27858 29552
rect 27908 29510 27936 32846
rect 28184 32570 28212 32914
rect 28172 32564 28224 32570
rect 28172 32506 28224 32512
rect 28276 30802 28304 42298
rect 28356 41064 28408 41070
rect 28356 41006 28408 41012
rect 28368 40730 28396 41006
rect 28356 40724 28408 40730
rect 28356 40666 28408 40672
rect 28356 33516 28408 33522
rect 28356 33458 28408 33464
rect 28368 32774 28396 33458
rect 28356 32768 28408 32774
rect 28356 32710 28408 32716
rect 28368 32230 28396 32710
rect 28356 32224 28408 32230
rect 28356 32166 28408 32172
rect 28264 30796 28316 30802
rect 28264 30738 28316 30744
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 27988 29776 28040 29782
rect 27988 29718 28040 29724
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 27896 29504 27948 29510
rect 27896 29446 27948 29452
rect 27580 29124 27660 29152
rect 27724 29152 27752 29446
rect 27804 29164 27856 29170
rect 27724 29124 27804 29152
rect 27528 29106 27580 29112
rect 27620 29028 27672 29034
rect 27620 28970 27672 28976
rect 26976 28620 27028 28626
rect 26976 28562 27028 28568
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 27356 28422 27384 28494
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27344 28416 27396 28422
rect 27344 28358 27396 28364
rect 26884 27872 26936 27878
rect 26884 27814 26936 27820
rect 26896 27470 26924 27814
rect 26608 27464 26660 27470
rect 26608 27406 26660 27412
rect 26884 27464 26936 27470
rect 26884 27406 26936 27412
rect 26516 27328 26568 27334
rect 26516 27270 26568 27276
rect 26528 27062 26556 27270
rect 26516 27056 26568 27062
rect 26516 26998 26568 27004
rect 26384 25860 26464 25888
rect 26332 25842 26384 25848
rect 25596 25832 25648 25838
rect 25410 25800 25466 25809
rect 25596 25774 25648 25780
rect 25780 25832 25832 25838
rect 25780 25774 25832 25780
rect 25410 25735 25466 25744
rect 25608 25430 25636 25774
rect 25884 25498 25912 25842
rect 25976 25702 26004 25842
rect 25964 25696 26016 25702
rect 25964 25638 26016 25644
rect 25872 25492 25924 25498
rect 25872 25434 25924 25440
rect 25596 25424 25648 25430
rect 25596 25366 25648 25372
rect 25976 25362 26004 25638
rect 26160 25498 26188 25842
rect 26148 25492 26200 25498
rect 26148 25434 26200 25440
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25228 25220 25280 25226
rect 25228 25162 25280 25168
rect 25042 24848 25098 24857
rect 25042 24783 25098 24792
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 21536 24900 23462
rect 24964 21894 24992 24142
rect 24952 21888 25004 21894
rect 24950 21856 24952 21865
rect 25004 21856 25006 21865
rect 24950 21791 25006 21800
rect 25056 21622 25084 24783
rect 25240 24206 25268 25162
rect 25792 25158 25820 25230
rect 25780 25152 25832 25158
rect 25780 25094 25832 25100
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25332 24206 25360 24550
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25332 23798 25360 24142
rect 25320 23792 25372 23798
rect 25516 23769 25544 24754
rect 25792 24750 25820 25094
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 26056 24744 26108 24750
rect 26056 24686 26108 24692
rect 26068 24206 26096 24686
rect 25964 24200 26016 24206
rect 25964 24142 26016 24148
rect 26056 24200 26108 24206
rect 26056 24142 26108 24148
rect 25976 23866 26004 24142
rect 25964 23860 26016 23866
rect 25964 23802 26016 23808
rect 25320 23734 25372 23740
rect 25502 23760 25558 23769
rect 25502 23695 25558 23704
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 25872 23656 25924 23662
rect 25872 23598 25924 23604
rect 25792 22982 25820 23598
rect 25884 22982 25912 23598
rect 25976 23050 26004 23802
rect 26344 23746 26372 25842
rect 26424 25220 26476 25226
rect 26424 25162 26476 25168
rect 26436 24954 26464 25162
rect 26424 24948 26476 24954
rect 26424 24890 26476 24896
rect 26252 23718 26372 23746
rect 26424 23724 26476 23730
rect 25964 23044 26016 23050
rect 25964 22986 26016 22992
rect 25780 22976 25832 22982
rect 25778 22944 25780 22953
rect 25872 22976 25924 22982
rect 25832 22944 25834 22953
rect 25872 22918 25924 22924
rect 25778 22879 25834 22888
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24952 21548 25004 21554
rect 24872 21508 24952 21536
rect 24952 21490 25004 21496
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 24964 20806 24992 21490
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 25056 20398 25084 21422
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 25240 21010 25268 21286
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25608 20806 25636 21490
rect 25700 21078 25728 21830
rect 25688 21072 25740 21078
rect 25688 21014 25740 21020
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25412 20528 25464 20534
rect 25412 20470 25464 20476
rect 25044 20392 25096 20398
rect 25044 20334 25096 20340
rect 25056 19922 25084 20334
rect 25044 19916 25096 19922
rect 25044 19858 25096 19864
rect 25424 19446 25452 20470
rect 25596 19780 25648 19786
rect 25596 19722 25648 19728
rect 25608 19514 25636 19722
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25044 19440 25096 19446
rect 25044 19382 25096 19388
rect 25412 19440 25464 19446
rect 25412 19382 25464 19388
rect 25056 18358 25084 19382
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 25044 18352 25096 18358
rect 25044 18294 25096 18300
rect 24872 17882 24900 18294
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24032 17060 24084 17066
rect 24032 17002 24084 17008
rect 24136 17054 24256 17082
rect 24320 17734 24808 17762
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 24044 16522 24072 17002
rect 24032 16516 24084 16522
rect 24032 16458 24084 16464
rect 24044 16250 24072 16458
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23940 16176 23992 16182
rect 23940 16118 23992 16124
rect 23664 15972 23716 15978
rect 23664 15914 23716 15920
rect 23676 15706 23704 15914
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 23572 14884 23624 14890
rect 23572 14826 23624 14832
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12986 24072 13126
rect 24136 12986 24164 17054
rect 24320 15502 24348 17734
rect 24964 17678 24992 17750
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17202 24440 17478
rect 24596 17338 24624 17614
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24688 17292 24900 17320
rect 24504 17218 24532 17274
rect 24688 17218 24716 17292
rect 24400 17196 24452 17202
rect 24504 17190 24716 17218
rect 24768 17196 24820 17202
rect 24400 17138 24452 17144
rect 24768 17138 24820 17144
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24688 16998 24716 17070
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24780 16658 24808 17138
rect 24872 17134 24900 17292
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24964 17066 24992 17138
rect 24952 17060 25004 17066
rect 24952 17002 25004 17008
rect 24964 16794 24992 17002
rect 24952 16788 25004 16794
rect 24952 16730 25004 16736
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24872 16538 24900 16594
rect 24780 16510 24900 16538
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 24320 14618 24348 15438
rect 24688 15434 24716 16118
rect 24780 16046 24808 16510
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24872 16182 24900 16390
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 24768 16040 24820 16046
rect 24768 15982 24820 15988
rect 24676 15428 24728 15434
rect 24676 15370 24728 15376
rect 24492 15088 24544 15094
rect 24492 15030 24544 15036
rect 24504 14958 24532 15030
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24504 14550 24532 14894
rect 24596 14618 24624 14894
rect 24780 14822 24808 15982
rect 25056 15858 25084 18294
rect 25148 17746 25176 18770
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 17338 25176 17546
rect 25332 17542 25360 18158
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25608 17954 25636 18022
rect 25516 17926 25636 17954
rect 25516 17678 25544 17926
rect 25700 17814 25728 18022
rect 25688 17808 25740 17814
rect 25688 17750 25740 17756
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25240 16250 25268 16526
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25516 16114 25544 17614
rect 25700 17270 25728 17750
rect 25688 17264 25740 17270
rect 25688 17206 25740 17212
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25056 15830 25176 15858
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24872 14958 24900 15506
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24964 14958 24992 15438
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 24952 14952 25004 14958
rect 24952 14894 25004 14900
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24492 14544 24544 14550
rect 24492 14486 24544 14492
rect 24780 14414 24808 14758
rect 24872 14482 24900 14894
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24412 14074 24440 14350
rect 24964 14074 24992 14894
rect 25148 14482 25176 15830
rect 25608 15706 25636 16526
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25148 14006 25176 14214
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 25504 13932 25556 13938
rect 25608 13920 25636 15642
rect 25700 15638 25728 15982
rect 25688 15632 25740 15638
rect 25688 15574 25740 15580
rect 25688 14612 25740 14618
rect 25688 14554 25740 14560
rect 25556 13892 25636 13920
rect 25504 13874 25556 13880
rect 24688 13190 24716 13874
rect 25700 13870 25728 14554
rect 25792 13920 25820 21966
rect 25884 14074 25912 22918
rect 25964 22432 26016 22438
rect 25964 22374 26016 22380
rect 25976 22030 26004 22374
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 26056 19304 26108 19310
rect 26108 19264 26188 19292
rect 26056 19246 26108 19252
rect 26160 18154 26188 19264
rect 26148 18148 26200 18154
rect 26148 18090 26200 18096
rect 26056 17740 26108 17746
rect 26160 17728 26188 18090
rect 26108 17700 26188 17728
rect 26056 17682 26108 17688
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 25976 16590 26004 16934
rect 26160 16590 26188 17700
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 25964 16448 26016 16454
rect 25962 16416 25964 16425
rect 26016 16416 26018 16425
rect 25962 16351 26018 16360
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25872 13932 25924 13938
rect 25792 13892 25872 13920
rect 25872 13874 25924 13880
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 25688 13728 25740 13734
rect 25042 13696 25098 13705
rect 25042 13631 25098 13640
rect 25686 13696 25688 13705
rect 25740 13696 25742 13705
rect 25686 13631 25742 13640
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24676 13184 24728 13190
rect 24676 13126 24728 13132
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 23572 12844 23624 12850
rect 23572 12786 23624 12792
rect 23584 12753 23612 12786
rect 23570 12744 23626 12753
rect 23570 12679 23626 12688
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 23296 12368 23348 12374
rect 23296 12310 23348 12316
rect 23480 12232 23532 12238
rect 23478 12200 23480 12209
rect 23532 12200 23534 12209
rect 23216 12170 23428 12186
rect 23216 12164 23440 12170
rect 23216 12158 23388 12164
rect 23478 12135 23534 12144
rect 23388 12106 23440 12112
rect 23400 11898 23428 12106
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23584 11830 23612 12582
rect 24688 12442 24716 12582
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24780 12306 24808 13262
rect 25056 12986 25084 13631
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 23676 11558 23704 12038
rect 24320 11898 24348 12038
rect 24308 11892 24360 11898
rect 24308 11834 24360 11840
rect 24400 11756 24452 11762
rect 24596 11744 24624 12106
rect 24452 11716 24624 11744
rect 24400 11698 24452 11704
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23664 11552 23716 11558
rect 23664 11494 23716 11500
rect 23400 11150 23428 11494
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 22928 10056 22980 10062
rect 22928 9998 22980 10004
rect 22940 9518 22968 9998
rect 23400 9518 23428 11086
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22376 9376 22428 9382
rect 22376 9318 22428 9324
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22388 9042 22416 9318
rect 22376 9036 22428 9042
rect 22376 8978 22428 8984
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22664 8498 22692 8910
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22652 8492 22704 8498
rect 22652 8434 22704 8440
rect 22388 7954 22416 8434
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22112 7546 22140 7754
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 22848 7410 22876 9318
rect 23400 7954 23428 9454
rect 23676 9178 23704 11494
rect 24412 11082 24440 11698
rect 24780 11694 24808 12242
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24872 11150 24900 12038
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23676 8566 23704 9114
rect 23768 9042 23796 10066
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23860 8838 23888 10542
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23952 9654 23980 10406
rect 24228 10266 24256 10610
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24412 10130 24440 11018
rect 24872 10742 24900 11086
rect 25516 10810 25544 11698
rect 25792 11150 25820 12786
rect 25884 12306 25912 13738
rect 25976 13190 26004 16351
rect 26252 16250 26280 23718
rect 26424 23666 26476 23672
rect 26436 23118 26464 23666
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26344 22098 26372 22646
rect 26436 22642 26464 23054
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26332 22092 26384 22098
rect 26332 22034 26384 22040
rect 26436 21622 26464 22578
rect 26528 22574 26556 26998
rect 26620 26926 26648 27406
rect 26700 27396 26752 27402
rect 26700 27338 26752 27344
rect 27068 27396 27120 27402
rect 27068 27338 27120 27344
rect 26712 27130 26740 27338
rect 27080 27130 27108 27338
rect 26700 27124 26752 27130
rect 26700 27066 26752 27072
rect 27068 27124 27120 27130
rect 27068 27066 27120 27072
rect 27264 26994 27292 28358
rect 27632 28082 27660 28970
rect 27620 28076 27672 28082
rect 27620 28018 27672 28024
rect 27632 27878 27660 28018
rect 27620 27872 27672 27878
rect 27620 27814 27672 27820
rect 27344 27396 27396 27402
rect 27344 27338 27396 27344
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 26608 26920 26660 26926
rect 26608 26862 26660 26868
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 26608 26240 26660 26246
rect 26608 26182 26660 26188
rect 26620 25838 26648 26182
rect 26988 25906 27016 26250
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 26608 25832 26660 25838
rect 26608 25774 26660 25780
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26620 24818 26648 25638
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 26884 24336 26936 24342
rect 26884 24278 26936 24284
rect 26700 24200 26752 24206
rect 26700 24142 26752 24148
rect 26712 23526 26740 24142
rect 26792 23860 26844 23866
rect 26792 23802 26844 23808
rect 26700 23520 26752 23526
rect 26700 23462 26752 23468
rect 26516 22568 26568 22574
rect 26516 22510 26568 22516
rect 26424 21616 26476 21622
rect 26424 21558 26476 21564
rect 26516 17604 26568 17610
rect 26516 17546 26568 17552
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26436 17202 26464 17478
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26056 15904 26108 15910
rect 26056 15846 26108 15852
rect 26068 15434 26096 15846
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 26056 15428 26108 15434
rect 26056 15370 26108 15376
rect 26160 15094 26188 15506
rect 26148 15088 26200 15094
rect 26148 15030 26200 15036
rect 26160 14482 26188 15030
rect 26344 14770 26372 16594
rect 26424 15972 26476 15978
rect 26424 15914 26476 15920
rect 26436 14958 26464 15914
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26344 14742 26464 14770
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26160 14074 26188 14418
rect 26332 14408 26384 14414
rect 26332 14350 26384 14356
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26344 13938 26372 14350
rect 26436 13938 26464 14742
rect 26528 14550 26556 17546
rect 26516 14544 26568 14550
rect 26516 14486 26568 14492
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26068 13394 26096 13670
rect 26252 13462 26280 13670
rect 26344 13530 26372 13874
rect 26528 13530 26556 14214
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26516 13524 26568 13530
rect 26516 13466 26568 13472
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26436 13190 26464 13262
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26424 12912 26476 12918
rect 26424 12854 26476 12860
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 26252 12442 26280 12718
rect 26240 12436 26292 12442
rect 26292 12396 26372 12424
rect 26240 12378 26292 12384
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 26148 11212 26200 11218
rect 26252 11200 26280 12038
rect 26344 11898 26372 12396
rect 26436 12374 26464 12854
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26712 12306 26740 23462
rect 26804 22658 26832 23802
rect 26896 22760 26924 24278
rect 26976 24064 27028 24070
rect 26976 24006 27028 24012
rect 26988 23118 27016 24006
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 26896 22732 27016 22760
rect 26804 22630 26924 22658
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26804 20942 26832 22510
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26792 20460 26844 20466
rect 26792 20402 26844 20408
rect 26804 13870 26832 20402
rect 26896 14618 26924 22630
rect 26988 22098 27016 22732
rect 26976 22092 27028 22098
rect 26976 22034 27028 22040
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26988 20602 27016 20878
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 27080 20058 27108 26318
rect 27160 26240 27212 26246
rect 27160 26182 27212 26188
rect 27172 26042 27200 26182
rect 27160 26036 27212 26042
rect 27160 25978 27212 25984
rect 27172 24682 27200 25978
rect 27356 25158 27384 27338
rect 27448 27130 27476 27338
rect 27436 27124 27488 27130
rect 27436 27066 27488 27072
rect 27344 25152 27396 25158
rect 27724 25106 27752 29124
rect 27804 29106 27856 29112
rect 27804 29028 27856 29034
rect 27804 28970 27856 28976
rect 27816 28082 27844 28970
rect 27804 28076 27856 28082
rect 27804 28018 27856 28024
rect 27816 27946 27844 28018
rect 27804 27940 27856 27946
rect 27804 27882 27856 27888
rect 27908 27554 27936 29446
rect 28000 29034 28028 29718
rect 27988 29028 28040 29034
rect 27988 28970 28040 28976
rect 28092 28422 28120 30670
rect 28356 30592 28408 30598
rect 28356 30534 28408 30540
rect 28368 30433 28396 30534
rect 28354 30424 28410 30433
rect 28354 30359 28410 30368
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28368 28490 28396 30194
rect 28460 29306 28488 43318
rect 29552 43308 29604 43314
rect 29552 43250 29604 43256
rect 29564 42702 29592 43250
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 29644 42764 29696 42770
rect 29644 42706 29696 42712
rect 37280 42764 37332 42770
rect 37280 42706 37332 42712
rect 29552 42696 29604 42702
rect 29552 42638 29604 42644
rect 28540 42628 28592 42634
rect 28540 42570 28592 42576
rect 28816 42628 28868 42634
rect 28816 42570 28868 42576
rect 28552 42294 28580 42570
rect 28540 42288 28592 42294
rect 28828 42242 28856 42570
rect 29564 42362 29592 42638
rect 29552 42356 29604 42362
rect 29552 42298 29604 42304
rect 29656 42294 29684 42706
rect 35440 42628 35492 42634
rect 35440 42570 35492 42576
rect 36820 42628 36872 42634
rect 36820 42570 36872 42576
rect 35452 42362 35480 42570
rect 35594 42460 35902 42469
rect 35594 42458 35600 42460
rect 35656 42458 35680 42460
rect 35736 42458 35760 42460
rect 35816 42458 35840 42460
rect 35896 42458 35902 42460
rect 35656 42406 35658 42458
rect 35838 42406 35840 42458
rect 35594 42404 35600 42406
rect 35656 42404 35680 42406
rect 35736 42404 35760 42406
rect 35816 42404 35840 42406
rect 35896 42404 35902 42406
rect 35594 42395 35902 42404
rect 35440 42356 35492 42362
rect 35440 42298 35492 42304
rect 36832 42294 36860 42570
rect 37004 42560 37056 42566
rect 37004 42502 37056 42508
rect 28540 42230 28592 42236
rect 28736 42214 28856 42242
rect 29644 42288 29696 42294
rect 29644 42230 29696 42236
rect 36820 42288 36872 42294
rect 36820 42230 36872 42236
rect 28736 42158 28764 42214
rect 28724 42152 28776 42158
rect 28724 42094 28776 42100
rect 28816 42152 28868 42158
rect 28816 42094 28868 42100
rect 28540 41812 28592 41818
rect 28540 41754 28592 41760
rect 28552 41546 28580 41754
rect 28724 41744 28776 41750
rect 28724 41686 28776 41692
rect 28736 41614 28764 41686
rect 28724 41608 28776 41614
rect 28724 41550 28776 41556
rect 28540 41540 28592 41546
rect 28540 41482 28592 41488
rect 28828 41414 28856 42094
rect 29092 41472 29144 41478
rect 29092 41414 29144 41420
rect 28828 41386 28948 41414
rect 28920 41206 28948 41386
rect 28908 41200 28960 41206
rect 28908 41142 28960 41148
rect 28920 41070 28948 41142
rect 28908 41064 28960 41070
rect 28908 41006 28960 41012
rect 28540 39568 28592 39574
rect 28540 39510 28592 39516
rect 28552 38962 28580 39510
rect 28540 38956 28592 38962
rect 28540 38898 28592 38904
rect 28552 38554 28580 38898
rect 28540 38548 28592 38554
rect 28540 38490 28592 38496
rect 28920 38486 28948 41006
rect 29104 40594 29132 41414
rect 29656 41206 29684 42230
rect 34796 42220 34848 42226
rect 34796 42162 34848 42168
rect 35624 42220 35676 42226
rect 35624 42162 35676 42168
rect 36452 42220 36504 42226
rect 36452 42162 36504 42168
rect 30840 42152 30892 42158
rect 30840 42094 30892 42100
rect 30932 42152 30984 42158
rect 30932 42094 30984 42100
rect 32036 42152 32088 42158
rect 32036 42094 32088 42100
rect 30852 41818 30880 42094
rect 30944 42022 30972 42094
rect 31576 42084 31628 42090
rect 31576 42026 31628 42032
rect 30932 42016 30984 42022
rect 30932 41958 30984 41964
rect 31208 42016 31260 42022
rect 31208 41958 31260 41964
rect 30840 41812 30892 41818
rect 30840 41754 30892 41760
rect 30932 41812 30984 41818
rect 30932 41754 30984 41760
rect 30944 41614 30972 41754
rect 31116 41744 31168 41750
rect 31116 41686 31168 41692
rect 31128 41614 31156 41686
rect 31220 41614 31248 41958
rect 31588 41614 31616 42026
rect 32048 41614 32076 42094
rect 32956 42016 33008 42022
rect 32956 41958 33008 41964
rect 32220 41812 32272 41818
rect 32220 41754 32272 41760
rect 32864 41812 32916 41818
rect 32864 41754 32916 41760
rect 32128 41676 32180 41682
rect 32128 41618 32180 41624
rect 30472 41608 30524 41614
rect 30472 41550 30524 41556
rect 30932 41608 30984 41614
rect 30932 41550 30984 41556
rect 31116 41608 31168 41614
rect 31116 41550 31168 41556
rect 31208 41608 31260 41614
rect 31208 41550 31260 41556
rect 31576 41608 31628 41614
rect 31576 41550 31628 41556
rect 31852 41608 31904 41614
rect 31852 41550 31904 41556
rect 31944 41608 31996 41614
rect 31944 41550 31996 41556
rect 32036 41608 32088 41614
rect 32036 41550 32088 41556
rect 29644 41200 29696 41206
rect 29644 41142 29696 41148
rect 29092 40588 29144 40594
rect 29092 40530 29144 40536
rect 29184 39568 29236 39574
rect 29184 39510 29236 39516
rect 29196 39370 29224 39510
rect 29184 39364 29236 39370
rect 29184 39306 29236 39312
rect 29196 38554 29224 39306
rect 29184 38548 29236 38554
rect 29184 38490 29236 38496
rect 28908 38480 28960 38486
rect 28908 38422 28960 38428
rect 28908 38344 28960 38350
rect 28908 38286 28960 38292
rect 28632 38276 28684 38282
rect 28632 38218 28684 38224
rect 28644 38010 28672 38218
rect 28920 38010 28948 38286
rect 29184 38276 29236 38282
rect 29184 38218 29236 38224
rect 29552 38276 29604 38282
rect 29552 38218 29604 38224
rect 28632 38004 28684 38010
rect 28632 37946 28684 37952
rect 28908 38004 28960 38010
rect 28908 37946 28960 37952
rect 28908 37868 28960 37874
rect 28908 37810 28960 37816
rect 28920 37670 28948 37810
rect 28908 37664 28960 37670
rect 28908 37606 28960 37612
rect 28920 37398 28948 37606
rect 28908 37392 28960 37398
rect 28908 37334 28960 37340
rect 28920 36786 28948 37334
rect 29196 36786 29224 38218
rect 29564 38010 29592 38218
rect 29552 38004 29604 38010
rect 29552 37946 29604 37952
rect 29276 37868 29328 37874
rect 29276 37810 29328 37816
rect 28908 36780 28960 36786
rect 28908 36722 28960 36728
rect 29184 36780 29236 36786
rect 29184 36722 29236 36728
rect 29092 36576 29144 36582
rect 29092 36518 29144 36524
rect 29104 35834 29132 36518
rect 29196 36378 29224 36722
rect 29184 36372 29236 36378
rect 29184 36314 29236 36320
rect 29288 36258 29316 37810
rect 29656 37346 29684 41142
rect 30484 41052 30512 41550
rect 30748 41540 30800 41546
rect 30748 41482 30800 41488
rect 30760 41138 30788 41482
rect 30748 41132 30800 41138
rect 30748 41074 30800 41080
rect 31116 41132 31168 41138
rect 31116 41074 31168 41080
rect 30564 41064 30616 41070
rect 30484 41024 30564 41052
rect 30484 40662 30512 41024
rect 30564 41006 30616 41012
rect 30564 40928 30616 40934
rect 30564 40870 30616 40876
rect 30472 40656 30524 40662
rect 30472 40598 30524 40604
rect 30288 40044 30340 40050
rect 30288 39986 30340 39992
rect 30300 39574 30328 39986
rect 30288 39568 30340 39574
rect 30288 39510 30340 39516
rect 30576 39522 30604 40870
rect 31128 40662 31156 41074
rect 31116 40656 31168 40662
rect 31116 40598 31168 40604
rect 30656 40588 30708 40594
rect 30656 40530 30708 40536
rect 30668 39642 30696 40530
rect 30748 40520 30800 40526
rect 30748 40462 30800 40468
rect 30760 40186 30788 40462
rect 30748 40180 30800 40186
rect 30748 40122 30800 40128
rect 30656 39636 30708 39642
rect 30656 39578 30708 39584
rect 31024 39636 31076 39642
rect 31024 39578 31076 39584
rect 30838 39536 30894 39545
rect 30576 39494 30696 39522
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 30564 38956 30616 38962
rect 30564 38898 30616 38904
rect 30208 37874 30236 38898
rect 30576 37874 30604 38898
rect 30196 37868 30248 37874
rect 30196 37810 30248 37816
rect 30564 37868 30616 37874
rect 30564 37810 30616 37816
rect 30012 37800 30064 37806
rect 30012 37742 30064 37748
rect 30104 37800 30156 37806
rect 30104 37742 30156 37748
rect 29472 37318 29684 37346
rect 29472 37262 29500 37318
rect 29460 37256 29512 37262
rect 29460 37198 29512 37204
rect 29552 37256 29604 37262
rect 29552 37198 29604 37204
rect 29656 37210 29684 37318
rect 29564 36378 29592 37198
rect 29656 37182 29776 37210
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29552 36372 29604 36378
rect 29552 36314 29604 36320
rect 29196 36230 29316 36258
rect 29092 35828 29144 35834
rect 29092 35770 29144 35776
rect 28724 35624 28776 35630
rect 28724 35566 28776 35572
rect 29000 35624 29052 35630
rect 29000 35566 29052 35572
rect 28736 34202 28764 35566
rect 29012 35154 29040 35566
rect 29000 35148 29052 35154
rect 29000 35090 29052 35096
rect 29196 35086 29224 36230
rect 29276 36100 29328 36106
rect 29276 36042 29328 36048
rect 29288 35154 29316 36042
rect 29656 35834 29684 37062
rect 29748 36718 29776 37182
rect 29736 36712 29788 36718
rect 29736 36654 29788 36660
rect 29748 36106 29776 36654
rect 29736 36100 29788 36106
rect 29736 36042 29788 36048
rect 29644 35828 29696 35834
rect 29644 35770 29696 35776
rect 29276 35148 29328 35154
rect 29276 35090 29328 35096
rect 29184 35080 29236 35086
rect 29184 35022 29236 35028
rect 29196 34746 29224 35022
rect 29184 34740 29236 34746
rect 29184 34682 29236 34688
rect 29288 34678 29316 35090
rect 29460 34944 29512 34950
rect 29460 34886 29512 34892
rect 29276 34672 29328 34678
rect 29276 34614 29328 34620
rect 29184 34604 29236 34610
rect 29184 34546 29236 34552
rect 28724 34196 28776 34202
rect 28724 34138 28776 34144
rect 29196 34066 29224 34546
rect 29472 34202 29500 34886
rect 30024 34746 30052 37742
rect 30116 37330 30144 37742
rect 30104 37324 30156 37330
rect 30104 37266 30156 37272
rect 30116 35698 30144 37266
rect 30208 37262 30236 37810
rect 30576 37398 30604 37810
rect 30564 37392 30616 37398
rect 30564 37334 30616 37340
rect 30196 37256 30248 37262
rect 30196 37198 30248 37204
rect 30472 37120 30524 37126
rect 30472 37062 30524 37068
rect 30484 36854 30512 37062
rect 30472 36848 30524 36854
rect 30472 36790 30524 36796
rect 30104 35692 30156 35698
rect 30104 35634 30156 35640
rect 30668 35578 30696 39494
rect 30838 39471 30840 39480
rect 30892 39471 30894 39480
rect 30840 39442 30892 39448
rect 31036 39438 31064 39578
rect 31024 39432 31076 39438
rect 31024 39374 31076 39380
rect 31036 39080 31064 39374
rect 30944 39052 31064 39080
rect 30746 38992 30802 39001
rect 30746 38927 30748 38936
rect 30800 38927 30802 38936
rect 30748 38898 30800 38904
rect 30760 37942 30788 38898
rect 30944 38826 30972 39052
rect 31024 38956 31076 38962
rect 31024 38898 31076 38904
rect 30932 38820 30984 38826
rect 30932 38762 30984 38768
rect 31036 38554 31064 38898
rect 31220 38654 31248 41550
rect 31668 41540 31720 41546
rect 31668 41482 31720 41488
rect 31680 41206 31708 41482
rect 31864 41478 31892 41550
rect 31852 41472 31904 41478
rect 31852 41414 31904 41420
rect 31864 41206 31892 41414
rect 31668 41200 31720 41206
rect 31668 41142 31720 41148
rect 31852 41200 31904 41206
rect 31852 41142 31904 41148
rect 31956 40390 31984 41550
rect 31944 40384 31996 40390
rect 31944 40326 31996 40332
rect 31392 40044 31444 40050
rect 31392 39986 31444 39992
rect 32036 40044 32088 40050
rect 32036 39986 32088 39992
rect 31404 39506 31432 39986
rect 32048 39642 32076 39986
rect 31944 39636 31996 39642
rect 31944 39578 31996 39584
rect 32036 39636 32088 39642
rect 32036 39578 32088 39584
rect 31392 39500 31444 39506
rect 31392 39442 31444 39448
rect 31404 39409 31432 39442
rect 31956 39438 31984 39578
rect 31668 39432 31720 39438
rect 31390 39400 31446 39409
rect 31760 39432 31812 39438
rect 31668 39374 31720 39380
rect 31758 39400 31760 39409
rect 31944 39432 31996 39438
rect 31812 39400 31814 39409
rect 31390 39335 31446 39344
rect 31404 38758 31432 39335
rect 31680 39302 31708 39374
rect 31944 39374 31996 39380
rect 31758 39335 31814 39344
rect 31668 39296 31720 39302
rect 31668 39238 31720 39244
rect 31944 38956 31996 38962
rect 31944 38898 31996 38904
rect 31392 38752 31444 38758
rect 31392 38694 31444 38700
rect 31128 38626 31248 38654
rect 31024 38548 31076 38554
rect 31024 38490 31076 38496
rect 30748 37936 30800 37942
rect 30748 37878 30800 37884
rect 31024 36100 31076 36106
rect 31024 36042 31076 36048
rect 30748 36032 30800 36038
rect 30748 35974 30800 35980
rect 30760 35766 30788 35974
rect 30748 35760 30800 35766
rect 30748 35702 30800 35708
rect 30840 35624 30892 35630
rect 30668 35550 30788 35578
rect 30840 35566 30892 35572
rect 30012 34740 30064 34746
rect 30012 34682 30064 34688
rect 30196 34468 30248 34474
rect 30196 34410 30248 34416
rect 29460 34196 29512 34202
rect 29460 34138 29512 34144
rect 30208 34066 30236 34410
rect 29184 34060 29236 34066
rect 29184 34002 29236 34008
rect 30196 34060 30248 34066
rect 30196 34002 30248 34008
rect 28632 33992 28684 33998
rect 28632 33934 28684 33940
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 28644 33862 28672 33934
rect 30024 33862 30052 33934
rect 28632 33856 28684 33862
rect 28632 33798 28684 33804
rect 29920 33856 29972 33862
rect 29920 33798 29972 33804
rect 30012 33856 30064 33862
rect 30012 33798 30064 33804
rect 28540 32428 28592 32434
rect 28540 32370 28592 32376
rect 28552 32026 28580 32370
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28644 31958 28672 33798
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29472 32842 29500 33390
rect 29748 33114 29776 33458
rect 29736 33108 29788 33114
rect 29736 33050 29788 33056
rect 29460 32836 29512 32842
rect 29460 32778 29512 32784
rect 28816 32768 28868 32774
rect 28816 32710 28868 32716
rect 28828 32502 28856 32710
rect 28816 32496 28868 32502
rect 28816 32438 28868 32444
rect 29472 32230 29500 32778
rect 29932 32434 29960 33798
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29920 32428 29972 32434
rect 29920 32370 29972 32376
rect 29460 32224 29512 32230
rect 29460 32166 29512 32172
rect 28632 31952 28684 31958
rect 28632 31894 28684 31900
rect 28644 30258 28672 31894
rect 29472 31890 29500 32166
rect 29460 31884 29512 31890
rect 29512 31844 29592 31872
rect 29460 31826 29512 31832
rect 29564 31346 29592 31844
rect 29656 31482 29684 32370
rect 30024 32366 30052 33798
rect 30564 33380 30616 33386
rect 30564 33322 30616 33328
rect 30196 33312 30248 33318
rect 30196 33254 30248 33260
rect 30208 32978 30236 33254
rect 30196 32972 30248 32978
rect 30196 32914 30248 32920
rect 30012 32360 30064 32366
rect 30012 32302 30064 32308
rect 30208 31754 30236 32914
rect 30576 32910 30604 33322
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 30564 32224 30616 32230
rect 30564 32166 30616 32172
rect 30656 32224 30708 32230
rect 30656 32166 30708 32172
rect 30380 31816 30432 31822
rect 30380 31758 30432 31764
rect 30196 31748 30248 31754
rect 30248 31708 30328 31736
rect 30196 31690 30248 31696
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 29644 31476 29696 31482
rect 29644 31418 29696 31424
rect 28816 31340 28868 31346
rect 28816 31282 28868 31288
rect 29552 31340 29604 31346
rect 29552 31282 29604 31288
rect 28828 30326 28856 31282
rect 28908 30728 28960 30734
rect 29736 30728 29788 30734
rect 28908 30670 28960 30676
rect 29182 30696 29238 30705
rect 28816 30320 28868 30326
rect 28816 30262 28868 30268
rect 28632 30252 28684 30258
rect 28632 30194 28684 30200
rect 28920 29850 28948 30670
rect 29736 30670 29788 30676
rect 29182 30631 29184 30640
rect 29236 30631 29238 30640
rect 29184 30602 29236 30608
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 28908 29844 28960 29850
rect 29104 29832 29132 30534
rect 29748 30258 29776 30670
rect 29552 30252 29604 30258
rect 29552 30194 29604 30200
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29828 30252 29880 30258
rect 29828 30194 29880 30200
rect 29460 30116 29512 30122
rect 29460 30058 29512 30064
rect 29104 29804 29224 29832
rect 28908 29786 28960 29792
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 29012 29578 29040 29650
rect 29000 29572 29052 29578
rect 29000 29514 29052 29520
rect 29012 29345 29040 29514
rect 28998 29336 29054 29345
rect 28448 29300 28500 29306
rect 28998 29271 29054 29280
rect 28448 29242 28500 29248
rect 29196 29238 29224 29804
rect 29472 29782 29500 30058
rect 29564 30025 29592 30194
rect 29550 30016 29606 30025
rect 29550 29951 29606 29960
rect 29460 29776 29512 29782
rect 29460 29718 29512 29724
rect 29644 29708 29696 29714
rect 29644 29650 29696 29656
rect 29368 29640 29420 29646
rect 29368 29582 29420 29588
rect 29184 29232 29236 29238
rect 29184 29174 29236 29180
rect 28906 28656 28962 28665
rect 28906 28591 28962 28600
rect 28356 28484 28408 28490
rect 28356 28426 28408 28432
rect 28080 28416 28132 28422
rect 28080 28358 28132 28364
rect 28092 28082 28120 28358
rect 28368 28218 28396 28426
rect 28920 28218 28948 28591
rect 28356 28212 28408 28218
rect 28356 28154 28408 28160
rect 28908 28212 28960 28218
rect 28908 28154 28960 28160
rect 28080 28076 28132 28082
rect 28080 28018 28132 28024
rect 28368 27946 28396 28154
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 28356 27940 28408 27946
rect 28356 27882 28408 27888
rect 27816 27526 27936 27554
rect 27816 25158 27844 27526
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 25294 27936 27338
rect 28000 26926 28028 27882
rect 28828 27849 28856 28018
rect 28814 27840 28870 27849
rect 28814 27775 28870 27784
rect 28920 27606 28948 28154
rect 29196 27606 29224 29174
rect 29380 28694 29408 29582
rect 29460 29504 29512 29510
rect 29460 29446 29512 29452
rect 29472 29170 29500 29446
rect 29656 29170 29684 29650
rect 29748 29510 29776 30194
rect 29840 29646 29868 30194
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29736 29504 29788 29510
rect 29736 29446 29788 29452
rect 29460 29164 29512 29170
rect 29460 29106 29512 29112
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29644 29028 29696 29034
rect 29644 28970 29696 28976
rect 29368 28688 29420 28694
rect 29368 28630 29420 28636
rect 29368 28484 29420 28490
rect 29368 28426 29420 28432
rect 29276 28416 29328 28422
rect 29276 28358 29328 28364
rect 29288 28150 29316 28358
rect 29380 28218 29408 28426
rect 29368 28212 29420 28218
rect 29368 28154 29420 28160
rect 29656 28150 29684 28970
rect 29736 28960 29788 28966
rect 29736 28902 29788 28908
rect 29748 28558 29776 28902
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29840 28218 29868 28494
rect 29920 28484 29972 28490
rect 29920 28426 29972 28432
rect 29828 28212 29880 28218
rect 29828 28154 29880 28160
rect 29932 28150 29960 28426
rect 29276 28144 29328 28150
rect 29276 28086 29328 28092
rect 29644 28144 29696 28150
rect 29644 28086 29696 28092
rect 29920 28144 29972 28150
rect 29920 28086 29972 28092
rect 29276 28008 29328 28014
rect 29276 27950 29328 27956
rect 28908 27600 28960 27606
rect 28908 27542 28960 27548
rect 29184 27600 29236 27606
rect 29184 27542 29236 27548
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 28080 27328 28132 27334
rect 28080 27270 28132 27276
rect 28092 27130 28120 27270
rect 28080 27124 28132 27130
rect 28080 27066 28132 27072
rect 27988 26920 28040 26926
rect 27988 26862 28040 26868
rect 28724 26308 28776 26314
rect 28724 26250 28776 26256
rect 28736 25906 28764 26250
rect 28724 25900 28776 25906
rect 28724 25842 28776 25848
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28908 25900 28960 25906
rect 28908 25842 28960 25848
rect 28722 25800 28778 25809
rect 28722 25735 28778 25744
rect 28736 25702 28764 25735
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28724 25696 28776 25702
rect 28724 25638 28776 25644
rect 28552 25362 28580 25638
rect 28736 25362 28764 25638
rect 28828 25498 28856 25842
rect 28816 25492 28868 25498
rect 28816 25434 28868 25440
rect 28920 25362 28948 25842
rect 29092 25764 29144 25770
rect 29092 25706 29144 25712
rect 29104 25430 29132 25706
rect 29000 25424 29052 25430
rect 29000 25366 29052 25372
rect 29092 25424 29144 25430
rect 29092 25366 29144 25372
rect 28540 25356 28592 25362
rect 28540 25298 28592 25304
rect 28724 25356 28776 25362
rect 28724 25298 28776 25304
rect 28908 25356 28960 25362
rect 28908 25298 28960 25304
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 27344 25094 27396 25100
rect 27356 24732 27384 25094
rect 27540 25078 27752 25106
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27540 24834 27568 25078
rect 27620 24948 27672 24954
rect 27816 24936 27844 25094
rect 27908 24954 27936 25230
rect 29012 25158 29040 25366
rect 29196 25226 29224 27406
rect 29288 26994 29316 27950
rect 29828 27600 29880 27606
rect 29828 27542 29880 27548
rect 29840 27062 29868 27542
rect 30024 27470 30052 31622
rect 30104 31340 30156 31346
rect 30104 31282 30156 31288
rect 30116 30326 30144 31282
rect 30300 31278 30328 31708
rect 30392 31482 30420 31758
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 30576 31346 30604 32166
rect 30668 32026 30696 32166
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 30760 31754 30788 35550
rect 30852 34406 30880 35566
rect 31036 35494 31064 36042
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 30932 34672 30984 34678
rect 30932 34614 30984 34620
rect 30840 34400 30892 34406
rect 30840 34342 30892 34348
rect 30944 33658 30972 34614
rect 30932 33652 30984 33658
rect 30932 33594 30984 33600
rect 31024 32768 31076 32774
rect 31024 32710 31076 32716
rect 31036 32230 31064 32710
rect 31024 32224 31076 32230
rect 31024 32166 31076 32172
rect 30668 31726 30788 31754
rect 30564 31340 30616 31346
rect 30564 31282 30616 31288
rect 30288 31272 30340 31278
rect 30288 31214 30340 31220
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 30104 30320 30156 30326
rect 30156 30280 30236 30308
rect 30104 30262 30156 30268
rect 30208 30190 30236 30280
rect 30392 30190 30420 30670
rect 30576 30394 30604 30670
rect 30564 30388 30616 30394
rect 30564 30330 30616 30336
rect 30196 30184 30248 30190
rect 30196 30126 30248 30132
rect 30380 30184 30432 30190
rect 30380 30126 30432 30132
rect 30208 29646 30236 30126
rect 30288 30048 30340 30054
rect 30288 29990 30340 29996
rect 30300 29646 30328 29990
rect 30196 29640 30248 29646
rect 30196 29582 30248 29588
rect 30288 29640 30340 29646
rect 30576 29628 30604 30330
rect 30668 29730 30696 31726
rect 30748 31340 30800 31346
rect 30748 31282 30800 31288
rect 30760 30258 30788 31282
rect 31024 31272 31076 31278
rect 31024 31214 31076 31220
rect 31036 30938 31064 31214
rect 31024 30932 31076 30938
rect 31024 30874 31076 30880
rect 30840 30864 30892 30870
rect 30840 30806 30892 30812
rect 30852 30394 30880 30806
rect 30840 30388 30892 30394
rect 30840 30330 30892 30336
rect 30748 30252 30800 30258
rect 30748 30194 30800 30200
rect 30760 29850 30788 30194
rect 31128 30138 31156 38626
rect 31392 38208 31444 38214
rect 31392 38150 31444 38156
rect 31404 38010 31432 38150
rect 31392 38004 31444 38010
rect 31392 37946 31444 37952
rect 31300 37868 31352 37874
rect 31300 37810 31352 37816
rect 31312 36922 31340 37810
rect 31956 37262 31984 38898
rect 32140 37874 32168 41618
rect 32232 41138 32260 41754
rect 32876 41614 32904 41754
rect 32968 41614 32996 41958
rect 34808 41818 34836 42162
rect 35348 42152 35400 42158
rect 35348 42094 35400 42100
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 35360 41818 35388 42094
rect 33048 41812 33100 41818
rect 33048 41754 33100 41760
rect 34796 41812 34848 41818
rect 34796 41754 34848 41760
rect 35348 41812 35400 41818
rect 35348 41754 35400 41760
rect 32404 41608 32456 41614
rect 32404 41550 32456 41556
rect 32772 41608 32824 41614
rect 32772 41550 32824 41556
rect 32864 41608 32916 41614
rect 32864 41550 32916 41556
rect 32956 41608 33008 41614
rect 32956 41550 33008 41556
rect 32416 41138 32444 41550
rect 32680 41472 32732 41478
rect 32680 41414 32732 41420
rect 32220 41132 32272 41138
rect 32220 41074 32272 41080
rect 32404 41132 32456 41138
rect 32404 41074 32456 41080
rect 32416 40186 32444 41074
rect 32496 41064 32548 41070
rect 32496 41006 32548 41012
rect 32404 40180 32456 40186
rect 32404 40122 32456 40128
rect 32220 39976 32272 39982
rect 32220 39918 32272 39924
rect 32404 39976 32456 39982
rect 32508 39964 32536 41006
rect 32692 40594 32720 41414
rect 32784 41206 32812 41550
rect 32772 41200 32824 41206
rect 32772 41142 32824 41148
rect 32864 41064 32916 41070
rect 32864 41006 32916 41012
rect 32772 40928 32824 40934
rect 32772 40870 32824 40876
rect 32680 40588 32732 40594
rect 32680 40530 32732 40536
rect 32784 40526 32812 40870
rect 32876 40730 32904 41006
rect 32864 40724 32916 40730
rect 32864 40666 32916 40672
rect 32968 40594 32996 41550
rect 33060 41018 33088 41754
rect 35636 41750 35664 42162
rect 36084 42016 36136 42022
rect 36084 41958 36136 41964
rect 35624 41744 35676 41750
rect 35624 41686 35676 41692
rect 34520 41608 34572 41614
rect 35716 41608 35768 41614
rect 34520 41550 34572 41556
rect 35452 41568 35716 41596
rect 33232 41200 33284 41206
rect 33232 41142 33284 41148
rect 34152 41200 34204 41206
rect 34152 41142 34204 41148
rect 33140 41064 33192 41070
rect 33060 41012 33140 41018
rect 33060 41006 33192 41012
rect 33060 40990 33180 41006
rect 33244 40730 33272 41142
rect 33324 40928 33376 40934
rect 33324 40870 33376 40876
rect 33232 40724 33284 40730
rect 33232 40666 33284 40672
rect 32956 40588 33008 40594
rect 32956 40530 33008 40536
rect 32772 40520 32824 40526
rect 32772 40462 32824 40468
rect 32456 39936 32536 39964
rect 32404 39918 32456 39924
rect 32232 39642 32260 39918
rect 32220 39636 32272 39642
rect 32220 39578 32272 39584
rect 32312 39568 32364 39574
rect 32312 39510 32364 39516
rect 32324 39098 32352 39510
rect 32312 39092 32364 39098
rect 32312 39034 32364 39040
rect 32416 38350 32444 39918
rect 32496 39500 32548 39506
rect 32496 39442 32548 39448
rect 32508 39098 32536 39442
rect 32772 39296 32824 39302
rect 32772 39238 32824 39244
rect 32784 39098 32812 39238
rect 32496 39092 32548 39098
rect 32496 39034 32548 39040
rect 32772 39092 32824 39098
rect 32772 39034 32824 39040
rect 33046 38992 33102 39001
rect 32496 38956 32548 38962
rect 32496 38898 32548 38904
rect 32772 38946 32824 38952
rect 32404 38344 32456 38350
rect 32404 38286 32456 38292
rect 32312 38276 32364 38282
rect 32312 38218 32364 38224
rect 32128 37868 32180 37874
rect 32128 37810 32180 37816
rect 31852 37256 31904 37262
rect 31852 37198 31904 37204
rect 31944 37256 31996 37262
rect 31944 37198 31996 37204
rect 31392 37188 31444 37194
rect 31392 37130 31444 37136
rect 31404 36922 31432 37130
rect 31668 37120 31720 37126
rect 31668 37062 31720 37068
rect 31300 36916 31352 36922
rect 31300 36858 31352 36864
rect 31392 36916 31444 36922
rect 31392 36858 31444 36864
rect 31312 36242 31340 36858
rect 31576 36780 31628 36786
rect 31576 36722 31628 36728
rect 31588 36582 31616 36722
rect 31576 36576 31628 36582
rect 31576 36518 31628 36524
rect 31300 36236 31352 36242
rect 31220 36196 31300 36224
rect 31220 35834 31248 36196
rect 31300 36178 31352 36184
rect 31484 36236 31536 36242
rect 31484 36178 31536 36184
rect 31208 35828 31260 35834
rect 31208 35770 31260 35776
rect 31220 35630 31248 35770
rect 31208 35624 31260 35630
rect 31208 35566 31260 35572
rect 31496 34202 31524 36178
rect 31588 35698 31616 36518
rect 31576 35692 31628 35698
rect 31576 35634 31628 35640
rect 31680 35290 31708 37062
rect 31864 36258 31892 37198
rect 31956 36922 31984 37198
rect 31944 36916 31996 36922
rect 31944 36858 31996 36864
rect 31864 36242 31984 36258
rect 31864 36236 31996 36242
rect 31864 36230 31944 36236
rect 31944 36178 31996 36184
rect 31668 35284 31720 35290
rect 31668 35226 31720 35232
rect 31944 35148 31996 35154
rect 31944 35090 31996 35096
rect 31760 34944 31812 34950
rect 31760 34886 31812 34892
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 31484 34196 31536 34202
rect 31484 34138 31536 34144
rect 31300 32836 31352 32842
rect 31300 32778 31352 32784
rect 31312 32298 31340 32778
rect 31300 32292 31352 32298
rect 31300 32234 31352 32240
rect 31208 31816 31260 31822
rect 31208 31758 31260 31764
rect 30840 30116 30892 30122
rect 30840 30058 30892 30064
rect 30944 30110 31156 30138
rect 30748 29844 30800 29850
rect 30748 29786 30800 29792
rect 30668 29702 30788 29730
rect 30656 29640 30708 29646
rect 30576 29600 30656 29628
rect 30288 29582 30340 29588
rect 30656 29582 30708 29588
rect 30208 28558 30236 29582
rect 30564 29504 30616 29510
rect 30564 29446 30616 29452
rect 30472 29164 30524 29170
rect 30576 29152 30604 29446
rect 30524 29124 30604 29152
rect 30472 29106 30524 29112
rect 30472 29028 30524 29034
rect 30472 28970 30524 28976
rect 30656 29028 30708 29034
rect 30656 28970 30708 28976
rect 30196 28552 30248 28558
rect 30196 28494 30248 28500
rect 30104 28144 30156 28150
rect 30104 28086 30156 28092
rect 30116 27946 30144 28086
rect 30104 27940 30156 27946
rect 30104 27882 30156 27888
rect 30208 27538 30236 28494
rect 30484 28014 30512 28970
rect 30668 28762 30696 28970
rect 30656 28756 30708 28762
rect 30656 28698 30708 28704
rect 30760 28422 30788 29702
rect 30852 28966 30880 30058
rect 30944 29238 30972 30110
rect 31024 30048 31076 30054
rect 31024 29990 31076 29996
rect 31036 29510 31064 29990
rect 31116 29640 31168 29646
rect 31220 29628 31248 31758
rect 31168 29600 31248 29628
rect 31116 29582 31168 29588
rect 31024 29504 31076 29510
rect 31024 29446 31076 29452
rect 30932 29232 30984 29238
rect 30932 29174 30984 29180
rect 30944 29073 30972 29174
rect 31024 29164 31076 29170
rect 31024 29106 31076 29112
rect 30930 29064 30986 29073
rect 30930 28999 30986 29008
rect 30840 28960 30892 28966
rect 30840 28902 30892 28908
rect 31036 28422 31064 29106
rect 31128 28558 31156 29582
rect 31208 28688 31260 28694
rect 31208 28630 31260 28636
rect 31116 28552 31168 28558
rect 31116 28494 31168 28500
rect 30748 28416 30800 28422
rect 30748 28358 30800 28364
rect 31024 28416 31076 28422
rect 31024 28358 31076 28364
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 29920 27328 29972 27334
rect 29920 27270 29972 27276
rect 29828 27056 29880 27062
rect 29828 26998 29880 27004
rect 29932 26994 29960 27270
rect 30760 27062 30788 28358
rect 31128 28218 31156 28494
rect 31116 28212 31168 28218
rect 31116 28154 31168 28160
rect 30932 28144 30984 28150
rect 30932 28086 30984 28092
rect 30944 28014 30972 28086
rect 30932 28008 30984 28014
rect 30932 27950 30984 27956
rect 30840 27872 30892 27878
rect 30840 27814 30892 27820
rect 30852 27577 30880 27814
rect 30838 27568 30894 27577
rect 30838 27503 30894 27512
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30748 27056 30800 27062
rect 30748 26998 30800 27004
rect 29276 26988 29328 26994
rect 29276 26930 29328 26936
rect 29920 26988 29972 26994
rect 29920 26930 29972 26936
rect 29288 25838 29316 26930
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 29564 25838 29592 26318
rect 29276 25832 29328 25838
rect 29276 25774 29328 25780
rect 29552 25832 29604 25838
rect 29552 25774 29604 25780
rect 29184 25220 29236 25226
rect 29184 25162 29236 25168
rect 28080 25152 28132 25158
rect 28080 25094 28132 25100
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 27672 24908 27844 24936
rect 27896 24948 27948 24954
rect 27620 24890 27672 24896
rect 27896 24890 27948 24896
rect 28092 24886 28120 25094
rect 28080 24880 28132 24886
rect 27540 24806 27752 24834
rect 28080 24822 28132 24828
rect 27528 24744 27580 24750
rect 27356 24704 27528 24732
rect 27160 24676 27212 24682
rect 27160 24618 27212 24624
rect 27448 23526 27476 24704
rect 27528 24686 27580 24692
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27448 23186 27476 23462
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27448 22710 27476 23122
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27264 22234 27292 22578
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 27724 22030 27752 24806
rect 29012 24206 29040 25094
rect 29196 24682 29224 25162
rect 29184 24676 29236 24682
rect 29184 24618 29236 24624
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28276 23322 28304 23666
rect 28264 23316 28316 23322
rect 28264 23258 28316 23264
rect 28264 23044 28316 23050
rect 28264 22986 28316 22992
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 28184 21690 28212 21830
rect 28172 21684 28224 21690
rect 28172 21626 28224 21632
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 27264 21350 27292 21422
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27264 20398 27292 21286
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 27448 20466 27476 20946
rect 27540 20806 27568 21286
rect 27724 20874 27752 21286
rect 27712 20868 27764 20874
rect 27712 20810 27764 20816
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27540 20602 27568 20742
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27252 20392 27304 20398
rect 27252 20334 27304 20340
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 27080 19514 27108 19994
rect 27172 19854 27200 20198
rect 27356 20058 27384 20402
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 27448 19922 27476 20402
rect 27436 19916 27488 19922
rect 27436 19858 27488 19864
rect 28080 19916 28132 19922
rect 28080 19858 28132 19864
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27172 18426 27200 19790
rect 27448 19378 27476 19858
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27160 18420 27212 18426
rect 27160 18362 27212 18368
rect 27068 18284 27120 18290
rect 26988 18244 27068 18272
rect 26988 17542 27016 18244
rect 27068 18226 27120 18232
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 27080 16794 27108 17546
rect 27172 17134 27200 18362
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27264 17270 27292 18226
rect 27712 17672 27764 17678
rect 27712 17614 27764 17620
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27528 17536 27580 17542
rect 27528 17478 27580 17484
rect 27356 17338 27384 17478
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27252 17264 27304 17270
rect 27540 17241 27568 17478
rect 27252 17206 27304 17212
rect 27526 17232 27582 17241
rect 27724 17202 27752 17614
rect 27896 17604 27948 17610
rect 27896 17546 27948 17552
rect 27908 17202 27936 17546
rect 27526 17167 27582 17176
rect 27712 17196 27764 17202
rect 27712 17138 27764 17144
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 27160 17128 27212 17134
rect 27160 17070 27212 17076
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 27344 16244 27396 16250
rect 27344 16186 27396 16192
rect 27356 15706 27384 16186
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27724 15570 27752 17138
rect 28092 16114 28120 19858
rect 28172 19712 28224 19718
rect 28172 19654 28224 19660
rect 28184 19446 28212 19654
rect 28172 19440 28224 19446
rect 28172 19382 28224 19388
rect 28172 19304 28224 19310
rect 28172 19246 28224 19252
rect 28184 18970 28212 19246
rect 28172 18964 28224 18970
rect 28172 18906 28224 18912
rect 28080 16108 28132 16114
rect 28000 16068 28080 16096
rect 27712 15564 27764 15570
rect 27712 15506 27764 15512
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27540 15026 27568 15370
rect 27724 15178 27752 15506
rect 27632 15150 27752 15178
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27632 14958 27660 15150
rect 27620 14952 27672 14958
rect 27620 14894 27672 14900
rect 28000 14770 28028 16068
rect 28080 16050 28132 16056
rect 28080 14816 28132 14822
rect 28000 14764 28080 14770
rect 28000 14758 28132 14764
rect 28000 14742 28120 14758
rect 26884 14612 26936 14618
rect 26884 14554 26936 14560
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27252 14544 27304 14550
rect 27252 14486 27304 14492
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26804 12918 26832 13806
rect 26792 12912 26844 12918
rect 26792 12854 26844 12860
rect 26884 12368 26936 12374
rect 26882 12336 26884 12345
rect 26936 12336 26938 12345
rect 26700 12300 26752 12306
rect 26882 12271 26938 12280
rect 26700 12242 26752 12248
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26200 11172 26280 11200
rect 26148 11154 26200 11160
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 24860 10736 24912 10742
rect 25596 10736 25648 10742
rect 24860 10678 24912 10684
rect 25594 10704 25596 10713
rect 25648 10704 25650 10713
rect 25594 10639 25650 10648
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 23940 9648 23992 9654
rect 23940 9590 23992 9596
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 23848 8832 23900 8838
rect 23848 8774 23900 8780
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23860 8430 23888 8774
rect 24044 8430 24072 9318
rect 24136 9178 24164 10066
rect 24228 9654 24256 10066
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24228 9058 24256 9590
rect 24688 9382 24716 10542
rect 25700 9722 25728 10542
rect 25792 10130 25820 11086
rect 27080 10962 27108 14350
rect 27264 14006 27292 14486
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 27436 13184 27488 13190
rect 27436 13126 27488 13132
rect 27448 12918 27476 13126
rect 27436 12912 27488 12918
rect 27436 12854 27488 12860
rect 27724 12238 27752 14554
rect 28000 13870 28028 14742
rect 28276 14618 28304 22986
rect 28356 22432 28408 22438
rect 28356 22374 28408 22380
rect 28368 22098 28396 22374
rect 28356 22092 28408 22098
rect 28356 22034 28408 22040
rect 28736 21078 28764 24142
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28828 23662 28856 24006
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 29012 23730 29040 23802
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28828 22982 28856 23598
rect 29000 23588 29052 23594
rect 29000 23530 29052 23536
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28920 23118 28948 23462
rect 29012 23118 29040 23530
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29196 23050 29224 24618
rect 29184 23044 29236 23050
rect 29184 22986 29236 22992
rect 28816 22976 28868 22982
rect 28816 22918 28868 22924
rect 28828 22166 28856 22918
rect 28816 22160 28868 22166
rect 28816 22102 28868 22108
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28920 21146 28948 21422
rect 28908 21140 28960 21146
rect 28908 21082 28960 21088
rect 28724 21072 28776 21078
rect 28724 21014 28776 21020
rect 28448 20392 28500 20398
rect 28448 20334 28500 20340
rect 28460 20058 28488 20334
rect 28448 20052 28500 20058
rect 28448 19994 28500 20000
rect 28724 19780 28776 19786
rect 28724 19722 28776 19728
rect 28736 19514 28764 19722
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 28736 18766 28764 19450
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 28368 17882 28396 18702
rect 28448 18692 28500 18698
rect 28448 18634 28500 18640
rect 28460 18426 28488 18634
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28356 17876 28408 17882
rect 28356 17818 28408 17824
rect 28552 17814 28580 18702
rect 28632 18624 28684 18630
rect 28632 18566 28684 18572
rect 28644 18426 28672 18566
rect 28632 18420 28684 18426
rect 28632 18362 28684 18368
rect 28920 18306 28948 21082
rect 29288 20584 29316 25774
rect 29564 24410 29592 25774
rect 29736 25696 29788 25702
rect 29736 25638 29788 25644
rect 29748 24886 29776 25638
rect 29736 24880 29788 24886
rect 29736 24822 29788 24828
rect 29828 24608 29880 24614
rect 29828 24550 29880 24556
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 29840 24206 29868 24550
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29840 24070 29868 24142
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29932 23866 29960 26930
rect 30012 25900 30064 25906
rect 30380 25900 30432 25906
rect 30064 25860 30380 25888
rect 30012 25842 30064 25848
rect 30380 25842 30432 25848
rect 30012 25764 30064 25770
rect 30012 25706 30064 25712
rect 30380 25764 30432 25770
rect 30380 25706 30432 25712
rect 30024 25294 30052 25706
rect 30392 25498 30420 25706
rect 30380 25492 30432 25498
rect 30380 25434 30432 25440
rect 30012 25288 30064 25294
rect 30748 25288 30800 25294
rect 30012 25230 30064 25236
rect 30746 25256 30748 25265
rect 30800 25256 30802 25265
rect 30852 25226 30880 27406
rect 31128 25362 31156 28154
rect 31220 27849 31248 28630
rect 31312 28558 31340 32234
rect 31392 32224 31444 32230
rect 31392 32166 31444 32172
rect 31300 28552 31352 28558
rect 31300 28494 31352 28500
rect 31312 28218 31340 28494
rect 31300 28212 31352 28218
rect 31300 28154 31352 28160
rect 31206 27840 31262 27849
rect 31206 27775 31262 27784
rect 31404 27334 31432 32166
rect 31588 31686 31616 34546
rect 31772 34066 31800 34886
rect 31956 34474 31984 35090
rect 32140 34950 32168 37810
rect 32324 36854 32352 38218
rect 32416 37942 32444 38286
rect 32404 37936 32456 37942
rect 32404 37878 32456 37884
rect 32508 37126 32536 38898
rect 33046 38927 33048 38936
rect 33100 38927 33102 38936
rect 33048 38898 33100 38904
rect 32680 38888 32732 38894
rect 32772 38888 32824 38894
rect 32680 38830 32732 38836
rect 32692 38758 32720 38830
rect 32680 38752 32732 38758
rect 32680 38694 32732 38700
rect 32784 38418 32812 38888
rect 32956 38752 33008 38758
rect 32956 38694 33008 38700
rect 32772 38412 32824 38418
rect 32772 38354 32824 38360
rect 32680 38276 32732 38282
rect 32680 38218 32732 38224
rect 32692 38010 32720 38218
rect 32680 38004 32732 38010
rect 32680 37946 32732 37952
rect 32968 37942 32996 38694
rect 33244 38282 33272 40666
rect 33336 40458 33364 40870
rect 34164 40730 34192 41142
rect 34152 40724 34204 40730
rect 34152 40666 34204 40672
rect 33324 40452 33376 40458
rect 33324 40394 33376 40400
rect 33232 38276 33284 38282
rect 33232 38218 33284 38224
rect 32956 37936 33008 37942
rect 32956 37878 33008 37884
rect 33140 37868 33192 37874
rect 33140 37810 33192 37816
rect 33152 37262 33180 37810
rect 32772 37256 32824 37262
rect 32772 37198 32824 37204
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32312 36848 32364 36854
rect 32312 36790 32364 36796
rect 32496 36848 32548 36854
rect 32496 36790 32548 36796
rect 32404 35624 32456 35630
rect 32404 35566 32456 35572
rect 32220 35012 32272 35018
rect 32220 34954 32272 34960
rect 32036 34944 32088 34950
rect 32036 34886 32088 34892
rect 32128 34944 32180 34950
rect 32128 34886 32180 34892
rect 31944 34468 31996 34474
rect 31944 34410 31996 34416
rect 31760 34060 31812 34066
rect 31760 34002 31812 34008
rect 32048 33862 32076 34886
rect 32128 34468 32180 34474
rect 32128 34410 32180 34416
rect 32140 34066 32168 34410
rect 32128 34060 32180 34066
rect 32128 34002 32180 34008
rect 32232 33930 32260 34954
rect 32416 34610 32444 35566
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32312 33992 32364 33998
rect 32312 33934 32364 33940
rect 32220 33924 32272 33930
rect 32220 33866 32272 33872
rect 32036 33856 32088 33862
rect 32036 33798 32088 33804
rect 32048 32756 32076 33798
rect 32128 33312 32180 33318
rect 32128 33254 32180 33260
rect 32140 32910 32168 33254
rect 32324 33114 32352 33934
rect 32312 33108 32364 33114
rect 32312 33050 32364 33056
rect 32128 32904 32180 32910
rect 32128 32846 32180 32852
rect 32048 32728 32168 32756
rect 32140 32366 32168 32728
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 32140 32026 32168 32302
rect 32128 32020 32180 32026
rect 32128 31962 32180 31968
rect 32128 31748 32180 31754
rect 32128 31690 32180 31696
rect 31576 31680 31628 31686
rect 31576 31622 31628 31628
rect 31588 30802 31616 31622
rect 32140 30938 32168 31690
rect 32508 31498 32536 36790
rect 32784 36174 32812 37198
rect 32772 36168 32824 36174
rect 32772 36110 32824 36116
rect 32680 36032 32732 36038
rect 32680 35974 32732 35980
rect 32692 34678 32720 35974
rect 32784 35834 32812 36110
rect 32772 35828 32824 35834
rect 32772 35770 32824 35776
rect 33244 35494 33272 38218
rect 33232 35488 33284 35494
rect 33232 35430 33284 35436
rect 33048 34944 33100 34950
rect 33048 34886 33100 34892
rect 32680 34672 32732 34678
rect 32680 34614 32732 34620
rect 32588 33856 32640 33862
rect 32588 33798 32640 33804
rect 32600 33658 32628 33798
rect 32588 33652 32640 33658
rect 32588 33594 32640 33600
rect 32588 33516 32640 33522
rect 32588 33458 32640 33464
rect 32600 31686 32628 33458
rect 32680 33380 32732 33386
rect 32680 33322 32732 33328
rect 32588 31680 32640 31686
rect 32588 31622 32640 31628
rect 32508 31470 32628 31498
rect 32496 31340 32548 31346
rect 32496 31282 32548 31288
rect 32128 30932 32180 30938
rect 32128 30874 32180 30880
rect 32508 30870 32536 31282
rect 32496 30864 32548 30870
rect 32496 30806 32548 30812
rect 31576 30796 31628 30802
rect 31576 30738 31628 30744
rect 31576 30592 31628 30598
rect 31576 30534 31628 30540
rect 31588 30258 31616 30534
rect 32508 30326 32536 30806
rect 32496 30320 32548 30326
rect 32496 30262 32548 30268
rect 31484 30252 31536 30258
rect 31484 30194 31536 30200
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31668 30252 31720 30258
rect 31668 30194 31720 30200
rect 31496 30138 31524 30194
rect 31496 30110 31616 30138
rect 31484 30048 31536 30054
rect 31484 29990 31536 29996
rect 31496 29714 31524 29990
rect 31484 29708 31536 29714
rect 31484 29650 31536 29656
rect 31484 29164 31536 29170
rect 31484 29106 31536 29112
rect 31496 27470 31524 29106
rect 31588 29034 31616 30110
rect 31680 29850 31708 30194
rect 32220 30184 32272 30190
rect 32218 30152 32220 30161
rect 32272 30152 32274 30161
rect 32218 30087 32274 30096
rect 31668 29844 31720 29850
rect 31668 29786 31720 29792
rect 32508 29782 32536 30262
rect 32496 29776 32548 29782
rect 32496 29718 32548 29724
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31668 29164 31720 29170
rect 31668 29106 31720 29112
rect 31576 29028 31628 29034
rect 31576 28970 31628 28976
rect 31588 27860 31616 28970
rect 31680 28694 31708 29106
rect 31772 29102 31800 29446
rect 32508 29306 32536 29718
rect 32496 29300 32548 29306
rect 32496 29242 32548 29248
rect 32312 29232 32364 29238
rect 32312 29174 32364 29180
rect 31760 29096 31812 29102
rect 31760 29038 31812 29044
rect 31668 28688 31720 28694
rect 31668 28630 31720 28636
rect 31668 28416 31720 28422
rect 31668 28358 31720 28364
rect 31680 28014 31708 28358
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31760 27872 31812 27878
rect 31588 27832 31760 27860
rect 31760 27814 31812 27820
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31772 27334 31800 27814
rect 31300 27328 31352 27334
rect 31300 27270 31352 27276
rect 31392 27328 31444 27334
rect 31392 27270 31444 27276
rect 31760 27328 31812 27334
rect 31760 27270 31812 27276
rect 31208 25696 31260 25702
rect 31208 25638 31260 25644
rect 31116 25356 31168 25362
rect 31116 25298 31168 25304
rect 31220 25226 31248 25638
rect 30746 25191 30802 25200
rect 30840 25220 30892 25226
rect 30840 25162 30892 25168
rect 31208 25220 31260 25226
rect 31208 25162 31260 25168
rect 30196 25152 30248 25158
rect 30196 25094 30248 25100
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 31024 25152 31076 25158
rect 31024 25094 31076 25100
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 29920 23588 29972 23594
rect 29920 23530 29972 23536
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29472 22234 29500 22510
rect 29460 22228 29512 22234
rect 29460 22170 29512 22176
rect 29932 22094 29960 23530
rect 30012 23520 30064 23526
rect 30012 23462 30064 23468
rect 30024 23050 30052 23462
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 30116 22574 30144 23054
rect 30104 22568 30156 22574
rect 30104 22510 30156 22516
rect 30116 22438 30144 22510
rect 30104 22432 30156 22438
rect 30104 22374 30156 22380
rect 30012 22094 30064 22098
rect 29932 22092 30064 22094
rect 29932 22066 30012 22092
rect 30012 22034 30064 22040
rect 29920 21888 29972 21894
rect 29920 21830 29972 21836
rect 29932 21690 29960 21830
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 30116 21010 30144 22374
rect 30104 21004 30156 21010
rect 30104 20946 30156 20952
rect 29460 20868 29512 20874
rect 29460 20810 29512 20816
rect 29368 20596 29420 20602
rect 29288 20556 29368 20584
rect 29288 19854 29316 20556
rect 29368 20538 29420 20544
rect 29472 20534 29500 20810
rect 29460 20528 29512 20534
rect 29460 20470 29512 20476
rect 29276 19848 29328 19854
rect 29276 19790 29328 19796
rect 29276 18828 29328 18834
rect 29276 18770 29328 18776
rect 29184 18624 29236 18630
rect 29184 18566 29236 18572
rect 29196 18426 29224 18566
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 28828 18278 28948 18306
rect 28540 17808 28592 17814
rect 28540 17750 28592 17756
rect 28356 17740 28408 17746
rect 28356 17682 28408 17688
rect 28632 17740 28684 17746
rect 28632 17682 28684 17688
rect 28368 16114 28396 17682
rect 28446 17232 28502 17241
rect 28446 17167 28448 17176
rect 28500 17167 28502 17176
rect 28540 17196 28592 17202
rect 28448 17138 28500 17144
rect 28540 17138 28592 17144
rect 28552 16998 28580 17138
rect 28644 16998 28672 17682
rect 28828 17678 28856 18278
rect 29092 18216 29144 18222
rect 29092 18158 29144 18164
rect 28908 18080 28960 18086
rect 28908 18022 28960 18028
rect 28920 17678 28948 18022
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28908 17672 28960 17678
rect 28908 17614 28960 17620
rect 28920 16998 28948 17614
rect 29104 17542 29132 18158
rect 29196 17678 29224 18362
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 29092 17536 29144 17542
rect 29092 17478 29144 17484
rect 29012 17202 29040 17478
rect 29196 17338 29224 17614
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 29012 17066 29040 17138
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 29092 17060 29144 17066
rect 29092 17002 29144 17008
rect 28540 16992 28592 16998
rect 28540 16934 28592 16940
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28446 16824 28502 16833
rect 28906 16824 28962 16833
rect 28446 16759 28502 16768
rect 28644 16782 28856 16810
rect 28460 16658 28488 16759
rect 28644 16726 28672 16782
rect 28828 16726 28856 16782
rect 29104 16794 29132 17002
rect 28906 16759 28908 16768
rect 28960 16759 28962 16768
rect 29092 16788 29144 16794
rect 28908 16730 28960 16736
rect 29092 16730 29144 16736
rect 29196 16726 29224 17070
rect 28632 16720 28684 16726
rect 28632 16662 28684 16668
rect 28724 16720 28776 16726
rect 28724 16662 28776 16668
rect 28816 16720 28868 16726
rect 28816 16662 28868 16668
rect 29184 16720 29236 16726
rect 29184 16662 29236 16668
rect 28448 16652 28500 16658
rect 28448 16594 28500 16600
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28368 15570 28396 16050
rect 28736 15910 28764 16662
rect 28908 16586 28960 16592
rect 28960 16534 28994 16538
rect 28908 16528 28994 16534
rect 28920 16510 28994 16528
rect 28966 16504 28994 16510
rect 29184 16516 29236 16522
rect 28966 16476 29132 16504
rect 28998 16280 29054 16289
rect 28920 16250 28998 16266
rect 28908 16244 28998 16250
rect 28960 16238 28998 16244
rect 28998 16215 29054 16224
rect 28908 16186 28960 16192
rect 28724 15904 28776 15910
rect 28724 15846 28776 15852
rect 29012 15706 29040 16215
rect 29104 16046 29132 16476
rect 29184 16458 29236 16464
rect 29196 16289 29224 16458
rect 29182 16280 29238 16289
rect 29182 16215 29238 16224
rect 29092 16040 29144 16046
rect 29092 15982 29144 15988
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 29104 15502 29132 15642
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29196 15366 29224 15846
rect 28448 15360 28500 15366
rect 28448 15302 28500 15308
rect 29184 15360 29236 15366
rect 29184 15302 29236 15308
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 28276 14414 28304 14554
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 28184 12442 28212 13262
rect 28172 12436 28224 12442
rect 28172 12378 28224 12384
rect 27712 12232 27764 12238
rect 27712 12174 27764 12180
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27172 11830 27200 12038
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27448 11082 27476 11698
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27540 11354 27568 11630
rect 27908 11354 27936 11698
rect 27988 11688 28040 11694
rect 27988 11630 28040 11636
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 28000 11150 28028 11630
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 27436 11076 27488 11082
rect 27436 11018 27488 11024
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 27080 10934 27292 10962
rect 27264 10656 27292 10934
rect 27344 10668 27396 10674
rect 27264 10628 27344 10656
rect 27344 10610 27396 10616
rect 26516 10600 26568 10606
rect 26516 10542 26568 10548
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25884 9722 25912 10202
rect 26424 9988 26476 9994
rect 26424 9930 26476 9936
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25872 9716 25924 9722
rect 25872 9658 25924 9664
rect 26240 9512 26292 9518
rect 26238 9480 26240 9489
rect 26292 9480 26294 9489
rect 26238 9415 26294 9424
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24688 9178 24716 9318
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24136 9030 24256 9058
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 24136 8906 24164 9030
rect 24412 8974 24440 9046
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23492 7750 23520 8230
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23204 7472 23256 7478
rect 23202 7440 23204 7449
rect 23256 7440 23258 7449
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 22836 7404 22888 7410
rect 23860 7410 23888 8366
rect 24044 7478 24072 8366
rect 24136 7818 24164 8842
rect 24412 8498 24440 8910
rect 26436 8634 26464 9930
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 26436 8498 26464 8570
rect 26528 8566 26556 10542
rect 27356 10470 27384 10610
rect 26976 10464 27028 10470
rect 26976 10406 27028 10412
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 26988 10266 27016 10406
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 27356 9994 27384 10406
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27344 9648 27396 9654
rect 26606 9616 26662 9625
rect 27342 9616 27344 9625
rect 27396 9616 27398 9625
rect 26606 9551 26608 9560
rect 26660 9551 26662 9560
rect 26896 9586 27200 9602
rect 26896 9580 27212 9586
rect 26896 9574 27160 9580
rect 26608 9522 26660 9528
rect 26620 8974 26648 9522
rect 26896 9518 26924 9574
rect 27342 9551 27398 9560
rect 27160 9522 27212 9528
rect 26884 9512 26936 9518
rect 27068 9512 27120 9518
rect 26884 9454 26936 9460
rect 27066 9480 27068 9489
rect 27120 9480 27122 9489
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26712 8974 26740 9318
rect 26896 9110 26924 9454
rect 27066 9415 27122 9424
rect 26884 9104 26936 9110
rect 26884 9046 26936 9052
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 27080 8498 27108 9415
rect 27448 8838 27476 11018
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27540 9722 27568 10610
rect 27620 10600 27672 10606
rect 27620 10542 27672 10548
rect 27528 9716 27580 9722
rect 27528 9658 27580 9664
rect 27632 9382 27660 10542
rect 27908 10266 27936 11018
rect 28092 10810 28120 11086
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 27896 10260 27948 10266
rect 27896 10202 27948 10208
rect 27908 9994 27936 10202
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27896 9988 27948 9994
rect 27896 9930 27948 9936
rect 27724 9722 27752 9930
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 28092 9654 28120 10746
rect 28184 10470 28212 10746
rect 28276 10713 28304 14350
rect 28368 13394 28396 14350
rect 28356 13388 28408 13394
rect 28356 13330 28408 13336
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28368 11082 28396 11494
rect 28356 11076 28408 11082
rect 28356 11018 28408 11024
rect 28262 10704 28318 10713
rect 28262 10639 28318 10648
rect 28172 10464 28224 10470
rect 28172 10406 28224 10412
rect 28276 9722 28304 10639
rect 28264 9716 28316 9722
rect 28264 9658 28316 9664
rect 28080 9648 28132 9654
rect 28080 9590 28132 9596
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27632 9042 27660 9318
rect 27620 9036 27672 9042
rect 27620 8978 27672 8984
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27160 8832 27212 8838
rect 27160 8774 27212 8780
rect 27436 8832 27488 8838
rect 27436 8774 27488 8780
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 24124 7812 24176 7818
rect 24124 7754 24176 7760
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 24136 7426 24164 7754
rect 24412 7546 24440 8434
rect 25240 8090 25268 8434
rect 27172 8430 27200 8774
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 27160 8424 27212 8430
rect 27160 8366 27212 8372
rect 26332 8356 26384 8362
rect 26332 8298 26384 8304
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 24504 7426 24532 7482
rect 25424 7478 25452 8230
rect 26344 7954 26372 8298
rect 27448 7954 27476 8434
rect 27540 8090 27568 8910
rect 28092 8906 28120 9454
rect 28460 8974 28488 15302
rect 29182 15192 29238 15201
rect 29182 15127 29238 15136
rect 29196 15026 29224 15127
rect 29184 15020 29236 15026
rect 29184 14962 29236 14968
rect 29092 14952 29144 14958
rect 29092 14894 29144 14900
rect 29104 14362 29132 14894
rect 29012 14346 29132 14362
rect 29000 14340 29132 14346
rect 29052 14334 29132 14340
rect 29000 14282 29052 14288
rect 29012 14006 29040 14282
rect 29000 14000 29052 14006
rect 29000 13942 29052 13948
rect 28816 13728 28868 13734
rect 28816 13670 28868 13676
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 28828 13326 28856 13670
rect 28920 13530 28948 13670
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 29012 13394 29040 13942
rect 29000 13388 29052 13394
rect 29000 13330 29052 13336
rect 28816 13320 28868 13326
rect 28816 13262 28868 13268
rect 28908 12912 28960 12918
rect 28908 12854 28960 12860
rect 28816 12640 28868 12646
rect 28816 12582 28868 12588
rect 28828 12238 28856 12582
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28828 11762 28856 12174
rect 28920 11778 28948 12854
rect 29012 12306 29040 13330
rect 29196 13002 29224 14962
rect 29288 13138 29316 18770
rect 29472 18358 29500 20470
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29736 19304 29788 19310
rect 29736 19246 29788 19252
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 29460 18352 29512 18358
rect 29460 18294 29512 18300
rect 29368 17808 29420 17814
rect 29368 17750 29420 17756
rect 29380 16590 29408 17750
rect 29472 17320 29500 18294
rect 29564 17882 29592 18702
rect 29552 17876 29604 17882
rect 29552 17818 29604 17824
rect 29748 17678 29776 19246
rect 29932 17678 29960 19314
rect 30104 18624 30156 18630
rect 30104 18566 30156 18572
rect 30116 18358 30144 18566
rect 30104 18352 30156 18358
rect 30104 18294 30156 18300
rect 30208 17762 30236 25094
rect 30576 24954 30604 25094
rect 30564 24948 30616 24954
rect 30564 24890 30616 24896
rect 31036 24886 31064 25094
rect 31024 24880 31076 24886
rect 31024 24822 31076 24828
rect 30932 23656 30984 23662
rect 30932 23598 30984 23604
rect 30944 23322 30972 23598
rect 30932 23316 30984 23322
rect 30932 23258 30984 23264
rect 31208 23044 31260 23050
rect 31208 22986 31260 22992
rect 30840 22704 30892 22710
rect 30840 22646 30892 22652
rect 30656 22432 30708 22438
rect 30656 22374 30708 22380
rect 30668 21554 30696 22374
rect 30656 21548 30708 21554
rect 30576 21508 30656 21536
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30392 21010 30420 21286
rect 30380 21004 30432 21010
rect 30380 20946 30432 20952
rect 30380 20868 30432 20874
rect 30380 20810 30432 20816
rect 30392 19718 30420 20810
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30392 18986 30420 19654
rect 30392 18958 30512 18986
rect 30380 18828 30432 18834
rect 30380 18770 30432 18776
rect 30392 18290 30420 18770
rect 30484 18630 30512 18958
rect 30576 18902 30604 21508
rect 30656 21490 30708 21496
rect 30852 20874 30880 22646
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30944 22234 30972 22578
rect 30932 22228 30984 22234
rect 30932 22170 30984 22176
rect 31220 22166 31248 22986
rect 31208 22160 31260 22166
rect 31208 22102 31260 22108
rect 31312 22030 31340 27270
rect 31404 25906 31432 27270
rect 31760 26444 31812 26450
rect 31760 26386 31812 26392
rect 31772 26246 31800 26386
rect 31760 26240 31812 26246
rect 31760 26182 31812 26188
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31404 24750 31432 25842
rect 31772 25838 31800 26182
rect 31760 25832 31812 25838
rect 31760 25774 31812 25780
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 31668 25356 31720 25362
rect 31668 25298 31720 25304
rect 31392 24744 31444 24750
rect 31392 24686 31444 24692
rect 31404 24206 31432 24686
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31404 22982 31432 24142
rect 31680 23186 31708 25298
rect 31864 24818 31892 25434
rect 31956 24886 31984 28018
rect 32324 27402 32352 29174
rect 32404 28484 32456 28490
rect 32404 28426 32456 28432
rect 32416 27674 32444 28426
rect 32600 28150 32628 31470
rect 32692 31278 32720 33322
rect 33060 32298 33088 34886
rect 33140 32836 33192 32842
rect 33140 32778 33192 32784
rect 33152 32570 33180 32778
rect 33140 32564 33192 32570
rect 33140 32506 33192 32512
rect 33048 32292 33100 32298
rect 33048 32234 33100 32240
rect 32772 32224 32824 32230
rect 32772 32166 32824 32172
rect 32784 31482 32812 32166
rect 33336 31906 33364 40394
rect 34428 40384 34480 40390
rect 34428 40326 34480 40332
rect 34440 38962 34468 40326
rect 34428 38956 34480 38962
rect 34428 38898 34480 38904
rect 33692 38208 33744 38214
rect 33692 38150 33744 38156
rect 33416 37868 33468 37874
rect 33416 37810 33468 37816
rect 33428 37126 33456 37810
rect 33416 37120 33468 37126
rect 33416 37062 33468 37068
rect 33416 36032 33468 36038
rect 33416 35974 33468 35980
rect 33428 33658 33456 35974
rect 33416 33652 33468 33658
rect 33416 33594 33468 33600
rect 33416 32496 33468 32502
rect 33416 32438 33468 32444
rect 32968 31878 33364 31906
rect 32864 31680 32916 31686
rect 32864 31622 32916 31628
rect 32772 31476 32824 31482
rect 32772 31418 32824 31424
rect 32680 31272 32732 31278
rect 32680 31214 32732 31220
rect 32772 31136 32824 31142
rect 32772 31078 32824 31084
rect 32784 30802 32812 31078
rect 32772 30796 32824 30802
rect 32772 30738 32824 30744
rect 32876 29306 32904 31622
rect 32968 30297 32996 31878
rect 33428 31822 33456 32438
rect 33508 32428 33560 32434
rect 33508 32370 33560 32376
rect 33324 31816 33376 31822
rect 33324 31758 33376 31764
rect 33416 31816 33468 31822
rect 33416 31758 33468 31764
rect 33336 31482 33364 31758
rect 33324 31476 33376 31482
rect 33324 31418 33376 31424
rect 32954 30288 33010 30297
rect 32954 30223 33010 30232
rect 32968 29510 32996 30223
rect 33416 30184 33468 30190
rect 33416 30126 33468 30132
rect 33428 29714 33456 30126
rect 33416 29708 33468 29714
rect 33416 29650 33468 29656
rect 33060 29578 33456 29594
rect 33048 29572 33456 29578
rect 33100 29566 33456 29572
rect 33048 29514 33100 29520
rect 32956 29504 33008 29510
rect 32956 29446 33008 29452
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 32772 29164 32824 29170
rect 32772 29106 32824 29112
rect 32784 28762 32812 29106
rect 32772 28756 32824 28762
rect 32772 28698 32824 28704
rect 32680 28688 32732 28694
rect 32680 28630 32732 28636
rect 32692 28150 32720 28630
rect 32770 28248 32826 28257
rect 32770 28183 32826 28192
rect 32588 28144 32640 28150
rect 32588 28086 32640 28092
rect 32680 28144 32732 28150
rect 32680 28086 32732 28092
rect 32784 28082 32812 28183
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32404 27668 32456 27674
rect 32404 27610 32456 27616
rect 32312 27396 32364 27402
rect 32312 27338 32364 27344
rect 32324 26994 32352 27338
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 32220 26036 32272 26042
rect 32220 25978 32272 25984
rect 32036 25900 32088 25906
rect 32036 25842 32088 25848
rect 31944 24880 31996 24886
rect 31944 24822 31996 24828
rect 32048 24818 32076 25842
rect 32232 25498 32260 25978
rect 32496 25696 32548 25702
rect 32496 25638 32548 25644
rect 32772 25696 32824 25702
rect 32772 25638 32824 25644
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32508 25226 32536 25638
rect 32678 25392 32734 25401
rect 32678 25327 32680 25336
rect 32732 25327 32734 25336
rect 32680 25298 32732 25304
rect 32784 25294 32812 25638
rect 32876 25498 32904 29242
rect 32956 29232 33008 29238
rect 33140 29232 33192 29238
rect 33008 29192 33140 29220
rect 32956 29174 33008 29180
rect 33140 29174 33192 29180
rect 33244 29170 33272 29446
rect 33232 29164 33284 29170
rect 33232 29106 33284 29112
rect 33048 29096 33100 29102
rect 33048 29038 33100 29044
rect 32956 28960 33008 28966
rect 33060 28937 33088 29038
rect 33140 29028 33192 29034
rect 33140 28970 33192 28976
rect 32956 28902 33008 28908
rect 33046 28928 33102 28937
rect 32968 27402 32996 28902
rect 33046 28863 33102 28872
rect 33048 28756 33100 28762
rect 33048 28698 33100 28704
rect 33060 28082 33088 28698
rect 33048 28076 33100 28082
rect 33048 28018 33100 28024
rect 33048 27940 33100 27946
rect 33048 27882 33100 27888
rect 33060 27674 33088 27882
rect 33048 27668 33100 27674
rect 33048 27610 33100 27616
rect 32956 27396 33008 27402
rect 32956 27338 33008 27344
rect 32956 26240 33008 26246
rect 32956 26182 33008 26188
rect 32968 25974 32996 26182
rect 32956 25968 33008 25974
rect 32956 25910 33008 25916
rect 32864 25492 32916 25498
rect 32864 25434 32916 25440
rect 32772 25288 32824 25294
rect 32772 25230 32824 25236
rect 32496 25220 32548 25226
rect 32496 25162 32548 25168
rect 32508 24970 32536 25162
rect 32508 24942 32628 24970
rect 32600 24886 32628 24942
rect 32588 24880 32640 24886
rect 32588 24822 32640 24828
rect 31852 24812 31904 24818
rect 31852 24754 31904 24760
rect 32036 24812 32088 24818
rect 32036 24754 32088 24760
rect 33048 24812 33100 24818
rect 33048 24754 33100 24760
rect 31760 24744 31812 24750
rect 31760 24686 31812 24692
rect 31772 24138 31800 24686
rect 31864 24426 31892 24754
rect 32680 24744 32732 24750
rect 32680 24686 32732 24692
rect 31864 24398 31984 24426
rect 31956 24342 31984 24398
rect 31944 24336 31996 24342
rect 31944 24278 31996 24284
rect 32404 24336 32456 24342
rect 32404 24278 32456 24284
rect 31760 24132 31812 24138
rect 31760 24074 31812 24080
rect 32312 23860 32364 23866
rect 32312 23802 32364 23808
rect 32324 23730 32352 23802
rect 32416 23730 32444 24278
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32404 23724 32456 23730
rect 32404 23666 32456 23672
rect 32496 23724 32548 23730
rect 32496 23666 32548 23672
rect 32036 23316 32088 23322
rect 32036 23258 32088 23264
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 32048 22778 32076 23258
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32048 22624 32076 22714
rect 32048 22596 32168 22624
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 32048 22098 32076 22374
rect 31392 22092 31444 22098
rect 31392 22034 31444 22040
rect 32036 22092 32088 22098
rect 32036 22034 32088 22040
rect 31300 22024 31352 22030
rect 31300 21966 31352 21972
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 31312 21690 31340 21830
rect 31300 21684 31352 21690
rect 31300 21626 31352 21632
rect 31404 21486 31432 22034
rect 32140 21570 32168 22596
rect 32324 21962 32352 23666
rect 32404 23588 32456 23594
rect 32404 23530 32456 23536
rect 32312 21956 32364 21962
rect 32312 21898 32364 21904
rect 31944 21548 31996 21554
rect 31944 21490 31996 21496
rect 32048 21542 32168 21570
rect 31392 21480 31444 21486
rect 31444 21440 31524 21468
rect 31392 21422 31444 21428
rect 31496 21078 31524 21440
rect 31956 21146 31984 21490
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31484 21072 31536 21078
rect 31484 21014 31536 21020
rect 30840 20868 30892 20874
rect 30840 20810 30892 20816
rect 31208 20392 31260 20398
rect 31208 20334 31260 20340
rect 31220 20058 31248 20334
rect 31208 20052 31260 20058
rect 31208 19994 31260 20000
rect 30656 19304 30708 19310
rect 30656 19246 30708 19252
rect 31496 19258 31524 21014
rect 31760 20800 31812 20806
rect 31760 20742 31812 20748
rect 31668 19712 31720 19718
rect 31668 19654 31720 19660
rect 30564 18896 30616 18902
rect 30564 18838 30616 18844
rect 30472 18624 30524 18630
rect 30472 18566 30524 18572
rect 30576 18358 30604 18838
rect 30668 18698 30696 19246
rect 31496 19230 31616 19258
rect 31484 19168 31536 19174
rect 31484 19110 31536 19116
rect 30656 18692 30708 18698
rect 30656 18634 30708 18640
rect 31208 18692 31260 18698
rect 31208 18634 31260 18640
rect 30668 18358 30696 18634
rect 31024 18624 31076 18630
rect 31024 18566 31076 18572
rect 30564 18352 30616 18358
rect 30564 18294 30616 18300
rect 30656 18352 30708 18358
rect 30656 18294 30708 18300
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30024 17734 30236 17762
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 29828 17604 29880 17610
rect 29828 17546 29880 17552
rect 29472 17292 29684 17320
rect 29460 17196 29512 17202
rect 29460 17138 29512 17144
rect 29472 16658 29500 17138
rect 29460 16652 29512 16658
rect 29460 16594 29512 16600
rect 29368 16584 29420 16590
rect 29368 16526 29420 16532
rect 29460 16516 29512 16522
rect 29460 16458 29512 16464
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29380 14550 29408 15982
rect 29472 15434 29500 16458
rect 29656 16182 29684 17292
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29644 16176 29696 16182
rect 29644 16118 29696 16124
rect 29460 15428 29512 15434
rect 29460 15370 29512 15376
rect 29472 14822 29500 15370
rect 29552 15360 29604 15366
rect 29552 15302 29604 15308
rect 29564 15094 29592 15302
rect 29656 15094 29684 16118
rect 29552 15088 29604 15094
rect 29552 15030 29604 15036
rect 29644 15088 29696 15094
rect 29644 15030 29696 15036
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29368 14544 29420 14550
rect 29368 14486 29420 14492
rect 29472 14414 29500 14758
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29460 14068 29512 14074
rect 29460 14010 29512 14016
rect 29472 13326 29500 14010
rect 29564 14006 29592 14894
rect 29748 14498 29776 16526
rect 29840 16522 29868 17546
rect 29828 16516 29880 16522
rect 29828 16458 29880 16464
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29932 15586 29960 16186
rect 29656 14470 29776 14498
rect 29840 15558 29960 15586
rect 29552 14000 29604 14006
rect 29552 13942 29604 13948
rect 29564 13870 29592 13942
rect 29552 13864 29604 13870
rect 29552 13806 29604 13812
rect 29564 13462 29592 13806
rect 29552 13456 29604 13462
rect 29552 13398 29604 13404
rect 29460 13320 29512 13326
rect 29460 13262 29512 13268
rect 29656 13190 29684 14470
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29644 13184 29696 13190
rect 29288 13110 29592 13138
rect 29644 13126 29696 13132
rect 29196 12974 29316 13002
rect 29184 12640 29236 12646
rect 29184 12582 29236 12588
rect 29196 12374 29224 12582
rect 29184 12368 29236 12374
rect 29184 12310 29236 12316
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 29000 11824 29052 11830
rect 28920 11772 29000 11778
rect 28920 11766 29052 11772
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 28920 11750 29040 11766
rect 28736 11150 28764 11698
rect 28724 11144 28776 11150
rect 28724 11086 28776 11092
rect 28920 11098 28948 11750
rect 28920 11070 29040 11098
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28736 10062 28764 10542
rect 28828 10198 28856 10610
rect 28908 10464 28960 10470
rect 28908 10406 28960 10412
rect 28816 10192 28868 10198
rect 28816 10134 28868 10140
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28828 9654 28856 10134
rect 28920 9654 28948 10406
rect 29012 10266 29040 11070
rect 29288 11014 29316 12974
rect 29276 11008 29328 11014
rect 29276 10950 29328 10956
rect 29092 10804 29144 10810
rect 29092 10746 29144 10752
rect 29104 10674 29132 10746
rect 29092 10668 29144 10674
rect 29092 10610 29144 10616
rect 29092 10532 29144 10538
rect 29092 10474 29144 10480
rect 29000 10260 29052 10266
rect 29000 10202 29052 10208
rect 29104 9926 29132 10474
rect 29288 10062 29316 10950
rect 29564 10810 29592 13110
rect 29656 12646 29684 13126
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29368 10260 29420 10266
rect 29368 10202 29420 10208
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29276 10056 29328 10062
rect 29276 9998 29328 10004
rect 29196 9926 29224 9998
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29184 9920 29236 9926
rect 29184 9862 29236 9868
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28908 9648 28960 9654
rect 28908 9590 28960 9596
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28632 9512 28684 9518
rect 28632 9454 28684 9460
rect 28552 9178 28580 9454
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28080 8900 28132 8906
rect 28080 8842 28132 8848
rect 28092 8362 28120 8842
rect 28172 8832 28224 8838
rect 28172 8774 28224 8780
rect 28356 8832 28408 8838
rect 28356 8774 28408 8780
rect 28184 8566 28212 8774
rect 28368 8566 28396 8774
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 28356 8560 28408 8566
rect 28356 8502 28408 8508
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 28264 8288 28316 8294
rect 28264 8230 28316 8236
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 25688 7948 25740 7954
rect 25688 7890 25740 7896
rect 26332 7948 26384 7954
rect 26332 7890 26384 7896
rect 27436 7948 27488 7954
rect 27436 7890 27488 7896
rect 23202 7375 23258 7384
rect 23848 7404 23900 7410
rect 22836 7346 22888 7352
rect 24136 7398 24532 7426
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 25700 7410 25728 7890
rect 27344 7812 27396 7818
rect 27344 7754 27396 7760
rect 27356 7546 27384 7754
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 25688 7404 25740 7410
rect 23848 7346 23900 7352
rect 25688 7346 25740 7352
rect 28276 7342 28304 8230
rect 28644 8090 28672 9454
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 29012 8974 29040 9318
rect 29104 8974 29132 9862
rect 29380 9654 29408 10202
rect 29368 9648 29420 9654
rect 29368 9590 29420 9596
rect 29276 9512 29328 9518
rect 29276 9454 29328 9460
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 29184 8968 29236 8974
rect 29184 8910 29236 8916
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28644 7546 28672 8026
rect 28920 7954 28948 8570
rect 29196 8430 29224 8910
rect 29288 8838 29316 9454
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29288 8430 29316 8774
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 28908 7948 28960 7954
rect 28908 7890 28960 7896
rect 29196 7546 29224 8366
rect 29380 7818 29408 9590
rect 29564 9518 29592 10746
rect 29748 10674 29776 14282
rect 29840 13326 29868 15558
rect 29920 15496 29972 15502
rect 29918 15464 29920 15473
rect 29972 15464 29974 15473
rect 29918 15399 29974 15408
rect 30024 15178 30052 17734
rect 30300 17678 30328 18022
rect 30840 17808 30892 17814
rect 30840 17750 30892 17756
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 30116 16266 30144 17614
rect 30852 17134 30880 17750
rect 30840 17128 30892 17134
rect 30840 17070 30892 17076
rect 30932 16584 30984 16590
rect 30930 16552 30932 16561
rect 30984 16552 30986 16561
rect 30930 16487 30986 16496
rect 30562 16280 30618 16289
rect 30116 16238 30236 16266
rect 30208 15706 30236 16238
rect 30562 16215 30618 16224
rect 30576 16114 30604 16215
rect 30288 16108 30340 16114
rect 30288 16050 30340 16056
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30300 16017 30328 16050
rect 30286 16008 30342 16017
rect 30286 15943 30342 15952
rect 30472 15904 30524 15910
rect 30472 15846 30524 15852
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30484 15502 30512 15846
rect 30472 15496 30524 15502
rect 30470 15464 30472 15473
rect 30524 15464 30526 15473
rect 30470 15399 30526 15408
rect 30196 15360 30248 15366
rect 30380 15360 30432 15366
rect 30248 15320 30380 15348
rect 30196 15302 30248 15308
rect 30380 15302 30432 15308
rect 30576 15201 30604 16050
rect 30656 15632 30708 15638
rect 30656 15574 30708 15580
rect 30668 15502 30696 15574
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 29932 15150 30052 15178
rect 30562 15192 30618 15201
rect 29932 14890 29960 15150
rect 30562 15127 30618 15136
rect 29920 14884 29972 14890
rect 29920 14826 29972 14832
rect 29932 14278 29960 14826
rect 30944 14346 30972 16487
rect 30932 14340 30984 14346
rect 30932 14282 30984 14288
rect 29920 14272 29972 14278
rect 29920 14214 29972 14220
rect 31036 14006 31064 18566
rect 31220 18426 31248 18634
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31496 18358 31524 19110
rect 31484 18352 31536 18358
rect 31484 18294 31536 18300
rect 31484 18216 31536 18222
rect 31404 18164 31484 18170
rect 31404 18158 31536 18164
rect 31404 18142 31524 18158
rect 31116 16448 31168 16454
rect 31116 16390 31168 16396
rect 31128 14346 31156 16390
rect 31404 16250 31432 18142
rect 31484 17060 31536 17066
rect 31484 17002 31536 17008
rect 31496 16522 31524 17002
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31392 16244 31444 16250
rect 31392 16186 31444 16192
rect 31208 16040 31260 16046
rect 31208 15982 31260 15988
rect 31220 15570 31248 15982
rect 31484 15904 31536 15910
rect 31484 15846 31536 15852
rect 31208 15564 31260 15570
rect 31208 15506 31260 15512
rect 31220 15094 31248 15506
rect 31496 15434 31524 15846
rect 31484 15428 31536 15434
rect 31484 15370 31536 15376
rect 31588 15314 31616 19230
rect 31680 18630 31708 19654
rect 31772 18986 31800 20742
rect 31944 20596 31996 20602
rect 31944 20538 31996 20544
rect 31956 19854 31984 20538
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31772 18958 31892 18986
rect 31668 18624 31720 18630
rect 31668 18566 31720 18572
rect 31680 18358 31708 18566
rect 31668 18352 31720 18358
rect 31668 18294 31720 18300
rect 31668 17672 31720 17678
rect 31668 17614 31720 17620
rect 31680 17134 31708 17614
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31760 17060 31812 17066
rect 31760 17002 31812 17008
rect 31772 16794 31800 17002
rect 31760 16788 31812 16794
rect 31760 16730 31812 16736
rect 31864 16658 31892 18958
rect 31944 18148 31996 18154
rect 31944 18090 31996 18096
rect 31956 17338 31984 18090
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 31852 16652 31904 16658
rect 31852 16594 31904 16600
rect 31668 16584 31720 16590
rect 31668 16526 31720 16532
rect 31680 16425 31708 16526
rect 31666 16416 31722 16425
rect 31666 16351 31722 16360
rect 31680 16250 31708 16351
rect 31668 16244 31720 16250
rect 31668 16186 31720 16192
rect 31496 15286 31616 15314
rect 31852 15360 31904 15366
rect 31852 15302 31904 15308
rect 31208 15088 31260 15094
rect 31208 15030 31260 15036
rect 31220 14482 31248 15030
rect 31208 14476 31260 14482
rect 31208 14418 31260 14424
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 31496 14006 31524 15286
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 31588 14074 31616 14962
rect 31576 14068 31628 14074
rect 31576 14010 31628 14016
rect 31024 14000 31076 14006
rect 31024 13942 31076 13948
rect 31484 14000 31536 14006
rect 31484 13942 31536 13948
rect 31036 13410 31064 13942
rect 30944 13382 31064 13410
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29840 12850 29868 13262
rect 30944 13258 30972 13382
rect 30932 13252 30984 13258
rect 30932 13194 30984 13200
rect 31024 13252 31076 13258
rect 31024 13194 31076 13200
rect 30564 13184 30616 13190
rect 30564 13126 30616 13132
rect 30576 12850 30604 13126
rect 31036 12986 31064 13194
rect 31024 12980 31076 12986
rect 31024 12922 31076 12928
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 30564 12844 30616 12850
rect 30564 12786 30616 12792
rect 31024 12844 31076 12850
rect 31024 12786 31076 12792
rect 30840 12776 30892 12782
rect 30840 12718 30892 12724
rect 30564 12640 30616 12646
rect 30564 12582 30616 12588
rect 30576 12306 30604 12582
rect 30564 12300 30616 12306
rect 30564 12242 30616 12248
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 29932 11830 29960 12106
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 29920 11824 29972 11830
rect 29920 11766 29972 11772
rect 30392 11218 30420 11834
rect 30852 11558 30880 12718
rect 31036 12434 31064 12786
rect 31496 12782 31524 13942
rect 31484 12776 31536 12782
rect 31484 12718 31536 12724
rect 31036 12406 31156 12434
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30380 11212 30432 11218
rect 30380 11154 30432 11160
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 30392 9382 30420 11154
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 30668 10266 30696 10610
rect 30656 10260 30708 10266
rect 30576 10220 30656 10248
rect 30472 9988 30524 9994
rect 30472 9930 30524 9936
rect 30484 9518 30512 9930
rect 30576 9722 30604 10220
rect 30656 10202 30708 10208
rect 31024 10260 31076 10266
rect 31024 10202 31076 10208
rect 31036 10062 31064 10202
rect 31024 10056 31076 10062
rect 31024 9998 31076 10004
rect 31128 9926 31156 12406
rect 31496 12306 31524 12718
rect 31760 12640 31812 12646
rect 31760 12582 31812 12588
rect 31484 12300 31536 12306
rect 31484 12242 31536 12248
rect 31772 12238 31800 12582
rect 31864 12442 31892 15302
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31956 12918 31984 13874
rect 31944 12912 31996 12918
rect 31944 12854 31996 12860
rect 31852 12436 31904 12442
rect 31852 12378 31904 12384
rect 32048 12238 32076 21542
rect 32128 21480 32180 21486
rect 32128 21422 32180 21428
rect 32140 20262 32168 21422
rect 32128 20256 32180 20262
rect 32128 20198 32180 20204
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32140 17814 32168 19314
rect 32220 18284 32272 18290
rect 32220 18226 32272 18232
rect 32232 17814 32260 18226
rect 32312 18148 32364 18154
rect 32312 18090 32364 18096
rect 32128 17808 32180 17814
rect 32128 17750 32180 17756
rect 32220 17808 32272 17814
rect 32220 17750 32272 17756
rect 32140 17202 32168 17750
rect 32220 17604 32272 17610
rect 32220 17546 32272 17552
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32140 16561 32168 16730
rect 32126 16552 32182 16561
rect 32126 16487 32182 16496
rect 32232 16114 32260 17546
rect 32324 17066 32352 18090
rect 32312 17060 32364 17066
rect 32312 17002 32364 17008
rect 32324 16794 32352 17002
rect 32312 16788 32364 16794
rect 32312 16730 32364 16736
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32220 16108 32272 16114
rect 32220 16050 32272 16056
rect 32232 15162 32260 16050
rect 32324 15978 32352 16594
rect 32312 15972 32364 15978
rect 32312 15914 32364 15920
rect 32220 15156 32272 15162
rect 32220 15098 32272 15104
rect 32232 14618 32260 15098
rect 32324 14618 32352 15914
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32416 14226 32444 23530
rect 32508 23118 32536 23666
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32588 21888 32640 21894
rect 32588 21830 32640 21836
rect 32600 21622 32628 21830
rect 32588 21616 32640 21622
rect 32588 21558 32640 21564
rect 32692 20602 32720 24686
rect 33060 24410 33088 24754
rect 33048 24404 33100 24410
rect 33048 24346 33100 24352
rect 32772 22976 32824 22982
rect 32772 22918 32824 22924
rect 32784 22574 32812 22918
rect 32772 22568 32824 22574
rect 32770 22536 32772 22545
rect 32824 22536 32826 22545
rect 32770 22471 32826 22480
rect 33152 22166 33180 28970
rect 33244 24750 33272 29106
rect 33324 28960 33376 28966
rect 33324 28902 33376 28908
rect 33336 28490 33364 28902
rect 33428 28529 33456 29566
rect 33520 28762 33548 32370
rect 33600 29640 33652 29646
rect 33600 29582 33652 29588
rect 33612 29510 33640 29582
rect 33600 29504 33652 29510
rect 33600 29446 33652 29452
rect 33508 28756 33560 28762
rect 33560 28716 33640 28744
rect 33508 28698 33560 28704
rect 33414 28520 33470 28529
rect 33324 28484 33376 28490
rect 33414 28455 33470 28464
rect 33324 28426 33376 28432
rect 33416 28416 33468 28422
rect 33336 28364 33416 28370
rect 33336 28358 33468 28364
rect 33336 28342 33456 28358
rect 33336 28082 33364 28342
rect 33324 28076 33376 28082
rect 33324 28018 33376 28024
rect 33508 28076 33560 28082
rect 33508 28018 33560 28024
rect 33336 26586 33364 28018
rect 33520 27402 33548 28018
rect 33612 27470 33640 28716
rect 33704 28257 33732 38150
rect 34244 37800 34296 37806
rect 34244 37742 34296 37748
rect 34256 37466 34284 37742
rect 34532 37738 34560 41550
rect 35452 41478 35480 41568
rect 35716 41550 35768 41556
rect 35900 41608 35952 41614
rect 36096 41596 36124 41958
rect 36360 41812 36412 41818
rect 36360 41754 36412 41760
rect 36268 41676 36320 41682
rect 36268 41618 36320 41624
rect 35952 41568 36124 41596
rect 35900 41550 35952 41556
rect 35072 41472 35124 41478
rect 35072 41414 35124 41420
rect 35440 41472 35492 41478
rect 35440 41414 35492 41420
rect 35084 41070 35112 41414
rect 35594 41372 35902 41381
rect 35594 41370 35600 41372
rect 35656 41370 35680 41372
rect 35736 41370 35760 41372
rect 35816 41370 35840 41372
rect 35896 41370 35902 41372
rect 35656 41318 35658 41370
rect 35838 41318 35840 41370
rect 35594 41316 35600 41318
rect 35656 41316 35680 41318
rect 35736 41316 35760 41318
rect 35816 41316 35840 41318
rect 35896 41316 35902 41318
rect 35594 41307 35902 41316
rect 34704 41064 34756 41070
rect 34704 41006 34756 41012
rect 35072 41064 35124 41070
rect 35072 41006 35124 41012
rect 34716 40526 34744 41006
rect 35348 40928 35400 40934
rect 35348 40870 35400 40876
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34796 40656 34848 40662
rect 35360 40610 35388 40870
rect 34796 40598 34848 40604
rect 34704 40520 34756 40526
rect 34704 40462 34756 40468
rect 34704 39976 34756 39982
rect 34704 39918 34756 39924
rect 34716 39642 34744 39918
rect 34704 39636 34756 39642
rect 34704 39578 34756 39584
rect 34808 39506 34836 40598
rect 35268 40582 35388 40610
rect 35268 40526 35296 40582
rect 35256 40520 35308 40526
rect 35256 40462 35308 40468
rect 35348 40520 35400 40526
rect 35348 40462 35400 40468
rect 35268 40032 35296 40462
rect 35360 40186 35388 40462
rect 35440 40452 35492 40458
rect 35440 40394 35492 40400
rect 35348 40180 35400 40186
rect 35348 40122 35400 40128
rect 35348 40044 35400 40050
rect 35268 40004 35348 40032
rect 35348 39986 35400 39992
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34796 39500 34848 39506
rect 34796 39442 34848 39448
rect 34612 39296 34664 39302
rect 34612 39238 34664 39244
rect 34520 37732 34572 37738
rect 34520 37674 34572 37680
rect 34244 37460 34296 37466
rect 34244 37402 34296 37408
rect 33968 37256 34020 37262
rect 33966 37224 33968 37233
rect 34152 37256 34204 37262
rect 34020 37224 34022 37233
rect 34152 37198 34204 37204
rect 33966 37159 34022 37168
rect 34164 36650 34192 37198
rect 34520 37188 34572 37194
rect 34520 37130 34572 37136
rect 34336 36780 34388 36786
rect 34336 36722 34388 36728
rect 34428 36780 34480 36786
rect 34428 36722 34480 36728
rect 34152 36644 34204 36650
rect 34152 36586 34204 36592
rect 34348 36582 34376 36722
rect 34336 36576 34388 36582
rect 34336 36518 34388 36524
rect 34348 36378 34376 36518
rect 34336 36372 34388 36378
rect 34336 36314 34388 36320
rect 34060 36100 34112 36106
rect 34060 36042 34112 36048
rect 33784 36032 33836 36038
rect 33784 35974 33836 35980
rect 33796 35630 33824 35974
rect 34072 35766 34100 36042
rect 34440 36038 34468 36722
rect 34532 36650 34560 37130
rect 34520 36644 34572 36650
rect 34520 36586 34572 36592
rect 34244 36032 34296 36038
rect 34244 35974 34296 35980
rect 34428 36032 34480 36038
rect 34428 35974 34480 35980
rect 34060 35760 34112 35766
rect 34060 35702 34112 35708
rect 33876 35692 33928 35698
rect 33876 35634 33928 35640
rect 33784 35624 33836 35630
rect 33784 35566 33836 35572
rect 33888 35494 33916 35634
rect 33876 35488 33928 35494
rect 33876 35430 33928 35436
rect 33888 34542 33916 35430
rect 33876 34536 33928 34542
rect 33876 34478 33928 34484
rect 34256 34202 34284 35974
rect 34440 35834 34468 35974
rect 34428 35828 34480 35834
rect 34428 35770 34480 35776
rect 34244 34196 34296 34202
rect 34244 34138 34296 34144
rect 33784 33992 33836 33998
rect 33784 33934 33836 33940
rect 33796 33522 33824 33934
rect 33968 33924 34020 33930
rect 33968 33866 34020 33872
rect 33784 33516 33836 33522
rect 33784 33458 33836 33464
rect 33796 31958 33824 33458
rect 33980 33454 34008 33866
rect 34060 33856 34112 33862
rect 34060 33798 34112 33804
rect 34072 33522 34100 33798
rect 34060 33516 34112 33522
rect 34060 33458 34112 33464
rect 33968 33448 34020 33454
rect 33968 33390 34020 33396
rect 34072 32774 34100 33458
rect 34060 32768 34112 32774
rect 34060 32710 34112 32716
rect 34072 32434 34100 32710
rect 34624 32552 34652 39238
rect 35360 39098 35388 39986
rect 35452 39982 35480 40394
rect 35992 40384 36044 40390
rect 35992 40326 36044 40332
rect 35594 40284 35902 40293
rect 35594 40282 35600 40284
rect 35656 40282 35680 40284
rect 35736 40282 35760 40284
rect 35816 40282 35840 40284
rect 35896 40282 35902 40284
rect 35656 40230 35658 40282
rect 35838 40230 35840 40282
rect 35594 40228 35600 40230
rect 35656 40228 35680 40230
rect 35736 40228 35760 40230
rect 35816 40228 35840 40230
rect 35896 40228 35902 40230
rect 35594 40219 35902 40228
rect 36004 40050 36032 40326
rect 35992 40044 36044 40050
rect 35992 39986 36044 39992
rect 36096 39982 36124 41568
rect 36176 41200 36228 41206
rect 36176 41142 36228 41148
rect 36188 40118 36216 41142
rect 36280 41138 36308 41618
rect 36268 41132 36320 41138
rect 36268 41074 36320 41080
rect 36372 41070 36400 41754
rect 36360 41064 36412 41070
rect 36360 41006 36412 41012
rect 36464 40882 36492 42162
rect 36544 42152 36596 42158
rect 36544 42094 36596 42100
rect 36636 42152 36688 42158
rect 36636 42094 36688 42100
rect 36556 41002 36584 42094
rect 36648 41818 36676 42094
rect 36636 41812 36688 41818
rect 36636 41754 36688 41760
rect 36832 41698 36860 42230
rect 37016 42090 37044 42502
rect 37292 42226 37320 42706
rect 37280 42220 37332 42226
rect 37280 42162 37332 42168
rect 37004 42084 37056 42090
rect 37004 42026 37056 42032
rect 36740 41670 36860 41698
rect 36740 41206 36768 41670
rect 36820 41608 36872 41614
rect 36820 41550 36872 41556
rect 36912 41608 36964 41614
rect 36912 41550 36964 41556
rect 36832 41478 36860 41550
rect 36820 41472 36872 41478
rect 36820 41414 36872 41420
rect 36728 41200 36780 41206
rect 36728 41142 36780 41148
rect 36544 40996 36596 41002
rect 36544 40938 36596 40944
rect 36832 40934 36860 41414
rect 36924 41070 36952 41550
rect 36912 41064 36964 41070
rect 36912 41006 36964 41012
rect 36820 40928 36872 40934
rect 36464 40854 36676 40882
rect 37016 40882 37044 42026
rect 37292 41138 37320 42162
rect 37188 41132 37240 41138
rect 37188 41074 37240 41080
rect 37280 41132 37332 41138
rect 37280 41074 37332 41080
rect 38200 41132 38252 41138
rect 38200 41074 38252 41080
rect 36820 40870 36872 40876
rect 36176 40112 36228 40118
rect 36176 40054 36228 40060
rect 35440 39976 35492 39982
rect 35440 39918 35492 39924
rect 36084 39976 36136 39982
rect 36084 39918 36136 39924
rect 35348 39092 35400 39098
rect 35348 39034 35400 39040
rect 35348 38956 35400 38962
rect 35348 38898 35400 38904
rect 35360 38758 35388 38898
rect 35452 38842 35480 39918
rect 35992 39908 36044 39914
rect 35992 39850 36044 39856
rect 35532 39840 35584 39846
rect 35532 39782 35584 39788
rect 35624 39840 35676 39846
rect 35624 39782 35676 39788
rect 35716 39840 35768 39846
rect 35716 39782 35768 39788
rect 35544 39370 35572 39782
rect 35636 39438 35664 39782
rect 35728 39545 35756 39782
rect 36004 39642 36032 39850
rect 36096 39642 36124 39918
rect 35992 39636 36044 39642
rect 35992 39578 36044 39584
rect 36084 39636 36136 39642
rect 36084 39578 36136 39584
rect 35714 39536 35770 39545
rect 35714 39471 35770 39480
rect 36084 39500 36136 39506
rect 36084 39442 36136 39448
rect 35624 39432 35676 39438
rect 35624 39374 35676 39380
rect 35992 39432 36044 39438
rect 35992 39374 36044 39380
rect 35532 39364 35584 39370
rect 35532 39306 35584 39312
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 36004 39098 36032 39374
rect 35808 39092 35860 39098
rect 35808 39034 35860 39040
rect 35992 39092 36044 39098
rect 35992 39034 36044 39040
rect 35530 38856 35586 38865
rect 35452 38814 35530 38842
rect 35530 38791 35532 38800
rect 35584 38791 35586 38800
rect 35532 38762 35584 38768
rect 35348 38752 35400 38758
rect 35348 38694 35400 38700
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34796 38412 34848 38418
rect 34796 38354 34848 38360
rect 34704 38208 34756 38214
rect 34704 38150 34756 38156
rect 34716 38010 34744 38150
rect 34808 38010 34836 38354
rect 34704 38004 34756 38010
rect 34704 37946 34756 37952
rect 34796 38004 34848 38010
rect 34796 37946 34848 37952
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35360 37482 35388 38694
rect 35820 38350 35848 39034
rect 35992 38956 36044 38962
rect 36096 38944 36124 39442
rect 36188 39438 36216 40054
rect 36176 39432 36228 39438
rect 36176 39374 36228 39380
rect 36176 39296 36228 39302
rect 36176 39238 36228 39244
rect 36188 39098 36216 39238
rect 36176 39092 36228 39098
rect 36176 39034 36228 39040
rect 36044 38916 36124 38944
rect 35992 38898 36044 38904
rect 35900 38888 35952 38894
rect 35900 38830 35952 38836
rect 35912 38758 35940 38830
rect 35900 38752 35952 38758
rect 35900 38694 35952 38700
rect 35808 38344 35860 38350
rect 35808 38286 35860 38292
rect 35440 38208 35492 38214
rect 35440 38150 35492 38156
rect 35452 37942 35480 38150
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 36004 38010 36032 38898
rect 36082 38856 36138 38865
rect 36082 38791 36138 38800
rect 36096 38758 36124 38791
rect 36084 38752 36136 38758
rect 36084 38694 36136 38700
rect 35992 38004 36044 38010
rect 35992 37946 36044 37952
rect 35440 37936 35492 37942
rect 35440 37878 35492 37884
rect 35440 37800 35492 37806
rect 35440 37742 35492 37748
rect 36452 37800 36504 37806
rect 36452 37742 36504 37748
rect 35268 37454 35388 37482
rect 35268 37262 35296 37454
rect 35348 37392 35400 37398
rect 35348 37334 35400 37340
rect 35360 37262 35388 37334
rect 35452 37262 35480 37742
rect 36464 37466 36492 37742
rect 36452 37460 36504 37466
rect 36452 37402 36504 37408
rect 35256 37256 35308 37262
rect 35256 37198 35308 37204
rect 35348 37256 35400 37262
rect 35348 37198 35400 37204
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 35992 37188 36044 37194
rect 35992 37130 36044 37136
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 35716 36780 35768 36786
rect 35716 36722 35768 36728
rect 35624 36576 35676 36582
rect 35624 36518 35676 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35440 36168 35492 36174
rect 35440 36110 35492 36116
rect 35452 35630 35480 36110
rect 35636 36106 35664 36518
rect 35728 36242 35756 36722
rect 36004 36650 36032 37130
rect 36268 37120 36320 37126
rect 36268 37062 36320 37068
rect 36280 36786 36308 37062
rect 36268 36780 36320 36786
rect 36268 36722 36320 36728
rect 36544 36780 36596 36786
rect 36544 36722 36596 36728
rect 36280 36666 36308 36722
rect 35992 36644 36044 36650
rect 36280 36638 36492 36666
rect 36556 36650 36584 36722
rect 35992 36586 36044 36592
rect 36464 36242 36492 36638
rect 36544 36644 36596 36650
rect 36544 36586 36596 36592
rect 35716 36236 35768 36242
rect 35716 36178 35768 36184
rect 36452 36236 36504 36242
rect 36452 36178 36504 36184
rect 35624 36100 35676 36106
rect 35624 36042 35676 36048
rect 36452 36100 36504 36106
rect 36452 36042 36504 36048
rect 36084 36032 36136 36038
rect 36084 35974 36136 35980
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 36096 35630 36124 35974
rect 34704 35624 34756 35630
rect 34704 35566 34756 35572
rect 35440 35624 35492 35630
rect 35440 35566 35492 35572
rect 35992 35624 36044 35630
rect 35992 35566 36044 35572
rect 36084 35624 36136 35630
rect 36084 35566 36136 35572
rect 34716 34746 34744 35566
rect 35532 35488 35584 35494
rect 35532 35430 35584 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 35148 34848 35154
rect 34796 35090 34848 35096
rect 34704 34740 34756 34746
rect 34704 34682 34756 34688
rect 34808 34610 34836 35090
rect 35544 35018 35572 35430
rect 35532 35012 35584 35018
rect 35532 34954 35584 34960
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34796 34604 34848 34610
rect 34796 34546 34848 34552
rect 34796 34400 34848 34406
rect 34796 34342 34848 34348
rect 34808 34202 34836 34342
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 36004 34202 36032 35566
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 35992 34196 36044 34202
rect 35992 34138 36044 34144
rect 36096 34066 36124 35566
rect 36360 35488 36412 35494
rect 36360 35430 36412 35436
rect 36372 35086 36400 35430
rect 36464 35222 36492 36042
rect 36544 36032 36596 36038
rect 36544 35974 36596 35980
rect 36556 35630 36584 35974
rect 36544 35624 36596 35630
rect 36544 35566 36596 35572
rect 36452 35216 36504 35222
rect 36452 35158 36504 35164
rect 36360 35080 36412 35086
rect 36360 35022 36412 35028
rect 36372 34678 36400 35022
rect 36360 34672 36412 34678
rect 36360 34614 36412 34620
rect 36464 34542 36492 35158
rect 36452 34536 36504 34542
rect 36452 34478 36504 34484
rect 36084 34060 36136 34066
rect 36084 34002 36136 34008
rect 36176 33856 36228 33862
rect 36176 33798 36228 33804
rect 36452 33856 36504 33862
rect 36452 33798 36504 33804
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 36188 33658 36216 33798
rect 36176 33652 36228 33658
rect 36176 33594 36228 33600
rect 36464 33454 36492 33798
rect 36544 33584 36596 33590
rect 36544 33526 36596 33532
rect 35808 33448 35860 33454
rect 35808 33390 35860 33396
rect 36452 33448 36504 33454
rect 36452 33390 36504 33396
rect 35440 33312 35492 33318
rect 35440 33254 35492 33260
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35072 32904 35124 32910
rect 35072 32846 35124 32852
rect 34624 32524 34836 32552
rect 34060 32428 34112 32434
rect 34060 32370 34112 32376
rect 34704 32428 34756 32434
rect 34704 32370 34756 32376
rect 34244 32360 34296 32366
rect 34244 32302 34296 32308
rect 34256 31958 34284 32302
rect 33784 31952 33836 31958
rect 33784 31894 33836 31900
rect 34244 31952 34296 31958
rect 34244 31894 34296 31900
rect 34152 31340 34204 31346
rect 34152 31282 34204 31288
rect 33784 30660 33836 30666
rect 33784 30602 33836 30608
rect 33796 29102 33824 30602
rect 34060 30320 34112 30326
rect 34060 30262 34112 30268
rect 33876 30048 33928 30054
rect 33876 29990 33928 29996
rect 33888 29170 33916 29990
rect 33966 29608 34022 29617
rect 33966 29543 34022 29552
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33784 29096 33836 29102
rect 33784 29038 33836 29044
rect 33980 29034 34008 29543
rect 34072 29209 34100 30262
rect 34164 30190 34192 31282
rect 34256 31278 34284 31894
rect 34520 31680 34572 31686
rect 34520 31622 34572 31628
rect 34532 31482 34560 31622
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 34244 31272 34296 31278
rect 34244 31214 34296 31220
rect 34520 31272 34572 31278
rect 34520 31214 34572 31220
rect 34336 31204 34388 31210
rect 34336 31146 34388 31152
rect 34348 30666 34376 31146
rect 34336 30660 34388 30666
rect 34336 30602 34388 30608
rect 34152 30184 34204 30190
rect 34152 30126 34204 30132
rect 34336 30184 34388 30190
rect 34336 30126 34388 30132
rect 34426 30152 34482 30161
rect 34244 30116 34296 30122
rect 34244 30058 34296 30064
rect 34152 29572 34204 29578
rect 34152 29514 34204 29520
rect 34164 29306 34192 29514
rect 34152 29300 34204 29306
rect 34152 29242 34204 29248
rect 34058 29200 34114 29209
rect 34058 29135 34114 29144
rect 34152 29164 34204 29170
rect 34152 29106 34204 29112
rect 33968 29028 34020 29034
rect 33968 28970 34020 28976
rect 33874 28928 33930 28937
rect 33874 28863 33930 28872
rect 33690 28248 33746 28257
rect 33690 28183 33746 28192
rect 33704 28064 33732 28183
rect 33784 28076 33836 28082
rect 33704 28036 33784 28064
rect 33784 28018 33836 28024
rect 33888 27538 33916 28863
rect 34058 28520 34114 28529
rect 34058 28455 34060 28464
rect 34112 28455 34114 28464
rect 34060 28426 34112 28432
rect 33968 28076 34020 28082
rect 33968 28018 34020 28024
rect 33980 27674 34008 28018
rect 33968 27668 34020 27674
rect 33968 27610 34020 27616
rect 33876 27532 33928 27538
rect 33876 27474 33928 27480
rect 33600 27464 33652 27470
rect 33600 27406 33652 27412
rect 34072 27418 34100 28426
rect 34164 27946 34192 29106
rect 34256 29034 34284 30058
rect 34348 29170 34376 30126
rect 34426 30087 34428 30096
rect 34480 30087 34482 30096
rect 34428 30058 34480 30064
rect 34440 29889 34468 30058
rect 34426 29880 34482 29889
rect 34426 29815 34482 29824
rect 34532 29730 34560 31214
rect 34624 29850 34652 31282
rect 34716 30802 34744 32370
rect 34808 31278 34836 32524
rect 35084 32434 35112 32846
rect 35348 32836 35400 32842
rect 35348 32778 35400 32784
rect 35072 32428 35124 32434
rect 35072 32370 35124 32376
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35360 32026 35388 32778
rect 35452 32502 35480 33254
rect 35820 32756 35848 33390
rect 35820 32728 36032 32756
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 36004 32552 36032 32728
rect 36464 32570 36492 33390
rect 35820 32524 36032 32552
rect 36452 32564 36504 32570
rect 35440 32496 35492 32502
rect 35440 32438 35492 32444
rect 35348 32020 35400 32026
rect 35348 31962 35400 31968
rect 35820 31890 35848 32524
rect 36452 32506 36504 32512
rect 35808 31884 35860 31890
rect 35808 31826 35860 31832
rect 36556 31754 36584 33526
rect 36464 31726 36584 31754
rect 35992 31680 36044 31686
rect 35992 31622 36044 31628
rect 36084 31680 36136 31686
rect 36084 31622 36136 31628
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 35348 31408 35400 31414
rect 35348 31350 35400 31356
rect 34796 31272 34848 31278
rect 34796 31214 34848 31220
rect 34796 31136 34848 31142
rect 34796 31078 34848 31084
rect 34808 30938 34836 31078
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30932 34848 30938
rect 34796 30874 34848 30880
rect 34704 30796 34756 30802
rect 34704 30738 34756 30744
rect 34796 30388 34848 30394
rect 34796 30330 34848 30336
rect 34808 30190 34836 30330
rect 34796 30184 34848 30190
rect 34796 30126 34848 30132
rect 34888 30184 34940 30190
rect 34888 30126 34940 30132
rect 35162 30152 35218 30161
rect 34900 30036 34928 30126
rect 35162 30087 35164 30096
rect 35216 30087 35218 30096
rect 35164 30058 35216 30064
rect 34808 30008 34928 30036
rect 34612 29844 34664 29850
rect 34808 29832 34836 30008
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34980 29844 35032 29850
rect 34808 29804 34928 29832
rect 34612 29786 34664 29792
rect 34532 29702 34836 29730
rect 34900 29714 34928 29804
rect 34980 29786 35032 29792
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34428 29300 34480 29306
rect 34428 29242 34480 29248
rect 34336 29164 34388 29170
rect 34336 29106 34388 29112
rect 34244 29028 34296 29034
rect 34244 28970 34296 28976
rect 34440 28966 34468 29242
rect 34612 29232 34664 29238
rect 34610 29200 34612 29209
rect 34664 29200 34666 29209
rect 34520 29164 34572 29170
rect 34610 29135 34666 29144
rect 34520 29106 34572 29112
rect 34428 28960 34480 28966
rect 34428 28902 34480 28908
rect 34440 28150 34468 28902
rect 34532 28762 34560 29106
rect 34716 28762 34744 29582
rect 34520 28756 34572 28762
rect 34704 28756 34756 28762
rect 34572 28716 34652 28744
rect 34520 28698 34572 28704
rect 34520 28212 34572 28218
rect 34520 28154 34572 28160
rect 34428 28144 34480 28150
rect 34334 28112 34390 28121
rect 34428 28086 34480 28092
rect 34334 28047 34336 28056
rect 34388 28047 34390 28056
rect 34336 28018 34388 28024
rect 34152 27940 34204 27946
rect 34152 27882 34204 27888
rect 34428 27532 34480 27538
rect 34428 27474 34480 27480
rect 33508 27396 33560 27402
rect 33508 27338 33560 27344
rect 33324 26580 33376 26586
rect 33324 26522 33376 26528
rect 33612 26382 33640 27406
rect 33968 27396 34020 27402
rect 34072 27390 34192 27418
rect 33968 27338 34020 27344
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33416 26240 33468 26246
rect 33416 26182 33468 26188
rect 33428 25498 33456 26182
rect 33612 25922 33640 26318
rect 33612 25894 33732 25922
rect 33704 25838 33732 25894
rect 33692 25832 33744 25838
rect 33692 25774 33744 25780
rect 33416 25492 33468 25498
rect 33416 25434 33468 25440
rect 33416 25288 33468 25294
rect 33416 25230 33468 25236
rect 33428 24886 33456 25230
rect 33704 24886 33732 25774
rect 33980 25294 34008 27338
rect 34060 27328 34112 27334
rect 34060 27270 34112 27276
rect 33784 25288 33836 25294
rect 33784 25230 33836 25236
rect 33876 25288 33928 25294
rect 33876 25230 33928 25236
rect 33968 25288 34020 25294
rect 33968 25230 34020 25236
rect 33416 24880 33468 24886
rect 33416 24822 33468 24828
rect 33692 24880 33744 24886
rect 33692 24822 33744 24828
rect 33428 24750 33456 24822
rect 33232 24744 33284 24750
rect 33232 24686 33284 24692
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 33796 24614 33824 25230
rect 33888 24954 33916 25230
rect 33876 24948 33928 24954
rect 33876 24890 33928 24896
rect 33784 24608 33836 24614
rect 33784 24550 33836 24556
rect 33796 24274 33824 24550
rect 33784 24268 33836 24274
rect 33784 24210 33836 24216
rect 33784 23792 33836 23798
rect 33784 23734 33836 23740
rect 33324 23520 33376 23526
rect 33324 23462 33376 23468
rect 33336 23050 33364 23462
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 33232 21888 33284 21894
rect 33232 21830 33284 21836
rect 32680 20596 32732 20602
rect 32680 20538 32732 20544
rect 32588 20392 32640 20398
rect 32588 20334 32640 20340
rect 32600 20058 32628 20334
rect 32772 20256 32824 20262
rect 32772 20198 32824 20204
rect 32588 20052 32640 20058
rect 32588 19994 32640 20000
rect 32784 19360 32812 20198
rect 33244 19922 33272 21830
rect 33520 21690 33548 21966
rect 33600 21888 33652 21894
rect 33600 21830 33652 21836
rect 33508 21684 33560 21690
rect 33508 21626 33560 21632
rect 33612 21078 33640 21830
rect 33796 21622 33824 23734
rect 33876 22092 33928 22098
rect 33876 22034 33928 22040
rect 33888 21690 33916 22034
rect 33876 21684 33928 21690
rect 33876 21626 33928 21632
rect 33784 21616 33836 21622
rect 33704 21576 33784 21604
rect 33600 21072 33652 21078
rect 33600 21014 33652 21020
rect 33612 20890 33640 21014
rect 33520 20862 33640 20890
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 33232 19916 33284 19922
rect 33232 19858 33284 19864
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 32864 19372 32916 19378
rect 32784 19332 32864 19360
rect 32680 19236 32732 19242
rect 32680 19178 32732 19184
rect 32496 18624 32548 18630
rect 32496 18566 32548 18572
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32508 18290 32536 18566
rect 32600 18358 32628 18566
rect 32588 18352 32640 18358
rect 32588 18294 32640 18300
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32496 17808 32548 17814
rect 32496 17750 32548 17756
rect 32508 16017 32536 17750
rect 32588 17740 32640 17746
rect 32588 17682 32640 17688
rect 32600 16998 32628 17682
rect 32692 17338 32720 19178
rect 32784 18834 32812 19332
rect 32864 19314 32916 19320
rect 32772 18828 32824 18834
rect 32772 18770 32824 18776
rect 32784 18222 32812 18770
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32784 17610 32812 18158
rect 32772 17604 32824 17610
rect 32772 17546 32824 17552
rect 32680 17332 32732 17338
rect 32680 17274 32732 17280
rect 32588 16992 32640 16998
rect 32588 16934 32640 16940
rect 32680 16516 32732 16522
rect 32680 16458 32732 16464
rect 32588 16176 32640 16182
rect 32588 16118 32640 16124
rect 32494 16008 32550 16017
rect 32494 15943 32550 15952
rect 32600 15706 32628 16118
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32692 15638 32720 16458
rect 32784 16046 32812 17546
rect 33060 17542 33088 19450
rect 33428 19378 33456 20538
rect 33520 19922 33548 20862
rect 33600 20800 33652 20806
rect 33600 20742 33652 20748
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33612 19854 33640 20742
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 33704 19514 33732 21576
rect 33784 21558 33836 21564
rect 33784 20936 33836 20942
rect 33784 20878 33836 20884
rect 33796 19922 33824 20878
rect 33888 20466 33916 21626
rect 33876 20460 33928 20466
rect 33876 20402 33928 20408
rect 33784 19916 33836 19922
rect 33784 19858 33836 19864
rect 33692 19508 33744 19514
rect 33692 19450 33744 19456
rect 33416 19372 33468 19378
rect 33416 19314 33468 19320
rect 33140 18080 33192 18086
rect 33140 18022 33192 18028
rect 33048 17536 33100 17542
rect 33048 17478 33100 17484
rect 33060 17202 33088 17478
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 33152 16658 33180 18022
rect 33428 17678 33456 19314
rect 33692 19304 33744 19310
rect 33692 19246 33744 19252
rect 33508 19236 33560 19242
rect 33508 19178 33560 19184
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33428 17202 33456 17614
rect 33416 17196 33468 17202
rect 33416 17138 33468 17144
rect 33232 17128 33284 17134
rect 33232 17070 33284 17076
rect 33244 16794 33272 17070
rect 33232 16788 33284 16794
rect 33232 16730 33284 16736
rect 33140 16652 33192 16658
rect 33140 16594 33192 16600
rect 32956 16516 33008 16522
rect 32956 16458 33008 16464
rect 32772 16040 32824 16046
rect 32772 15982 32824 15988
rect 32680 15632 32732 15638
rect 32680 15574 32732 15580
rect 32496 15428 32548 15434
rect 32496 15370 32548 15376
rect 32508 14414 32536 15370
rect 32968 15366 32996 16458
rect 33152 16289 33180 16594
rect 33232 16448 33284 16454
rect 33324 16448 33376 16454
rect 33232 16390 33284 16396
rect 33322 16416 33324 16425
rect 33376 16416 33378 16425
rect 33138 16280 33194 16289
rect 33138 16215 33194 16224
rect 32956 15360 33008 15366
rect 32956 15302 33008 15308
rect 33152 14958 33180 16215
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 33140 14952 33192 14958
rect 33140 14894 33192 14900
rect 32784 14618 32812 14894
rect 32772 14612 32824 14618
rect 32772 14554 32824 14560
rect 33244 14482 33272 16390
rect 33322 16351 33378 16360
rect 33324 16176 33376 16182
rect 33324 16118 33376 16124
rect 33336 15892 33364 16118
rect 33416 15904 33468 15910
rect 33336 15864 33416 15892
rect 33336 15434 33364 15864
rect 33416 15846 33468 15852
rect 33416 15564 33468 15570
rect 33416 15506 33468 15512
rect 33324 15428 33376 15434
rect 33324 15370 33376 15376
rect 33428 14890 33456 15506
rect 33416 14884 33468 14890
rect 33416 14826 33468 14832
rect 33428 14482 33456 14826
rect 33232 14476 33284 14482
rect 33232 14418 33284 14424
rect 33416 14476 33468 14482
rect 33416 14418 33468 14424
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 33416 14340 33468 14346
rect 33416 14282 33468 14288
rect 32416 14198 32536 14226
rect 32312 13864 32364 13870
rect 32312 13806 32364 13812
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32128 13320 32180 13326
rect 32128 13262 32180 13268
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 32036 12232 32088 12238
rect 32036 12174 32088 12180
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11830 31432 12038
rect 31392 11824 31444 11830
rect 31392 11766 31444 11772
rect 31852 11756 31904 11762
rect 31852 11698 31904 11704
rect 31576 11688 31628 11694
rect 31576 11630 31628 11636
rect 31300 11552 31352 11558
rect 31300 11494 31352 11500
rect 31312 11150 31340 11494
rect 31300 11144 31352 11150
rect 31300 11086 31352 11092
rect 31484 10192 31536 10198
rect 31484 10134 31536 10140
rect 31208 9988 31260 9994
rect 31208 9930 31260 9936
rect 31116 9920 31168 9926
rect 31116 9862 31168 9868
rect 30564 9716 30616 9722
rect 30564 9658 30616 9664
rect 30748 9648 30800 9654
rect 30748 9590 30800 9596
rect 30472 9512 30524 9518
rect 30472 9454 30524 9460
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 29460 8832 29512 8838
rect 29460 8774 29512 8780
rect 29472 8498 29500 8774
rect 30392 8634 30420 9318
rect 30484 9110 30512 9454
rect 30472 9104 30524 9110
rect 30472 9046 30524 9052
rect 30760 9042 30788 9590
rect 31220 9518 31248 9930
rect 31496 9586 31524 10134
rect 31588 9654 31616 11630
rect 31760 11144 31812 11150
rect 31864 11132 31892 11698
rect 31812 11104 31892 11132
rect 31760 11086 31812 11092
rect 31668 10056 31720 10062
rect 31668 9998 31720 10004
rect 31760 10056 31812 10062
rect 31760 9998 31812 10004
rect 31680 9654 31708 9998
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 31208 9512 31260 9518
rect 31208 9454 31260 9460
rect 31300 9512 31352 9518
rect 31300 9454 31352 9460
rect 30748 9036 30800 9042
rect 30748 8978 30800 8984
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30760 8566 30788 8978
rect 30748 8560 30800 8566
rect 30748 8502 30800 8508
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29564 7954 29592 8434
rect 30472 8424 30524 8430
rect 30472 8366 30524 8372
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 29840 7954 29868 8230
rect 30484 8090 30512 8366
rect 30564 8288 30616 8294
rect 30564 8230 30616 8236
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30576 7954 30604 8230
rect 31220 8022 31248 9454
rect 31312 9382 31340 9454
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 31680 8838 31708 9590
rect 31772 9178 31800 9998
rect 31864 9382 31892 11104
rect 32140 10810 32168 13262
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 32232 11150 32260 11494
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 31944 9920 31996 9926
rect 31944 9862 31996 9868
rect 31956 9654 31984 9862
rect 31944 9648 31996 9654
rect 31944 9590 31996 9596
rect 31852 9376 31904 9382
rect 31852 9318 31904 9324
rect 31760 9172 31812 9178
rect 31760 9114 31812 9120
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31208 8016 31260 8022
rect 31208 7958 31260 7964
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29828 7948 29880 7954
rect 29828 7890 29880 7896
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 29368 7812 29420 7818
rect 29368 7754 29420 7760
rect 28632 7540 28684 7546
rect 28632 7482 28684 7488
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 29380 7410 29408 7754
rect 31588 7750 31616 8434
rect 31864 7954 31892 9318
rect 32140 8974 32168 10746
rect 32324 9926 32352 13806
rect 32416 13394 32444 13806
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 32416 11830 32444 13330
rect 32508 12850 32536 14198
rect 33428 14074 33456 14282
rect 33520 14074 33548 19178
rect 33704 18766 33732 19246
rect 33692 18760 33744 18766
rect 33692 18702 33744 18708
rect 33704 18086 33732 18702
rect 33692 18080 33744 18086
rect 33692 18022 33744 18028
rect 33704 17678 33732 18022
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 33704 17270 33732 17614
rect 33692 17264 33744 17270
rect 33692 17206 33744 17212
rect 33980 16250 34008 25230
rect 34072 22094 34100 27270
rect 34164 25974 34192 27390
rect 34440 26926 34468 27474
rect 34428 26920 34480 26926
rect 34428 26862 34480 26868
rect 34152 25968 34204 25974
rect 34152 25910 34204 25916
rect 34152 25832 34204 25838
rect 34152 25774 34204 25780
rect 34164 24818 34192 25774
rect 34532 25294 34560 28154
rect 34624 27470 34652 28716
rect 34704 28698 34756 28704
rect 34808 28694 34836 29702
rect 34888 29708 34940 29714
rect 34888 29650 34940 29656
rect 34888 29572 34940 29578
rect 34888 29514 34940 29520
rect 34900 29306 34928 29514
rect 34992 29345 35020 29786
rect 35360 29782 35388 31350
rect 36004 31346 36032 31622
rect 35992 31340 36044 31346
rect 35992 31282 36044 31288
rect 36004 30938 36032 31282
rect 35992 30932 36044 30938
rect 35992 30874 36044 30880
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 36004 30326 36032 30874
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 35624 30252 35676 30258
rect 35624 30194 35676 30200
rect 35532 30184 35584 30190
rect 35532 30126 35584 30132
rect 35544 29850 35572 30126
rect 35532 29844 35584 29850
rect 35532 29786 35584 29792
rect 35348 29776 35400 29782
rect 35070 29744 35126 29753
rect 35348 29718 35400 29724
rect 35070 29679 35126 29688
rect 35084 29646 35112 29679
rect 35072 29640 35124 29646
rect 35072 29582 35124 29588
rect 34978 29336 35034 29345
rect 34888 29300 34940 29306
rect 34978 29271 35034 29280
rect 34888 29242 34940 29248
rect 34992 29102 35020 29271
rect 35084 29170 35112 29582
rect 35072 29164 35124 29170
rect 35072 29106 35124 29112
rect 34980 29096 35032 29102
rect 34980 29038 35032 29044
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28688 34848 28694
rect 34796 28630 34848 28636
rect 35256 28620 35308 28626
rect 35256 28562 35308 28568
rect 35070 28520 35126 28529
rect 35070 28455 35072 28464
rect 35124 28455 35126 28464
rect 35164 28484 35216 28490
rect 35072 28426 35124 28432
rect 35164 28426 35216 28432
rect 34796 28212 34848 28218
rect 34796 28154 34848 28160
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 34716 27470 34744 27814
rect 34808 27674 34836 28154
rect 35176 28014 35204 28426
rect 35268 28082 35296 28562
rect 35360 28218 35388 29718
rect 35544 29714 35572 29786
rect 35636 29753 35664 30194
rect 35900 30184 35952 30190
rect 35900 30126 35952 30132
rect 35622 29744 35678 29753
rect 35532 29708 35584 29714
rect 35622 29679 35678 29688
rect 35532 29650 35584 29656
rect 35808 29640 35860 29646
rect 35912 29628 35940 30126
rect 36004 29714 36032 30262
rect 36096 30190 36124 31622
rect 36268 31272 36320 31278
rect 36268 31214 36320 31220
rect 36176 30796 36228 30802
rect 36176 30738 36228 30744
rect 36188 30190 36216 30738
rect 36280 30394 36308 31214
rect 36360 30796 36412 30802
rect 36360 30738 36412 30744
rect 36268 30388 36320 30394
rect 36268 30330 36320 30336
rect 36372 30258 36400 30738
rect 36360 30252 36412 30258
rect 36360 30194 36412 30200
rect 36084 30184 36136 30190
rect 36084 30126 36136 30132
rect 36176 30184 36228 30190
rect 36176 30126 36228 30132
rect 35992 29708 36044 29714
rect 35992 29650 36044 29656
rect 35860 29600 35940 29628
rect 35808 29582 35860 29588
rect 36004 29578 36032 29650
rect 35992 29572 36044 29578
rect 35992 29514 36044 29520
rect 35440 29504 35492 29510
rect 35440 29446 35492 29452
rect 35452 29170 35480 29446
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 36004 29238 36032 29514
rect 35992 29232 36044 29238
rect 35992 29174 36044 29180
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35716 28960 35768 28966
rect 35716 28902 35768 28908
rect 35440 28756 35492 28762
rect 35440 28698 35492 28704
rect 35452 28558 35480 28698
rect 35532 28688 35584 28694
rect 35532 28630 35584 28636
rect 35440 28552 35492 28558
rect 35440 28494 35492 28500
rect 35544 28506 35572 28630
rect 35728 28558 35756 28902
rect 35716 28552 35768 28558
rect 35544 28478 35664 28506
rect 35716 28494 35768 28500
rect 35808 28552 35860 28558
rect 35808 28494 35860 28500
rect 35440 28416 35492 28422
rect 35636 28404 35664 28478
rect 35820 28404 35848 28494
rect 35636 28376 35848 28404
rect 35992 28416 36044 28422
rect 35440 28358 35492 28364
rect 35992 28358 36044 28364
rect 35348 28212 35400 28218
rect 35348 28154 35400 28160
rect 35256 28076 35308 28082
rect 35256 28018 35308 28024
rect 35164 28008 35216 28014
rect 35164 27950 35216 27956
rect 35268 27826 35296 28018
rect 35268 27798 35388 27826
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27668 34848 27674
rect 34796 27610 34848 27616
rect 35072 27600 35124 27606
rect 35256 27600 35308 27606
rect 35124 27560 35256 27588
rect 35072 27542 35124 27548
rect 35256 27542 35308 27548
rect 34612 27464 34664 27470
rect 34612 27406 34664 27412
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 35164 27464 35216 27470
rect 35164 27406 35216 27412
rect 35176 27130 35204 27406
rect 35164 27124 35216 27130
rect 35164 27066 35216 27072
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35256 26444 35308 26450
rect 35256 26386 35308 26392
rect 34796 26036 34848 26042
rect 34796 25978 34848 25984
rect 34612 25832 34664 25838
rect 34612 25774 34664 25780
rect 34520 25288 34572 25294
rect 34520 25230 34572 25236
rect 34624 24954 34652 25774
rect 34808 25362 34836 25978
rect 35268 25650 35296 26386
rect 35360 26382 35388 27798
rect 35452 27538 35480 28358
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 35624 27872 35676 27878
rect 35624 27814 35676 27820
rect 35440 27532 35492 27538
rect 35440 27474 35492 27480
rect 35636 27402 35664 27814
rect 36004 27470 36032 28358
rect 36096 27538 36124 30126
rect 36188 28762 36216 30126
rect 36372 29306 36400 30194
rect 36464 29646 36492 31726
rect 36648 31414 36676 40854
rect 36832 40662 36860 40870
rect 36924 40854 37044 40882
rect 36820 40656 36872 40662
rect 36820 40598 36872 40604
rect 36924 38554 36952 40854
rect 37200 40050 37228 41074
rect 37372 40996 37424 41002
rect 37372 40938 37424 40944
rect 37188 40044 37240 40050
rect 37188 39986 37240 39992
rect 37280 39976 37332 39982
rect 37108 39924 37280 39930
rect 37108 39918 37332 39924
rect 37004 39908 37056 39914
rect 37004 39850 37056 39856
rect 37108 39902 37320 39918
rect 37016 39642 37044 39850
rect 37004 39636 37056 39642
rect 37004 39578 37056 39584
rect 37108 39302 37136 39902
rect 37096 39296 37148 39302
rect 37096 39238 37148 39244
rect 36912 38548 36964 38554
rect 36912 38490 36964 38496
rect 36912 37392 36964 37398
rect 36912 37334 36964 37340
rect 36924 37194 36952 37334
rect 36912 37188 36964 37194
rect 36912 37130 36964 37136
rect 36924 36922 36952 37130
rect 36912 36916 36964 36922
rect 36912 36858 36964 36864
rect 36820 36780 36872 36786
rect 36820 36722 36872 36728
rect 36832 36378 36860 36722
rect 36912 36712 36964 36718
rect 36912 36654 36964 36660
rect 37004 36712 37056 36718
rect 37004 36654 37056 36660
rect 36820 36372 36872 36378
rect 36820 36314 36872 36320
rect 36924 36174 36952 36654
rect 36912 36168 36964 36174
rect 36912 36110 36964 36116
rect 37016 35986 37044 36654
rect 36924 35958 37044 35986
rect 36924 35698 36952 35958
rect 36912 35692 36964 35698
rect 36912 35634 36964 35640
rect 36924 35290 36952 35634
rect 36912 35284 36964 35290
rect 36912 35226 36964 35232
rect 36820 34944 36872 34950
rect 36820 34886 36872 34892
rect 36832 34134 36860 34886
rect 36820 34128 36872 34134
rect 36820 34070 36872 34076
rect 36820 33856 36872 33862
rect 36820 33798 36872 33804
rect 36832 33658 36860 33798
rect 36820 33652 36872 33658
rect 36820 33594 36872 33600
rect 36832 32774 36860 33594
rect 36820 32768 36872 32774
rect 36820 32710 36872 32716
rect 36832 31890 36860 32710
rect 36820 31884 36872 31890
rect 36820 31826 36872 31832
rect 36636 31408 36688 31414
rect 36636 31350 36688 31356
rect 37004 31408 37056 31414
rect 37004 31350 37056 31356
rect 37016 30734 37044 31350
rect 37004 30728 37056 30734
rect 37004 30670 37056 30676
rect 36912 30660 36964 30666
rect 36912 30602 36964 30608
rect 36636 30592 36688 30598
rect 36636 30534 36688 30540
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 36556 29782 36584 30194
rect 36544 29776 36596 29782
rect 36544 29718 36596 29724
rect 36452 29640 36504 29646
rect 36452 29582 36504 29588
rect 36360 29300 36412 29306
rect 36360 29242 36412 29248
rect 36360 29028 36412 29034
rect 36360 28970 36412 28976
rect 36176 28756 36228 28762
rect 36228 28716 36308 28744
rect 36176 28698 36228 28704
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36188 28218 36216 28358
rect 36280 28218 36308 28716
rect 36372 28558 36400 28970
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 36360 28416 36412 28422
rect 36360 28358 36412 28364
rect 36176 28212 36228 28218
rect 36176 28154 36228 28160
rect 36268 28212 36320 28218
rect 36268 28154 36320 28160
rect 36268 28008 36320 28014
rect 36372 27996 36400 28358
rect 36320 27968 36400 27996
rect 36268 27950 36320 27956
rect 36084 27532 36136 27538
rect 36084 27474 36136 27480
rect 35992 27464 36044 27470
rect 35992 27406 36044 27412
rect 36268 27464 36320 27470
rect 36268 27406 36320 27412
rect 35624 27396 35676 27402
rect 35624 27338 35676 27344
rect 35440 27328 35492 27334
rect 35440 27270 35492 27276
rect 35452 26586 35480 27270
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 36004 27010 36032 27406
rect 36280 27130 36308 27406
rect 36372 27334 36400 27968
rect 36464 27554 36492 29582
rect 36544 29300 36596 29306
rect 36544 29242 36596 29248
rect 36556 28694 36584 29242
rect 36544 28688 36596 28694
rect 36544 28630 36596 28636
rect 36542 28520 36598 28529
rect 36542 28455 36598 28464
rect 36556 27962 36584 28455
rect 36648 28082 36676 30534
rect 36924 30394 36952 30602
rect 36912 30388 36964 30394
rect 36912 30330 36964 30336
rect 36728 30252 36780 30258
rect 36780 30212 36860 30240
rect 36728 30194 36780 30200
rect 36728 28688 36780 28694
rect 36728 28630 36780 28636
rect 36740 28422 36768 28630
rect 36728 28416 36780 28422
rect 36728 28358 36780 28364
rect 36636 28076 36688 28082
rect 36636 28018 36688 28024
rect 36556 27934 36676 27962
rect 36464 27526 36584 27554
rect 36452 27464 36504 27470
rect 36452 27406 36504 27412
rect 36360 27328 36412 27334
rect 36360 27270 36412 27276
rect 36268 27124 36320 27130
rect 36268 27066 36320 27072
rect 36464 27062 36492 27406
rect 36452 27056 36504 27062
rect 36004 26982 36400 27010
rect 36452 26998 36504 27004
rect 35440 26580 35492 26586
rect 35440 26522 35492 26528
rect 35440 26444 35492 26450
rect 35440 26386 35492 26392
rect 35348 26376 35400 26382
rect 35348 26318 35400 26324
rect 35360 26042 35388 26318
rect 35348 26036 35400 26042
rect 35348 25978 35400 25984
rect 35268 25622 35388 25650
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35164 25492 35216 25498
rect 35164 25434 35216 25440
rect 34796 25356 34848 25362
rect 34796 25298 34848 25304
rect 34612 24948 34664 24954
rect 34612 24890 34664 24896
rect 34704 24880 34756 24886
rect 34624 24828 34704 24834
rect 34624 24822 34756 24828
rect 34152 24812 34204 24818
rect 34520 24812 34572 24818
rect 34204 24772 34284 24800
rect 34152 24754 34204 24760
rect 34072 22066 34192 22094
rect 34060 20936 34112 20942
rect 34060 20878 34112 20884
rect 34072 20602 34100 20878
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34060 20460 34112 20466
rect 34060 20402 34112 20408
rect 34072 19378 34100 20402
rect 34164 19854 34192 22066
rect 34152 19848 34204 19854
rect 34152 19790 34204 19796
rect 34256 19378 34284 24772
rect 34520 24754 34572 24760
rect 34624 24806 34744 24822
rect 34532 24342 34560 24754
rect 34520 24336 34572 24342
rect 34520 24278 34572 24284
rect 34334 24168 34390 24177
rect 34334 24103 34390 24112
rect 34348 21622 34376 24103
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34532 22982 34560 23598
rect 34520 22976 34572 22982
rect 34520 22918 34572 22924
rect 34336 21616 34388 21622
rect 34336 21558 34388 21564
rect 34336 21344 34388 21350
rect 34336 21286 34388 21292
rect 34348 19938 34376 21286
rect 34428 20460 34480 20466
rect 34428 20402 34480 20408
rect 34440 20058 34468 20402
rect 34428 20052 34480 20058
rect 34428 19994 34480 20000
rect 34348 19910 34468 19938
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 34348 19378 34376 19450
rect 34060 19372 34112 19378
rect 34060 19314 34112 19320
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34336 19372 34388 19378
rect 34336 19314 34388 19320
rect 34060 18624 34112 18630
rect 34060 18566 34112 18572
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 33600 16040 33652 16046
rect 33600 15982 33652 15988
rect 33612 15706 33640 15982
rect 33600 15700 33652 15706
rect 33600 15642 33652 15648
rect 33980 15502 34008 16186
rect 33968 15496 34020 15502
rect 33968 15438 34020 15444
rect 33968 14408 34020 14414
rect 33968 14350 34020 14356
rect 33416 14068 33468 14074
rect 33416 14010 33468 14016
rect 33508 14068 33560 14074
rect 33508 14010 33560 14016
rect 32864 13796 32916 13802
rect 32864 13738 32916 13744
rect 33140 13796 33192 13802
rect 33140 13738 33192 13744
rect 32876 13394 32904 13738
rect 32956 13728 33008 13734
rect 32956 13670 33008 13676
rect 32864 13388 32916 13394
rect 32864 13330 32916 13336
rect 32864 13252 32916 13258
rect 32864 13194 32916 13200
rect 32496 12844 32548 12850
rect 32496 12786 32548 12792
rect 32876 12782 32904 13194
rect 32968 12986 32996 13670
rect 32956 12980 33008 12986
rect 32956 12922 33008 12928
rect 33152 12866 33180 13738
rect 33416 13728 33468 13734
rect 33416 13670 33468 13676
rect 33428 12918 33456 13670
rect 32968 12850 33180 12866
rect 33416 12912 33468 12918
rect 33416 12854 33468 12860
rect 32956 12844 33180 12850
rect 33008 12838 33180 12844
rect 32956 12786 33008 12792
rect 33980 12782 34008 14350
rect 34072 13938 34100 18566
rect 34336 16720 34388 16726
rect 34336 16662 34388 16668
rect 34242 16008 34298 16017
rect 34242 15943 34298 15952
rect 34256 15638 34284 15943
rect 34244 15632 34296 15638
rect 34244 15574 34296 15580
rect 34256 15026 34284 15574
rect 34244 15020 34296 15026
rect 34244 14962 34296 14968
rect 34348 14906 34376 16662
rect 34164 14878 34376 14906
rect 34060 13932 34112 13938
rect 34060 13874 34112 13880
rect 34164 13326 34192 14878
rect 34336 14408 34388 14414
rect 34336 14350 34388 14356
rect 34244 14272 34296 14278
rect 34244 14214 34296 14220
rect 34256 14074 34284 14214
rect 34244 14068 34296 14074
rect 34244 14010 34296 14016
rect 34348 13462 34376 14350
rect 34440 14074 34468 19910
rect 34532 19258 34560 22918
rect 34624 21049 34652 24806
rect 34704 23520 34756 23526
rect 34704 23462 34756 23468
rect 34716 22710 34744 23462
rect 34808 23322 34836 25298
rect 35176 24954 35204 25434
rect 35360 25430 35388 25622
rect 35348 25424 35400 25430
rect 35348 25366 35400 25372
rect 35256 25152 35308 25158
rect 35256 25094 35308 25100
rect 35268 24954 35296 25094
rect 35164 24948 35216 24954
rect 35164 24890 35216 24896
rect 35256 24948 35308 24954
rect 35256 24890 35308 24896
rect 34886 24848 34942 24857
rect 34886 24783 34942 24792
rect 35164 24812 35216 24818
rect 34900 24750 34928 24783
rect 35164 24754 35216 24760
rect 34888 24744 34940 24750
rect 34888 24686 34940 24692
rect 35176 24596 35204 24754
rect 35360 24750 35388 25366
rect 35452 24857 35480 26386
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 36004 25294 36032 26250
rect 36096 25702 36124 26318
rect 36176 26240 36228 26246
rect 36176 26182 36228 26188
rect 36084 25696 36136 25702
rect 36084 25638 36136 25644
rect 36096 25498 36124 25638
rect 36084 25492 36136 25498
rect 36084 25434 36136 25440
rect 36188 25362 36216 26182
rect 36268 25696 36320 25702
rect 36268 25638 36320 25644
rect 36176 25356 36228 25362
rect 36176 25298 36228 25304
rect 35992 25288 36044 25294
rect 35898 25256 35954 25265
rect 35992 25230 36044 25236
rect 35898 25191 35954 25200
rect 36084 25220 36136 25226
rect 35912 25140 35940 25191
rect 36084 25162 36136 25168
rect 35912 25112 36032 25140
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 36004 24954 36032 25112
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 35624 24880 35676 24886
rect 35438 24848 35494 24857
rect 35624 24822 35676 24828
rect 35438 24783 35440 24792
rect 35492 24783 35494 24792
rect 35440 24754 35492 24760
rect 35348 24744 35400 24750
rect 35346 24712 35348 24721
rect 35400 24712 35402 24721
rect 35346 24647 35402 24656
rect 35176 24568 35480 24596
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35452 24410 35480 24568
rect 35256 24404 35308 24410
rect 35256 24346 35308 24352
rect 35440 24404 35492 24410
rect 35440 24346 35492 24352
rect 35268 24290 35296 24346
rect 35176 24262 35296 24290
rect 35636 24274 35664 24822
rect 36096 24750 36124 25162
rect 36084 24744 36136 24750
rect 36084 24686 36136 24692
rect 36188 24682 36216 25298
rect 36280 24886 36308 25638
rect 36268 24880 36320 24886
rect 36268 24822 36320 24828
rect 36176 24676 36228 24682
rect 36176 24618 36228 24624
rect 36174 24576 36230 24585
rect 36174 24511 36230 24520
rect 36188 24274 36216 24511
rect 35624 24268 35676 24274
rect 35176 23798 35204 24262
rect 35624 24210 35676 24216
rect 36176 24268 36228 24274
rect 36176 24210 36228 24216
rect 36280 24206 36308 24822
rect 36372 24750 36400 26982
rect 36556 26314 36584 27526
rect 36648 27062 36676 27934
rect 36636 27056 36688 27062
rect 36636 26998 36688 27004
rect 36648 26586 36676 26998
rect 36636 26580 36688 26586
rect 36636 26522 36688 26528
rect 36544 26308 36596 26314
rect 36544 26250 36596 26256
rect 36452 25492 36504 25498
rect 36452 25434 36504 25440
rect 36464 25362 36492 25434
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 36648 24970 36676 26522
rect 36728 26444 36780 26450
rect 36728 26386 36780 26392
rect 36740 26042 36768 26386
rect 36728 26036 36780 26042
rect 36728 25978 36780 25984
rect 36464 24942 36676 24970
rect 36360 24744 36412 24750
rect 36360 24686 36412 24692
rect 36464 24410 36492 24942
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 36556 24410 36584 24754
rect 36636 24676 36688 24682
rect 36636 24618 36688 24624
rect 36452 24404 36504 24410
rect 36452 24346 36504 24352
rect 36544 24404 36596 24410
rect 36544 24346 36596 24352
rect 36268 24200 36320 24206
rect 35530 24168 35586 24177
rect 36268 24142 36320 24148
rect 36464 24188 36492 24346
rect 36544 24200 36596 24206
rect 36464 24160 36544 24188
rect 35530 24103 35532 24112
rect 35584 24103 35586 24112
rect 35532 24074 35584 24080
rect 36464 24070 36492 24160
rect 36544 24142 36596 24148
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 36452 24064 36504 24070
rect 36452 24006 36504 24012
rect 35164 23792 35216 23798
rect 35164 23734 35216 23740
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 23316 34848 23322
rect 34796 23258 34848 23264
rect 34888 23112 34940 23118
rect 34888 23054 34940 23060
rect 34900 22778 34928 23054
rect 35360 22982 35388 23666
rect 35452 23050 35480 24006
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 36464 23322 36492 24006
rect 36084 23316 36136 23322
rect 36084 23258 36136 23264
rect 36452 23316 36504 23322
rect 36452 23258 36504 23264
rect 35440 23044 35492 23050
rect 35440 22986 35492 22992
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 34888 22772 34940 22778
rect 34888 22714 34940 22720
rect 34704 22704 34756 22710
rect 34704 22646 34756 22652
rect 34796 22432 34848 22438
rect 34716 22392 34796 22420
rect 34716 21486 34744 22392
rect 34796 22374 34848 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35360 22234 35388 22918
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 34796 22228 34848 22234
rect 34796 22170 34848 22176
rect 35348 22228 35400 22234
rect 35348 22170 35400 22176
rect 34704 21480 34756 21486
rect 34704 21422 34756 21428
rect 34610 21040 34666 21049
rect 34610 20975 34666 20984
rect 34532 19230 34652 19258
rect 34520 19168 34572 19174
rect 34520 19110 34572 19116
rect 34532 18834 34560 19110
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34624 18714 34652 19230
rect 34532 18686 34652 18714
rect 34428 14068 34480 14074
rect 34428 14010 34480 14016
rect 34532 14006 34560 18686
rect 34612 18216 34664 18222
rect 34612 18158 34664 18164
rect 34624 17610 34652 18158
rect 34612 17604 34664 17610
rect 34612 17546 34664 17552
rect 34624 16114 34652 17546
rect 34612 16108 34664 16114
rect 34612 16050 34664 16056
rect 34716 15994 34744 21422
rect 34808 19802 34836 22170
rect 35256 21956 35308 21962
rect 35256 21898 35308 21904
rect 35268 21690 35296 21898
rect 35256 21684 35308 21690
rect 35256 21626 35308 21632
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34888 21072 34940 21078
rect 34888 21014 34940 21020
rect 34978 21040 35034 21049
rect 34900 20874 34928 21014
rect 35360 21026 35388 21490
rect 34978 20975 35034 20984
rect 35268 20998 35388 21026
rect 34992 20942 35020 20975
rect 35268 20942 35296 20998
rect 34980 20936 35032 20942
rect 34980 20878 35032 20884
rect 35256 20936 35308 20942
rect 35256 20878 35308 20884
rect 35348 20936 35400 20942
rect 35348 20878 35400 20884
rect 34888 20868 34940 20874
rect 34888 20810 34940 20816
rect 35360 20330 35388 20878
rect 35348 20324 35400 20330
rect 35348 20266 35400 20272
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34808 19774 34928 19802
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34808 17270 34836 19654
rect 34900 19174 34928 19774
rect 34888 19168 34940 19174
rect 34888 19110 34940 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34980 17604 35032 17610
rect 34980 17546 35032 17552
rect 34992 17338 35020 17546
rect 34980 17332 35032 17338
rect 34980 17274 35032 17280
rect 34796 17264 34848 17270
rect 34796 17206 34848 17212
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16726 35388 20266
rect 35452 19394 35480 22714
rect 35532 22704 35584 22710
rect 35532 22646 35584 22652
rect 35544 22030 35572 22646
rect 36096 22094 36124 23258
rect 36004 22066 36124 22094
rect 35532 22024 35584 22030
rect 35532 21966 35584 21972
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 36004 21622 36032 22066
rect 36084 21888 36136 21894
rect 36084 21830 36136 21836
rect 36452 21888 36504 21894
rect 36452 21830 36504 21836
rect 35992 21616 36044 21622
rect 35992 21558 36044 21564
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 35636 21350 35664 21490
rect 36096 21468 36124 21830
rect 36464 21554 36492 21830
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36004 21440 36124 21468
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35636 21146 35664 21286
rect 35624 21140 35676 21146
rect 35624 21082 35676 21088
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35532 20256 35584 20262
rect 35532 20198 35584 20204
rect 35544 19922 35572 20198
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35452 19366 35572 19394
rect 35544 18630 35572 19366
rect 35624 19372 35676 19378
rect 35624 19314 35676 19320
rect 35636 18970 35664 19314
rect 35624 18964 35676 18970
rect 35624 18906 35676 18912
rect 35532 18624 35584 18630
rect 35532 18566 35584 18572
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35440 18420 35492 18426
rect 35440 18362 35492 18368
rect 35452 17610 35480 18362
rect 35440 17604 35492 17610
rect 35440 17546 35492 17552
rect 35348 16720 35400 16726
rect 35348 16662 35400 16668
rect 35348 16176 35400 16182
rect 35452 16164 35480 17546
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35400 16136 35480 16164
rect 35348 16118 35400 16124
rect 34624 15966 34744 15994
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35532 16040 35584 16046
rect 35532 15982 35584 15988
rect 34520 14000 34572 14006
rect 34520 13942 34572 13948
rect 34624 13870 34652 15966
rect 35348 15904 35400 15910
rect 35348 15846 35400 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34888 15496 34940 15502
rect 34888 15438 34940 15444
rect 34716 14890 34744 15438
rect 34900 14958 34928 15438
rect 35360 15094 35388 15846
rect 35452 15706 35480 15982
rect 35440 15700 35492 15706
rect 35440 15642 35492 15648
rect 35544 15502 35572 15982
rect 35532 15496 35584 15502
rect 35532 15438 35584 15444
rect 35440 15360 35492 15366
rect 35440 15302 35492 15308
rect 35348 15088 35400 15094
rect 35348 15030 35400 15036
rect 35452 15026 35480 15302
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 34888 14952 34940 14958
rect 34888 14894 34940 14900
rect 34704 14884 34756 14890
rect 34704 14826 34756 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 14476 34756 14482
rect 34704 14418 34756 14424
rect 34612 13864 34664 13870
rect 34612 13806 34664 13812
rect 34428 13796 34480 13802
rect 34428 13738 34480 13744
rect 34336 13456 34388 13462
rect 34440 13433 34468 13738
rect 34336 13398 34388 13404
rect 34426 13424 34482 13433
rect 34152 13320 34204 13326
rect 34152 13262 34204 13268
rect 32864 12776 32916 12782
rect 32864 12718 32916 12724
rect 33968 12776 34020 12782
rect 33968 12718 34020 12724
rect 32404 11824 32456 11830
rect 32404 11766 32456 11772
rect 32416 11218 32444 11766
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 32508 11218 32536 11698
rect 32588 11688 32640 11694
rect 32588 11630 32640 11636
rect 32600 11354 32628 11630
rect 32876 11626 32904 12718
rect 34348 11830 34376 13398
rect 34426 13359 34482 13368
rect 34428 13252 34480 13258
rect 34428 13194 34480 13200
rect 34440 12850 34468 13194
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34716 12714 34744 14418
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 35452 14074 35480 14214
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 35256 13864 35308 13870
rect 34886 13832 34942 13841
rect 35308 13812 35388 13818
rect 35256 13806 35388 13812
rect 35268 13790 35388 13806
rect 34886 13767 34942 13776
rect 34900 13734 34928 13767
rect 34888 13728 34940 13734
rect 34888 13670 34940 13676
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34980 13524 35032 13530
rect 34980 13466 35032 13472
rect 34992 13297 35020 13466
rect 35360 13394 35388 13790
rect 35532 13728 35584 13734
rect 35532 13670 35584 13676
rect 35348 13388 35400 13394
rect 35348 13330 35400 13336
rect 34978 13288 35034 13297
rect 35544 13258 35572 13670
rect 36004 13297 36032 21440
rect 36268 20800 36320 20806
rect 36268 20742 36320 20748
rect 36084 19168 36136 19174
rect 36084 19110 36136 19116
rect 36096 17762 36124 19110
rect 36176 18828 36228 18834
rect 36176 18770 36228 18776
rect 36188 17882 36216 18770
rect 36176 17876 36228 17882
rect 36176 17818 36228 17824
rect 36096 17734 36216 17762
rect 36084 16652 36136 16658
rect 36084 16594 36136 16600
rect 36096 15026 36124 16594
rect 36084 15020 36136 15026
rect 36084 14962 36136 14968
rect 36188 13530 36216 17734
rect 36280 14618 36308 20742
rect 36360 20256 36412 20262
rect 36360 20198 36412 20204
rect 36372 19786 36400 20198
rect 36360 19780 36412 19786
rect 36360 19722 36412 19728
rect 36452 17536 36504 17542
rect 36452 17478 36504 17484
rect 36544 17536 36596 17542
rect 36544 17478 36596 17484
rect 36464 16726 36492 17478
rect 36556 17338 36584 17478
rect 36648 17338 36676 24618
rect 36740 24614 36768 25978
rect 36832 25498 36860 30212
rect 36924 28966 36952 30330
rect 37108 29782 37136 39238
rect 37384 38894 37412 40938
rect 38212 40594 38240 41074
rect 38200 40588 38252 40594
rect 38200 40530 38252 40536
rect 37832 40520 37884 40526
rect 37832 40462 37884 40468
rect 37844 40186 37872 40462
rect 38108 40452 38160 40458
rect 38108 40394 38160 40400
rect 37832 40180 37884 40186
rect 37832 40122 37884 40128
rect 37740 39840 37792 39846
rect 37740 39782 37792 39788
rect 37924 39840 37976 39846
rect 37924 39782 37976 39788
rect 37752 39506 37780 39782
rect 37740 39500 37792 39506
rect 37740 39442 37792 39448
rect 37464 39364 37516 39370
rect 37464 39306 37516 39312
rect 37476 39098 37504 39306
rect 37936 39098 37964 39782
rect 37464 39092 37516 39098
rect 37464 39034 37516 39040
rect 37924 39092 37976 39098
rect 37924 39034 37976 39040
rect 37372 38888 37424 38894
rect 37372 38830 37424 38836
rect 37372 38752 37424 38758
rect 37372 38694 37424 38700
rect 37384 38418 37412 38694
rect 37556 38548 37608 38554
rect 37556 38490 37608 38496
rect 37372 38412 37424 38418
rect 37372 38354 37424 38360
rect 37372 37732 37424 37738
rect 37372 37674 37424 37680
rect 37384 37262 37412 37674
rect 37464 37664 37516 37670
rect 37464 37606 37516 37612
rect 37476 37398 37504 37606
rect 37464 37392 37516 37398
rect 37464 37334 37516 37340
rect 37372 37256 37424 37262
rect 37372 37198 37424 37204
rect 37372 36168 37424 36174
rect 37372 36110 37424 36116
rect 37280 35148 37332 35154
rect 37280 35090 37332 35096
rect 37292 35034 37320 35090
rect 37384 35034 37412 36110
rect 37292 35006 37412 35034
rect 37384 34542 37412 35006
rect 37372 34536 37424 34542
rect 37372 34478 37424 34484
rect 37384 33454 37412 34478
rect 37372 33448 37424 33454
rect 37372 33390 37424 33396
rect 37384 32910 37412 33390
rect 37372 32904 37424 32910
rect 37372 32846 37424 32852
rect 37384 32366 37412 32846
rect 37372 32360 37424 32366
rect 37372 32302 37424 32308
rect 37384 31822 37412 32302
rect 37372 31816 37424 31822
rect 37372 31758 37424 31764
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 37292 29850 37320 31282
rect 37384 30734 37412 31758
rect 37464 31340 37516 31346
rect 37464 31282 37516 31288
rect 37476 30938 37504 31282
rect 37464 30932 37516 30938
rect 37464 30874 37516 30880
rect 37372 30728 37424 30734
rect 37372 30670 37424 30676
rect 37280 29844 37332 29850
rect 37280 29786 37332 29792
rect 37096 29776 37148 29782
rect 37096 29718 37148 29724
rect 37280 29640 37332 29646
rect 37280 29582 37332 29588
rect 37188 29504 37240 29510
rect 37188 29446 37240 29452
rect 37200 29102 37228 29446
rect 37188 29096 37240 29102
rect 37188 29038 37240 29044
rect 36912 28960 36964 28966
rect 36912 28902 36964 28908
rect 36924 28014 36952 28902
rect 37004 28552 37056 28558
rect 37004 28494 37056 28500
rect 36912 28008 36964 28014
rect 36912 27950 36964 27956
rect 37016 27878 37044 28494
rect 36912 27872 36964 27878
rect 36912 27814 36964 27820
rect 37004 27872 37056 27878
rect 37004 27814 37056 27820
rect 36924 27010 36952 27814
rect 37016 27538 37044 27814
rect 37292 27538 37320 29582
rect 37384 28626 37412 30670
rect 37568 29322 37596 38490
rect 37924 38344 37976 38350
rect 37924 38286 37976 38292
rect 37936 38010 37964 38286
rect 37924 38004 37976 38010
rect 37924 37946 37976 37952
rect 37648 37868 37700 37874
rect 37648 37810 37700 37816
rect 37660 37262 37688 37810
rect 37740 37732 37792 37738
rect 37740 37674 37792 37680
rect 37752 37398 37780 37674
rect 37740 37392 37792 37398
rect 37740 37334 37792 37340
rect 37648 37256 37700 37262
rect 37648 37198 37700 37204
rect 37660 36922 37688 37198
rect 37648 36916 37700 36922
rect 37648 36858 37700 36864
rect 38120 36242 38148 40394
rect 38212 40118 38240 40530
rect 39304 40520 39356 40526
rect 39304 40462 39356 40468
rect 42156 40520 42208 40526
rect 42156 40462 42208 40468
rect 38200 40112 38252 40118
rect 38200 40054 38252 40060
rect 38212 39506 38240 40054
rect 39316 39982 39344 40462
rect 41052 40384 41104 40390
rect 41052 40326 41104 40332
rect 39580 40044 39632 40050
rect 39580 39986 39632 39992
rect 39672 40044 39724 40050
rect 39672 39986 39724 39992
rect 38476 39976 38528 39982
rect 38476 39918 38528 39924
rect 39304 39976 39356 39982
rect 39304 39918 39356 39924
rect 38200 39500 38252 39506
rect 38200 39442 38252 39448
rect 38292 39296 38344 39302
rect 38292 39238 38344 39244
rect 38304 38350 38332 39238
rect 38488 39098 38516 39918
rect 38936 39908 38988 39914
rect 38936 39850 38988 39856
rect 39028 39908 39080 39914
rect 39028 39850 39080 39856
rect 38948 39642 38976 39850
rect 38936 39636 38988 39642
rect 38936 39578 38988 39584
rect 39040 39574 39068 39850
rect 39592 39642 39620 39986
rect 39684 39914 39712 39986
rect 40316 39976 40368 39982
rect 40316 39918 40368 39924
rect 39672 39908 39724 39914
rect 39672 39850 39724 39856
rect 39580 39636 39632 39642
rect 39580 39578 39632 39584
rect 39028 39568 39080 39574
rect 39028 39510 39080 39516
rect 38936 39432 38988 39438
rect 38936 39374 38988 39380
rect 39396 39432 39448 39438
rect 39396 39374 39448 39380
rect 38476 39092 38528 39098
rect 38476 39034 38528 39040
rect 38948 38826 38976 39374
rect 39408 38962 39436 39374
rect 39580 39364 39632 39370
rect 39684 39352 39712 39850
rect 39948 39432 40000 39438
rect 39948 39374 40000 39380
rect 40224 39432 40276 39438
rect 40224 39374 40276 39380
rect 39632 39324 39712 39352
rect 39580 39306 39632 39312
rect 39396 38956 39448 38962
rect 39396 38898 39448 38904
rect 39120 38888 39172 38894
rect 39120 38830 39172 38836
rect 38936 38820 38988 38826
rect 38936 38762 38988 38768
rect 39132 38350 39160 38830
rect 39684 38826 39712 39324
rect 39960 39098 39988 39374
rect 40040 39364 40092 39370
rect 40040 39306 40092 39312
rect 40132 39364 40184 39370
rect 40132 39306 40184 39312
rect 40052 39098 40080 39306
rect 39948 39092 40000 39098
rect 39948 39034 40000 39040
rect 40040 39092 40092 39098
rect 40040 39034 40092 39040
rect 40144 38962 40172 39306
rect 40236 38962 40264 39374
rect 40132 38956 40184 38962
rect 40052 38916 40132 38944
rect 39672 38820 39724 38826
rect 39672 38762 39724 38768
rect 38292 38344 38344 38350
rect 38292 38286 38344 38292
rect 39120 38344 39172 38350
rect 39120 38286 39172 38292
rect 39396 38344 39448 38350
rect 39396 38286 39448 38292
rect 38304 37738 38332 38286
rect 38476 37868 38528 37874
rect 38476 37810 38528 37816
rect 38292 37732 38344 37738
rect 38292 37674 38344 37680
rect 38488 36922 38516 37810
rect 39408 37670 39436 38286
rect 39856 37936 39908 37942
rect 39856 37878 39908 37884
rect 39396 37664 39448 37670
rect 39396 37606 39448 37612
rect 39408 37466 39436 37606
rect 39868 37466 39896 37878
rect 40052 37874 40080 38916
rect 40132 38898 40184 38904
rect 40224 38956 40276 38962
rect 40224 38898 40276 38904
rect 40328 38554 40356 39918
rect 40776 39500 40828 39506
rect 40776 39442 40828 39448
rect 40684 39364 40736 39370
rect 40684 39306 40736 39312
rect 40696 39098 40724 39306
rect 40684 39092 40736 39098
rect 40684 39034 40736 39040
rect 40500 38752 40552 38758
rect 40500 38694 40552 38700
rect 40316 38548 40368 38554
rect 40316 38490 40368 38496
rect 40512 38010 40540 38694
rect 40592 38276 40644 38282
rect 40592 38218 40644 38224
rect 40500 38004 40552 38010
rect 40500 37946 40552 37952
rect 39948 37868 40000 37874
rect 39948 37810 40000 37816
rect 40040 37868 40092 37874
rect 40040 37810 40092 37816
rect 40316 37868 40368 37874
rect 40316 37810 40368 37816
rect 39396 37460 39448 37466
rect 39396 37402 39448 37408
rect 39856 37460 39908 37466
rect 39856 37402 39908 37408
rect 39960 37262 39988 37810
rect 40052 37262 40080 37810
rect 40328 37670 40356 37810
rect 40316 37664 40368 37670
rect 40316 37606 40368 37612
rect 39948 37256 40000 37262
rect 39948 37198 40000 37204
rect 40040 37256 40092 37262
rect 40040 37198 40092 37204
rect 39960 36922 39988 37198
rect 38476 36916 38528 36922
rect 38476 36858 38528 36864
rect 39948 36916 40000 36922
rect 39948 36858 40000 36864
rect 38200 36780 38252 36786
rect 38200 36722 38252 36728
rect 38292 36780 38344 36786
rect 38292 36722 38344 36728
rect 38936 36780 38988 36786
rect 38936 36722 38988 36728
rect 39120 36780 39172 36786
rect 39120 36722 39172 36728
rect 38212 36582 38240 36722
rect 38200 36576 38252 36582
rect 38200 36518 38252 36524
rect 38304 36378 38332 36722
rect 38948 36582 38976 36722
rect 38936 36576 38988 36582
rect 38936 36518 38988 36524
rect 39028 36576 39080 36582
rect 39028 36518 39080 36524
rect 38292 36372 38344 36378
rect 38292 36314 38344 36320
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 37648 36100 37700 36106
rect 37648 36042 37700 36048
rect 37660 35834 37688 36042
rect 37648 35828 37700 35834
rect 37648 35770 37700 35776
rect 38120 35018 38148 36178
rect 38752 36168 38804 36174
rect 38752 36110 38804 36116
rect 38476 35624 38528 35630
rect 38476 35566 38528 35572
rect 38488 35154 38516 35566
rect 38476 35148 38528 35154
rect 38476 35090 38528 35096
rect 38108 35012 38160 35018
rect 38108 34954 38160 34960
rect 37924 34944 37976 34950
rect 37924 34886 37976 34892
rect 37936 34678 37964 34886
rect 37924 34672 37976 34678
rect 37924 34614 37976 34620
rect 38120 33522 38148 34954
rect 38384 34944 38436 34950
rect 38384 34886 38436 34892
rect 38396 34202 38424 34886
rect 38764 34610 38792 36110
rect 38948 36038 38976 36518
rect 39040 36174 39068 36518
rect 39132 36378 39160 36722
rect 39212 36712 39264 36718
rect 40052 36666 40080 37198
rect 40328 37194 40356 37606
rect 40316 37188 40368 37194
rect 40316 37130 40368 37136
rect 40408 37188 40460 37194
rect 40408 37130 40460 37136
rect 40500 37188 40552 37194
rect 40500 37130 40552 37136
rect 39212 36654 39264 36660
rect 39120 36372 39172 36378
rect 39120 36314 39172 36320
rect 39224 36174 39252 36654
rect 39868 36650 40080 36666
rect 39396 36644 39448 36650
rect 39396 36586 39448 36592
rect 39856 36644 40080 36650
rect 39908 36638 40080 36644
rect 39856 36586 39908 36592
rect 39408 36174 39436 36586
rect 40040 36576 40092 36582
rect 40040 36518 40092 36524
rect 39028 36168 39080 36174
rect 39028 36110 39080 36116
rect 39212 36168 39264 36174
rect 39212 36110 39264 36116
rect 39396 36168 39448 36174
rect 39396 36110 39448 36116
rect 38936 36032 38988 36038
rect 38936 35974 38988 35980
rect 39120 35760 39172 35766
rect 39120 35702 39172 35708
rect 38936 35012 38988 35018
rect 38936 34954 38988 34960
rect 38948 34746 38976 34954
rect 38936 34740 38988 34746
rect 38936 34682 38988 34688
rect 38752 34604 38804 34610
rect 38752 34546 38804 34552
rect 38384 34196 38436 34202
rect 38384 34138 38436 34144
rect 38936 33924 38988 33930
rect 38936 33866 38988 33872
rect 38660 33856 38712 33862
rect 38660 33798 38712 33804
rect 38672 33674 38700 33798
rect 38672 33658 38792 33674
rect 38672 33652 38804 33658
rect 38672 33646 38752 33652
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 38568 33516 38620 33522
rect 38568 33458 38620 33464
rect 38384 33448 38436 33454
rect 38384 33390 38436 33396
rect 37648 33312 37700 33318
rect 37648 33254 37700 33260
rect 37660 32910 37688 33254
rect 37648 32904 37700 32910
rect 37648 32846 37700 32852
rect 37648 32428 37700 32434
rect 37648 32370 37700 32376
rect 37660 32026 37688 32370
rect 38292 32224 38344 32230
rect 38292 32166 38344 32172
rect 37648 32020 37700 32026
rect 37648 31962 37700 31968
rect 38304 31890 38332 32166
rect 38292 31884 38344 31890
rect 38292 31826 38344 31832
rect 38396 31754 38424 33390
rect 38580 32994 38608 33458
rect 38672 33114 38700 33646
rect 38752 33594 38804 33600
rect 38844 33312 38896 33318
rect 38844 33254 38896 33260
rect 38856 33114 38884 33254
rect 38660 33108 38712 33114
rect 38660 33050 38712 33056
rect 38844 33108 38896 33114
rect 38844 33050 38896 33056
rect 38580 32966 38792 32994
rect 38396 31726 38516 31754
rect 38292 31680 38344 31686
rect 38292 31622 38344 31628
rect 37832 31340 37884 31346
rect 37832 31282 37884 31288
rect 37740 31204 37792 31210
rect 37740 31146 37792 31152
rect 37648 31136 37700 31142
rect 37648 31078 37700 31084
rect 37660 30802 37688 31078
rect 37648 30796 37700 30802
rect 37648 30738 37700 30744
rect 37648 30320 37700 30326
rect 37648 30262 37700 30268
rect 37660 29714 37688 30262
rect 37648 29708 37700 29714
rect 37648 29650 37700 29656
rect 37476 29294 37596 29322
rect 37372 28620 37424 28626
rect 37372 28562 37424 28568
rect 37476 28218 37504 29294
rect 37556 29164 37608 29170
rect 37556 29106 37608 29112
rect 37568 28218 37596 29106
rect 37752 29034 37780 31146
rect 37844 30394 37872 31282
rect 38304 30598 38332 31622
rect 37924 30592 37976 30598
rect 37924 30534 37976 30540
rect 38292 30592 38344 30598
rect 38292 30534 38344 30540
rect 37936 30394 37964 30534
rect 37832 30388 37884 30394
rect 37832 30330 37884 30336
rect 37924 30388 37976 30394
rect 37924 30330 37976 30336
rect 38108 30252 38160 30258
rect 38304 30240 38332 30534
rect 38160 30212 38332 30240
rect 38108 30194 38160 30200
rect 37832 30184 37884 30190
rect 37832 30126 37884 30132
rect 37844 29646 37872 30126
rect 38120 29850 38148 30194
rect 38384 30116 38436 30122
rect 38384 30058 38436 30064
rect 38108 29844 38160 29850
rect 38108 29786 38160 29792
rect 38292 29844 38344 29850
rect 38292 29786 38344 29792
rect 37832 29640 37884 29646
rect 37832 29582 37884 29588
rect 38200 29640 38252 29646
rect 38200 29582 38252 29588
rect 37844 29102 37872 29582
rect 37924 29504 37976 29510
rect 37924 29446 37976 29452
rect 37936 29238 37964 29446
rect 37924 29232 37976 29238
rect 38108 29198 38160 29204
rect 37924 29174 37976 29180
rect 38028 29158 38108 29186
rect 37832 29096 37884 29102
rect 38028 29050 38056 29158
rect 38108 29140 38160 29146
rect 37884 29044 38056 29050
rect 37832 29038 38056 29044
rect 38108 29096 38160 29102
rect 38108 29038 38160 29044
rect 37740 29028 37792 29034
rect 37844 29022 38056 29038
rect 37740 28970 37792 28976
rect 37648 28960 37700 28966
rect 37648 28902 37700 28908
rect 37660 28626 37688 28902
rect 37752 28762 37780 28970
rect 37740 28756 37792 28762
rect 37740 28698 37792 28704
rect 37648 28620 37700 28626
rect 37648 28562 37700 28568
rect 37740 28416 37792 28422
rect 37740 28358 37792 28364
rect 37464 28212 37516 28218
rect 37464 28154 37516 28160
rect 37556 28212 37608 28218
rect 37556 28154 37608 28160
rect 37752 28082 37780 28358
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37740 28076 37792 28082
rect 37740 28018 37792 28024
rect 37004 27532 37056 27538
rect 37004 27474 37056 27480
rect 37280 27532 37332 27538
rect 37280 27474 37332 27480
rect 37016 27130 37044 27474
rect 37004 27124 37056 27130
rect 37004 27066 37056 27072
rect 36924 26982 37044 27010
rect 36912 26240 36964 26246
rect 36912 26182 36964 26188
rect 36924 25906 36952 26182
rect 36912 25900 36964 25906
rect 36912 25842 36964 25848
rect 36820 25492 36872 25498
rect 36820 25434 36872 25440
rect 36820 25152 36872 25158
rect 36820 25094 36872 25100
rect 36832 24818 36860 25094
rect 36820 24812 36872 24818
rect 36820 24754 36872 24760
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36740 24342 36768 24550
rect 36728 24336 36780 24342
rect 36728 24278 36780 24284
rect 36832 24138 36860 24754
rect 36924 24410 36952 25842
rect 37016 25838 37044 26982
rect 37476 26382 37504 28018
rect 37924 28008 37976 28014
rect 37924 27950 37976 27956
rect 37936 27577 37964 27950
rect 37922 27568 37978 27577
rect 37922 27503 37978 27512
rect 38120 27402 38148 29038
rect 38108 27396 38160 27402
rect 38108 27338 38160 27344
rect 37832 27328 37884 27334
rect 37832 27270 37884 27276
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 37844 26450 37872 27270
rect 37832 26444 37884 26450
rect 37832 26386 37884 26392
rect 38028 26382 38056 27270
rect 37464 26376 37516 26382
rect 37464 26318 37516 26324
rect 38016 26376 38068 26382
rect 38016 26318 38068 26324
rect 37372 25900 37424 25906
rect 37372 25842 37424 25848
rect 37004 25832 37056 25838
rect 37004 25774 37056 25780
rect 36912 24404 36964 24410
rect 36912 24346 36964 24352
rect 36820 24132 36872 24138
rect 36820 24074 36872 24080
rect 37016 23050 37044 25774
rect 37096 25696 37148 25702
rect 37096 25638 37148 25644
rect 37280 25696 37332 25702
rect 37280 25638 37332 25644
rect 37108 24206 37136 25638
rect 37292 25362 37320 25638
rect 37280 25356 37332 25362
rect 37280 25298 37332 25304
rect 37278 25256 37334 25265
rect 37278 25191 37334 25200
rect 37292 25158 37320 25191
rect 37280 25152 37332 25158
rect 37280 25094 37332 25100
rect 37384 24750 37412 25842
rect 37372 24744 37424 24750
rect 37372 24686 37424 24692
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37292 24206 37320 24550
rect 37096 24200 37148 24206
rect 37096 24142 37148 24148
rect 37280 24200 37332 24206
rect 37280 24142 37332 24148
rect 37476 24070 37504 26318
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37568 25294 37596 25774
rect 37648 25424 37700 25430
rect 37648 25366 37700 25372
rect 37740 25424 37792 25430
rect 37740 25366 37792 25372
rect 37556 25288 37608 25294
rect 37556 25230 37608 25236
rect 37568 24206 37596 25230
rect 37660 24750 37688 25366
rect 37752 25158 37780 25366
rect 37740 25152 37792 25158
rect 37740 25094 37792 25100
rect 37740 24880 37792 24886
rect 37740 24822 37792 24828
rect 37648 24744 37700 24750
rect 37648 24686 37700 24692
rect 37556 24200 37608 24206
rect 37556 24142 37608 24148
rect 37464 24064 37516 24070
rect 37464 24006 37516 24012
rect 37004 23044 37056 23050
rect 37004 22986 37056 22992
rect 37280 22636 37332 22642
rect 37280 22578 37332 22584
rect 36912 22568 36964 22574
rect 36912 22510 36964 22516
rect 36924 21418 36952 22510
rect 37292 21486 37320 22578
rect 37280 21480 37332 21486
rect 37332 21440 37412 21468
rect 37280 21422 37332 21428
rect 36912 21412 36964 21418
rect 36912 21354 36964 21360
rect 36728 21072 36780 21078
rect 36728 21014 36780 21020
rect 37280 21072 37332 21078
rect 37280 21014 37332 21020
rect 36740 20534 36768 21014
rect 36728 20528 36780 20534
rect 36728 20470 36780 20476
rect 36728 19372 36780 19378
rect 37292 19334 37320 21014
rect 37384 20398 37412 21440
rect 37476 20534 37504 24006
rect 37752 23798 37780 24822
rect 37832 24744 37884 24750
rect 37832 24686 37884 24692
rect 37844 24410 37872 24686
rect 37832 24404 37884 24410
rect 37832 24346 37884 24352
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37924 23520 37976 23526
rect 37924 23462 37976 23468
rect 37936 23118 37964 23462
rect 37924 23112 37976 23118
rect 37924 23054 37976 23060
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37568 22234 37596 22578
rect 37556 22228 37608 22234
rect 37556 22170 37608 22176
rect 38028 22030 38056 26318
rect 38120 26314 38148 27338
rect 38108 26308 38160 26314
rect 38108 26250 38160 26256
rect 38108 25832 38160 25838
rect 38108 25774 38160 25780
rect 38016 22024 38068 22030
rect 38016 21966 38068 21972
rect 37648 21888 37700 21894
rect 37648 21830 37700 21836
rect 37556 21480 37608 21486
rect 37556 21422 37608 21428
rect 37568 21146 37596 21422
rect 37556 21140 37608 21146
rect 37556 21082 37608 21088
rect 37660 21010 37688 21830
rect 37924 21480 37976 21486
rect 37924 21422 37976 21428
rect 37936 21350 37964 21422
rect 37924 21344 37976 21350
rect 37924 21286 37976 21292
rect 37648 21004 37700 21010
rect 37648 20946 37700 20952
rect 38016 20868 38068 20874
rect 38016 20810 38068 20816
rect 38028 20777 38056 20810
rect 38014 20768 38070 20777
rect 38014 20703 38070 20712
rect 37464 20528 37516 20534
rect 37464 20470 37516 20476
rect 37832 20528 37884 20534
rect 37832 20470 37884 20476
rect 37372 20392 37424 20398
rect 37372 20334 37424 20340
rect 37384 19922 37412 20334
rect 37476 20058 37504 20470
rect 37740 20392 37792 20398
rect 37740 20334 37792 20340
rect 37464 20052 37516 20058
rect 37464 19994 37516 20000
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 36728 19314 36780 19320
rect 36544 17332 36596 17338
rect 36544 17274 36596 17280
rect 36636 17332 36688 17338
rect 36636 17274 36688 17280
rect 36648 16794 36676 17274
rect 36636 16788 36688 16794
rect 36636 16730 36688 16736
rect 36452 16720 36504 16726
rect 36452 16662 36504 16668
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 36372 16250 36400 16526
rect 36360 16244 36412 16250
rect 36360 16186 36412 16192
rect 36544 15156 36596 15162
rect 36544 15098 36596 15104
rect 36452 14952 36504 14958
rect 36452 14894 36504 14900
rect 36268 14612 36320 14618
rect 36268 14554 36320 14560
rect 36360 14476 36412 14482
rect 36360 14418 36412 14424
rect 36268 14272 36320 14278
rect 36268 14214 36320 14220
rect 36176 13524 36228 13530
rect 36176 13466 36228 13472
rect 36280 13394 36308 14214
rect 36372 13433 36400 14418
rect 36464 14414 36492 14894
rect 36452 14408 36504 14414
rect 36452 14350 36504 14356
rect 36358 13424 36414 13433
rect 36268 13388 36320 13394
rect 36358 13359 36414 13368
rect 36268 13330 36320 13336
rect 35990 13288 36046 13297
rect 34978 13223 35034 13232
rect 35532 13252 35584 13258
rect 35990 13223 36046 13232
rect 35532 13194 35584 13200
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35164 12980 35216 12986
rect 35164 12922 35216 12928
rect 35176 12889 35204 12922
rect 35162 12880 35218 12889
rect 35162 12815 35218 12824
rect 35346 12880 35402 12889
rect 35346 12815 35402 12824
rect 35532 12844 35584 12850
rect 34704 12708 34756 12714
rect 34704 12650 34756 12656
rect 34716 12434 34744 12650
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34716 12406 34928 12434
rect 34704 12232 34756 12238
rect 34704 12174 34756 12180
rect 34520 12164 34572 12170
rect 34520 12106 34572 12112
rect 34336 11824 34388 11830
rect 34336 11766 34388 11772
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 32864 11620 32916 11626
rect 32864 11562 32916 11568
rect 33980 11354 34008 11698
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 33968 11348 34020 11354
rect 33968 11290 34020 11296
rect 33600 11280 33652 11286
rect 33600 11222 33652 11228
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32496 11212 32548 11218
rect 32496 11154 32548 11160
rect 32404 10600 32456 10606
rect 32404 10542 32456 10548
rect 32416 10266 32444 10542
rect 32404 10260 32456 10266
rect 32404 10202 32456 10208
rect 32508 10062 32536 11154
rect 32588 10464 32640 10470
rect 32588 10406 32640 10412
rect 32496 10056 32548 10062
rect 32496 9998 32548 10004
rect 32312 9920 32364 9926
rect 32312 9862 32364 9868
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31944 8288 31996 8294
rect 31944 8230 31996 8236
rect 31956 7954 31984 8230
rect 31852 7948 31904 7954
rect 31852 7890 31904 7896
rect 31944 7948 31996 7954
rect 31944 7890 31996 7896
rect 32324 7800 32352 9862
rect 32508 9518 32536 9998
rect 32496 9512 32548 9518
rect 32496 9454 32548 9460
rect 32600 7954 32628 10406
rect 33324 10056 33376 10062
rect 33324 9998 33376 10004
rect 32772 9988 32824 9994
rect 32772 9930 32824 9936
rect 32784 8378 32812 9930
rect 33336 9586 33364 9998
rect 33140 9580 33192 9586
rect 33140 9522 33192 9528
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 33152 9450 33180 9522
rect 33244 9466 33272 9522
rect 33612 9466 33640 11222
rect 34348 11218 34376 11766
rect 34532 11694 34560 12106
rect 34612 11892 34664 11898
rect 34612 11834 34664 11840
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 34428 11552 34480 11558
rect 34428 11494 34480 11500
rect 34336 11212 34388 11218
rect 34336 11154 34388 11160
rect 34244 11144 34296 11150
rect 34244 11086 34296 11092
rect 34256 11014 34284 11086
rect 34440 11082 34468 11494
rect 34520 11144 34572 11150
rect 34520 11086 34572 11092
rect 34428 11076 34480 11082
rect 34428 11018 34480 11024
rect 34244 11008 34296 11014
rect 34244 10950 34296 10956
rect 34152 10736 34204 10742
rect 34150 10704 34152 10713
rect 34204 10704 34206 10713
rect 34150 10639 34206 10648
rect 33876 10464 33928 10470
rect 33876 10406 33928 10412
rect 34152 10464 34204 10470
rect 34152 10406 34204 10412
rect 33888 10130 33916 10406
rect 33784 10124 33836 10130
rect 33784 10066 33836 10072
rect 33876 10124 33928 10130
rect 33876 10066 33928 10072
rect 33140 9444 33192 9450
rect 33140 9386 33192 9392
rect 33244 9438 33640 9466
rect 33152 9178 33180 9386
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 32956 9104 33008 9110
rect 32956 9046 33008 9052
rect 32864 8968 32916 8974
rect 32864 8910 32916 8916
rect 32876 8634 32904 8910
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 32968 8566 32996 9046
rect 33048 9036 33100 9042
rect 33048 8978 33100 8984
rect 32956 8560 33008 8566
rect 32956 8502 33008 8508
rect 32956 8424 33008 8430
rect 32784 8372 32956 8378
rect 32784 8366 33008 8372
rect 33060 8378 33088 8978
rect 33140 8492 33192 8498
rect 33244 8480 33272 9438
rect 33324 9172 33376 9178
rect 33324 9114 33376 9120
rect 33336 8498 33364 9114
rect 33612 9110 33640 9438
rect 33600 9104 33652 9110
rect 33600 9046 33652 9052
rect 33796 9058 33824 10066
rect 33876 9988 33928 9994
rect 33876 9930 33928 9936
rect 33888 9722 33916 9930
rect 34164 9926 34192 10406
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 33876 9716 33928 9722
rect 33876 9658 33928 9664
rect 33888 9518 33916 9658
rect 34164 9654 34192 9862
rect 34152 9648 34204 9654
rect 34152 9590 34204 9596
rect 34060 9580 34112 9586
rect 34060 9522 34112 9528
rect 33876 9512 33928 9518
rect 33876 9454 33928 9460
rect 33888 9178 33916 9454
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 33968 9172 34020 9178
rect 33968 9114 34020 9120
rect 33980 9058 34008 9114
rect 33796 9030 34008 9058
rect 33980 8566 34008 9030
rect 33968 8560 34020 8566
rect 33968 8502 34020 8508
rect 33192 8452 33272 8480
rect 33324 8492 33376 8498
rect 33140 8434 33192 8440
rect 33324 8434 33376 8440
rect 32784 8350 32996 8366
rect 33060 8350 33180 8378
rect 34072 8362 34100 9522
rect 34164 9382 34192 9590
rect 34152 9376 34204 9382
rect 34152 9318 34204 9324
rect 34256 9330 34284 10950
rect 34532 10810 34560 11086
rect 34520 10804 34572 10810
rect 34520 10746 34572 10752
rect 34624 10554 34652 11834
rect 34716 11354 34744 12174
rect 34796 12096 34848 12102
rect 34796 12038 34848 12044
rect 34808 11830 34836 12038
rect 34796 11824 34848 11830
rect 34796 11766 34848 11772
rect 34900 11676 34928 12406
rect 35360 12288 35388 12815
rect 35532 12786 35584 12792
rect 35900 12844 35952 12850
rect 35900 12786 35952 12792
rect 35440 12436 35492 12442
rect 35440 12378 35492 12384
rect 35268 12260 35388 12288
rect 35268 11694 35296 12260
rect 35348 12164 35400 12170
rect 35348 12106 35400 12112
rect 34808 11648 34928 11676
rect 35256 11688 35308 11694
rect 34704 11348 34756 11354
rect 34704 11290 34756 11296
rect 34808 11150 34836 11648
rect 35256 11630 35308 11636
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 35360 10742 35388 12106
rect 34980 10736 35032 10742
rect 34978 10704 34980 10713
rect 35348 10736 35400 10742
rect 35032 10704 35034 10713
rect 35348 10678 35400 10684
rect 34978 10639 35034 10648
rect 34796 10600 34848 10606
rect 34624 10526 34744 10554
rect 34796 10542 34848 10548
rect 34716 10470 34744 10526
rect 34704 10464 34756 10470
rect 34704 10406 34756 10412
rect 34704 10192 34756 10198
rect 34704 10134 34756 10140
rect 34336 9988 34388 9994
rect 34336 9930 34388 9936
rect 34348 9654 34376 9930
rect 34716 9654 34744 10134
rect 34336 9648 34388 9654
rect 34336 9590 34388 9596
rect 34704 9648 34756 9654
rect 34704 9590 34756 9596
rect 34808 9586 34836 10542
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 35348 9444 35400 9450
rect 35348 9386 35400 9392
rect 34520 9376 34572 9382
rect 34256 9324 34520 9330
rect 34256 9318 34572 9324
rect 34256 9302 34560 9318
rect 34256 8498 34284 9302
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34612 9172 34664 9178
rect 34612 9114 34664 9120
rect 35256 9172 35308 9178
rect 35256 9114 35308 9120
rect 34336 8968 34388 8974
rect 34336 8910 34388 8916
rect 34348 8634 34376 8910
rect 34624 8906 34652 9114
rect 34612 8900 34664 8906
rect 34612 8842 34664 8848
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34704 8832 34756 8838
rect 34704 8774 34756 8780
rect 35164 8832 35216 8838
rect 35164 8774 35216 8780
rect 34440 8634 34468 8774
rect 34336 8628 34388 8634
rect 34336 8570 34388 8576
rect 34428 8628 34480 8634
rect 34428 8570 34480 8576
rect 34244 8492 34296 8498
rect 34244 8434 34296 8440
rect 32968 8090 32996 8350
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 32496 7812 32548 7818
rect 32324 7772 32496 7800
rect 32496 7754 32548 7760
rect 31576 7744 31628 7750
rect 31576 7686 31628 7692
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 32508 7206 32536 7754
rect 33152 7750 33180 8350
rect 34060 8356 34112 8362
rect 34060 8298 34112 8304
rect 33232 8288 33284 8294
rect 33232 8230 33284 8236
rect 33244 7818 33272 8230
rect 33232 7812 33284 7818
rect 33232 7754 33284 7760
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 33152 7478 33180 7686
rect 34072 7546 34100 8298
rect 34060 7540 34112 7546
rect 34060 7482 34112 7488
rect 34716 7478 34744 8774
rect 35176 8498 35204 8774
rect 35164 8492 35216 8498
rect 35164 8434 35216 8440
rect 34796 8424 34848 8430
rect 34796 8366 34848 8372
rect 34808 8090 34836 8366
rect 35268 8276 35296 9114
rect 35360 8974 35388 9386
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 35360 8378 35388 8910
rect 35452 8566 35480 12378
rect 35544 12102 35572 12786
rect 35912 12442 35940 12786
rect 35900 12436 35952 12442
rect 35900 12378 35952 12384
rect 35532 12096 35584 12102
rect 35532 12038 35584 12044
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35532 11688 35584 11694
rect 35532 11630 35584 11636
rect 35544 11218 35572 11630
rect 36004 11354 36032 13223
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 36084 12912 36136 12918
rect 36084 12854 36136 12860
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 35532 11212 35584 11218
rect 35532 11154 35584 11160
rect 35992 11008 36044 11014
rect 35992 10950 36044 10956
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 36004 10742 36032 10950
rect 35992 10736 36044 10742
rect 35992 10678 36044 10684
rect 36096 10656 36124 12854
rect 36176 12096 36228 12102
rect 36176 12038 36228 12044
rect 36188 11898 36216 12038
rect 36176 11892 36228 11898
rect 36176 11834 36228 11840
rect 36188 10810 36216 11834
rect 36280 11354 36308 13126
rect 36556 12918 36584 15098
rect 36740 14414 36768 19314
rect 37108 19306 37320 19334
rect 37108 17134 37136 19306
rect 37556 19304 37608 19310
rect 37556 19246 37608 19252
rect 37188 19168 37240 19174
rect 37188 19110 37240 19116
rect 37280 19168 37332 19174
rect 37280 19110 37332 19116
rect 37200 18766 37228 19110
rect 37292 18834 37320 19110
rect 37568 18834 37596 19246
rect 37648 18896 37700 18902
rect 37648 18838 37700 18844
rect 37280 18828 37332 18834
rect 37280 18770 37332 18776
rect 37556 18828 37608 18834
rect 37556 18770 37608 18776
rect 37188 18760 37240 18766
rect 37188 18702 37240 18708
rect 37200 17814 37228 18702
rect 37556 18692 37608 18698
rect 37556 18634 37608 18640
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 37476 18358 37504 18566
rect 37464 18352 37516 18358
rect 37464 18294 37516 18300
rect 37280 18216 37332 18222
rect 37280 18158 37332 18164
rect 37292 17882 37320 18158
rect 37568 17882 37596 18634
rect 37280 17876 37332 17882
rect 37280 17818 37332 17824
rect 37556 17876 37608 17882
rect 37556 17818 37608 17824
rect 37188 17808 37240 17814
rect 37188 17750 37240 17756
rect 37660 17678 37688 18838
rect 37752 18426 37780 20334
rect 37844 19786 37872 20470
rect 38120 20398 38148 25774
rect 38212 23866 38240 29582
rect 38304 27538 38332 29786
rect 38396 29646 38424 30058
rect 38384 29640 38436 29646
rect 38384 29582 38436 29588
rect 38396 29209 38424 29582
rect 38382 29200 38438 29209
rect 38382 29135 38438 29144
rect 38292 27532 38344 27538
rect 38292 27474 38344 27480
rect 38304 26926 38332 27474
rect 38292 26920 38344 26926
rect 38292 26862 38344 26868
rect 38396 26314 38424 29135
rect 38488 27334 38516 31726
rect 38568 30388 38620 30394
rect 38568 30330 38620 30336
rect 38580 30258 38608 30330
rect 38568 30252 38620 30258
rect 38568 30194 38620 30200
rect 38476 27328 38528 27334
rect 38476 27270 38528 27276
rect 38384 26308 38436 26314
rect 38384 26250 38436 26256
rect 38488 25770 38516 27270
rect 38580 25838 38608 30194
rect 38660 29708 38712 29714
rect 38660 29650 38712 29656
rect 38672 27062 38700 29650
rect 38764 27577 38792 32966
rect 38844 32836 38896 32842
rect 38844 32778 38896 32784
rect 38856 30326 38884 32778
rect 38948 32570 38976 33866
rect 39028 33448 39080 33454
rect 39028 33390 39080 33396
rect 38936 32564 38988 32570
rect 38936 32506 38988 32512
rect 39040 31890 39068 33390
rect 39132 33386 39160 35702
rect 39224 35154 39252 36110
rect 40052 36106 40080 36518
rect 40132 36236 40184 36242
rect 40132 36178 40184 36184
rect 40040 36100 40092 36106
rect 40040 36042 40092 36048
rect 39304 36032 39356 36038
rect 39304 35974 39356 35980
rect 39316 35698 39344 35974
rect 39304 35692 39356 35698
rect 39304 35634 39356 35640
rect 40144 35630 40172 36178
rect 40420 35834 40448 37130
rect 40512 36786 40540 37130
rect 40500 36780 40552 36786
rect 40500 36722 40552 36728
rect 40604 35834 40632 38218
rect 40788 37874 40816 39442
rect 41064 39098 41092 40326
rect 41420 40044 41472 40050
rect 41420 39986 41472 39992
rect 41432 39370 41460 39986
rect 41788 39840 41840 39846
rect 41788 39782 41840 39788
rect 41420 39364 41472 39370
rect 41472 39324 41552 39352
rect 41420 39306 41472 39312
rect 41052 39092 41104 39098
rect 41052 39034 41104 39040
rect 41144 38888 41196 38894
rect 41144 38830 41196 38836
rect 41052 38820 41104 38826
rect 41052 38762 41104 38768
rect 40868 38752 40920 38758
rect 40868 38694 40920 38700
rect 40880 38350 40908 38694
rect 41064 38418 41092 38762
rect 41052 38412 41104 38418
rect 41052 38354 41104 38360
rect 40868 38344 40920 38350
rect 40868 38286 40920 38292
rect 40960 38208 41012 38214
rect 40960 38150 41012 38156
rect 40684 37868 40736 37874
rect 40684 37810 40736 37816
rect 40776 37868 40828 37874
rect 40776 37810 40828 37816
rect 40696 37126 40724 37810
rect 40788 37330 40816 37810
rect 40776 37324 40828 37330
rect 40776 37266 40828 37272
rect 40684 37120 40736 37126
rect 40684 37062 40736 37068
rect 40788 36922 40816 37266
rect 40776 36916 40828 36922
rect 40776 36858 40828 36864
rect 40408 35828 40460 35834
rect 40408 35770 40460 35776
rect 40592 35828 40644 35834
rect 40592 35770 40644 35776
rect 40132 35624 40184 35630
rect 40132 35566 40184 35572
rect 40408 35624 40460 35630
rect 40408 35566 40460 35572
rect 40420 35290 40448 35566
rect 40408 35284 40460 35290
rect 40408 35226 40460 35232
rect 39212 35148 39264 35154
rect 39212 35090 39264 35096
rect 40040 35148 40092 35154
rect 40040 35090 40092 35096
rect 39224 34746 39252 35090
rect 40052 34950 40080 35090
rect 40776 35012 40828 35018
rect 40776 34954 40828 34960
rect 40040 34944 40092 34950
rect 40040 34886 40092 34892
rect 39212 34740 39264 34746
rect 39212 34682 39264 34688
rect 39948 34604 40000 34610
rect 39948 34546 40000 34552
rect 39580 33924 39632 33930
rect 39580 33866 39632 33872
rect 39592 33658 39620 33866
rect 39672 33856 39724 33862
rect 39672 33798 39724 33804
rect 39580 33652 39632 33658
rect 39580 33594 39632 33600
rect 39684 33590 39712 33798
rect 39960 33658 39988 34546
rect 40052 33998 40080 34886
rect 40788 34746 40816 34954
rect 40972 34746 41000 38150
rect 41064 35630 41092 38354
rect 41156 35834 41184 38830
rect 41524 37738 41552 39324
rect 41800 38962 41828 39782
rect 42168 39642 42196 40462
rect 42156 39636 42208 39642
rect 42156 39578 42208 39584
rect 41788 38956 41840 38962
rect 41788 38898 41840 38904
rect 41880 38344 41932 38350
rect 41880 38286 41932 38292
rect 41696 37868 41748 37874
rect 41696 37810 41748 37816
rect 41512 37732 41564 37738
rect 41512 37674 41564 37680
rect 41328 36916 41380 36922
rect 41328 36858 41380 36864
rect 41340 36242 41368 36858
rect 41524 36718 41552 37674
rect 41512 36712 41564 36718
rect 41512 36654 41564 36660
rect 41604 36712 41656 36718
rect 41604 36654 41656 36660
rect 41616 36378 41644 36654
rect 41604 36372 41656 36378
rect 41604 36314 41656 36320
rect 41328 36236 41380 36242
rect 41328 36178 41380 36184
rect 41236 36032 41288 36038
rect 41236 35974 41288 35980
rect 41144 35828 41196 35834
rect 41144 35770 41196 35776
rect 41052 35624 41104 35630
rect 41052 35566 41104 35572
rect 41144 35556 41196 35562
rect 41144 35498 41196 35504
rect 41156 35154 41184 35498
rect 41248 35290 41276 35974
rect 41236 35284 41288 35290
rect 41236 35226 41288 35232
rect 41144 35148 41196 35154
rect 41144 35090 41196 35096
rect 40776 34740 40828 34746
rect 40776 34682 40828 34688
rect 40960 34740 41012 34746
rect 40960 34682 41012 34688
rect 40408 34604 40460 34610
rect 40408 34546 40460 34552
rect 40420 34066 40448 34546
rect 40788 34202 40816 34682
rect 41156 34542 41184 35090
rect 41236 34944 41288 34950
rect 41236 34886 41288 34892
rect 41144 34536 41196 34542
rect 41144 34478 41196 34484
rect 40776 34196 40828 34202
rect 40776 34138 40828 34144
rect 40408 34060 40460 34066
rect 40408 34002 40460 34008
rect 40040 33992 40092 33998
rect 40040 33934 40092 33940
rect 39948 33652 40000 33658
rect 39948 33594 40000 33600
rect 39304 33584 39356 33590
rect 39304 33526 39356 33532
rect 39672 33584 39724 33590
rect 39672 33526 39724 33532
rect 39120 33380 39172 33386
rect 39120 33322 39172 33328
rect 39028 31884 39080 31890
rect 39028 31826 39080 31832
rect 38936 30660 38988 30666
rect 38936 30602 38988 30608
rect 38844 30320 38896 30326
rect 38844 30262 38896 30268
rect 38856 29578 38884 30262
rect 38844 29572 38896 29578
rect 38844 29514 38896 29520
rect 38856 29306 38884 29514
rect 38844 29300 38896 29306
rect 38844 29242 38896 29248
rect 38856 28626 38884 29242
rect 38844 28620 38896 28626
rect 38844 28562 38896 28568
rect 38948 28490 38976 30602
rect 39212 30252 39264 30258
rect 39212 30194 39264 30200
rect 39224 29238 39252 30194
rect 39316 29714 39344 33526
rect 40052 33454 40080 33934
rect 40868 33924 40920 33930
rect 40868 33866 40920 33872
rect 40408 33856 40460 33862
rect 40408 33798 40460 33804
rect 40420 33658 40448 33798
rect 40880 33658 40908 33866
rect 40408 33652 40460 33658
rect 40408 33594 40460 33600
rect 40868 33652 40920 33658
rect 40868 33594 40920 33600
rect 40316 33516 40368 33522
rect 40316 33458 40368 33464
rect 40040 33448 40092 33454
rect 40040 33390 40092 33396
rect 40132 31340 40184 31346
rect 40132 31282 40184 31288
rect 40040 30660 40092 30666
rect 40040 30602 40092 30608
rect 39672 30592 39724 30598
rect 39672 30534 39724 30540
rect 39580 30320 39632 30326
rect 39580 30262 39632 30268
rect 39304 29708 39356 29714
rect 39304 29650 39356 29656
rect 39212 29232 39264 29238
rect 39212 29174 39264 29180
rect 39592 29170 39620 30262
rect 39684 30258 39712 30534
rect 39672 30252 39724 30258
rect 39672 30194 39724 30200
rect 39120 29164 39172 29170
rect 39120 29106 39172 29112
rect 39580 29164 39632 29170
rect 39580 29106 39632 29112
rect 39028 29028 39080 29034
rect 39028 28970 39080 28976
rect 38936 28484 38988 28490
rect 38936 28426 38988 28432
rect 38936 28076 38988 28082
rect 38936 28018 38988 28024
rect 38948 27985 38976 28018
rect 38934 27976 38990 27985
rect 38934 27911 38990 27920
rect 39040 27878 39068 28970
rect 39132 28948 39160 29106
rect 39132 28920 39344 28948
rect 39120 28620 39172 28626
rect 39120 28562 39172 28568
rect 39132 28422 39160 28562
rect 39120 28416 39172 28422
rect 39120 28358 39172 28364
rect 39028 27872 39080 27878
rect 39028 27814 39080 27820
rect 38750 27568 38806 27577
rect 38750 27503 38806 27512
rect 38936 27532 38988 27538
rect 38936 27474 38988 27480
rect 38948 27418 38976 27474
rect 38764 27390 38976 27418
rect 38764 27334 38792 27390
rect 38752 27328 38804 27334
rect 38752 27270 38804 27276
rect 38936 27328 38988 27334
rect 38936 27270 38988 27276
rect 38750 27160 38806 27169
rect 38750 27095 38806 27104
rect 38660 27056 38712 27062
rect 38660 26998 38712 27004
rect 38764 26382 38792 27095
rect 38948 26586 38976 27270
rect 38936 26580 38988 26586
rect 38936 26522 38988 26528
rect 38752 26376 38804 26382
rect 38752 26318 38804 26324
rect 39040 25906 39068 27814
rect 39132 27538 39160 28358
rect 39120 27532 39172 27538
rect 39120 27474 39172 27480
rect 39212 27396 39264 27402
rect 39212 27338 39264 27344
rect 39224 26042 39252 27338
rect 39212 26036 39264 26042
rect 39212 25978 39264 25984
rect 39316 25922 39344 28920
rect 39580 28484 39632 28490
rect 39580 28426 39632 28432
rect 39488 28144 39540 28150
rect 39488 28086 39540 28092
rect 39396 27328 39448 27334
rect 39396 27270 39448 27276
rect 39408 27062 39436 27270
rect 39396 27056 39448 27062
rect 39396 26998 39448 27004
rect 39500 25974 39528 28086
rect 39592 27062 39620 28426
rect 39580 27056 39632 27062
rect 39580 26998 39632 27004
rect 39028 25900 39080 25906
rect 39028 25842 39080 25848
rect 39224 25894 39344 25922
rect 39488 25968 39540 25974
rect 39488 25910 39540 25916
rect 38568 25832 38620 25838
rect 38568 25774 38620 25780
rect 38476 25764 38528 25770
rect 38476 25706 38528 25712
rect 38384 25356 38436 25362
rect 38384 25298 38436 25304
rect 38396 25265 38424 25298
rect 38382 25256 38438 25265
rect 38292 25220 38344 25226
rect 38382 25191 38438 25200
rect 38292 25162 38344 25168
rect 38304 24818 38332 25162
rect 38488 24970 38516 25706
rect 38488 24942 38608 24970
rect 38292 24812 38344 24818
rect 38292 24754 38344 24760
rect 38200 23860 38252 23866
rect 38200 23802 38252 23808
rect 38304 23730 38332 24754
rect 38488 24614 38516 24942
rect 38580 24886 38608 24942
rect 38568 24880 38620 24886
rect 38568 24822 38620 24828
rect 39040 24750 39068 25842
rect 39224 25498 39252 25894
rect 39212 25492 39264 25498
rect 39212 25434 39264 25440
rect 39028 24744 39080 24750
rect 39028 24686 39080 24692
rect 38476 24608 38528 24614
rect 38476 24550 38528 24556
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38304 23322 38332 23666
rect 38568 23656 38620 23662
rect 38568 23598 38620 23604
rect 38384 23588 38436 23594
rect 38384 23530 38436 23536
rect 38292 23316 38344 23322
rect 38292 23258 38344 23264
rect 38292 22092 38344 22098
rect 38292 22034 38344 22040
rect 38304 21486 38332 22034
rect 38292 21480 38344 21486
rect 38292 21422 38344 21428
rect 38108 20392 38160 20398
rect 38108 20334 38160 20340
rect 38120 19938 38148 20334
rect 38120 19922 38332 19938
rect 38120 19916 38344 19922
rect 38120 19910 38292 19916
rect 38292 19858 38344 19864
rect 38108 19848 38160 19854
rect 38108 19790 38160 19796
rect 37832 19780 37884 19786
rect 37832 19722 37884 19728
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 37648 17672 37700 17678
rect 37648 17614 37700 17620
rect 37752 17610 37780 18362
rect 37740 17604 37792 17610
rect 37740 17546 37792 17552
rect 37464 17536 37516 17542
rect 37464 17478 37516 17484
rect 37096 17128 37148 17134
rect 37096 17070 37148 17076
rect 37108 14464 37136 17070
rect 37476 16130 37504 17478
rect 37844 16522 37872 19722
rect 37924 19712 37976 19718
rect 37924 19654 37976 19660
rect 38016 19712 38068 19718
rect 38016 19654 38068 19660
rect 37936 19378 37964 19654
rect 37924 19372 37976 19378
rect 37924 19314 37976 19320
rect 37924 19168 37976 19174
rect 37924 19110 37976 19116
rect 37936 17746 37964 19110
rect 37924 17740 37976 17746
rect 37924 17682 37976 17688
rect 38028 17542 38056 19654
rect 38120 18290 38148 19790
rect 38292 19780 38344 19786
rect 38292 19722 38344 19728
rect 38304 19514 38332 19722
rect 38292 19508 38344 19514
rect 38292 19450 38344 19456
rect 38200 19168 38252 19174
rect 38200 19110 38252 19116
rect 38212 18834 38240 19110
rect 38200 18828 38252 18834
rect 38200 18770 38252 18776
rect 38396 18426 38424 23530
rect 38580 23168 38608 23598
rect 38660 23180 38712 23186
rect 38580 23140 38660 23168
rect 38580 22098 38608 23140
rect 38660 23122 38712 23128
rect 39028 22976 39080 22982
rect 39028 22918 39080 22924
rect 38660 22432 38712 22438
rect 38660 22374 38712 22380
rect 38672 22098 38700 22374
rect 38568 22092 38620 22098
rect 38568 22034 38620 22040
rect 38660 22092 38712 22098
rect 38660 22034 38712 22040
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38580 21010 38608 21286
rect 38568 21004 38620 21010
rect 38568 20946 38620 20952
rect 38476 20256 38528 20262
rect 38476 20198 38528 20204
rect 38384 18420 38436 18426
rect 38212 18380 38384 18408
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 38016 17536 38068 17542
rect 38016 17478 38068 17484
rect 38120 17270 38148 17614
rect 38108 17264 38160 17270
rect 38108 17206 38160 17212
rect 37832 16516 37884 16522
rect 37832 16458 37884 16464
rect 37740 16448 37792 16454
rect 37740 16390 37792 16396
rect 37384 16114 37504 16130
rect 37752 16114 37780 16390
rect 37844 16250 37872 16458
rect 38120 16454 38148 17206
rect 38108 16448 38160 16454
rect 38108 16390 38160 16396
rect 37832 16244 37884 16250
rect 37832 16186 37884 16192
rect 37384 16108 37516 16114
rect 37384 16102 37464 16108
rect 37188 15904 37240 15910
rect 37188 15846 37240 15852
rect 37200 15570 37228 15846
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37280 14952 37332 14958
rect 37280 14894 37332 14900
rect 37188 14476 37240 14482
rect 37108 14436 37188 14464
rect 36728 14408 36780 14414
rect 36728 14350 36780 14356
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 36636 13932 36688 13938
rect 36636 13874 36688 13880
rect 36648 13394 36676 13874
rect 36924 13530 36952 14214
rect 36912 13524 36964 13530
rect 36912 13466 36964 13472
rect 36636 13388 36688 13394
rect 36636 13330 36688 13336
rect 36544 12912 36596 12918
rect 36544 12854 36596 12860
rect 36544 12776 36596 12782
rect 36544 12718 36596 12724
rect 36556 12238 36584 12718
rect 36648 12714 36676 13330
rect 37004 13184 37056 13190
rect 37004 13126 37056 13132
rect 37016 12918 37044 13126
rect 37004 12912 37056 12918
rect 37108 12889 37136 14436
rect 37188 14418 37240 14424
rect 37292 14074 37320 14894
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 37188 12980 37240 12986
rect 37188 12922 37240 12928
rect 37004 12854 37056 12860
rect 37094 12880 37150 12889
rect 36636 12708 36688 12714
rect 36636 12650 36688 12656
rect 36544 12232 36596 12238
rect 36544 12174 36596 12180
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36360 11552 36412 11558
rect 36360 11494 36412 11500
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 36372 11218 36400 11494
rect 36360 11212 36412 11218
rect 36360 11154 36412 11160
rect 36176 10804 36228 10810
rect 36176 10746 36228 10752
rect 36464 10713 36492 11630
rect 37016 11218 37044 12854
rect 37094 12815 37150 12824
rect 37108 12306 37136 12815
rect 37096 12300 37148 12306
rect 37096 12242 37148 12248
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 37200 11150 37228 12922
rect 37384 12782 37412 16102
rect 37464 16050 37516 16056
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37740 16108 37792 16114
rect 37740 16050 37792 16056
rect 37464 15972 37516 15978
rect 37464 15914 37516 15920
rect 37476 15502 37504 15914
rect 37464 15496 37516 15502
rect 37464 15438 37516 15444
rect 37476 14414 37504 15438
rect 37660 14822 37688 16050
rect 37844 15434 37872 16186
rect 38120 15910 38148 16390
rect 38108 15904 38160 15910
rect 38108 15846 38160 15852
rect 37832 15428 37884 15434
rect 37832 15370 37884 15376
rect 37844 15094 37872 15370
rect 37832 15088 37884 15094
rect 37884 15036 37964 15042
rect 37832 15030 37964 15036
rect 37844 15014 37964 15030
rect 37832 14952 37884 14958
rect 37832 14894 37884 14900
rect 37648 14816 37700 14822
rect 37648 14758 37700 14764
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 37476 13870 37504 14350
rect 37844 14278 37872 14894
rect 37832 14272 37884 14278
rect 37832 14214 37884 14220
rect 37556 14068 37608 14074
rect 37556 14010 37608 14016
rect 37464 13864 37516 13870
rect 37464 13806 37516 13812
rect 37568 12850 37596 14010
rect 37936 14006 37964 15014
rect 38212 14482 38240 18380
rect 38384 18362 38436 18368
rect 38488 17202 38516 20198
rect 38580 19446 38608 20946
rect 38936 19848 38988 19854
rect 38936 19790 38988 19796
rect 38948 19514 38976 19790
rect 38936 19508 38988 19514
rect 38936 19450 38988 19456
rect 38568 19440 38620 19446
rect 38568 19382 38620 19388
rect 39040 18290 39068 22918
rect 39224 22094 39252 25434
rect 39592 25294 39620 26998
rect 39304 25288 39356 25294
rect 39304 25230 39356 25236
rect 39580 25288 39632 25294
rect 39580 25230 39632 25236
rect 39316 24886 39344 25230
rect 39580 25152 39632 25158
rect 39580 25094 39632 25100
rect 39592 24954 39620 25094
rect 39580 24948 39632 24954
rect 39580 24890 39632 24896
rect 39304 24880 39356 24886
rect 39304 24822 39356 24828
rect 39684 24698 39712 30194
rect 40052 30122 40080 30602
rect 40144 30326 40172 31282
rect 40328 30598 40356 33458
rect 40960 33448 41012 33454
rect 40960 33390 41012 33396
rect 40972 32978 41000 33390
rect 40960 32972 41012 32978
rect 40960 32914 41012 32920
rect 40592 32768 40644 32774
rect 40592 32710 40644 32716
rect 40604 32502 40632 32710
rect 40592 32496 40644 32502
rect 40592 32438 40644 32444
rect 40408 32428 40460 32434
rect 40408 32370 40460 32376
rect 40420 31822 40448 32370
rect 41248 31958 41276 34886
rect 41340 34746 41368 36178
rect 41708 35766 41736 37810
rect 41892 37126 41920 38286
rect 41880 37120 41932 37126
rect 41880 37062 41932 37068
rect 41696 35760 41748 35766
rect 41696 35702 41748 35708
rect 41420 35692 41472 35698
rect 41420 35634 41472 35640
rect 41432 34746 41460 35634
rect 41512 35624 41564 35630
rect 41512 35566 41564 35572
rect 41328 34740 41380 34746
rect 41328 34682 41380 34688
rect 41420 34740 41472 34746
rect 41420 34682 41472 34688
rect 41340 33998 41368 34682
rect 41328 33992 41380 33998
rect 41328 33934 41380 33940
rect 41432 32978 41460 34682
rect 41524 34678 41552 35566
rect 41512 34672 41564 34678
rect 41512 34614 41564 34620
rect 41420 32972 41472 32978
rect 41420 32914 41472 32920
rect 41432 32570 41460 32914
rect 41420 32564 41472 32570
rect 41420 32506 41472 32512
rect 41236 31952 41288 31958
rect 41236 31894 41288 31900
rect 40408 31816 40460 31822
rect 40408 31758 40460 31764
rect 40420 31346 40448 31758
rect 41708 31754 41736 35702
rect 41972 34604 42024 34610
rect 41972 34546 42024 34552
rect 41984 34202 42012 34546
rect 41972 34196 42024 34202
rect 41972 34138 42024 34144
rect 41972 32428 42024 32434
rect 41972 32370 42024 32376
rect 41708 31726 41828 31754
rect 41800 31346 41828 31726
rect 41984 31482 42012 32370
rect 42064 32224 42116 32230
rect 42064 32166 42116 32172
rect 41972 31476 42024 31482
rect 41972 31418 42024 31424
rect 42076 31385 42104 32166
rect 42062 31376 42118 31385
rect 40408 31340 40460 31346
rect 40408 31282 40460 31288
rect 41788 31340 41840 31346
rect 42062 31311 42118 31320
rect 41788 31282 41840 31288
rect 41052 31272 41104 31278
rect 41052 31214 41104 31220
rect 40868 31136 40920 31142
rect 40868 31078 40920 31084
rect 40408 30796 40460 30802
rect 40408 30738 40460 30744
rect 40316 30592 40368 30598
rect 40316 30534 40368 30540
rect 40132 30320 40184 30326
rect 40132 30262 40184 30268
rect 40224 30252 40276 30258
rect 40224 30194 40276 30200
rect 40040 30116 40092 30122
rect 40040 30058 40092 30064
rect 40236 29646 40264 30194
rect 40420 29850 40448 30738
rect 40880 30734 40908 31078
rect 41064 30938 41092 31214
rect 41052 30932 41104 30938
rect 41052 30874 41104 30880
rect 40868 30728 40920 30734
rect 40868 30670 40920 30676
rect 40592 30592 40644 30598
rect 40592 30534 40644 30540
rect 40498 30288 40554 30297
rect 40498 30223 40500 30232
rect 40552 30223 40554 30232
rect 40500 30194 40552 30200
rect 40408 29844 40460 29850
rect 40408 29786 40460 29792
rect 40224 29640 40276 29646
rect 40408 29640 40460 29646
rect 40276 29588 40356 29594
rect 40224 29582 40356 29588
rect 40408 29582 40460 29588
rect 40040 29572 40092 29578
rect 40236 29566 40356 29582
rect 40040 29514 40092 29520
rect 40052 29306 40080 29514
rect 40224 29504 40276 29510
rect 40224 29446 40276 29452
rect 40040 29300 40092 29306
rect 40040 29242 40092 29248
rect 40236 29238 40264 29446
rect 39856 29232 39908 29238
rect 40224 29232 40276 29238
rect 39908 29180 39988 29186
rect 39856 29174 39988 29180
rect 40224 29174 40276 29180
rect 39868 29158 39988 29174
rect 39960 29102 39988 29158
rect 39948 29096 40000 29102
rect 39948 29038 40000 29044
rect 40038 28928 40094 28937
rect 40038 28863 40094 28872
rect 39856 28484 39908 28490
rect 39856 28426 39908 28432
rect 39764 28416 39816 28422
rect 39764 28358 39816 28364
rect 39776 28082 39804 28358
rect 39764 28076 39816 28082
rect 39764 28018 39816 28024
rect 39868 27606 39896 28426
rect 40052 28150 40080 28863
rect 40040 28144 40092 28150
rect 40328 28098 40356 29566
rect 40420 28966 40448 29582
rect 40408 28960 40460 28966
rect 40408 28902 40460 28908
rect 40040 28086 40092 28092
rect 40236 28082 40356 28098
rect 40224 28076 40356 28082
rect 40276 28070 40356 28076
rect 40224 28018 40276 28024
rect 40236 27946 40264 28018
rect 40420 28014 40448 28902
rect 40500 28484 40552 28490
rect 40500 28426 40552 28432
rect 40512 28218 40540 28426
rect 40500 28212 40552 28218
rect 40500 28154 40552 28160
rect 40316 28008 40368 28014
rect 40316 27950 40368 27956
rect 40408 28008 40460 28014
rect 40408 27950 40460 27956
rect 40224 27940 40276 27946
rect 40224 27882 40276 27888
rect 39856 27600 39908 27606
rect 39856 27542 39908 27548
rect 40236 27334 40264 27882
rect 40328 27402 40356 27950
rect 40316 27396 40368 27402
rect 40316 27338 40368 27344
rect 40224 27328 40276 27334
rect 40144 27288 40224 27316
rect 40040 27124 40092 27130
rect 40040 27066 40092 27072
rect 39948 25288 40000 25294
rect 39948 25230 40000 25236
rect 39684 24670 39804 24698
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39408 23730 39436 24142
rect 39396 23724 39448 23730
rect 39396 23666 39448 23672
rect 39672 23724 39724 23730
rect 39672 23666 39724 23672
rect 39684 23322 39712 23666
rect 39672 23316 39724 23322
rect 39672 23258 39724 23264
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39224 22066 39344 22094
rect 39212 21412 39264 21418
rect 39212 21354 39264 21360
rect 39224 20874 39252 21354
rect 39212 20868 39264 20874
rect 39212 20810 39264 20816
rect 39224 20262 39252 20810
rect 39120 20256 39172 20262
rect 39120 20198 39172 20204
rect 39212 20256 39264 20262
rect 39212 20198 39264 20204
rect 39132 19922 39160 20198
rect 39120 19916 39172 19922
rect 39120 19858 39172 19864
rect 39224 19310 39252 20198
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 39224 18766 39252 19246
rect 39212 18760 39264 18766
rect 39212 18702 39264 18708
rect 39028 18284 39080 18290
rect 39028 18226 39080 18232
rect 38476 17196 38528 17202
rect 38476 17138 38528 17144
rect 38384 16992 38436 16998
rect 38384 16934 38436 16940
rect 38396 16658 38424 16934
rect 38384 16652 38436 16658
rect 38384 16594 38436 16600
rect 38292 16516 38344 16522
rect 38292 16458 38344 16464
rect 38304 16046 38332 16458
rect 38292 16040 38344 16046
rect 38292 15982 38344 15988
rect 38290 15464 38346 15473
rect 38290 15399 38292 15408
rect 38344 15399 38346 15408
rect 38292 15370 38344 15376
rect 38304 15162 38332 15370
rect 38488 15366 38516 17138
rect 38752 17128 38804 17134
rect 38752 17070 38804 17076
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38672 16182 38700 16934
rect 38764 16794 38792 17070
rect 38844 17060 38896 17066
rect 38844 17002 38896 17008
rect 38752 16788 38804 16794
rect 38752 16730 38804 16736
rect 38660 16176 38712 16182
rect 38660 16118 38712 16124
rect 38568 15496 38620 15502
rect 38568 15438 38620 15444
rect 38476 15360 38528 15366
rect 38476 15302 38528 15308
rect 38292 15156 38344 15162
rect 38292 15098 38344 15104
rect 38488 15042 38516 15302
rect 38580 15162 38608 15438
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 38488 15014 38700 15042
rect 38200 14476 38252 14482
rect 38200 14418 38252 14424
rect 38384 14408 38436 14414
rect 38384 14350 38436 14356
rect 37924 14000 37976 14006
rect 37924 13942 37976 13948
rect 38396 13870 38424 14350
rect 37832 13864 37884 13870
rect 37832 13806 37884 13812
rect 38384 13864 38436 13870
rect 38384 13806 38436 13812
rect 37844 13530 37872 13806
rect 37832 13524 37884 13530
rect 37832 13466 37884 13472
rect 38672 13462 38700 15014
rect 38660 13456 38712 13462
rect 38660 13398 38712 13404
rect 37924 13388 37976 13394
rect 37924 13330 37976 13336
rect 37936 12918 37964 13330
rect 37924 12912 37976 12918
rect 37924 12854 37976 12860
rect 38660 12912 38712 12918
rect 38660 12854 38712 12860
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37372 12776 37424 12782
rect 37372 12718 37424 12724
rect 37372 12640 37424 12646
rect 37372 12582 37424 12588
rect 37280 12232 37332 12238
rect 37280 12174 37332 12180
rect 37292 11898 37320 12174
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 36450 10704 36506 10713
rect 36176 10668 36228 10674
rect 36096 10628 36176 10656
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 36096 9722 36124 10628
rect 37002 10704 37058 10713
rect 36450 10639 36506 10648
rect 36912 10668 36964 10674
rect 36176 10610 36228 10616
rect 37002 10639 37058 10648
rect 36912 10610 36964 10616
rect 36924 10130 36952 10610
rect 36912 10124 36964 10130
rect 36912 10066 36964 10072
rect 36924 9722 36952 10066
rect 37016 9722 37044 10639
rect 36084 9716 36136 9722
rect 36084 9658 36136 9664
rect 36912 9716 36964 9722
rect 36912 9658 36964 9664
rect 37004 9716 37056 9722
rect 37004 9658 37056 9664
rect 35532 9580 35584 9586
rect 35532 9522 35584 9528
rect 35544 9466 35572 9522
rect 35716 9512 35768 9518
rect 35544 9460 35716 9466
rect 35544 9454 35768 9460
rect 35544 9438 35756 9454
rect 35544 9178 35572 9438
rect 35532 9172 35584 9178
rect 35532 9114 35584 9120
rect 35728 9042 35756 9438
rect 35716 9036 35768 9042
rect 35716 8978 35768 8984
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 36096 8480 36124 9658
rect 37292 9586 37320 11834
rect 37384 11354 37412 12582
rect 37568 12434 37596 12786
rect 37648 12776 37700 12782
rect 37648 12718 37700 12724
rect 37476 12406 37596 12434
rect 37372 11348 37424 11354
rect 37372 11290 37424 11296
rect 37476 11150 37504 12406
rect 37556 12164 37608 12170
rect 37556 12106 37608 12112
rect 37568 11626 37596 12106
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37660 11150 37688 12718
rect 37924 12708 37976 12714
rect 37924 12650 37976 12656
rect 37832 12640 37884 12646
rect 37832 12582 37884 12588
rect 37844 11762 37872 12582
rect 37936 11762 37964 12650
rect 38672 12186 38700 12854
rect 38856 12850 38884 17002
rect 39224 16658 39252 18702
rect 39212 16652 39264 16658
rect 39212 16594 39264 16600
rect 39316 14074 39344 22066
rect 39592 21690 39620 22578
rect 39776 21690 39804 24670
rect 39960 24206 39988 25230
rect 39948 24200 40000 24206
rect 39948 24142 40000 24148
rect 40052 23118 40080 27066
rect 40144 25838 40172 27288
rect 40224 27270 40276 27276
rect 40420 26926 40448 27950
rect 40408 26920 40460 26926
rect 40408 26862 40460 26868
rect 40224 26852 40276 26858
rect 40224 26794 40276 26800
rect 40236 25906 40264 26794
rect 40420 26314 40448 26862
rect 40408 26308 40460 26314
rect 40408 26250 40460 26256
rect 40224 25900 40276 25906
rect 40224 25842 40276 25848
rect 40420 25838 40448 26250
rect 40132 25832 40184 25838
rect 40132 25774 40184 25780
rect 40408 25832 40460 25838
rect 40408 25774 40460 25780
rect 40132 25696 40184 25702
rect 40132 25638 40184 25644
rect 40144 25265 40172 25638
rect 40420 25294 40448 25774
rect 40604 25514 40632 30534
rect 40868 30252 40920 30258
rect 40868 30194 40920 30200
rect 40684 30048 40736 30054
rect 40684 29990 40736 29996
rect 40696 29714 40724 29990
rect 40684 29708 40736 29714
rect 40684 29650 40736 29656
rect 40880 29617 40908 30194
rect 40866 29608 40922 29617
rect 40866 29543 40922 29552
rect 41420 29572 41472 29578
rect 41420 29514 41472 29520
rect 41432 28558 41460 29514
rect 41420 28552 41472 28558
rect 41420 28494 41472 28500
rect 40684 28416 40736 28422
rect 40684 28358 40736 28364
rect 40696 28150 40724 28358
rect 41432 28150 41460 28494
rect 41696 28416 41748 28422
rect 41696 28358 41748 28364
rect 40684 28144 40736 28150
rect 40684 28086 40736 28092
rect 41420 28144 41472 28150
rect 41420 28086 41472 28092
rect 40776 27464 40828 27470
rect 40776 27406 40828 27412
rect 40788 26790 40816 27406
rect 41052 27396 41104 27402
rect 41052 27338 41104 27344
rect 41064 26858 41092 27338
rect 41144 27328 41196 27334
rect 41144 27270 41196 27276
rect 41052 26852 41104 26858
rect 41052 26794 41104 26800
rect 40776 26784 40828 26790
rect 40776 26726 40828 26732
rect 41052 26512 41104 26518
rect 41052 26454 41104 26460
rect 40512 25498 40632 25514
rect 40500 25492 40632 25498
rect 40552 25486 40632 25492
rect 40500 25434 40552 25440
rect 40408 25288 40460 25294
rect 40130 25256 40186 25265
rect 40408 25230 40460 25236
rect 40130 25191 40186 25200
rect 40684 25220 40736 25226
rect 40684 25162 40736 25168
rect 40696 24954 40724 25162
rect 41064 24954 41092 26454
rect 41156 25838 41184 27270
rect 41236 26988 41288 26994
rect 41236 26930 41288 26936
rect 41144 25832 41196 25838
rect 41144 25774 41196 25780
rect 40684 24948 40736 24954
rect 40684 24890 40736 24896
rect 41052 24948 41104 24954
rect 41052 24890 41104 24896
rect 40592 24608 40644 24614
rect 40590 24576 40592 24585
rect 40644 24576 40646 24585
rect 40590 24511 40646 24520
rect 40960 24132 41012 24138
rect 40960 24074 41012 24080
rect 40972 23866 41000 24074
rect 40960 23860 41012 23866
rect 40960 23802 41012 23808
rect 40776 23520 40828 23526
rect 40776 23462 40828 23468
rect 40788 23186 40816 23462
rect 40776 23180 40828 23186
rect 40776 23122 40828 23128
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 41052 22976 41104 22982
rect 41052 22918 41104 22924
rect 41064 22778 41092 22918
rect 41052 22772 41104 22778
rect 41052 22714 41104 22720
rect 39856 22704 39908 22710
rect 39856 22646 39908 22652
rect 39868 22030 39896 22646
rect 40776 22568 40828 22574
rect 40776 22510 40828 22516
rect 40684 22432 40736 22438
rect 40684 22374 40736 22380
rect 39856 22024 39908 22030
rect 39856 21966 39908 21972
rect 40224 22024 40276 22030
rect 40224 21966 40276 21972
rect 39580 21684 39632 21690
rect 39580 21626 39632 21632
rect 39764 21684 39816 21690
rect 39764 21626 39816 21632
rect 40132 21548 40184 21554
rect 40132 21490 40184 21496
rect 40144 20806 40172 21490
rect 40236 21486 40264 21966
rect 40592 21956 40644 21962
rect 40592 21898 40644 21904
rect 40604 21622 40632 21898
rect 40592 21616 40644 21622
rect 40592 21558 40644 21564
rect 40224 21480 40276 21486
rect 40224 21422 40276 21428
rect 40592 21480 40644 21486
rect 40592 21422 40644 21428
rect 40604 21146 40632 21422
rect 40592 21140 40644 21146
rect 40592 21082 40644 21088
rect 40132 20800 40184 20806
rect 40132 20742 40184 20748
rect 40144 20534 40172 20742
rect 40132 20528 40184 20534
rect 40132 20470 40184 20476
rect 40696 20466 40724 22374
rect 40788 21894 40816 22510
rect 41144 22092 41196 22098
rect 41144 22034 41196 22040
rect 40776 21888 40828 21894
rect 40776 21830 40828 21836
rect 41156 21146 41184 22034
rect 41144 21140 41196 21146
rect 41144 21082 41196 21088
rect 40684 20460 40736 20466
rect 40684 20402 40736 20408
rect 39580 20392 39632 20398
rect 39580 20334 39632 20340
rect 40316 20392 40368 20398
rect 40316 20334 40368 20340
rect 39592 20058 39620 20334
rect 40040 20324 40092 20330
rect 40040 20266 40092 20272
rect 39580 20052 39632 20058
rect 39580 19994 39632 20000
rect 39396 19848 39448 19854
rect 39396 19790 39448 19796
rect 39408 19718 39436 19790
rect 39396 19712 39448 19718
rect 39396 19654 39448 19660
rect 39488 19712 39540 19718
rect 39488 19654 39540 19660
rect 39500 19446 39528 19654
rect 39488 19440 39540 19446
rect 39488 19382 39540 19388
rect 39764 18896 39816 18902
rect 39764 18838 39816 18844
rect 39776 18222 39804 18838
rect 40052 18290 40080 20266
rect 40224 19780 40276 19786
rect 40224 19722 40276 19728
rect 40132 19440 40184 19446
rect 40132 19382 40184 19388
rect 40144 19310 40172 19382
rect 40132 19304 40184 19310
rect 40132 19246 40184 19252
rect 40144 18630 40172 19246
rect 40132 18624 40184 18630
rect 40132 18566 40184 18572
rect 40040 18284 40092 18290
rect 40040 18226 40092 18232
rect 40236 18222 40264 19722
rect 40328 18834 40356 20334
rect 40592 19848 40644 19854
rect 40592 19790 40644 19796
rect 41144 19848 41196 19854
rect 41144 19790 41196 19796
rect 40316 18828 40368 18834
rect 40316 18770 40368 18776
rect 40328 18714 40356 18770
rect 40328 18686 40448 18714
rect 40316 18624 40368 18630
rect 40316 18566 40368 18572
rect 39764 18216 39816 18222
rect 39764 18158 39816 18164
rect 40224 18216 40276 18222
rect 40224 18158 40276 18164
rect 40132 18148 40184 18154
rect 40132 18090 40184 18096
rect 39856 17264 39908 17270
rect 39856 17206 39908 17212
rect 39868 16590 39896 17206
rect 40040 16720 40092 16726
rect 40040 16662 40092 16668
rect 39856 16584 39908 16590
rect 39856 16526 39908 16532
rect 40052 16250 40080 16662
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 40052 16046 40080 16186
rect 40144 16130 40172 18090
rect 40328 17270 40356 18566
rect 40420 18154 40448 18686
rect 40500 18352 40552 18358
rect 40500 18294 40552 18300
rect 40408 18148 40460 18154
rect 40408 18090 40460 18096
rect 40316 17264 40368 17270
rect 40316 17206 40368 17212
rect 40224 17196 40276 17202
rect 40224 17138 40276 17144
rect 40236 16590 40264 17138
rect 40328 16590 40356 17206
rect 40224 16584 40276 16590
rect 40224 16526 40276 16532
rect 40316 16584 40368 16590
rect 40316 16526 40368 16532
rect 40512 16130 40540 18294
rect 40604 17678 40632 19790
rect 41156 19514 41184 19790
rect 40776 19508 40828 19514
rect 40776 19450 40828 19456
rect 41144 19508 41196 19514
rect 41144 19450 41196 19456
rect 40788 18222 40816 19450
rect 41052 19168 41104 19174
rect 41052 19110 41104 19116
rect 41064 18834 41092 19110
rect 41052 18828 41104 18834
rect 41052 18770 41104 18776
rect 41156 18290 41184 19450
rect 41144 18284 41196 18290
rect 41144 18226 41196 18232
rect 40776 18216 40828 18222
rect 40776 18158 40828 18164
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40776 17536 40828 17542
rect 40776 17478 40828 17484
rect 40788 17270 40816 17478
rect 40776 17264 40828 17270
rect 40776 17206 40828 17212
rect 41248 17116 41276 26930
rect 41328 26444 41380 26450
rect 41328 26386 41380 26392
rect 41340 23866 41368 26386
rect 41432 25974 41460 28086
rect 41708 27985 41736 28358
rect 41694 27976 41750 27985
rect 41694 27911 41750 27920
rect 41604 27464 41656 27470
rect 41604 27406 41656 27412
rect 41512 27328 41564 27334
rect 41510 27296 41512 27305
rect 41564 27296 41566 27305
rect 41510 27231 41566 27240
rect 41512 26784 41564 26790
rect 41512 26726 41564 26732
rect 41420 25968 41472 25974
rect 41420 25910 41472 25916
rect 41432 25226 41460 25910
rect 41420 25220 41472 25226
rect 41420 25162 41472 25168
rect 41432 24886 41460 25162
rect 41420 24880 41472 24886
rect 41420 24822 41472 24828
rect 41432 24138 41460 24822
rect 41524 24818 41552 26726
rect 41616 26042 41644 27406
rect 41696 26852 41748 26858
rect 41800 26840 41828 31282
rect 41880 30252 41932 30258
rect 41880 30194 41932 30200
rect 41892 29850 41920 30194
rect 42064 30048 42116 30054
rect 42064 29990 42116 29996
rect 41880 29844 41932 29850
rect 41880 29786 41932 29792
rect 42076 29345 42104 29990
rect 42062 29336 42118 29345
rect 42062 29271 42118 29280
rect 41972 29232 42024 29238
rect 41972 29174 42024 29180
rect 41878 28656 41934 28665
rect 41878 28591 41934 28600
rect 41892 28558 41920 28591
rect 41880 28552 41932 28558
rect 41880 28494 41932 28500
rect 41880 27328 41932 27334
rect 41880 27270 41932 27276
rect 41748 26812 41828 26840
rect 41696 26794 41748 26800
rect 41604 26036 41656 26042
rect 41604 25978 41656 25984
rect 41708 25922 41736 26794
rect 41892 26625 41920 27270
rect 41878 26616 41934 26625
rect 41878 26551 41934 26560
rect 41616 25894 41736 25922
rect 41616 25158 41644 25894
rect 41604 25152 41656 25158
rect 41604 25094 41656 25100
rect 41512 24812 41564 24818
rect 41512 24754 41564 24760
rect 41512 24676 41564 24682
rect 41512 24618 41564 24624
rect 41420 24132 41472 24138
rect 41420 24074 41472 24080
rect 41328 23860 41380 23866
rect 41328 23802 41380 23808
rect 41524 23662 41552 24618
rect 41420 23656 41472 23662
rect 41420 23598 41472 23604
rect 41512 23656 41564 23662
rect 41512 23598 41564 23604
rect 41432 23322 41460 23598
rect 41420 23316 41472 23322
rect 41420 23258 41472 23264
rect 41616 22710 41644 25094
rect 41984 24818 42012 29174
rect 42064 29028 42116 29034
rect 42064 28970 42116 28976
rect 42076 28665 42104 28970
rect 42062 28656 42118 28665
rect 42062 28591 42118 28600
rect 42064 28416 42116 28422
rect 42064 28358 42116 28364
rect 42076 25945 42104 28358
rect 42156 26920 42208 26926
rect 42156 26862 42208 26868
rect 42062 25936 42118 25945
rect 42062 25871 42118 25880
rect 42064 25696 42116 25702
rect 42168 25650 42196 26862
rect 42116 25644 42196 25650
rect 42064 25638 42196 25644
rect 42076 25622 42196 25638
rect 42168 25498 42196 25622
rect 42156 25492 42208 25498
rect 42156 25434 42208 25440
rect 41972 24812 42024 24818
rect 41972 24754 42024 24760
rect 41696 24608 41748 24614
rect 41696 24550 41748 24556
rect 41708 24410 41736 24550
rect 41696 24404 41748 24410
rect 41696 24346 41748 24352
rect 41984 23050 42012 24754
rect 42064 24404 42116 24410
rect 42064 24346 42116 24352
rect 42076 23186 42104 24346
rect 42064 23180 42116 23186
rect 42064 23122 42116 23128
rect 41972 23044 42024 23050
rect 41972 22986 42024 22992
rect 41984 22778 42012 22986
rect 41972 22772 42024 22778
rect 41972 22714 42024 22720
rect 41604 22704 41656 22710
rect 41604 22646 41656 22652
rect 41696 22636 41748 22642
rect 41696 22578 41748 22584
rect 41512 22432 41564 22438
rect 41512 22374 41564 22380
rect 41420 21888 41472 21894
rect 41420 21830 41472 21836
rect 41328 21616 41380 21622
rect 41432 21570 41460 21830
rect 41380 21564 41460 21570
rect 41328 21558 41460 21564
rect 41340 21542 41460 21558
rect 41328 19984 41380 19990
rect 41328 19926 41380 19932
rect 41340 18358 41368 19926
rect 41432 19242 41460 21542
rect 41524 21010 41552 22374
rect 41708 22098 41736 22578
rect 41696 22092 41748 22098
rect 41696 22034 41748 22040
rect 41880 22092 41932 22098
rect 41880 22034 41932 22040
rect 41512 21004 41564 21010
rect 41512 20946 41564 20952
rect 41512 20868 41564 20874
rect 41512 20810 41564 20816
rect 41524 20602 41552 20810
rect 41512 20596 41564 20602
rect 41512 20538 41564 20544
rect 41696 20528 41748 20534
rect 41696 20470 41748 20476
rect 41512 19712 41564 19718
rect 41512 19654 41564 19660
rect 41420 19236 41472 19242
rect 41420 19178 41472 19184
rect 41432 18698 41460 19178
rect 41420 18692 41472 18698
rect 41420 18634 41472 18640
rect 41524 18358 41552 19654
rect 41708 19378 41736 20470
rect 41788 20460 41840 20466
rect 41788 20402 41840 20408
rect 41696 19372 41748 19378
rect 41696 19314 41748 19320
rect 41604 19304 41656 19310
rect 41604 19246 41656 19252
rect 41616 18426 41644 19246
rect 41604 18420 41656 18426
rect 41604 18362 41656 18368
rect 41328 18352 41380 18358
rect 41328 18294 41380 18300
rect 41512 18352 41564 18358
rect 41512 18294 41564 18300
rect 40788 17088 41276 17116
rect 40684 16516 40736 16522
rect 40684 16458 40736 16464
rect 40592 16448 40644 16454
rect 40592 16390 40644 16396
rect 40144 16114 40356 16130
rect 40420 16114 40540 16130
rect 40604 16114 40632 16390
rect 40696 16250 40724 16458
rect 40684 16244 40736 16250
rect 40684 16186 40736 16192
rect 40132 16108 40356 16114
rect 40184 16102 40356 16108
rect 40132 16050 40184 16056
rect 40040 16040 40092 16046
rect 40040 15982 40092 15988
rect 39764 15904 39816 15910
rect 39764 15846 39816 15852
rect 40224 15904 40276 15910
rect 40224 15846 40276 15852
rect 39304 14068 39356 14074
rect 39304 14010 39356 14016
rect 39316 13326 39344 14010
rect 39776 13394 39804 15846
rect 40236 15706 40264 15846
rect 40224 15700 40276 15706
rect 40224 15642 40276 15648
rect 40040 15156 40092 15162
rect 40040 15098 40092 15104
rect 39856 14884 39908 14890
rect 39856 14826 39908 14832
rect 39868 14414 39896 14826
rect 39856 14408 39908 14414
rect 40052 14362 40080 15098
rect 40236 15026 40264 15642
rect 40224 15020 40276 15026
rect 40224 14962 40276 14968
rect 40132 14952 40184 14958
rect 40132 14894 40184 14900
rect 40144 14618 40172 14894
rect 40132 14612 40184 14618
rect 40132 14554 40184 14560
rect 40236 14550 40264 14962
rect 40224 14544 40276 14550
rect 40224 14486 40276 14492
rect 39856 14350 39908 14356
rect 39960 14334 40080 14362
rect 39960 14278 39988 14334
rect 39948 14272 40000 14278
rect 39948 14214 40000 14220
rect 40040 14272 40092 14278
rect 40040 14214 40092 14220
rect 39948 13864 40000 13870
rect 39948 13806 40000 13812
rect 39960 13530 39988 13806
rect 39948 13524 40000 13530
rect 39948 13466 40000 13472
rect 39488 13388 39540 13394
rect 39488 13330 39540 13336
rect 39764 13388 39816 13394
rect 39764 13330 39816 13336
rect 39304 13320 39356 13326
rect 39304 13262 39356 13268
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 38856 12374 38884 12786
rect 38844 12368 38896 12374
rect 38844 12310 38896 12316
rect 39500 12238 39528 13330
rect 40052 13326 40080 14214
rect 40040 13320 40092 13326
rect 40040 13262 40092 13268
rect 39488 12232 39540 12238
rect 38672 12170 38884 12186
rect 39488 12174 39540 12180
rect 38672 12164 38896 12170
rect 38672 12158 38844 12164
rect 38844 12106 38896 12112
rect 38856 11830 38884 12106
rect 39488 12096 39540 12102
rect 39488 12038 39540 12044
rect 38844 11824 38896 11830
rect 38844 11766 38896 11772
rect 37832 11756 37884 11762
rect 37832 11698 37884 11704
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 37740 11688 37792 11694
rect 37740 11630 37792 11636
rect 37464 11144 37516 11150
rect 37464 11086 37516 11092
rect 37648 11144 37700 11150
rect 37648 11086 37700 11092
rect 37464 11008 37516 11014
rect 37464 10950 37516 10956
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 37384 10062 37412 10610
rect 37476 10062 37504 10950
rect 37556 10192 37608 10198
rect 37660 10180 37688 11086
rect 37752 11014 37780 11630
rect 37844 11354 37872 11698
rect 38200 11688 38252 11694
rect 38200 11630 38252 11636
rect 37832 11348 37884 11354
rect 37832 11290 37884 11296
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 37740 11008 37792 11014
rect 37740 10950 37792 10956
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 37936 10674 37964 10950
rect 38120 10810 38148 11154
rect 38108 10804 38160 10810
rect 38108 10746 38160 10752
rect 37740 10668 37792 10674
rect 37740 10610 37792 10616
rect 37924 10668 37976 10674
rect 37924 10610 37976 10616
rect 38016 10668 38068 10674
rect 38016 10610 38068 10616
rect 37752 10266 37780 10610
rect 37740 10260 37792 10266
rect 37740 10202 37792 10208
rect 37608 10152 37688 10180
rect 37556 10134 37608 10140
rect 37660 10062 37688 10152
rect 37372 10056 37424 10062
rect 37372 9998 37424 10004
rect 37464 10056 37516 10062
rect 37464 9998 37516 10004
rect 37648 10056 37700 10062
rect 37648 9998 37700 10004
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37372 9172 37424 9178
rect 37372 9114 37424 9120
rect 37384 9042 37412 9114
rect 37372 9036 37424 9042
rect 37372 8978 37424 8984
rect 37476 8922 37504 9998
rect 37556 9920 37608 9926
rect 37556 9862 37608 9868
rect 37648 9920 37700 9926
rect 37648 9862 37700 9868
rect 37568 9654 37596 9862
rect 37556 9648 37608 9654
rect 37556 9590 37608 9596
rect 37292 8906 37504 8922
rect 37280 8900 37504 8906
rect 37332 8894 37504 8900
rect 37280 8842 37332 8848
rect 36268 8492 36320 8498
rect 36096 8452 36268 8480
rect 36268 8434 36320 8440
rect 37476 8430 37504 8894
rect 37660 8838 37688 9862
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37648 8832 37700 8838
rect 37648 8774 37700 8780
rect 37740 8832 37792 8838
rect 37740 8774 37792 8780
rect 37660 8498 37688 8774
rect 37648 8492 37700 8498
rect 37648 8434 37700 8440
rect 35440 8424 35492 8430
rect 35360 8372 35440 8378
rect 35360 8366 35492 8372
rect 37464 8424 37516 8430
rect 37464 8366 37516 8372
rect 35360 8350 35480 8366
rect 35268 8248 35388 8276
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 8084 34848 8090
rect 34796 8026 34848 8032
rect 34980 7948 35032 7954
rect 34980 7890 35032 7896
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 34704 7472 34756 7478
rect 34704 7414 34756 7420
rect 34992 7410 35020 7890
rect 35360 7546 35388 8248
rect 35452 7954 35480 8350
rect 35900 8356 35952 8362
rect 35900 8298 35952 8304
rect 35912 8090 35940 8298
rect 35900 8084 35952 8090
rect 35900 8026 35952 8032
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 35452 7546 35480 7890
rect 35900 7812 35952 7818
rect 35952 7772 36032 7800
rect 35900 7754 35952 7760
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 36004 7562 36032 7772
rect 35348 7540 35400 7546
rect 35348 7482 35400 7488
rect 35440 7540 35492 7546
rect 36004 7534 36124 7562
rect 35440 7482 35492 7488
rect 36096 7478 36124 7534
rect 36084 7472 36136 7478
rect 36084 7414 36136 7420
rect 34980 7404 35032 7410
rect 34980 7346 35032 7352
rect 37752 7342 37780 8774
rect 37844 8566 37872 8910
rect 37936 8906 37964 10610
rect 38028 10130 38056 10610
rect 38108 10600 38160 10606
rect 38108 10542 38160 10548
rect 38120 10198 38148 10542
rect 38108 10192 38160 10198
rect 38108 10134 38160 10140
rect 38016 10124 38068 10130
rect 38016 10066 38068 10072
rect 38212 9994 38240 11630
rect 38844 11620 38896 11626
rect 38844 11562 38896 11568
rect 38384 11552 38436 11558
rect 38384 11494 38436 11500
rect 38396 11150 38424 11494
rect 38856 11354 38884 11562
rect 38844 11348 38896 11354
rect 38844 11290 38896 11296
rect 38384 11144 38436 11150
rect 38384 11086 38436 11092
rect 38396 10674 38424 11086
rect 38568 11008 38620 11014
rect 38568 10950 38620 10956
rect 38580 10674 38608 10950
rect 38856 10674 38884 11290
rect 39500 11218 39528 12038
rect 39488 11212 39540 11218
rect 39488 11154 39540 11160
rect 38384 10668 38436 10674
rect 38384 10610 38436 10616
rect 38476 10668 38528 10674
rect 38476 10610 38528 10616
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38844 10668 38896 10674
rect 38844 10610 38896 10616
rect 38488 10470 38516 10610
rect 39396 10532 39448 10538
rect 39396 10474 39448 10480
rect 38476 10464 38528 10470
rect 38476 10406 38528 10412
rect 38936 10464 38988 10470
rect 38936 10406 38988 10412
rect 38488 10180 38516 10406
rect 38568 10192 38620 10198
rect 38488 10152 38568 10180
rect 38200 9988 38252 9994
rect 38200 9930 38252 9936
rect 38488 9178 38516 10152
rect 38568 10134 38620 10140
rect 38948 10062 38976 10406
rect 38936 10056 38988 10062
rect 38936 9998 38988 10004
rect 39028 10056 39080 10062
rect 39028 9998 39080 10004
rect 38936 9920 38988 9926
rect 38936 9862 38988 9868
rect 38948 9722 38976 9862
rect 39040 9722 39068 9998
rect 39304 9988 39356 9994
rect 39304 9930 39356 9936
rect 38936 9716 38988 9722
rect 38936 9658 38988 9664
rect 39028 9716 39080 9722
rect 39028 9658 39080 9664
rect 39316 9654 39344 9930
rect 39408 9654 39436 10474
rect 40328 10198 40356 16102
rect 40408 16108 40540 16114
rect 40460 16102 40540 16108
rect 40408 16050 40460 16056
rect 40408 15496 40460 15502
rect 40408 15438 40460 15444
rect 40420 15162 40448 15438
rect 40512 15434 40540 16102
rect 40592 16108 40644 16114
rect 40592 16050 40644 16056
rect 40500 15428 40552 15434
rect 40500 15370 40552 15376
rect 40408 15156 40460 15162
rect 40408 15098 40460 15104
rect 40604 15026 40632 16050
rect 40592 15020 40644 15026
rect 40512 14980 40592 15008
rect 40512 14618 40540 14980
rect 40592 14962 40644 14968
rect 40684 14816 40736 14822
rect 40684 14758 40736 14764
rect 40500 14612 40552 14618
rect 40500 14554 40552 14560
rect 40696 14482 40724 14758
rect 40684 14476 40736 14482
rect 40684 14418 40736 14424
rect 40408 13864 40460 13870
rect 40408 13806 40460 13812
rect 40420 13462 40448 13806
rect 40408 13456 40460 13462
rect 40408 13398 40460 13404
rect 40500 13320 40552 13326
rect 40500 13262 40552 13268
rect 40512 12714 40540 13262
rect 40500 12708 40552 12714
rect 40500 12650 40552 12656
rect 40788 12434 40816 17088
rect 41236 16992 41288 16998
rect 41236 16934 41288 16940
rect 41248 16182 41276 16934
rect 41708 16574 41736 19314
rect 41800 18970 41828 20402
rect 41788 18964 41840 18970
rect 41788 18906 41840 18912
rect 41800 18426 41828 18906
rect 41788 18420 41840 18426
rect 41788 18362 41840 18368
rect 41788 17672 41840 17678
rect 41788 17614 41840 17620
rect 41800 17202 41828 17614
rect 41892 17610 41920 22034
rect 42064 21344 42116 21350
rect 42064 21286 42116 21292
rect 42076 20466 42104 21286
rect 42064 20460 42116 20466
rect 42064 20402 42116 20408
rect 42076 18290 42104 20402
rect 42156 19848 42208 19854
rect 42156 19790 42208 19796
rect 42168 18970 42196 19790
rect 42156 18964 42208 18970
rect 42156 18906 42208 18912
rect 42168 18290 42196 18906
rect 42064 18284 42116 18290
rect 42064 18226 42116 18232
rect 42156 18284 42208 18290
rect 42156 18226 42208 18232
rect 41880 17604 41932 17610
rect 41880 17546 41932 17552
rect 41892 17202 41920 17546
rect 41788 17196 41840 17202
rect 41788 17138 41840 17144
rect 41880 17196 41932 17202
rect 41880 17138 41932 17144
rect 42156 17196 42208 17202
rect 42156 17138 42208 17144
rect 42168 16794 42196 17138
rect 42156 16788 42208 16794
rect 42156 16730 42208 16736
rect 41708 16546 41828 16574
rect 41236 16176 41288 16182
rect 41236 16118 41288 16124
rect 41604 16040 41656 16046
rect 41604 15982 41656 15988
rect 40868 15428 40920 15434
rect 40868 15370 40920 15376
rect 41512 15428 41564 15434
rect 41512 15370 41564 15376
rect 40604 12406 40816 12434
rect 40316 10192 40368 10198
rect 40316 10134 40368 10140
rect 40604 10062 40632 12406
rect 40776 11688 40828 11694
rect 40776 11630 40828 11636
rect 40788 10810 40816 11630
rect 40880 11014 40908 15370
rect 41420 15360 41472 15366
rect 41420 15302 41472 15308
rect 41432 15026 41460 15302
rect 41420 15020 41472 15026
rect 41420 14962 41472 14968
rect 41524 14074 41552 15370
rect 41616 14890 41644 15982
rect 41696 15904 41748 15910
rect 41696 15846 41748 15852
rect 41604 14884 41656 14890
rect 41604 14826 41656 14832
rect 41512 14068 41564 14074
rect 41512 14010 41564 14016
rect 41708 13190 41736 15846
rect 41800 13326 41828 16546
rect 42064 16516 42116 16522
rect 42064 16458 42116 16464
rect 41972 15632 42024 15638
rect 41972 15574 42024 15580
rect 41984 15026 42012 15574
rect 41972 15020 42024 15026
rect 41972 14962 42024 14968
rect 41984 14618 42012 14962
rect 41972 14612 42024 14618
rect 41972 14554 42024 14560
rect 42076 14498 42104 16458
rect 41984 14470 42104 14498
rect 41984 14346 42012 14470
rect 41972 14340 42024 14346
rect 41972 14282 42024 14288
rect 41984 14006 42012 14282
rect 41972 14000 42024 14006
rect 41972 13942 42024 13948
rect 41984 13462 42012 13942
rect 41972 13456 42024 13462
rect 41972 13398 42024 13404
rect 41788 13320 41840 13326
rect 41788 13262 41840 13268
rect 41696 13184 41748 13190
rect 41696 13126 41748 13132
rect 41800 12918 41828 13262
rect 41788 12912 41840 12918
rect 41788 12854 41840 12860
rect 40868 11008 40920 11014
rect 40868 10950 40920 10956
rect 40776 10804 40828 10810
rect 40776 10746 40828 10752
rect 40684 10736 40736 10742
rect 40684 10678 40736 10684
rect 40696 10130 40724 10678
rect 41800 10266 41828 12854
rect 41880 10668 41932 10674
rect 41880 10610 41932 10616
rect 41788 10260 41840 10266
rect 41788 10202 41840 10208
rect 40684 10124 40736 10130
rect 40684 10066 40736 10072
rect 40592 10056 40644 10062
rect 40592 9998 40644 10004
rect 39856 9920 39908 9926
rect 39856 9862 39908 9868
rect 39868 9654 39896 9862
rect 40696 9722 40724 10066
rect 40684 9716 40736 9722
rect 40684 9658 40736 9664
rect 39304 9648 39356 9654
rect 39304 9590 39356 9596
rect 39396 9648 39448 9654
rect 39396 9590 39448 9596
rect 39856 9648 39908 9654
rect 39856 9590 39908 9596
rect 38476 9172 38528 9178
rect 38476 9114 38528 9120
rect 37924 8900 37976 8906
rect 37924 8842 37976 8848
rect 37832 8560 37884 8566
rect 37832 8502 37884 8508
rect 37844 8090 37872 8502
rect 37832 8084 37884 8090
rect 37832 8026 37884 8032
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 32496 7200 32548 7206
rect 32496 7142 32548 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 6186 13032 6734
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4622 12480 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11808 3670 11836 4490
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 41892 3602 41920 10610
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 11520 3528 11572 3534
rect 42156 3528 42208 3534
rect 11520 3470 11572 3476
rect 42154 3496 42156 3505
rect 42208 3496 42210 3505
rect 42154 3431 42210 3440
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10336 2854 10364 3062
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 11624 800 11652 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 11610 0 11666 800
<< via2 >>
rect 4880 43546 4936 43548
rect 4960 43546 5016 43548
rect 5040 43546 5096 43548
rect 5120 43546 5176 43548
rect 4880 43494 4926 43546
rect 4926 43494 4936 43546
rect 4960 43494 4990 43546
rect 4990 43494 5002 43546
rect 5002 43494 5016 43546
rect 5040 43494 5054 43546
rect 5054 43494 5066 43546
rect 5066 43494 5096 43546
rect 5120 43494 5130 43546
rect 5130 43494 5176 43546
rect 4880 43492 4936 43494
rect 4960 43492 5016 43494
rect 5040 43492 5096 43494
rect 5120 43492 5176 43494
rect 35600 43546 35656 43548
rect 35680 43546 35736 43548
rect 35760 43546 35816 43548
rect 35840 43546 35896 43548
rect 35600 43494 35646 43546
rect 35646 43494 35656 43546
rect 35680 43494 35710 43546
rect 35710 43494 35722 43546
rect 35722 43494 35736 43546
rect 35760 43494 35774 43546
rect 35774 43494 35786 43546
rect 35786 43494 35816 43546
rect 35840 43494 35850 43546
rect 35850 43494 35896 43546
rect 35600 43492 35656 43494
rect 35680 43492 35736 43494
rect 35760 43492 35816 43494
rect 35840 43492 35896 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4880 42458 4936 42460
rect 4960 42458 5016 42460
rect 5040 42458 5096 42460
rect 5120 42458 5176 42460
rect 4880 42406 4926 42458
rect 4926 42406 4936 42458
rect 4960 42406 4990 42458
rect 4990 42406 5002 42458
rect 5002 42406 5016 42458
rect 5040 42406 5054 42458
rect 5054 42406 5066 42458
rect 5066 42406 5096 42458
rect 5120 42406 5130 42458
rect 5130 42406 5176 42458
rect 4880 42404 4936 42406
rect 4960 42404 5016 42406
rect 5040 42404 5096 42406
rect 5120 42404 5176 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 1306 41520 1362 41576
rect 4880 41370 4936 41372
rect 4960 41370 5016 41372
rect 5040 41370 5096 41372
rect 5120 41370 5176 41372
rect 4880 41318 4926 41370
rect 4926 41318 4936 41370
rect 4960 41318 4990 41370
rect 4990 41318 5002 41370
rect 5002 41318 5016 41370
rect 5040 41318 5054 41370
rect 5054 41318 5066 41370
rect 5066 41318 5096 41370
rect 5120 41318 5130 41370
rect 5130 41318 5176 41370
rect 4880 41316 4936 41318
rect 4960 41316 5016 41318
rect 5040 41316 5096 41318
rect 5120 41316 5176 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4880 40282 4936 40284
rect 4960 40282 5016 40284
rect 5040 40282 5096 40284
rect 5120 40282 5176 40284
rect 4880 40230 4926 40282
rect 4926 40230 4936 40282
rect 4960 40230 4990 40282
rect 4990 40230 5002 40282
rect 5002 40230 5016 40282
rect 5040 40230 5054 40282
rect 5054 40230 5066 40282
rect 5066 40230 5096 40282
rect 5120 40230 5130 40282
rect 5130 40230 5176 40282
rect 4880 40228 4936 40230
rect 4960 40228 5016 40230
rect 5040 40228 5096 40230
rect 5120 40228 5176 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4342 36660 4344 36680
rect 4344 36660 4396 36680
rect 4396 36660 4398 36680
rect 4342 36624 4398 36660
rect 4710 36624 4766 36680
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4342 35012 4398 35048
rect 4342 34992 4344 35012
rect 4344 34992 4396 35012
rect 4396 34992 4398 35012
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4894 35572 4896 35592
rect 4896 35572 4948 35592
rect 4948 35572 4950 35592
rect 4894 35536 4950 35572
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 5170 34448 5226 34504
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 2686 30096 2742 30152
rect 2870 29588 2872 29608
rect 2872 29588 2924 29608
rect 2924 29588 2926 29608
rect 2870 29552 2926 29588
rect 3330 30252 3386 30288
rect 3330 30232 3332 30252
rect 3332 30232 3384 30252
rect 3384 30232 3386 30252
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 5630 35572 5632 35592
rect 5632 35572 5684 35592
rect 5684 35572 5686 35592
rect 5630 35536 5686 35572
rect 5906 34992 5962 35048
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4250 30252 4306 30288
rect 4250 30232 4252 30252
rect 4252 30232 4304 30252
rect 4304 30232 4306 30252
rect 4434 30096 4490 30152
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 846 26732 848 26752
rect 848 26732 900 26752
rect 900 26732 902 26752
rect 846 26696 902 26732
rect 4618 29552 4674 29608
rect 5446 30640 5502 30696
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 3974 26288 4030 26344
rect 846 22616 902 22672
rect 1306 21800 1362 21856
rect 1030 21120 1086 21176
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 5170 26324 5172 26344
rect 5172 26324 5224 26344
rect 5224 26324 5226 26344
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 5170 26288 5226 26324
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 1490 17720 1546 17776
rect 846 16904 902 16960
rect 846 15816 902 15872
rect 1674 15000 1730 15056
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4526 22072 4582 22128
rect 1490 12280 1546 12336
rect 846 11500 848 11520
rect 848 11500 900 11520
rect 900 11500 902 11520
rect 846 11464 902 11500
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 5078 22072 5134 22128
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 7378 36624 7434 36680
rect 7378 34448 7434 34504
rect 7562 24812 7618 24848
rect 7562 24792 7564 24812
rect 7564 24792 7616 24812
rect 7616 24792 7618 24812
rect 6826 23160 6882 23216
rect 9586 24812 9642 24848
rect 9586 24792 9588 24812
rect 9588 24792 9640 24812
rect 9640 24792 9642 24812
rect 8298 23196 8300 23216
rect 8300 23196 8352 23216
rect 8352 23196 8354 23216
rect 8298 23160 8354 23196
rect 11978 28076 12034 28112
rect 12254 28364 12256 28384
rect 12256 28364 12308 28384
rect 12308 28364 12310 28384
rect 12254 28328 12310 28364
rect 12530 29144 12586 29200
rect 12530 29028 12586 29064
rect 12530 29008 12532 29028
rect 12532 29008 12584 29028
rect 12584 29008 12586 29028
rect 12438 28192 12494 28248
rect 11978 28056 11980 28076
rect 11980 28056 12032 28076
rect 12032 28056 12034 28076
rect 12254 26424 12310 26480
rect 13174 29708 13230 29744
rect 13174 29688 13176 29708
rect 13176 29688 13228 29708
rect 13228 29688 13230 29708
rect 12990 27920 13046 27976
rect 12898 27784 12954 27840
rect 12714 27648 12770 27704
rect 12714 27512 12770 27568
rect 13358 28056 13414 28112
rect 13542 28192 13598 28248
rect 13450 27784 13506 27840
rect 13818 28328 13874 28384
rect 13358 23976 13414 24032
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4250 11736 4306 11792
rect 4434 11600 4490 11656
rect 4710 11756 4766 11792
rect 4710 11736 4712 11756
rect 4712 11736 4764 11756
rect 4764 11736 4766 11756
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5354 11736 5410 11792
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 9586 18708 9588 18728
rect 9588 18708 9640 18728
rect 9640 18708 9642 18728
rect 9586 18672 9642 18708
rect 13910 27920 13966 27976
rect 13910 27648 13966 27704
rect 15750 31084 15752 31104
rect 15752 31084 15804 31104
rect 15804 31084 15806 31104
rect 15750 31048 15806 31084
rect 17590 40976 17646 41032
rect 14554 27784 14610 27840
rect 15198 28076 15254 28112
rect 15198 28056 15200 28076
rect 15200 28056 15252 28076
rect 15252 28056 15254 28076
rect 6734 11636 6736 11656
rect 6736 11636 6788 11656
rect 6788 11636 6790 11656
rect 6734 11600 6790 11636
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3698 7928 3754 7984
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4526 7928 4582 7984
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 12530 18708 12532 18728
rect 12532 18708 12584 18728
rect 12584 18708 12586 18728
rect 12530 18672 12586 18708
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 9586 11464 9642 11520
rect 9586 11056 9642 11112
rect 7838 7964 7840 7984
rect 7840 7964 7892 7984
rect 7892 7964 7894 7984
rect 7838 7928 7894 7964
rect 7838 7828 7840 7848
rect 7840 7828 7892 7848
rect 7892 7828 7894 7848
rect 7838 7792 7894 7828
rect 8298 7828 8300 7848
rect 8300 7828 8352 7848
rect 8352 7828 8354 7848
rect 8298 7792 8354 7828
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9034 7948 9090 7984
rect 9034 7928 9036 7948
rect 9036 7928 9088 7948
rect 9088 7928 9090 7948
rect 15198 26444 15254 26480
rect 15198 26424 15200 26444
rect 15200 26424 15252 26444
rect 15252 26424 15254 26444
rect 15658 29044 15660 29064
rect 15660 29044 15712 29064
rect 15712 29044 15714 29064
rect 15658 29008 15714 29044
rect 15934 29960 15990 30016
rect 16578 31592 16634 31648
rect 16486 31320 16542 31376
rect 16210 30232 16266 30288
rect 16118 29824 16174 29880
rect 16854 31184 16910 31240
rect 16394 28056 16450 28112
rect 15474 25236 15476 25256
rect 15476 25236 15528 25256
rect 15528 25236 15530 25256
rect 15474 25200 15530 25236
rect 15566 24792 15622 24848
rect 16578 25336 16634 25392
rect 16394 23724 16450 23760
rect 16394 23704 16396 23724
rect 16396 23704 16448 23724
rect 16448 23704 16450 23724
rect 17130 30776 17186 30832
rect 17130 30096 17186 30152
rect 17130 29280 17186 29336
rect 16946 29008 17002 29064
rect 17038 24656 17094 24712
rect 17406 31592 17462 31648
rect 17314 31340 17370 31376
rect 17314 31320 17316 31340
rect 17316 31320 17368 31340
rect 17368 31320 17370 31340
rect 17314 31184 17370 31240
rect 17498 31340 17554 31376
rect 17498 31320 17500 31340
rect 17500 31320 17552 31340
rect 17552 31320 17554 31340
rect 17498 30776 17554 30832
rect 17498 29144 17554 29200
rect 18142 30232 18198 30288
rect 18970 37204 18972 37224
rect 18972 37204 19024 37224
rect 19024 37204 19026 37224
rect 18970 37168 19026 37204
rect 18602 31320 18658 31376
rect 18142 29960 18198 30016
rect 17682 29280 17738 29336
rect 17406 25372 17408 25392
rect 17408 25372 17460 25392
rect 17460 25372 17462 25392
rect 17406 25336 17462 25372
rect 18234 29280 18290 29336
rect 17958 25200 18014 25256
rect 17774 24792 17830 24848
rect 17682 24656 17738 24712
rect 18418 31048 18474 31104
rect 19246 41012 19248 41032
rect 19248 41012 19300 41032
rect 19300 41012 19302 41032
rect 19246 40976 19302 41012
rect 20994 42880 21050 42936
rect 20810 41520 20866 41576
rect 21362 38276 21418 38312
rect 21362 38256 21364 38276
rect 21364 38256 21416 38276
rect 21416 38256 21418 38276
rect 18602 30504 18658 30560
rect 18602 29996 18604 30016
rect 18604 29996 18656 30016
rect 18656 29996 18658 30016
rect 18602 29960 18658 29996
rect 19062 30504 19118 30560
rect 18234 24248 18290 24304
rect 18142 24112 18198 24168
rect 18694 25336 18750 25392
rect 18694 24812 18750 24848
rect 18694 24792 18696 24812
rect 18696 24792 18748 24812
rect 18748 24792 18750 24812
rect 18418 24112 18474 24168
rect 18326 23840 18382 23896
rect 19338 28056 19394 28112
rect 20718 31456 20774 31512
rect 20994 31456 21050 31512
rect 19706 28056 19762 28112
rect 20810 29572 20866 29608
rect 20810 29552 20812 29572
rect 20812 29552 20864 29572
rect 20864 29552 20866 29572
rect 19246 24248 19302 24304
rect 18602 21972 18604 21992
rect 18604 21972 18656 21992
rect 18656 21972 18658 21992
rect 18602 21936 18658 21972
rect 19292 24112 19348 24168
rect 19246 24012 19248 24032
rect 19248 24012 19300 24032
rect 19300 24012 19302 24032
rect 19246 23976 19302 24012
rect 19154 23840 19210 23896
rect 21178 31728 21234 31784
rect 20994 29688 21050 29744
rect 20994 28756 21050 28792
rect 20994 28736 20996 28756
rect 20996 28736 21048 28756
rect 21048 28736 21050 28756
rect 21638 38392 21694 38448
rect 21546 31764 21548 31784
rect 21548 31764 21600 31784
rect 21600 31764 21602 31784
rect 21546 31728 21602 31764
rect 22006 41556 22008 41576
rect 22008 41556 22060 41576
rect 22060 41556 22062 41576
rect 22006 41520 22062 41556
rect 22558 41132 22614 41168
rect 22558 41112 22560 41132
rect 22560 41112 22612 41132
rect 22612 41112 22614 41132
rect 21822 39344 21878 39400
rect 22282 38428 22284 38448
rect 22284 38428 22336 38448
rect 22336 38428 22338 38448
rect 22282 38392 22338 38428
rect 22374 38292 22376 38312
rect 22376 38292 22428 38312
rect 22428 38292 22430 38312
rect 22374 38256 22430 38292
rect 21822 38156 21824 38176
rect 21824 38156 21876 38176
rect 21876 38156 21878 38176
rect 21822 38120 21878 38156
rect 22558 38156 22560 38176
rect 22560 38156 22612 38176
rect 22612 38156 22614 38176
rect 22558 38120 22614 38156
rect 21454 30540 21456 30560
rect 21456 30540 21508 30560
rect 21508 30540 21510 30560
rect 21454 30504 21510 30540
rect 21178 27512 21234 27568
rect 21914 29164 21970 29200
rect 21914 29144 21916 29164
rect 21916 29144 21968 29164
rect 21968 29144 21970 29164
rect 18970 16088 19026 16144
rect 19154 17040 19210 17096
rect 19430 17040 19486 17096
rect 19522 15952 19578 16008
rect 20166 15952 20222 16008
rect 19706 12688 19762 12744
rect 20166 10920 20222 10976
rect 21638 21972 21640 21992
rect 21640 21972 21692 21992
rect 21692 21972 21694 21992
rect 21638 21936 21694 21972
rect 23754 41132 23810 41168
rect 23754 41112 23756 41132
rect 23756 41112 23808 41132
rect 23808 41112 23810 41132
rect 24030 34040 24086 34096
rect 23478 25780 23480 25800
rect 23480 25780 23532 25800
rect 23532 25780 23534 25800
rect 23478 25744 23534 25780
rect 23570 24812 23626 24848
rect 23570 24792 23572 24812
rect 23572 24792 23624 24812
rect 23624 24792 23626 24812
rect 23202 24656 23258 24712
rect 21362 12280 21418 12336
rect 20902 10920 20958 10976
rect 25962 40588 26018 40624
rect 25962 40568 25964 40588
rect 25964 40568 26016 40588
rect 26016 40568 26018 40588
rect 26238 40568 26294 40624
rect 24306 27940 24362 27976
rect 24306 27920 24308 27940
rect 24308 27920 24360 27940
rect 24360 27920 24362 27940
rect 27526 34060 27582 34096
rect 27526 34040 27528 34060
rect 27528 34040 27580 34060
rect 27580 34040 27582 34060
rect 26054 28600 26110 28656
rect 25042 25900 25098 25936
rect 25042 25880 25044 25900
rect 25044 25880 25096 25900
rect 25096 25880 25098 25900
rect 24490 24812 24546 24848
rect 24490 24792 24492 24812
rect 24492 24792 24544 24812
rect 24544 24792 24546 24812
rect 23570 16360 23626 16416
rect 22834 12144 22890 12200
rect 19798 7420 19800 7440
rect 19800 7420 19852 7440
rect 19852 7420 19854 7440
rect 19798 7384 19854 7420
rect 25686 25900 25742 25936
rect 25686 25880 25688 25900
rect 25688 25880 25740 25900
rect 25740 25880 25742 25900
rect 27802 29552 27858 29608
rect 25410 25744 25466 25800
rect 25042 24792 25098 24848
rect 24950 21836 24952 21856
rect 24952 21836 25004 21856
rect 25004 21836 25006 21856
rect 24950 21800 25006 21836
rect 25502 23704 25558 23760
rect 25778 22924 25780 22944
rect 25780 22924 25832 22944
rect 25832 22924 25834 22944
rect 25778 22888 25834 22924
rect 25962 16396 25964 16416
rect 25964 16396 26016 16416
rect 26016 16396 26018 16416
rect 25962 16360 26018 16396
rect 25042 13640 25098 13696
rect 25686 13676 25688 13696
rect 25688 13676 25740 13696
rect 25740 13676 25742 13696
rect 25686 13640 25742 13676
rect 23570 12688 23626 12744
rect 23478 12180 23480 12200
rect 23480 12180 23532 12200
rect 23532 12180 23534 12200
rect 23478 12144 23534 12180
rect 28354 30368 28410 30424
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35600 42458 35656 42460
rect 35680 42458 35736 42460
rect 35760 42458 35816 42460
rect 35840 42458 35896 42460
rect 35600 42406 35646 42458
rect 35646 42406 35656 42458
rect 35680 42406 35710 42458
rect 35710 42406 35722 42458
rect 35722 42406 35736 42458
rect 35760 42406 35774 42458
rect 35774 42406 35786 42458
rect 35786 42406 35816 42458
rect 35840 42406 35850 42458
rect 35850 42406 35896 42458
rect 35600 42404 35656 42406
rect 35680 42404 35736 42406
rect 35760 42404 35816 42406
rect 35840 42404 35896 42406
rect 30838 39500 30894 39536
rect 30838 39480 30840 39500
rect 30840 39480 30892 39500
rect 30892 39480 30894 39500
rect 30746 38956 30802 38992
rect 30746 38936 30748 38956
rect 30748 38936 30800 38956
rect 30800 38936 30802 38956
rect 31390 39344 31446 39400
rect 31758 39380 31760 39400
rect 31760 39380 31812 39400
rect 31812 39380 31814 39400
rect 31758 39344 31814 39380
rect 29182 30660 29238 30696
rect 29182 30640 29184 30660
rect 29184 30640 29236 30660
rect 29236 30640 29238 30660
rect 28998 29280 29054 29336
rect 29550 29960 29606 30016
rect 28906 28600 28962 28656
rect 28814 27784 28870 27840
rect 28722 25744 28778 25800
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 33046 38956 33102 38992
rect 30930 29008 30986 29064
rect 30838 27512 30894 27568
rect 27526 17176 27582 17232
rect 26882 12316 26884 12336
rect 26884 12316 26936 12336
rect 26936 12316 26938 12336
rect 26882 12280 26938 12316
rect 25594 10684 25596 10704
rect 25596 10684 25648 10704
rect 25648 10684 25650 10704
rect 25594 10648 25650 10684
rect 30746 25236 30748 25256
rect 30748 25236 30800 25256
rect 30800 25236 30802 25256
rect 30746 25200 30802 25236
rect 31206 27784 31262 27840
rect 33046 38936 33048 38956
rect 33048 38936 33100 38956
rect 33100 38936 33102 38956
rect 32218 30132 32220 30152
rect 32220 30132 32272 30152
rect 32272 30132 32274 30152
rect 32218 30096 32274 30132
rect 28446 17196 28502 17232
rect 28446 17176 28448 17196
rect 28448 17176 28500 17196
rect 28500 17176 28502 17196
rect 28446 16768 28502 16824
rect 28906 16788 28962 16824
rect 28906 16768 28908 16788
rect 28908 16768 28960 16788
rect 28960 16768 28962 16788
rect 28998 16224 29054 16280
rect 29182 16224 29238 16280
rect 26238 9460 26240 9480
rect 26240 9460 26292 9480
rect 26292 9460 26294 9480
rect 26238 9424 26294 9460
rect 23202 7420 23204 7440
rect 23204 7420 23256 7440
rect 23256 7420 23258 7440
rect 23202 7384 23258 7420
rect 26606 9580 26662 9616
rect 26606 9560 26608 9580
rect 26608 9560 26660 9580
rect 26660 9560 26662 9580
rect 27342 9596 27344 9616
rect 27344 9596 27396 9616
rect 27396 9596 27398 9616
rect 27342 9560 27398 9596
rect 27066 9460 27068 9480
rect 27068 9460 27120 9480
rect 27120 9460 27122 9480
rect 27066 9424 27122 9460
rect 28262 10648 28318 10704
rect 29182 15136 29238 15192
rect 32954 30232 33010 30288
rect 32770 28192 32826 28248
rect 32678 25356 32734 25392
rect 32678 25336 32680 25356
rect 32680 25336 32732 25356
rect 32732 25336 32734 25356
rect 33046 28872 33102 28928
rect 29918 15444 29920 15464
rect 29920 15444 29972 15464
rect 29972 15444 29974 15464
rect 29918 15408 29974 15444
rect 30930 16532 30932 16552
rect 30932 16532 30984 16552
rect 30984 16532 30986 16552
rect 30930 16496 30986 16532
rect 30562 16224 30618 16280
rect 30286 15952 30342 16008
rect 30470 15444 30472 15464
rect 30472 15444 30524 15464
rect 30524 15444 30526 15464
rect 30470 15408 30526 15444
rect 30562 15136 30618 15192
rect 31666 16360 31722 16416
rect 32126 16496 32182 16552
rect 32770 22516 32772 22536
rect 32772 22516 32824 22536
rect 32824 22516 32826 22536
rect 32770 22480 32826 22516
rect 33414 28464 33470 28520
rect 35600 41370 35656 41372
rect 35680 41370 35736 41372
rect 35760 41370 35816 41372
rect 35840 41370 35896 41372
rect 35600 41318 35646 41370
rect 35646 41318 35656 41370
rect 35680 41318 35710 41370
rect 35710 41318 35722 41370
rect 35722 41318 35736 41370
rect 35760 41318 35774 41370
rect 35774 41318 35786 41370
rect 35786 41318 35816 41370
rect 35840 41318 35850 41370
rect 35850 41318 35896 41370
rect 35600 41316 35656 41318
rect 35680 41316 35736 41318
rect 35760 41316 35816 41318
rect 35840 41316 35896 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 33966 37204 33968 37224
rect 33968 37204 34020 37224
rect 34020 37204 34022 37224
rect 33966 37168 34022 37204
rect 35600 40282 35656 40284
rect 35680 40282 35736 40284
rect 35760 40282 35816 40284
rect 35840 40282 35896 40284
rect 35600 40230 35646 40282
rect 35646 40230 35656 40282
rect 35680 40230 35710 40282
rect 35710 40230 35722 40282
rect 35722 40230 35736 40282
rect 35760 40230 35774 40282
rect 35774 40230 35786 40282
rect 35786 40230 35816 40282
rect 35840 40230 35850 40282
rect 35850 40230 35896 40282
rect 35600 40228 35656 40230
rect 35680 40228 35736 40230
rect 35760 40228 35816 40230
rect 35840 40228 35896 40230
rect 35714 39480 35770 39536
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 35530 38820 35586 38856
rect 35530 38800 35532 38820
rect 35532 38800 35584 38820
rect 35584 38800 35586 38820
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 36082 38800 36138 38856
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 33966 29552 34022 29608
rect 34058 29144 34114 29200
rect 33874 28872 33930 28928
rect 33690 28192 33746 28248
rect 34058 28484 34114 28520
rect 34058 28464 34060 28484
rect 34060 28464 34112 28484
rect 34112 28464 34114 28484
rect 34426 30116 34482 30152
rect 34426 30096 34428 30116
rect 34428 30096 34480 30116
rect 34480 30096 34482 30116
rect 34426 29824 34482 29880
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35162 30116 35218 30152
rect 35162 30096 35164 30116
rect 35164 30096 35216 30116
rect 35216 30096 35218 30116
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34610 29180 34612 29200
rect 34612 29180 34664 29200
rect 34664 29180 34666 29200
rect 34610 29144 34666 29180
rect 34334 28076 34390 28112
rect 34334 28056 34336 28076
rect 34336 28056 34388 28076
rect 34388 28056 34390 28076
rect 32494 15952 32550 16008
rect 33322 16396 33324 16416
rect 33324 16396 33376 16416
rect 33376 16396 33378 16416
rect 33138 16224 33194 16280
rect 33322 16360 33378 16396
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 35070 29688 35126 29744
rect 34978 29280 35034 29336
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35070 28484 35126 28520
rect 35070 28464 35072 28484
rect 35072 28464 35124 28484
rect 35124 28464 35126 28484
rect 35622 29688 35678 29744
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 36542 28464 36598 28520
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34334 24112 34390 24168
rect 34242 15952 34298 16008
rect 34886 24792 34942 24848
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 35898 25200 35954 25256
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 35438 24812 35494 24848
rect 35438 24792 35440 24812
rect 35440 24792 35492 24812
rect 35492 24792 35494 24812
rect 35346 24692 35348 24712
rect 35348 24692 35400 24712
rect 35400 24692 35402 24712
rect 35346 24656 35402 24692
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 36174 24520 36230 24576
rect 35530 24132 35586 24168
rect 35530 24112 35532 24132
rect 35532 24112 35584 24132
rect 35584 24112 35586 24132
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34610 20984 34666 21040
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34978 20984 35034 21040
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34426 13368 34482 13424
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34886 13776 34942 13832
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34978 13232 35034 13288
rect 37922 27512 37978 27568
rect 37278 25200 37334 25256
rect 38014 20712 38070 20768
rect 36358 13368 36414 13424
rect 35990 13232 36046 13288
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 35162 12824 35218 12880
rect 35346 12824 35402 12880
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34150 10684 34152 10704
rect 34152 10684 34204 10704
rect 34204 10684 34206 10704
rect 34150 10648 34206 10684
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34978 10684 34980 10704
rect 34980 10684 35032 10704
rect 35032 10684 35034 10704
rect 34978 10648 35034 10684
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 38382 29144 38438 29200
rect 38934 27920 38990 27976
rect 38750 27512 38806 27568
rect 38750 27104 38806 27160
rect 38382 25200 38438 25256
rect 37094 12824 37150 12880
rect 42062 31320 42118 31376
rect 40498 30252 40554 30288
rect 40498 30232 40500 30252
rect 40500 30232 40552 30252
rect 40552 30232 40554 30252
rect 40038 28872 40094 28928
rect 38290 15428 38346 15464
rect 38290 15408 38292 15428
rect 38292 15408 38344 15428
rect 38344 15408 38346 15428
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 36450 10648 36506 10704
rect 37002 10648 37058 10704
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 40866 29552 40922 29608
rect 40130 25200 40186 25256
rect 40590 24556 40592 24576
rect 40592 24556 40644 24576
rect 40644 24556 40646 24576
rect 40590 24520 40646 24556
rect 41694 27920 41750 27976
rect 41510 27276 41512 27296
rect 41512 27276 41564 27296
rect 41564 27276 41566 27296
rect 41510 27240 41566 27276
rect 42062 29280 42118 29336
rect 41878 28600 41934 28656
rect 41878 26560 41934 26616
rect 42062 28600 42118 28656
rect 42062 25880 42118 25936
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 42154 3476 42156 3496
rect 42156 3476 42208 3496
rect 42208 3476 42210 3496
rect 42154 3440 42210 3476
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4870 43552 5186 43553
rect 4870 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5186 43552
rect 4870 43487 5186 43488
rect 35590 43552 35906 43553
rect 35590 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35906 43552
rect 35590 43487 35906 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 20989 42940 21055 42941
rect 20989 42936 21036 42940
rect 21100 42938 21106 42940
rect 20989 42880 20994 42936
rect 20989 42876 21036 42880
rect 21100 42878 21146 42938
rect 21100 42876 21106 42878
rect 20989 42875 21055 42876
rect 4870 42464 5186 42465
rect 4870 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5186 42464
rect 4870 42399 5186 42400
rect 35590 42464 35906 42465
rect 35590 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35906 42464
rect 35590 42399 35906 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 0 41578 800 41608
rect 1301 41578 1367 41581
rect 20805 41580 20871 41581
rect 20805 41578 20852 41580
rect 0 41576 1367 41578
rect 0 41520 1306 41576
rect 1362 41520 1367 41576
rect 0 41518 1367 41520
rect 20724 41576 20852 41578
rect 20916 41578 20922 41580
rect 22001 41578 22067 41581
rect 20916 41576 22067 41578
rect 20724 41520 20810 41576
rect 20916 41520 22006 41576
rect 22062 41520 22067 41576
rect 20724 41518 20852 41520
rect 0 41488 800 41518
rect 1301 41515 1367 41518
rect 20805 41516 20852 41518
rect 20916 41518 22067 41520
rect 20916 41516 20922 41518
rect 20805 41515 20871 41516
rect 22001 41515 22067 41518
rect 4870 41376 5186 41377
rect 4870 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5186 41376
rect 4870 41311 5186 41312
rect 35590 41376 35906 41377
rect 35590 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35906 41376
rect 35590 41311 35906 41312
rect 22553 41170 22619 41173
rect 23749 41170 23815 41173
rect 22553 41168 23815 41170
rect 22553 41112 22558 41168
rect 22614 41112 23754 41168
rect 23810 41112 23815 41168
rect 22553 41110 23815 41112
rect 22553 41107 22619 41110
rect 23749 41107 23815 41110
rect 17585 41034 17651 41037
rect 19241 41034 19307 41037
rect 17585 41032 19307 41034
rect 17585 40976 17590 41032
rect 17646 40976 19246 41032
rect 19302 40976 19307 41032
rect 17585 40974 19307 40976
rect 17585 40971 17651 40974
rect 19241 40971 19307 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 25957 40628 26023 40629
rect 25957 40626 26004 40628
rect 25912 40624 26004 40626
rect 26068 40626 26074 40628
rect 26233 40626 26299 40629
rect 26068 40624 26299 40626
rect 25912 40568 25962 40624
rect 26068 40568 26238 40624
rect 26294 40568 26299 40624
rect 25912 40566 26004 40568
rect 25957 40564 26004 40566
rect 26068 40566 26299 40568
rect 26068 40564 26074 40566
rect 25957 40563 26023 40564
rect 26233 40563 26299 40566
rect 4870 40288 5186 40289
rect 4870 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5186 40288
rect 4870 40223 5186 40224
rect 35590 40288 35906 40289
rect 35590 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35906 40288
rect 35590 40223 35906 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 30833 39538 30899 39541
rect 35709 39538 35775 39541
rect 30833 39536 35775 39538
rect 30833 39480 30838 39536
rect 30894 39480 35714 39536
rect 35770 39480 35775 39536
rect 30833 39478 35775 39480
rect 30833 39475 30899 39478
rect 35709 39475 35775 39478
rect 21817 39402 21883 39405
rect 21950 39402 21956 39404
rect 21817 39400 21956 39402
rect 21817 39344 21822 39400
rect 21878 39344 21956 39400
rect 21817 39342 21956 39344
rect 21817 39339 21883 39342
rect 21950 39340 21956 39342
rect 22020 39340 22026 39404
rect 31385 39402 31451 39405
rect 31753 39402 31819 39405
rect 31385 39400 31819 39402
rect 31385 39344 31390 39400
rect 31446 39344 31758 39400
rect 31814 39344 31819 39400
rect 31385 39342 31819 39344
rect 31385 39339 31451 39342
rect 31753 39339 31819 39342
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 30741 38994 30807 38997
rect 33041 38994 33107 38997
rect 30741 38992 33107 38994
rect 30741 38936 30746 38992
rect 30802 38936 33046 38992
rect 33102 38936 33107 38992
rect 30741 38934 33107 38936
rect 30741 38931 30807 38934
rect 33041 38931 33107 38934
rect 35525 38858 35591 38861
rect 36077 38858 36143 38861
rect 35525 38856 36143 38858
rect 35525 38800 35530 38856
rect 35586 38800 36082 38856
rect 36138 38800 36143 38856
rect 35525 38798 36143 38800
rect 35525 38795 35591 38798
rect 36077 38795 36143 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 21633 38450 21699 38453
rect 22277 38450 22343 38453
rect 21633 38448 22343 38450
rect 21633 38392 21638 38448
rect 21694 38392 22282 38448
rect 22338 38392 22343 38448
rect 21633 38390 22343 38392
rect 21633 38387 21699 38390
rect 22277 38387 22343 38390
rect 21357 38314 21423 38317
rect 22369 38314 22435 38317
rect 21357 38312 22435 38314
rect 21357 38256 21362 38312
rect 21418 38256 22374 38312
rect 22430 38256 22435 38312
rect 21357 38254 22435 38256
rect 21357 38251 21423 38254
rect 22369 38251 22435 38254
rect 21817 38178 21883 38181
rect 22553 38178 22619 38181
rect 21817 38176 22619 38178
rect 21817 38120 21822 38176
rect 21878 38120 22558 38176
rect 22614 38120 22619 38176
rect 21817 38118 22619 38120
rect 21817 38115 21883 38118
rect 22553 38115 22619 38118
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 18965 37226 19031 37229
rect 33961 37226 34027 37229
rect 18965 37224 34027 37226
rect 18965 37168 18970 37224
rect 19026 37168 33966 37224
rect 34022 37168 34027 37224
rect 18965 37166 34027 37168
rect 18965 37163 19031 37166
rect 33961 37163 34027 37166
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4337 36682 4403 36685
rect 4705 36682 4771 36685
rect 7373 36682 7439 36685
rect 4337 36680 7439 36682
rect 4337 36624 4342 36680
rect 4398 36624 4710 36680
rect 4766 36624 7378 36680
rect 7434 36624 7439 36680
rect 4337 36622 7439 36624
rect 4337 36619 4403 36622
rect 4705 36619 4771 36622
rect 7373 36619 7439 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4889 35594 4955 35597
rect 5625 35594 5691 35597
rect 4889 35592 5691 35594
rect 4889 35536 4894 35592
rect 4950 35536 5630 35592
rect 5686 35536 5691 35592
rect 4889 35534 5691 35536
rect 4889 35531 4955 35534
rect 5625 35531 5691 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4337 35050 4403 35053
rect 5901 35050 5967 35053
rect 4337 35048 5967 35050
rect 4337 34992 4342 35048
rect 4398 34992 5906 35048
rect 5962 34992 5967 35048
rect 4337 34990 5967 34992
rect 4337 34987 4403 34990
rect 5901 34987 5967 34990
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 5165 34506 5231 34509
rect 5390 34506 5396 34508
rect 5165 34504 5396 34506
rect 5165 34448 5170 34504
rect 5226 34448 5396 34504
rect 5165 34446 5396 34448
rect 5165 34443 5231 34446
rect 5390 34444 5396 34446
rect 5460 34506 5466 34508
rect 7373 34506 7439 34509
rect 5460 34504 7439 34506
rect 5460 34448 7378 34504
rect 7434 34448 7439 34504
rect 5460 34446 7439 34448
rect 5460 34444 5466 34446
rect 7373 34443 7439 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 24025 34098 24091 34101
rect 27521 34098 27587 34101
rect 24025 34096 27587 34098
rect 24025 34040 24030 34096
rect 24086 34040 27526 34096
rect 27582 34040 27587 34096
rect 24025 34038 27587 34040
rect 24025 34035 24091 34038
rect 27521 34035 27587 34038
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 21173 31786 21239 31789
rect 21541 31786 21607 31789
rect 21173 31784 21607 31786
rect 21173 31728 21178 31784
rect 21234 31728 21546 31784
rect 21602 31728 21607 31784
rect 21173 31726 21607 31728
rect 21173 31723 21239 31726
rect 21541 31723 21607 31726
rect 16573 31650 16639 31653
rect 17401 31650 17467 31653
rect 16573 31648 17467 31650
rect 16573 31592 16578 31648
rect 16634 31592 17406 31648
rect 17462 31592 17467 31648
rect 16573 31590 17467 31592
rect 16573 31587 16639 31590
rect 17401 31587 17467 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 20713 31514 20779 31517
rect 20989 31514 21055 31517
rect 20713 31512 21055 31514
rect 20713 31456 20718 31512
rect 20774 31456 20994 31512
rect 21050 31456 21055 31512
rect 20713 31454 21055 31456
rect 20713 31451 20779 31454
rect 20989 31451 21055 31454
rect 16481 31378 16547 31381
rect 17309 31378 17375 31381
rect 16481 31376 17375 31378
rect 16481 31320 16486 31376
rect 16542 31320 17314 31376
rect 17370 31320 17375 31376
rect 16481 31318 17375 31320
rect 16481 31315 16547 31318
rect 17309 31315 17375 31318
rect 17493 31378 17559 31381
rect 18597 31378 18663 31381
rect 17493 31376 18663 31378
rect 17493 31320 17498 31376
rect 17554 31320 18602 31376
rect 18658 31320 18663 31376
rect 17493 31318 18663 31320
rect 17493 31315 17559 31318
rect 18597 31315 18663 31318
rect 42057 31378 42123 31381
rect 42843 31378 43643 31408
rect 42057 31376 43643 31378
rect 42057 31320 42062 31376
rect 42118 31320 43643 31376
rect 42057 31318 43643 31320
rect 42057 31315 42123 31318
rect 42843 31288 43643 31318
rect 16849 31242 16915 31245
rect 17309 31242 17375 31245
rect 16849 31240 17375 31242
rect 16849 31184 16854 31240
rect 16910 31184 17314 31240
rect 17370 31184 17375 31240
rect 16849 31182 17375 31184
rect 16849 31179 16915 31182
rect 17309 31179 17375 31182
rect 15745 31108 15811 31109
rect 15694 31044 15700 31108
rect 15764 31106 15811 31108
rect 18413 31106 18479 31109
rect 15764 31104 18479 31106
rect 15806 31048 18418 31104
rect 18474 31048 18479 31104
rect 15764 31046 18479 31048
rect 15764 31044 15811 31046
rect 15745 31043 15811 31044
rect 18413 31043 18479 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 17125 30834 17191 30837
rect 17493 30834 17559 30837
rect 17125 30832 17559 30834
rect 17125 30776 17130 30832
rect 17186 30776 17498 30832
rect 17554 30776 17559 30832
rect 17125 30774 17559 30776
rect 17125 30771 17191 30774
rect 17493 30771 17559 30774
rect 5441 30700 5507 30701
rect 5390 30698 5396 30700
rect 5350 30638 5396 30698
rect 5460 30696 5507 30700
rect 5502 30640 5507 30696
rect 5390 30636 5396 30638
rect 5460 30636 5507 30640
rect 17902 30636 17908 30700
rect 17972 30698 17978 30700
rect 29177 30698 29243 30701
rect 17972 30696 29243 30698
rect 17972 30640 29182 30696
rect 29238 30640 29243 30696
rect 17972 30638 29243 30640
rect 17972 30636 17978 30638
rect 5441 30635 5507 30636
rect 29177 30635 29243 30638
rect 18597 30562 18663 30565
rect 19057 30562 19123 30565
rect 18597 30560 19123 30562
rect 18597 30504 18602 30560
rect 18658 30504 19062 30560
rect 19118 30504 19123 30560
rect 18597 30502 19123 30504
rect 18597 30499 18663 30502
rect 19057 30499 19123 30502
rect 21449 30562 21515 30565
rect 21766 30562 21772 30564
rect 21449 30560 21772 30562
rect 21449 30504 21454 30560
rect 21510 30504 21772 30560
rect 21449 30502 21772 30504
rect 21449 30499 21515 30502
rect 21766 30500 21772 30502
rect 21836 30500 21842 30564
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 28349 30426 28415 30429
rect 17910 30424 28415 30426
rect 17910 30368 28354 30424
rect 28410 30368 28415 30424
rect 17910 30366 28415 30368
rect 3325 30290 3391 30293
rect 4245 30290 4311 30293
rect 3325 30288 4311 30290
rect 3325 30232 3330 30288
rect 3386 30232 4250 30288
rect 4306 30232 4311 30288
rect 3325 30230 4311 30232
rect 3325 30227 3391 30230
rect 4245 30227 4311 30230
rect 16205 30290 16271 30293
rect 17910 30290 17970 30366
rect 28349 30363 28415 30366
rect 16205 30288 17970 30290
rect 16205 30232 16210 30288
rect 16266 30232 17970 30288
rect 16205 30230 17970 30232
rect 18137 30290 18203 30293
rect 32949 30290 33015 30293
rect 40493 30290 40559 30293
rect 18137 30288 22110 30290
rect 18137 30232 18142 30288
rect 18198 30232 22110 30288
rect 18137 30230 22110 30232
rect 16205 30227 16271 30230
rect 18137 30227 18203 30230
rect 2681 30154 2747 30157
rect 4429 30154 4495 30157
rect 2681 30152 4495 30154
rect 2681 30096 2686 30152
rect 2742 30096 4434 30152
rect 4490 30096 4495 30152
rect 2681 30094 4495 30096
rect 2681 30091 2747 30094
rect 4429 30091 4495 30094
rect 17125 30154 17191 30157
rect 22050 30154 22110 30230
rect 32949 30288 40559 30290
rect 32949 30232 32954 30288
rect 33010 30232 40498 30288
rect 40554 30232 40559 30288
rect 32949 30230 40559 30232
rect 32949 30227 33015 30230
rect 40493 30227 40559 30230
rect 32213 30154 32279 30157
rect 17125 30152 18890 30154
rect 17125 30096 17130 30152
rect 17186 30096 18890 30152
rect 17125 30094 18890 30096
rect 22050 30152 32279 30154
rect 22050 30096 32218 30152
rect 32274 30096 32279 30152
rect 22050 30094 32279 30096
rect 17125 30091 17191 30094
rect 15929 30018 15995 30021
rect 18137 30018 18203 30021
rect 18597 30020 18663 30021
rect 18597 30018 18644 30020
rect 15929 30016 18203 30018
rect 15929 29960 15934 30016
rect 15990 29960 18142 30016
rect 18198 29960 18203 30016
rect 15929 29958 18203 29960
rect 18552 30016 18644 30018
rect 18552 29960 18602 30016
rect 18552 29958 18644 29960
rect 15929 29955 15995 29958
rect 18137 29955 18203 29958
rect 18597 29956 18644 29958
rect 18708 29956 18714 30020
rect 18830 30018 18890 30094
rect 32213 30091 32279 30094
rect 34421 30154 34487 30157
rect 35157 30154 35223 30157
rect 34421 30152 35223 30154
rect 34421 30096 34426 30152
rect 34482 30096 35162 30152
rect 35218 30096 35223 30152
rect 34421 30094 35223 30096
rect 34421 30091 34487 30094
rect 35157 30091 35223 30094
rect 29545 30018 29611 30021
rect 18830 30016 29611 30018
rect 18830 29960 29550 30016
rect 29606 29960 29611 30016
rect 18830 29958 29611 29960
rect 18597 29955 18663 29956
rect 29545 29955 29611 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 16113 29882 16179 29885
rect 34421 29882 34487 29885
rect 16113 29880 34487 29882
rect 16113 29824 16118 29880
rect 16174 29824 34426 29880
rect 34482 29824 34487 29880
rect 16113 29822 34487 29824
rect 16113 29819 16179 29822
rect 34421 29819 34487 29822
rect 13169 29746 13235 29749
rect 17902 29746 17908 29748
rect 13169 29744 17908 29746
rect 13169 29688 13174 29744
rect 13230 29688 17908 29744
rect 13169 29686 17908 29688
rect 13169 29683 13235 29686
rect 17902 29684 17908 29686
rect 17972 29684 17978 29748
rect 20846 29684 20852 29748
rect 20916 29746 20922 29748
rect 20989 29746 21055 29749
rect 20916 29744 21055 29746
rect 20916 29688 20994 29744
rect 21050 29688 21055 29744
rect 20916 29686 21055 29688
rect 20916 29684 20922 29686
rect 20989 29683 21055 29686
rect 35065 29746 35131 29749
rect 35617 29746 35683 29749
rect 35065 29744 35683 29746
rect 35065 29688 35070 29744
rect 35126 29688 35622 29744
rect 35678 29688 35683 29744
rect 35065 29686 35683 29688
rect 35065 29683 35131 29686
rect 35617 29683 35683 29686
rect 2865 29610 2931 29613
rect 4613 29610 4679 29613
rect 2865 29608 4679 29610
rect 2865 29552 2870 29608
rect 2926 29552 4618 29608
rect 4674 29552 4679 29608
rect 2865 29550 4679 29552
rect 2865 29547 2931 29550
rect 4613 29547 4679 29550
rect 20805 29610 20871 29613
rect 27797 29610 27863 29613
rect 20805 29608 27863 29610
rect 20805 29552 20810 29608
rect 20866 29552 27802 29608
rect 27858 29552 27863 29608
rect 20805 29550 27863 29552
rect 20805 29547 20871 29550
rect 27797 29547 27863 29550
rect 33961 29610 34027 29613
rect 40861 29610 40927 29613
rect 33961 29608 40927 29610
rect 33961 29552 33966 29608
rect 34022 29552 40866 29608
rect 40922 29552 40927 29608
rect 33961 29550 40927 29552
rect 33961 29547 34027 29550
rect 40861 29547 40927 29550
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 17125 29338 17191 29341
rect 17677 29338 17743 29341
rect 17125 29336 17743 29338
rect 17125 29280 17130 29336
rect 17186 29280 17682 29336
rect 17738 29280 17743 29336
rect 17125 29278 17743 29280
rect 17125 29275 17191 29278
rect 17677 29275 17743 29278
rect 18229 29340 18295 29341
rect 18229 29336 18276 29340
rect 18340 29338 18346 29340
rect 28993 29338 29059 29341
rect 34973 29338 35039 29341
rect 18229 29280 18234 29336
rect 18229 29276 18276 29280
rect 18340 29278 18386 29338
rect 28993 29336 35039 29338
rect 28993 29280 28998 29336
rect 29054 29280 34978 29336
rect 35034 29280 35039 29336
rect 28993 29278 35039 29280
rect 18340 29276 18346 29278
rect 18229 29275 18295 29276
rect 28993 29275 29059 29278
rect 34973 29275 35039 29278
rect 42057 29338 42123 29341
rect 42843 29338 43643 29368
rect 42057 29336 43643 29338
rect 42057 29280 42062 29336
rect 42118 29280 43643 29336
rect 42057 29278 43643 29280
rect 42057 29275 42123 29278
rect 42843 29248 43643 29278
rect 12525 29204 12591 29205
rect 12525 29200 12572 29204
rect 12636 29202 12642 29204
rect 17493 29202 17559 29205
rect 21909 29204 21975 29205
rect 21909 29202 21956 29204
rect 12525 29144 12530 29200
rect 12525 29140 12572 29144
rect 12636 29142 12682 29202
rect 17493 29200 17602 29202
rect 17493 29144 17498 29200
rect 17554 29144 17602 29200
rect 12636 29140 12642 29142
rect 12525 29139 12591 29140
rect 17493 29139 17602 29144
rect 21864 29200 21956 29202
rect 21864 29144 21914 29200
rect 21864 29142 21956 29144
rect 21909 29140 21956 29142
rect 22020 29140 22026 29204
rect 34053 29202 34119 29205
rect 26926 29200 34119 29202
rect 26926 29144 34058 29200
rect 34114 29144 34119 29200
rect 26926 29142 34119 29144
rect 21909 29139 21975 29140
rect 12525 29066 12591 29069
rect 15653 29066 15719 29069
rect 12525 29064 15719 29066
rect 12525 29008 12530 29064
rect 12586 29008 15658 29064
rect 15714 29008 15719 29064
rect 12525 29006 15719 29008
rect 12525 29003 12591 29006
rect 15653 29003 15719 29006
rect 16941 29066 17007 29069
rect 17542 29066 17602 29139
rect 26926 29066 26986 29142
rect 34053 29139 34119 29142
rect 34605 29202 34671 29205
rect 38377 29202 38443 29205
rect 34605 29200 38443 29202
rect 34605 29144 34610 29200
rect 34666 29144 38382 29200
rect 38438 29144 38443 29200
rect 34605 29142 38443 29144
rect 34605 29139 34671 29142
rect 38377 29139 38443 29142
rect 16941 29064 26986 29066
rect 16941 29008 16946 29064
rect 17002 29008 26986 29064
rect 16941 29006 26986 29008
rect 30925 29066 30991 29069
rect 30925 29064 35450 29066
rect 30925 29008 30930 29064
rect 30986 29008 35450 29064
rect 30925 29006 35450 29008
rect 16941 29003 17007 29006
rect 30925 29003 30991 29006
rect 33041 28930 33107 28933
rect 33869 28930 33935 28933
rect 33041 28928 33935 28930
rect 33041 28872 33046 28928
rect 33102 28872 33874 28928
rect 33930 28872 33935 28928
rect 33041 28870 33935 28872
rect 35390 28930 35450 29006
rect 40033 28930 40099 28933
rect 35390 28928 40099 28930
rect 35390 28872 40038 28928
rect 40094 28872 40099 28928
rect 35390 28870 40099 28872
rect 33041 28867 33107 28870
rect 33869 28867 33935 28870
rect 40033 28867 40099 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 20989 28796 21055 28797
rect 20989 28794 21036 28796
rect 20944 28792 21036 28794
rect 20944 28736 20994 28792
rect 20944 28734 21036 28736
rect 20989 28732 21036 28734
rect 21100 28732 21106 28796
rect 20989 28731 21055 28732
rect 26049 28660 26115 28661
rect 25998 28596 26004 28660
rect 26068 28658 26115 28660
rect 28901 28658 28967 28661
rect 41873 28658 41939 28661
rect 26068 28656 26160 28658
rect 26110 28600 26160 28656
rect 26068 28598 26160 28600
rect 28901 28656 41939 28658
rect 28901 28600 28906 28656
rect 28962 28600 41878 28656
rect 41934 28600 41939 28656
rect 28901 28598 41939 28600
rect 26068 28596 26115 28598
rect 26049 28595 26115 28596
rect 28901 28595 28967 28598
rect 41873 28595 41939 28598
rect 42057 28658 42123 28661
rect 42843 28658 43643 28688
rect 42057 28656 43643 28658
rect 42057 28600 42062 28656
rect 42118 28600 43643 28656
rect 42057 28598 43643 28600
rect 42057 28595 42123 28598
rect 42843 28568 43643 28598
rect 33409 28522 33475 28525
rect 34053 28522 34119 28525
rect 33409 28520 34119 28522
rect 33409 28464 33414 28520
rect 33470 28464 34058 28520
rect 34114 28464 34119 28520
rect 33409 28462 34119 28464
rect 33409 28459 33475 28462
rect 34053 28459 34119 28462
rect 35065 28522 35131 28525
rect 36537 28522 36603 28525
rect 35065 28520 36603 28522
rect 35065 28464 35070 28520
rect 35126 28464 36542 28520
rect 36598 28464 36603 28520
rect 35065 28462 36603 28464
rect 35065 28459 35131 28462
rect 36537 28459 36603 28462
rect 12249 28386 12315 28389
rect 13813 28386 13879 28389
rect 12249 28384 13879 28386
rect 12249 28328 12254 28384
rect 12310 28328 13818 28384
rect 13874 28328 13879 28384
rect 12249 28326 13879 28328
rect 12249 28323 12315 28326
rect 13813 28323 13879 28326
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 12433 28250 12499 28253
rect 13537 28250 13603 28253
rect 12433 28248 13603 28250
rect 12433 28192 12438 28248
rect 12494 28192 13542 28248
rect 13598 28192 13603 28248
rect 12433 28190 13603 28192
rect 12433 28187 12499 28190
rect 13537 28187 13603 28190
rect 32765 28250 32831 28253
rect 33685 28250 33751 28253
rect 32765 28248 33751 28250
rect 32765 28192 32770 28248
rect 32826 28192 33690 28248
rect 33746 28192 33751 28248
rect 32765 28190 33751 28192
rect 32765 28187 32831 28190
rect 33685 28187 33751 28190
rect 11973 28114 12039 28117
rect 13353 28114 13419 28117
rect 11973 28112 13419 28114
rect 11973 28056 11978 28112
rect 12034 28056 13358 28112
rect 13414 28056 13419 28112
rect 11973 28054 13419 28056
rect 11973 28051 12039 28054
rect 13353 28051 13419 28054
rect 15193 28114 15259 28117
rect 16389 28114 16455 28117
rect 15193 28112 16455 28114
rect 15193 28056 15198 28112
rect 15254 28056 16394 28112
rect 16450 28056 16455 28112
rect 15193 28054 16455 28056
rect 15193 28051 15259 28054
rect 16389 28051 16455 28054
rect 19333 28114 19399 28117
rect 19701 28114 19767 28117
rect 34329 28114 34395 28117
rect 19333 28112 34395 28114
rect 19333 28056 19338 28112
rect 19394 28056 19706 28112
rect 19762 28056 34334 28112
rect 34390 28056 34395 28112
rect 19333 28054 34395 28056
rect 19333 28051 19399 28054
rect 19701 28051 19767 28054
rect 34329 28051 34395 28054
rect 12985 27978 13051 27981
rect 13905 27978 13971 27981
rect 12985 27976 13971 27978
rect 12985 27920 12990 27976
rect 13046 27920 13910 27976
rect 13966 27920 13971 27976
rect 12985 27918 13971 27920
rect 12985 27915 13051 27918
rect 13905 27915 13971 27918
rect 24301 27978 24367 27981
rect 38929 27978 38995 27981
rect 24301 27976 38995 27978
rect 24301 27920 24306 27976
rect 24362 27920 38934 27976
rect 38990 27920 38995 27976
rect 24301 27918 38995 27920
rect 24301 27915 24367 27918
rect 38929 27915 38995 27918
rect 41689 27978 41755 27981
rect 42843 27978 43643 28008
rect 41689 27976 43643 27978
rect 41689 27920 41694 27976
rect 41750 27920 43643 27976
rect 41689 27918 43643 27920
rect 41689 27915 41755 27918
rect 42843 27888 43643 27918
rect 12893 27842 12959 27845
rect 13445 27842 13511 27845
rect 14549 27842 14615 27845
rect 12893 27840 14615 27842
rect 12893 27784 12898 27840
rect 12954 27784 13450 27840
rect 13506 27784 14554 27840
rect 14610 27784 14615 27840
rect 12893 27782 14615 27784
rect 12893 27779 12959 27782
rect 13445 27779 13511 27782
rect 14549 27779 14615 27782
rect 28809 27842 28875 27845
rect 31201 27842 31267 27845
rect 28809 27840 31267 27842
rect 28809 27784 28814 27840
rect 28870 27784 31206 27840
rect 31262 27784 31267 27840
rect 28809 27782 31267 27784
rect 28809 27779 28875 27782
rect 31201 27779 31267 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 12709 27706 12775 27709
rect 13905 27706 13971 27709
rect 12709 27704 13971 27706
rect 12709 27648 12714 27704
rect 12770 27648 13910 27704
rect 13966 27648 13971 27704
rect 12709 27646 13971 27648
rect 12709 27643 12775 27646
rect 13905 27643 13971 27646
rect 12566 27508 12572 27572
rect 12636 27570 12642 27572
rect 12709 27570 12775 27573
rect 21173 27570 21239 27573
rect 12636 27568 21239 27570
rect 12636 27512 12714 27568
rect 12770 27512 21178 27568
rect 21234 27512 21239 27568
rect 12636 27510 21239 27512
rect 12636 27508 12642 27510
rect 12709 27507 12775 27510
rect 21173 27507 21239 27510
rect 30833 27570 30899 27573
rect 37917 27570 37983 27573
rect 38745 27570 38811 27573
rect 30833 27568 37983 27570
rect 30833 27512 30838 27568
rect 30894 27512 37922 27568
rect 37978 27512 37983 27568
rect 30833 27510 37983 27512
rect 30833 27507 30899 27510
rect 37917 27507 37983 27510
rect 38702 27568 38811 27570
rect 38702 27512 38750 27568
rect 38806 27512 38811 27568
rect 38702 27507 38811 27512
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 38702 27165 38762 27507
rect 41505 27298 41571 27301
rect 42843 27298 43643 27328
rect 41505 27296 43643 27298
rect 41505 27240 41510 27296
rect 41566 27240 43643 27296
rect 41505 27238 43643 27240
rect 41505 27235 41571 27238
rect 42843 27208 43643 27238
rect 38702 27160 38811 27165
rect 38702 27104 38750 27160
rect 38806 27104 38811 27160
rect 38702 27102 38811 27104
rect 38745 27099 38811 27102
rect 841 26754 907 26757
rect 798 26752 907 26754
rect 798 26696 846 26752
rect 902 26696 907 26752
rect 798 26691 907 26696
rect 798 26648 858 26691
rect 0 26558 858 26648
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 41873 26618 41939 26621
rect 42843 26618 43643 26648
rect 41873 26616 43643 26618
rect 41873 26560 41878 26616
rect 41934 26560 43643 26616
rect 41873 26558 43643 26560
rect 0 26528 800 26558
rect 41873 26555 41939 26558
rect 42843 26528 43643 26558
rect 12249 26482 12315 26485
rect 15193 26482 15259 26485
rect 12249 26480 15259 26482
rect 12249 26424 12254 26480
rect 12310 26424 15198 26480
rect 15254 26424 15259 26480
rect 12249 26422 15259 26424
rect 12249 26419 12315 26422
rect 15193 26419 15259 26422
rect 3969 26346 4035 26349
rect 5165 26346 5231 26349
rect 3969 26344 5231 26346
rect 3969 26288 3974 26344
rect 4030 26288 5170 26344
rect 5226 26288 5231 26344
rect 3969 26286 5231 26288
rect 3969 26283 4035 26286
rect 5165 26283 5231 26286
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 25037 25938 25103 25941
rect 25681 25938 25747 25941
rect 25037 25936 25747 25938
rect 25037 25880 25042 25936
rect 25098 25880 25686 25936
rect 25742 25880 25747 25936
rect 25037 25878 25747 25880
rect 25037 25875 25103 25878
rect 25681 25875 25747 25878
rect 42057 25938 42123 25941
rect 42843 25938 43643 25968
rect 42057 25936 43643 25938
rect 42057 25880 42062 25936
rect 42118 25880 43643 25936
rect 42057 25878 43643 25880
rect 42057 25875 42123 25878
rect 42843 25848 43643 25878
rect 23473 25802 23539 25805
rect 25405 25802 25471 25805
rect 28717 25802 28783 25805
rect 23473 25800 28783 25802
rect 23473 25744 23478 25800
rect 23534 25744 25410 25800
rect 25466 25744 28722 25800
rect 28778 25744 28783 25800
rect 23473 25742 28783 25744
rect 23473 25739 23539 25742
rect 25405 25739 25471 25742
rect 28717 25739 28783 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 16573 25394 16639 25397
rect 17401 25394 17467 25397
rect 16573 25392 17467 25394
rect 16573 25336 16578 25392
rect 16634 25336 17406 25392
rect 17462 25336 17467 25392
rect 16573 25334 17467 25336
rect 16573 25331 16639 25334
rect 17401 25331 17467 25334
rect 18689 25394 18755 25397
rect 32673 25394 32739 25397
rect 18689 25392 32739 25394
rect 18689 25336 18694 25392
rect 18750 25336 32678 25392
rect 32734 25336 32739 25392
rect 18689 25334 32739 25336
rect 18689 25331 18755 25334
rect 32673 25331 32739 25334
rect 15469 25258 15535 25261
rect 17953 25258 18019 25261
rect 15469 25256 18019 25258
rect 15469 25200 15474 25256
rect 15530 25200 17958 25256
rect 18014 25200 18019 25256
rect 15469 25198 18019 25200
rect 15469 25195 15535 25198
rect 17953 25195 18019 25198
rect 30741 25258 30807 25261
rect 35893 25258 35959 25261
rect 30741 25256 35959 25258
rect 30741 25200 30746 25256
rect 30802 25200 35898 25256
rect 35954 25200 35959 25256
rect 30741 25198 35959 25200
rect 30741 25195 30807 25198
rect 35893 25195 35959 25198
rect 37273 25258 37339 25261
rect 38377 25258 38443 25261
rect 37273 25256 38443 25258
rect 37273 25200 37278 25256
rect 37334 25200 38382 25256
rect 38438 25200 38443 25256
rect 37273 25198 38443 25200
rect 37273 25195 37339 25198
rect 38377 25195 38443 25198
rect 40125 25258 40191 25261
rect 42843 25258 43643 25288
rect 40125 25256 43643 25258
rect 40125 25200 40130 25256
rect 40186 25200 43643 25256
rect 40125 25198 43643 25200
rect 40125 25195 40191 25198
rect 42843 25168 43643 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 7557 24850 7623 24853
rect 9581 24850 9647 24853
rect 7557 24848 9647 24850
rect 7557 24792 7562 24848
rect 7618 24792 9586 24848
rect 9642 24792 9647 24848
rect 7557 24790 9647 24792
rect 7557 24787 7623 24790
rect 9581 24787 9647 24790
rect 15561 24850 15627 24853
rect 15694 24850 15700 24852
rect 15561 24848 15700 24850
rect 15561 24792 15566 24848
rect 15622 24792 15700 24848
rect 15561 24790 15700 24792
rect 15561 24787 15627 24790
rect 15694 24788 15700 24790
rect 15764 24788 15770 24852
rect 17769 24850 17835 24853
rect 18270 24850 18276 24852
rect 17769 24848 18276 24850
rect 17769 24792 17774 24848
rect 17830 24792 18276 24848
rect 17769 24790 18276 24792
rect 17769 24787 17835 24790
rect 18270 24788 18276 24790
rect 18340 24850 18346 24852
rect 18689 24850 18755 24853
rect 18340 24848 18755 24850
rect 18340 24792 18694 24848
rect 18750 24792 18755 24848
rect 18340 24790 18755 24792
rect 18340 24788 18346 24790
rect 18689 24787 18755 24790
rect 23565 24850 23631 24853
rect 24485 24850 24551 24853
rect 25037 24850 25103 24853
rect 23565 24848 25103 24850
rect 23565 24792 23570 24848
rect 23626 24792 24490 24848
rect 24546 24792 25042 24848
rect 25098 24792 25103 24848
rect 23565 24790 25103 24792
rect 23565 24787 23631 24790
rect 24485 24787 24551 24790
rect 25037 24787 25103 24790
rect 34881 24850 34947 24853
rect 35433 24850 35499 24853
rect 34881 24848 35499 24850
rect 34881 24792 34886 24848
rect 34942 24792 35438 24848
rect 35494 24792 35499 24848
rect 34881 24790 35499 24792
rect 34881 24787 34947 24790
rect 35433 24787 35499 24790
rect 17033 24714 17099 24717
rect 17677 24714 17743 24717
rect 23197 24714 23263 24717
rect 17033 24712 23263 24714
rect 17033 24656 17038 24712
rect 17094 24656 17682 24712
rect 17738 24656 23202 24712
rect 23258 24656 23263 24712
rect 17033 24654 23263 24656
rect 17033 24651 17099 24654
rect 17677 24651 17743 24654
rect 23197 24651 23263 24654
rect 35341 24712 35407 24717
rect 35341 24656 35346 24712
rect 35402 24656 35407 24712
rect 35341 24651 35407 24656
rect 35344 24578 35404 24651
rect 36169 24578 36235 24581
rect 35344 24576 36235 24578
rect 35344 24520 36174 24576
rect 36230 24520 36235 24576
rect 35344 24518 36235 24520
rect 36169 24515 36235 24518
rect 40585 24578 40651 24581
rect 42843 24578 43643 24608
rect 40585 24576 43643 24578
rect 40585 24520 40590 24576
rect 40646 24520 43643 24576
rect 40585 24518 43643 24520
rect 40585 24515 40651 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 42843 24488 43643 24518
rect 34930 24447 35246 24448
rect 18229 24306 18295 24309
rect 19241 24306 19307 24309
rect 18229 24304 19307 24306
rect 18229 24248 18234 24304
rect 18290 24248 19246 24304
rect 19302 24248 19307 24304
rect 18229 24246 19307 24248
rect 18229 24243 18295 24246
rect 19241 24243 19307 24246
rect 18137 24170 18203 24173
rect 18413 24170 18479 24173
rect 19287 24170 19353 24173
rect 18137 24168 19353 24170
rect 18137 24112 18142 24168
rect 18198 24112 18418 24168
rect 18474 24112 19292 24168
rect 19348 24112 19353 24168
rect 18137 24110 19353 24112
rect 18137 24107 18203 24110
rect 18413 24107 18479 24110
rect 19287 24107 19353 24110
rect 34329 24170 34395 24173
rect 35525 24170 35591 24173
rect 34329 24168 35591 24170
rect 34329 24112 34334 24168
rect 34390 24112 35530 24168
rect 35586 24112 35591 24168
rect 34329 24110 35591 24112
rect 34329 24107 34395 24110
rect 35525 24107 35591 24110
rect 13353 24034 13419 24037
rect 19241 24034 19307 24037
rect 13353 24032 19307 24034
rect 13353 23976 13358 24032
rect 13414 23976 19246 24032
rect 19302 23976 19307 24032
rect 13353 23974 19307 23976
rect 13353 23971 13419 23974
rect 19241 23971 19307 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 18321 23898 18387 23901
rect 19149 23898 19215 23901
rect 18321 23896 19215 23898
rect 18321 23840 18326 23896
rect 18382 23840 19154 23896
rect 19210 23840 19215 23896
rect 18321 23838 19215 23840
rect 18321 23835 18387 23838
rect 19149 23835 19215 23838
rect 16389 23762 16455 23765
rect 25497 23762 25563 23765
rect 16389 23760 25563 23762
rect 16389 23704 16394 23760
rect 16450 23704 25502 23760
rect 25558 23704 25563 23760
rect 16389 23702 25563 23704
rect 16389 23699 16455 23702
rect 25497 23699 25563 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 6821 23218 6887 23221
rect 8293 23218 8359 23221
rect 6821 23216 8359 23218
rect 6821 23160 6826 23216
rect 6882 23160 8298 23216
rect 8354 23160 8359 23216
rect 6821 23158 8359 23160
rect 6821 23155 6887 23158
rect 8293 23155 8359 23158
rect 25630 22884 25636 22948
rect 25700 22946 25706 22948
rect 25773 22946 25839 22949
rect 25700 22944 25839 22946
rect 25700 22888 25778 22944
rect 25834 22888 25839 22944
rect 25700 22886 25839 22888
rect 25700 22884 25706 22886
rect 25773 22883 25839 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 841 22674 907 22677
rect 798 22672 907 22674
rect 798 22616 846 22672
rect 902 22616 907 22672
rect 798 22611 907 22616
rect 798 22568 858 22611
rect 0 22478 858 22568
rect 32765 22540 32831 22541
rect 32765 22538 32812 22540
rect 32720 22536 32812 22538
rect 32720 22480 32770 22536
rect 32720 22478 32812 22480
rect 0 22448 800 22478
rect 32765 22476 32812 22478
rect 32876 22476 32882 22540
rect 32765 22475 32831 22476
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 4521 22130 4587 22133
rect 5073 22130 5139 22133
rect 4521 22128 5139 22130
rect 4521 22072 4526 22128
rect 4582 22072 5078 22128
rect 5134 22072 5139 22128
rect 4521 22070 5139 22072
rect 4521 22067 4587 22070
rect 5073 22067 5139 22070
rect 18597 21996 18663 21997
rect 18597 21994 18644 21996
rect 18552 21992 18644 21994
rect 18552 21936 18602 21992
rect 18552 21934 18644 21936
rect 18597 21932 18644 21934
rect 18708 21932 18714 21996
rect 21633 21994 21699 21997
rect 21766 21994 21772 21996
rect 21633 21992 21772 21994
rect 21633 21936 21638 21992
rect 21694 21936 21772 21992
rect 21633 21934 21772 21936
rect 18597 21931 18663 21932
rect 21633 21931 21699 21934
rect 21766 21932 21772 21934
rect 21836 21932 21842 21996
rect 0 21858 800 21888
rect 1301 21858 1367 21861
rect 24945 21860 25011 21861
rect 0 21856 1367 21858
rect 0 21800 1306 21856
rect 1362 21800 1367 21856
rect 0 21798 1367 21800
rect 0 21768 800 21798
rect 1301 21795 1367 21798
rect 24894 21796 24900 21860
rect 24964 21858 25011 21860
rect 24964 21856 25056 21858
rect 25006 21800 25056 21856
rect 24964 21798 25056 21800
rect 24964 21796 25011 21798
rect 24945 21795 25011 21796
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 1025 21178 1091 21181
rect 0 21176 1091 21178
rect 0 21120 1030 21176
rect 1086 21120 1091 21176
rect 0 21118 1091 21120
rect 0 21088 800 21118
rect 1025 21115 1091 21118
rect 34605 21042 34671 21045
rect 34973 21042 35039 21045
rect 34605 21040 35039 21042
rect 34605 20984 34610 21040
rect 34666 20984 34978 21040
rect 35034 20984 35039 21040
rect 34605 20982 35039 20984
rect 34605 20979 34671 20982
rect 34973 20979 35039 20982
rect 38009 20770 38075 20773
rect 38142 20770 38148 20772
rect 38009 20768 38148 20770
rect 38009 20712 38014 20768
rect 38070 20712 38148 20768
rect 38009 20710 38148 20712
rect 38009 20707 38075 20710
rect 38142 20708 38148 20710
rect 38212 20708 38218 20772
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 9581 18730 9647 18733
rect 12525 18730 12591 18733
rect 9581 18728 12591 18730
rect 9581 18672 9586 18728
rect 9642 18672 12530 18728
rect 12586 18672 12591 18728
rect 9581 18670 12591 18672
rect 9581 18667 9647 18670
rect 12525 18667 12591 18670
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 27521 17234 27587 17237
rect 28441 17234 28507 17237
rect 27521 17232 28507 17234
rect 27521 17176 27526 17232
rect 27582 17176 28446 17232
rect 28502 17176 28507 17232
rect 27521 17174 28507 17176
rect 27521 17171 27587 17174
rect 28441 17171 28507 17174
rect 0 17098 800 17128
rect 19149 17098 19215 17101
rect 19425 17098 19491 17101
rect 0 17008 858 17098
rect 19149 17096 19491 17098
rect 19149 17040 19154 17096
rect 19210 17040 19430 17096
rect 19486 17040 19491 17096
rect 19149 17038 19491 17040
rect 19149 17035 19215 17038
rect 19425 17035 19491 17038
rect 798 16965 858 17008
rect 798 16960 907 16965
rect 798 16904 846 16960
rect 902 16904 907 16960
rect 798 16902 907 16904
rect 841 16899 907 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 28441 16826 28507 16829
rect 28901 16826 28967 16829
rect 28441 16824 28967 16826
rect 28441 16768 28446 16824
rect 28502 16768 28906 16824
rect 28962 16768 28967 16824
rect 28441 16766 28967 16768
rect 28441 16763 28507 16766
rect 28901 16763 28967 16766
rect 30925 16554 30991 16557
rect 32121 16554 32187 16557
rect 30925 16552 32187 16554
rect 30925 16496 30930 16552
rect 30986 16496 32126 16552
rect 32182 16496 32187 16552
rect 30925 16494 32187 16496
rect 30925 16491 30991 16494
rect 32121 16491 32187 16494
rect 23565 16418 23631 16421
rect 25957 16418 26023 16421
rect 23565 16416 26023 16418
rect 23565 16360 23570 16416
rect 23626 16360 25962 16416
rect 26018 16360 26023 16416
rect 23565 16358 26023 16360
rect 23565 16355 23631 16358
rect 25957 16355 26023 16358
rect 31661 16418 31727 16421
rect 33317 16418 33383 16421
rect 31661 16416 33383 16418
rect 31661 16360 31666 16416
rect 31722 16360 33322 16416
rect 33378 16360 33383 16416
rect 31661 16358 33383 16360
rect 31661 16355 31727 16358
rect 33317 16355 33383 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 28993 16282 29059 16285
rect 29177 16282 29243 16285
rect 28993 16280 29243 16282
rect 28993 16224 28998 16280
rect 29054 16224 29182 16280
rect 29238 16224 29243 16280
rect 28993 16222 29243 16224
rect 28993 16219 29059 16222
rect 29177 16219 29243 16222
rect 30557 16282 30623 16285
rect 33133 16282 33199 16285
rect 30557 16280 33199 16282
rect 30557 16224 30562 16280
rect 30618 16224 33138 16280
rect 33194 16224 33199 16280
rect 30557 16222 33199 16224
rect 30557 16219 30623 16222
rect 33133 16219 33199 16222
rect 18965 16146 19031 16149
rect 18965 16144 19350 16146
rect 18965 16088 18970 16144
rect 19026 16088 19350 16144
rect 18965 16086 19350 16088
rect 18965 16083 19031 16086
rect 19290 16010 19350 16086
rect 19517 16010 19583 16013
rect 20161 16010 20227 16013
rect 19290 16008 20227 16010
rect 19290 15952 19522 16008
rect 19578 15952 20166 16008
rect 20222 15952 20227 16008
rect 19290 15950 20227 15952
rect 19517 15947 19583 15950
rect 20161 15947 20227 15950
rect 30281 16010 30347 16013
rect 32489 16010 32555 16013
rect 34237 16010 34303 16013
rect 30281 16008 34303 16010
rect 30281 15952 30286 16008
rect 30342 15952 32494 16008
rect 32550 15952 34242 16008
rect 34298 15952 34303 16008
rect 30281 15950 34303 15952
rect 30281 15947 30347 15950
rect 32489 15947 32555 15950
rect 34237 15947 34303 15950
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 0 15648 800 15678
rect 29913 15466 29979 15469
rect 30465 15466 30531 15469
rect 29913 15464 30531 15466
rect 29913 15408 29918 15464
rect 29974 15408 30470 15464
rect 30526 15408 30531 15464
rect 29913 15406 30531 15408
rect 29913 15403 29979 15406
rect 30465 15403 30531 15406
rect 38142 15404 38148 15468
rect 38212 15466 38218 15468
rect 38285 15466 38351 15469
rect 38212 15464 38351 15466
rect 38212 15408 38290 15464
rect 38346 15408 38351 15464
rect 38212 15406 38351 15408
rect 38212 15404 38218 15406
rect 38285 15403 38351 15406
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 29177 15194 29243 15197
rect 30557 15194 30623 15197
rect 29177 15192 30623 15194
rect 29177 15136 29182 15192
rect 29238 15136 30562 15192
rect 30618 15136 30623 15192
rect 29177 15134 30623 15136
rect 29177 15131 29243 15134
rect 30557 15131 30623 15134
rect 0 15058 800 15088
rect 1669 15058 1735 15061
rect 0 15056 1735 15058
rect 0 15000 1674 15056
rect 1730 15000 1735 15056
rect 0 14998 1735 15000
rect 0 14968 800 14998
rect 1669 14995 1735 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 32806 13772 32812 13836
rect 32876 13834 32882 13836
rect 34881 13834 34947 13837
rect 32876 13832 34947 13834
rect 32876 13776 34886 13832
rect 34942 13776 34947 13832
rect 32876 13774 34947 13776
rect 32876 13772 32882 13774
rect 34881 13771 34947 13774
rect 24894 13636 24900 13700
rect 24964 13698 24970 13700
rect 25037 13698 25103 13701
rect 25681 13700 25747 13701
rect 25630 13698 25636 13700
rect 24964 13696 25103 13698
rect 24964 13640 25042 13696
rect 25098 13640 25103 13696
rect 24964 13638 25103 13640
rect 25590 13638 25636 13698
rect 25700 13696 25747 13700
rect 25742 13640 25747 13696
rect 24964 13636 24970 13638
rect 25037 13635 25103 13638
rect 25630 13636 25636 13638
rect 25700 13636 25747 13640
rect 25681 13635 25747 13636
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 34421 13426 34487 13429
rect 36353 13426 36419 13429
rect 34421 13424 36419 13426
rect 34421 13368 34426 13424
rect 34482 13368 36358 13424
rect 36414 13368 36419 13424
rect 34421 13366 36419 13368
rect 34421 13363 34487 13366
rect 36353 13363 36419 13366
rect 34973 13290 35039 13293
rect 35985 13290 36051 13293
rect 34973 13288 36051 13290
rect 34973 13232 34978 13288
rect 35034 13232 35990 13288
rect 36046 13232 36051 13288
rect 34973 13230 36051 13232
rect 34973 13227 35039 13230
rect 35985 13227 36051 13230
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 35157 12882 35223 12885
rect 35341 12882 35407 12885
rect 37089 12882 37155 12885
rect 35157 12880 37155 12882
rect 35157 12824 35162 12880
rect 35218 12824 35346 12880
rect 35402 12824 37094 12880
rect 37150 12824 37155 12880
rect 35157 12822 37155 12824
rect 35157 12819 35223 12822
rect 35341 12819 35407 12822
rect 37089 12819 37155 12822
rect 19701 12746 19767 12749
rect 23565 12746 23631 12749
rect 19701 12744 23631 12746
rect 19701 12688 19706 12744
rect 19762 12688 23570 12744
rect 23626 12688 23631 12744
rect 19701 12686 23631 12688
rect 19701 12683 19767 12686
rect 23565 12683 23631 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 21357 12338 21423 12341
rect 26877 12338 26943 12341
rect 21357 12336 26943 12338
rect 21357 12280 21362 12336
rect 21418 12280 26882 12336
rect 26938 12280 26943 12336
rect 21357 12278 26943 12280
rect 21357 12275 21423 12278
rect 26877 12275 26943 12278
rect 22829 12202 22895 12205
rect 23473 12202 23539 12205
rect 22829 12200 23539 12202
rect 22829 12144 22834 12200
rect 22890 12144 23478 12200
rect 23534 12144 23539 12200
rect 22829 12142 23539 12144
rect 22829 12139 22895 12142
rect 23473 12139 23539 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 4245 11794 4311 11797
rect 4705 11794 4771 11797
rect 5349 11794 5415 11797
rect 4245 11792 5415 11794
rect 4245 11736 4250 11792
rect 4306 11736 4710 11792
rect 4766 11736 5354 11792
rect 5410 11736 5415 11792
rect 4245 11734 5415 11736
rect 4245 11731 4311 11734
rect 4705 11731 4771 11734
rect 5349 11731 5415 11734
rect 0 11658 800 11688
rect 4429 11658 4495 11661
rect 6729 11658 6795 11661
rect 0 11568 858 11658
rect 4429 11656 6795 11658
rect 4429 11600 4434 11656
rect 4490 11600 6734 11656
rect 6790 11600 6795 11656
rect 4429 11598 6795 11600
rect 4429 11595 4495 11598
rect 6729 11595 6795 11598
rect 798 11525 858 11568
rect 798 11520 907 11525
rect 798 11464 846 11520
rect 902 11464 907 11520
rect 798 11462 907 11464
rect 841 11459 907 11462
rect 9581 11520 9647 11525
rect 9581 11464 9586 11520
rect 9642 11464 9647 11520
rect 9581 11459 9647 11464
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 9584 11117 9644 11459
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 9581 11112 9647 11117
rect 9581 11056 9586 11112
rect 9642 11056 9647 11112
rect 9581 11051 9647 11056
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 20161 10978 20227 10981
rect 20897 10978 20963 10981
rect 20161 10976 20963 10978
rect 20161 10920 20166 10976
rect 20222 10920 20902 10976
rect 20958 10920 20963 10976
rect 20161 10918 20963 10920
rect 20161 10915 20227 10918
rect 20897 10915 20963 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 25589 10706 25655 10709
rect 28257 10706 28323 10709
rect 25589 10704 28323 10706
rect 25589 10648 25594 10704
rect 25650 10648 28262 10704
rect 28318 10648 28323 10704
rect 25589 10646 28323 10648
rect 25589 10643 25655 10646
rect 28257 10643 28323 10646
rect 34145 10706 34211 10709
rect 34973 10706 35039 10709
rect 36445 10706 36511 10709
rect 36997 10706 37063 10709
rect 34145 10704 37063 10706
rect 34145 10648 34150 10704
rect 34206 10648 34978 10704
rect 35034 10648 36450 10704
rect 36506 10648 37002 10704
rect 37058 10648 37063 10704
rect 34145 10646 37063 10648
rect 34145 10643 34211 10646
rect 34973 10643 35039 10646
rect 36445 10643 36511 10646
rect 36997 10643 37063 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 26601 9618 26667 9621
rect 27337 9618 27403 9621
rect 26601 9616 27403 9618
rect 26601 9560 26606 9616
rect 26662 9560 27342 9616
rect 27398 9560 27403 9616
rect 26601 9558 27403 9560
rect 26601 9555 26667 9558
rect 27337 9555 27403 9558
rect 26233 9482 26299 9485
rect 27061 9482 27127 9485
rect 26233 9480 27127 9482
rect 26233 9424 26238 9480
rect 26294 9424 27066 9480
rect 27122 9424 27127 9480
rect 26233 9422 27127 9424
rect 26233 9419 26299 9422
rect 27061 9419 27127 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 3693 7986 3759 7989
rect 4521 7986 4587 7989
rect 3693 7984 4587 7986
rect 3693 7928 3698 7984
rect 3754 7928 4526 7984
rect 4582 7928 4587 7984
rect 3693 7926 4587 7928
rect 3693 7923 3759 7926
rect 4521 7923 4587 7926
rect 7833 7986 7899 7989
rect 9029 7986 9095 7989
rect 7833 7984 9095 7986
rect 7833 7928 7838 7984
rect 7894 7928 9034 7984
rect 9090 7928 9095 7984
rect 7833 7926 9095 7928
rect 7833 7923 7899 7926
rect 9029 7923 9095 7926
rect 7833 7850 7899 7853
rect 8293 7850 8359 7853
rect 7833 7848 8359 7850
rect 7833 7792 7838 7848
rect 7894 7792 8298 7848
rect 8354 7792 8359 7848
rect 7833 7790 8359 7792
rect 7833 7787 7899 7790
rect 8293 7787 8359 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 19793 7442 19859 7445
rect 23197 7442 23263 7445
rect 19793 7440 23263 7442
rect 19793 7384 19798 7440
rect 19854 7384 23202 7440
rect 23258 7384 23263 7440
rect 19793 7382 23263 7384
rect 19793 7379 19859 7382
rect 23197 7379 23263 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 42149 3498 42215 3501
rect 42843 3498 43643 3528
rect 42149 3496 43643 3498
rect 42149 3440 42154 3496
rect 42210 3440 43643 3496
rect 42149 3438 43643 3440
rect 42149 3435 42215 3438
rect 42843 3408 43643 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4876 43548 4940 43552
rect 4876 43492 4880 43548
rect 4880 43492 4936 43548
rect 4936 43492 4940 43548
rect 4876 43488 4940 43492
rect 4956 43548 5020 43552
rect 4956 43492 4960 43548
rect 4960 43492 5016 43548
rect 5016 43492 5020 43548
rect 4956 43488 5020 43492
rect 5036 43548 5100 43552
rect 5036 43492 5040 43548
rect 5040 43492 5096 43548
rect 5096 43492 5100 43548
rect 5036 43488 5100 43492
rect 5116 43548 5180 43552
rect 5116 43492 5120 43548
rect 5120 43492 5176 43548
rect 5176 43492 5180 43548
rect 5116 43488 5180 43492
rect 35596 43548 35660 43552
rect 35596 43492 35600 43548
rect 35600 43492 35656 43548
rect 35656 43492 35660 43548
rect 35596 43488 35660 43492
rect 35676 43548 35740 43552
rect 35676 43492 35680 43548
rect 35680 43492 35736 43548
rect 35736 43492 35740 43548
rect 35676 43488 35740 43492
rect 35756 43548 35820 43552
rect 35756 43492 35760 43548
rect 35760 43492 35816 43548
rect 35816 43492 35820 43548
rect 35756 43488 35820 43492
rect 35836 43548 35900 43552
rect 35836 43492 35840 43548
rect 35840 43492 35896 43548
rect 35896 43492 35900 43548
rect 35836 43488 35900 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 21036 42936 21100 42940
rect 21036 42880 21050 42936
rect 21050 42880 21100 42936
rect 21036 42876 21100 42880
rect 4876 42460 4940 42464
rect 4876 42404 4880 42460
rect 4880 42404 4936 42460
rect 4936 42404 4940 42460
rect 4876 42400 4940 42404
rect 4956 42460 5020 42464
rect 4956 42404 4960 42460
rect 4960 42404 5016 42460
rect 5016 42404 5020 42460
rect 4956 42400 5020 42404
rect 5036 42460 5100 42464
rect 5036 42404 5040 42460
rect 5040 42404 5096 42460
rect 5096 42404 5100 42460
rect 5036 42400 5100 42404
rect 5116 42460 5180 42464
rect 5116 42404 5120 42460
rect 5120 42404 5176 42460
rect 5176 42404 5180 42460
rect 5116 42400 5180 42404
rect 35596 42460 35660 42464
rect 35596 42404 35600 42460
rect 35600 42404 35656 42460
rect 35656 42404 35660 42460
rect 35596 42400 35660 42404
rect 35676 42460 35740 42464
rect 35676 42404 35680 42460
rect 35680 42404 35736 42460
rect 35736 42404 35740 42460
rect 35676 42400 35740 42404
rect 35756 42460 35820 42464
rect 35756 42404 35760 42460
rect 35760 42404 35816 42460
rect 35816 42404 35820 42460
rect 35756 42400 35820 42404
rect 35836 42460 35900 42464
rect 35836 42404 35840 42460
rect 35840 42404 35896 42460
rect 35896 42404 35900 42460
rect 35836 42400 35900 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 20852 41576 20916 41580
rect 20852 41520 20866 41576
rect 20866 41520 20916 41576
rect 20852 41516 20916 41520
rect 4876 41372 4940 41376
rect 4876 41316 4880 41372
rect 4880 41316 4936 41372
rect 4936 41316 4940 41372
rect 4876 41312 4940 41316
rect 4956 41372 5020 41376
rect 4956 41316 4960 41372
rect 4960 41316 5016 41372
rect 5016 41316 5020 41372
rect 4956 41312 5020 41316
rect 5036 41372 5100 41376
rect 5036 41316 5040 41372
rect 5040 41316 5096 41372
rect 5096 41316 5100 41372
rect 5036 41312 5100 41316
rect 5116 41372 5180 41376
rect 5116 41316 5120 41372
rect 5120 41316 5176 41372
rect 5176 41316 5180 41372
rect 5116 41312 5180 41316
rect 35596 41372 35660 41376
rect 35596 41316 35600 41372
rect 35600 41316 35656 41372
rect 35656 41316 35660 41372
rect 35596 41312 35660 41316
rect 35676 41372 35740 41376
rect 35676 41316 35680 41372
rect 35680 41316 35736 41372
rect 35736 41316 35740 41372
rect 35676 41312 35740 41316
rect 35756 41372 35820 41376
rect 35756 41316 35760 41372
rect 35760 41316 35816 41372
rect 35816 41316 35820 41372
rect 35756 41312 35820 41316
rect 35836 41372 35900 41376
rect 35836 41316 35840 41372
rect 35840 41316 35896 41372
rect 35896 41316 35900 41372
rect 35836 41312 35900 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 26004 40624 26068 40628
rect 26004 40568 26018 40624
rect 26018 40568 26068 40624
rect 26004 40564 26068 40568
rect 4876 40284 4940 40288
rect 4876 40228 4880 40284
rect 4880 40228 4936 40284
rect 4936 40228 4940 40284
rect 4876 40224 4940 40228
rect 4956 40284 5020 40288
rect 4956 40228 4960 40284
rect 4960 40228 5016 40284
rect 5016 40228 5020 40284
rect 4956 40224 5020 40228
rect 5036 40284 5100 40288
rect 5036 40228 5040 40284
rect 5040 40228 5096 40284
rect 5096 40228 5100 40284
rect 5036 40224 5100 40228
rect 5116 40284 5180 40288
rect 5116 40228 5120 40284
rect 5120 40228 5176 40284
rect 5176 40228 5180 40284
rect 5116 40224 5180 40228
rect 35596 40284 35660 40288
rect 35596 40228 35600 40284
rect 35600 40228 35656 40284
rect 35656 40228 35660 40284
rect 35596 40224 35660 40228
rect 35676 40284 35740 40288
rect 35676 40228 35680 40284
rect 35680 40228 35736 40284
rect 35736 40228 35740 40284
rect 35676 40224 35740 40228
rect 35756 40284 35820 40288
rect 35756 40228 35760 40284
rect 35760 40228 35816 40284
rect 35816 40228 35820 40284
rect 35756 40224 35820 40228
rect 35836 40284 35900 40288
rect 35836 40228 35840 40284
rect 35840 40228 35896 40284
rect 35896 40228 35900 40284
rect 35836 40224 35900 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 21956 39340 22020 39404
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 5396 34444 5460 34508
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 15700 31104 15764 31108
rect 15700 31048 15750 31104
rect 15750 31048 15764 31104
rect 15700 31044 15764 31048
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 5396 30696 5460 30700
rect 5396 30640 5446 30696
rect 5446 30640 5460 30696
rect 5396 30636 5460 30640
rect 17908 30636 17972 30700
rect 21772 30500 21836 30564
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 18644 30016 18708 30020
rect 18644 29960 18658 30016
rect 18658 29960 18708 30016
rect 18644 29956 18708 29960
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 17908 29684 17972 29748
rect 20852 29684 20916 29748
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 18276 29336 18340 29340
rect 18276 29280 18290 29336
rect 18290 29280 18340 29336
rect 18276 29276 18340 29280
rect 12572 29200 12636 29204
rect 12572 29144 12586 29200
rect 12586 29144 12636 29200
rect 12572 29140 12636 29144
rect 21956 29200 22020 29204
rect 21956 29144 21970 29200
rect 21970 29144 22020 29200
rect 21956 29140 22020 29144
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 21036 28792 21100 28796
rect 21036 28736 21050 28792
rect 21050 28736 21100 28792
rect 21036 28732 21100 28736
rect 26004 28656 26068 28660
rect 26004 28600 26054 28656
rect 26054 28600 26068 28656
rect 26004 28596 26068 28600
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 12572 27508 12636 27572
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 15700 24788 15764 24852
rect 18276 24788 18340 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 25636 22884 25700 22948
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 32812 22536 32876 22540
rect 32812 22480 32826 22536
rect 32826 22480 32876 22536
rect 32812 22476 32876 22480
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 18644 21992 18708 21996
rect 18644 21936 18658 21992
rect 18658 21936 18708 21992
rect 18644 21932 18708 21936
rect 21772 21932 21836 21996
rect 24900 21856 24964 21860
rect 24900 21800 24950 21856
rect 24950 21800 24964 21856
rect 24900 21796 24964 21800
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 38148 20708 38212 20772
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 38148 15404 38212 15468
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 32812 13772 32876 13836
rect 24900 13636 24964 13700
rect 25636 13696 25700 13700
rect 25636 13640 25686 13696
rect 25686 13640 25700 13696
rect 25636 13636 25700 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 43008 4528 43568
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 43552 5188 43568
rect 4868 43488 4876 43552
rect 4940 43488 4956 43552
rect 5020 43488 5036 43552
rect 5100 43488 5116 43552
rect 5180 43488 5188 43552
rect 4868 42464 5188 43488
rect 34928 43008 35248 43568
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 21035 42940 21101 42941
rect 21035 42876 21036 42940
rect 21100 42876 21101 42940
rect 21035 42875 21101 42876
rect 4868 42400 4876 42464
rect 4940 42400 4956 42464
rect 5020 42400 5036 42464
rect 5100 42400 5116 42464
rect 5180 42400 5188 42464
rect 4868 41376 5188 42400
rect 20851 41580 20917 41581
rect 20851 41516 20852 41580
rect 20916 41516 20917 41580
rect 20851 41515 20917 41516
rect 4868 41312 4876 41376
rect 4940 41312 4956 41376
rect 5020 41312 5036 41376
rect 5100 41312 5116 41376
rect 5180 41312 5188 41376
rect 4868 40288 5188 41312
rect 4868 40224 4876 40288
rect 4940 40224 4956 40288
rect 5020 40224 5036 40288
rect 5100 40224 5116 40288
rect 5180 40224 5188 40288
rect 4868 39200 5188 40224
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 5395 34508 5461 34509
rect 5395 34444 5396 34508
rect 5460 34444 5461 34508
rect 5395 34443 5461 34444
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 5398 30701 5458 34443
rect 15699 31108 15765 31109
rect 15699 31044 15700 31108
rect 15764 31044 15765 31108
rect 15699 31043 15765 31044
rect 5395 30700 5461 30701
rect 5395 30636 5396 30700
rect 5460 30636 5461 30700
rect 5395 30635 5461 30636
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 12571 29204 12637 29205
rect 12571 29140 12572 29204
rect 12636 29140 12637 29204
rect 12571 29139 12637 29140
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 12574 27573 12634 29139
rect 12571 27572 12637 27573
rect 12571 27508 12572 27572
rect 12636 27508 12637 27572
rect 12571 27507 12637 27508
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 15702 24853 15762 31043
rect 17907 30700 17973 30701
rect 17907 30636 17908 30700
rect 17972 30636 17973 30700
rect 17907 30635 17973 30636
rect 17910 29749 17970 30635
rect 18643 30020 18709 30021
rect 18643 29956 18644 30020
rect 18708 29956 18709 30020
rect 18643 29955 18709 29956
rect 17907 29748 17973 29749
rect 17907 29684 17908 29748
rect 17972 29684 17973 29748
rect 17907 29683 17973 29684
rect 18275 29340 18341 29341
rect 18275 29276 18276 29340
rect 18340 29276 18341 29340
rect 18275 29275 18341 29276
rect 18278 24853 18338 29275
rect 15699 24852 15765 24853
rect 15699 24788 15700 24852
rect 15764 24788 15765 24852
rect 15699 24787 15765 24788
rect 18275 24852 18341 24853
rect 18275 24788 18276 24852
rect 18340 24788 18341 24852
rect 18275 24787 18341 24788
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 18646 21997 18706 29955
rect 20854 29749 20914 41515
rect 20851 29748 20917 29749
rect 20851 29684 20852 29748
rect 20916 29684 20917 29748
rect 20851 29683 20917 29684
rect 21038 28797 21098 42875
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 26003 40628 26069 40629
rect 26003 40564 26004 40628
rect 26068 40564 26069 40628
rect 26003 40563 26069 40564
rect 21955 39404 22021 39405
rect 21955 39340 21956 39404
rect 22020 39340 22021 39404
rect 21955 39339 22021 39340
rect 21771 30564 21837 30565
rect 21771 30500 21772 30564
rect 21836 30500 21837 30564
rect 21771 30499 21837 30500
rect 21035 28796 21101 28797
rect 21035 28732 21036 28796
rect 21100 28732 21101 28796
rect 21035 28731 21101 28732
rect 21774 21997 21834 30499
rect 21958 29205 22018 39339
rect 21955 29204 22021 29205
rect 21955 29140 21956 29204
rect 22020 29140 22021 29204
rect 21955 29139 22021 29140
rect 26006 28661 26066 40563
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 26003 28660 26069 28661
rect 26003 28596 26004 28660
rect 26068 28596 26069 28660
rect 26003 28595 26069 28596
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 25635 22948 25701 22949
rect 25635 22884 25636 22948
rect 25700 22884 25701 22948
rect 25635 22883 25701 22884
rect 18643 21996 18709 21997
rect 18643 21932 18644 21996
rect 18708 21932 18709 21996
rect 18643 21931 18709 21932
rect 21771 21996 21837 21997
rect 21771 21932 21772 21996
rect 21836 21932 21837 21996
rect 21771 21931 21837 21932
rect 24899 21860 24965 21861
rect 24899 21796 24900 21860
rect 24964 21796 24965 21860
rect 24899 21795 24965 21796
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 24902 13701 24962 21795
rect 25638 13701 25698 22883
rect 32811 22540 32877 22541
rect 32811 22476 32812 22540
rect 32876 22476 32877 22540
rect 32811 22475 32877 22476
rect 32814 13837 32874 22475
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 32811 13836 32877 13837
rect 32811 13772 32812 13836
rect 32876 13772 32877 13836
rect 32811 13771 32877 13772
rect 24899 13700 24965 13701
rect 24899 13636 24900 13700
rect 24964 13636 24965 13700
rect 24899 13635 24965 13636
rect 25635 13700 25701 13701
rect 25635 13636 25636 13700
rect 25700 13636 25701 13700
rect 25635 13635 25701 13636
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 43552 35908 43568
rect 35588 43488 35596 43552
rect 35660 43488 35676 43552
rect 35740 43488 35756 43552
rect 35820 43488 35836 43552
rect 35900 43488 35908 43552
rect 35588 42464 35908 43488
rect 35588 42400 35596 42464
rect 35660 42400 35676 42464
rect 35740 42400 35756 42464
rect 35820 42400 35836 42464
rect 35900 42400 35908 42464
rect 35588 41376 35908 42400
rect 35588 41312 35596 41376
rect 35660 41312 35676 41376
rect 35740 41312 35756 41376
rect 35820 41312 35836 41376
rect 35900 41312 35908 41376
rect 35588 40288 35908 41312
rect 35588 40224 35596 40288
rect 35660 40224 35676 40288
rect 35740 40224 35756 40288
rect 35820 40224 35836 40288
rect 35900 40224 35908 40288
rect 35588 39200 35908 40224
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 38147 20772 38213 20773
rect 38147 20708 38148 20772
rect 38212 20708 38213 20772
rect 38147 20707 38213 20708
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 38150 15469 38210 20707
rect 38147 15468 38213 15469
rect 38147 15404 38148 15468
rect 38212 15404 38213 15468
rect 38147 15403 38213 15404
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 42552 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 42552 36920
rect 1056 36642 42552 36684
rect 1056 36260 42552 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 42552 36260
rect 1056 35982 42552 36024
rect 1056 6284 42552 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 42552 6284
rect 1056 6006 42552 6048
rect 1056 5624 42552 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 42552 5624
rect 1056 5346 42552 5388
use sky130_fd_sc_hd__a21o_1  _1211_
timestamp 18001
transform -1 0 15732 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1212_
timestamp 18001
transform -1 0 17572 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1213_
timestamp 18001
transform -1 0 17756 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1214_
timestamp 18001
transform 1 0 16100 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 18001
transform -1 0 16928 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1216_
timestamp 18001
transform 1 0 15640 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1217_
timestamp 18001
transform 1 0 19320 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1218_
timestamp 18001
transform -1 0 19320 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1219_
timestamp 18001
transform -1 0 19504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1220_
timestamp 18001
transform -1 0 18124 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1221_
timestamp 18001
transform 1 0 18768 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1222_
timestamp 18001
transform -1 0 18768 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1223_
timestamp 18001
transform 1 0 17756 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1224_
timestamp 18001
transform 1 0 20884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 18001
transform 1 0 21528 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 18001
transform 1 0 19504 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1227_
timestamp 18001
transform -1 0 20608 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1228_
timestamp 18001
transform -1 0 20700 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1229_
timestamp 18001
transform 1 0 20240 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1230_
timestamp 18001
transform 1 0 20700 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1231_
timestamp 18001
transform 1 0 21344 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1232_
timestamp 18001
transform 1 0 23184 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 18001
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 18001
transform -1 0 22264 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 18001
transform -1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1236_
timestamp 18001
transform -1 0 22264 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1237_
timestamp 18001
transform -1 0 23184 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1238_
timestamp 18001
transform -1 0 22356 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1239_
timestamp 18001
transform -1 0 22356 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1240_
timestamp 18001
transform 1 0 25024 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1241_
timestamp 18001
transform 1 0 24656 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1242_
timestamp 18001
transform 1 0 24380 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1243_
timestamp 18001
transform -1 0 25392 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1244_
timestamp 18001
transform 1 0 23552 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1245_
timestamp 18001
transform 1 0 25300 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1246_
timestamp 18001
transform 1 0 25760 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1247_
timestamp 18001
transform -1 0 26496 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1248_
timestamp 18001
transform 1 0 25116 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1249_
timestamp 18001
transform -1 0 25760 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1250_
timestamp 18001
transform -1 0 26496 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1251_
timestamp 18001
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1252_
timestamp 18001
transform -1 0 27876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1253_
timestamp 18001
transform 1 0 26864 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 18001
transform -1 0 30084 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1255_
timestamp 18001
transform -1 0 29440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1256_
timestamp 18001
transform 1 0 29440 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1257_
timestamp 18001
transform 1 0 28888 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1258_
timestamp 18001
transform 1 0 29532 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1259_
timestamp 18001
transform 1 0 30084 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 18001
transform 1 0 30820 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1261_
timestamp 18001
transform -1 0 30820 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1262_
timestamp 18001
transform -1 0 31648 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1263_
timestamp 18001
transform 1 0 30268 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1264_
timestamp 18001
transform 1 0 30544 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1265_
timestamp 18001
transform -1 0 30084 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1266_
timestamp 18001
transform -1 0 31004 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1267_
timestamp 18001
transform -1 0 33764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1268_
timestamp 18001
transform 1 0 31372 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1269_
timestamp 18001
transform -1 0 37996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1270_
timestamp 18001
transform 1 0 37904 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1271_
timestamp 18001
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1272_
timestamp 18001
transform -1 0 37904 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1273_
timestamp 18001
transform -1 0 37628 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1274_
timestamp 18001
transform 1 0 37904 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1275_
timestamp 18001
transform 1 0 37260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1276_
timestamp 18001
transform 1 0 36616 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1277_
timestamp 18001
transform -1 0 37904 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1278_
timestamp 18001
transform -1 0 36064 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1279_
timestamp 18001
transform 1 0 35328 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1280_
timestamp 18001
transform -1 0 35604 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1281_
timestamp 18001
transform 1 0 35420 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1282_
timestamp 18001
transform 1 0 36156 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1283_
timestamp 18001
transform -1 0 35236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1284_
timestamp 18001
transform 1 0 34776 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1285_
timestamp 18001
transform -1 0 36984 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1286_
timestamp 18001
transform 1 0 34868 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1287_
timestamp 18001
transform -1 0 35604 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1288_
timestamp 18001
transform 1 0 34500 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1289_
timestamp 18001
transform -1 0 34500 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1290_
timestamp 18001
transform 1 0 33396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1291_
timestamp 18001
transform 1 0 33856 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1292_
timestamp 18001
transform -1 0 23368 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1293_
timestamp 18001
transform -1 0 19044 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1294_
timestamp 18001
transform 1 0 19228 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 18001
transform 1 0 17388 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1296_
timestamp 18001
transform -1 0 18400 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1297_
timestamp 18001
transform 1 0 17848 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1298_
timestamp 18001
transform 1 0 17388 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1299_
timestamp 18001
transform 1 0 18584 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1300_
timestamp 18001
transform 1 0 18584 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1301_
timestamp 18001
transform -1 0 19872 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1302_
timestamp 18001
transform -1 0 18584 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1303_
timestamp 18001
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1304_
timestamp 18001
transform 1 0 16652 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1305_
timestamp 18001
transform 1 0 20056 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1306_
timestamp 18001
transform -1 0 19780 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1307_
timestamp 18001
transform 1 0 20516 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1308_
timestamp 18001
transform -1 0 20516 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1309_
timestamp 18001
transform 1 0 20240 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1310_
timestamp 18001
transform 1 0 20148 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1311_
timestamp 18001
transform -1 0 20884 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1312_
timestamp 18001
transform 1 0 22816 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 18001
transform -1 0 21896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1314_
timestamp 18001
transform 1 0 21160 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1315_
timestamp 18001
transform -1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1316_
timestamp 18001
transform -1 0 22540 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1317_
timestamp 18001
transform -1 0 21712 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1318_
timestamp 18001
transform 1 0 21528 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1319_
timestamp 18001
transform 1 0 21804 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1320_
timestamp 18001
transform -1 0 24748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1321_
timestamp 18001
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1322_
timestamp 18001
transform -1 0 24012 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1323_
timestamp 18001
transform 1 0 23644 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1324_
timestamp 18001
transform -1 0 24196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1325_
timestamp 18001
transform -1 0 25944 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1326_
timestamp 18001
transform 1 0 25116 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1327_
timestamp 18001
transform -1 0 25116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1328_
timestamp 18001
transform 1 0 24564 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1329_
timestamp 18001
transform -1 0 26036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1330_
timestamp 18001
transform -1 0 25392 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1331_
timestamp 18001
transform -1 0 25944 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1332_
timestamp 18001
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1333_
timestamp 18001
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 18001
transform -1 0 29348 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1335_
timestamp 18001
transform -1 0 29992 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1336_
timestamp 18001
transform -1 0 29808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1337_
timestamp 18001
transform 1 0 28520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1338_
timestamp 18001
transform 1 0 28060 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1339_
timestamp 18001
transform 1 0 29256 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1340_
timestamp 18001
transform 1 0 29716 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1341_
timestamp 18001
transform 1 0 29900 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1342_
timestamp 18001
transform 1 0 31280 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1343_
timestamp 18001
transform -1 0 33120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1344_
timestamp 18001
transform -1 0 32016 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1345_
timestamp 18001
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1346_
timestamp 18001
transform 1 0 31188 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 18001
transform 1 0 37260 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1348_
timestamp 18001
transform -1 0 36892 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1349_
timestamp 18001
transform 1 0 37076 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1350_
timestamp 18001
transform -1 0 38364 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1351_
timestamp 18001
transform -1 0 35604 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 18001
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 18001
transform -1 0 37168 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1354_
timestamp 18001
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1355_
timestamp 18001
transform -1 0 37720 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1356_
timestamp 18001
transform 1 0 34316 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1357_
timestamp 18001
transform -1 0 36800 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1358_
timestamp 18001
transform 1 0 35696 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1359_
timestamp 18001
transform 1 0 35604 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1360_
timestamp 18001
transform -1 0 36616 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1361_
timestamp 18001
transform 1 0 35512 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1362_
timestamp 18001
transform 1 0 35696 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1363_
timestamp 18001
transform 1 0 34776 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1364_
timestamp 18001
transform 1 0 33396 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1365_
timestamp 18001
transform -1 0 34224 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1366_
timestamp 18001
transform 1 0 33580 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1367_
timestamp 18001
transform 1 0 32936 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1368_
timestamp 18001
transform 1 0 8004 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 18001
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1370_
timestamp 18001
transform 1 0 19228 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1371_
timestamp 18001
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1372_
timestamp 18001
transform 1 0 21068 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1373_
timestamp 18001
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1374_
timestamp 18001
transform 1 0 23460 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1375_
timestamp 18001
transform 1 0 23920 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1376_
timestamp 18001
transform 1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1377_
timestamp 18001
transform 1 0 27876 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1378_
timestamp 18001
transform 1 0 28612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1379_
timestamp 18001
transform 1 0 31372 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1380_
timestamp 18001
transform 1 0 32108 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1381_
timestamp 18001
transform 1 0 33488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1382_
timestamp 18001
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1383_
timestamp 18001
transform 1 0 37260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1384_
timestamp 18001
transform 1 0 37536 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1385_
timestamp 18001
transform 1 0 13340 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1386_
timestamp 18001
transform -1 0 14720 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1387_
timestamp 18001
transform -1 0 13984 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1388_
timestamp 18001
transform 1 0 14076 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1389_
timestamp 18001
transform 1 0 14536 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1390_
timestamp 18001
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1391_
timestamp 18001
transform 1 0 16652 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1392_
timestamp 18001
transform 1 0 17204 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1393_
timestamp 18001
transform 1 0 20240 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1394_
timestamp 18001
transform 1 0 21896 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1395_
timestamp 18001
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1396_
timestamp 18001
transform 1 0 25576 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1397_
timestamp 18001
transform 1 0 26956 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1398_
timestamp 18001
transform 1 0 28428 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1399_
timestamp 18001
transform 1 0 32752 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1400_
timestamp 18001
transform 1 0 31188 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1401_
timestamp 18001
transform 1 0 37260 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1402_
timestamp 18001
transform 1 0 38640 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1403_
timestamp 18001
transform -1 0 38640 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1404_
timestamp 18001
transform 1 0 38272 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1405_
timestamp 18001
transform 1 0 33580 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1406_
timestamp 18001
transform 1 0 15640 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 18001
transform -1 0 19872 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1408_
timestamp 18001
transform -1 0 19320 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1409_
timestamp 18001
transform 1 0 20056 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 18001
transform -1 0 23920 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1411_
timestamp 18001
transform -1 0 25024 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1412_
timestamp 18001
transform 1 0 25760 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1413_
timestamp 18001
transform -1 0 30912 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 18001
transform -1 0 30176 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1415_
timestamp 18001
transform 1 0 30268 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1416_
timestamp 18001
transform 1 0 32108 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1417_
timestamp 18001
transform -1 0 38548 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1418_
timestamp 18001
transform -1 0 41676 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1419_
timestamp 18001
transform 1 0 40112 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1420_
timestamp 18001
transform 1 0 40756 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 18001
transform 1 0 34224 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1422_
timestamp 18001
transform -1 0 17664 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1423_
timestamp 18001
transform 1 0 16744 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1424_
timestamp 18001
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1425_
timestamp 18001
transform 1 0 17664 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1426_
timestamp 18001
transform 1 0 20424 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1427_
timestamp 18001
transform -1 0 23000 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1428_
timestamp 18001
transform 1 0 24380 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1429_
timestamp 18001
transform 1 0 26956 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1430_
timestamp 18001
transform 1 0 27692 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1431_
timestamp 18001
transform 1 0 29532 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1432_
timestamp 18001
transform 1 0 30820 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1433_
timestamp 18001
transform 1 0 32752 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1434_
timestamp 18001
transform 1 0 37168 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1435_
timestamp 18001
transform 1 0 40480 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1436_
timestamp 18001
transform -1 0 41584 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1437_
timestamp 18001
transform -1 0 38272 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1438_
timestamp 18001
transform 1 0 34684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1439_
timestamp 18001
transform 1 0 18952 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 18001
transform 1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1441_
timestamp 18001
transform 1 0 20608 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1442_
timestamp 18001
transform 1 0 21804 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1443_
timestamp 18001
transform 1 0 23644 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 18001
transform 1 0 24564 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1445_
timestamp 18001
transform 1 0 26220 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1446_
timestamp 18001
transform 1 0 27692 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1447_
timestamp 18001
transform 1 0 31372 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1448_
timestamp 18001
transform 1 0 32108 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1449_
timestamp 18001
transform 1 0 33028 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1450_
timestamp 18001
transform 1 0 33856 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1451_
timestamp 18001
transform 1 0 34960 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 18001
transform 1 0 35696 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1453_
timestamp 18001
transform 1 0 36524 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1454_
timestamp 18001
transform -1 0 19044 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1455_
timestamp 18001
transform -1 0 19688 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1456_
timestamp 18001
transform 1 0 18216 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1457_
timestamp 18001
transform 1 0 19228 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1458_
timestamp 18001
transform -1 0 19964 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1459_
timestamp 18001
transform -1 0 20424 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1460_
timestamp 18001
transform -1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1461_
timestamp 18001
transform 1 0 18676 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1462_
timestamp 18001
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1463_
timestamp 18001
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1464_
timestamp 18001
transform -1 0 21436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _1465_
timestamp 18001
transform -1 0 19964 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1466_
timestamp 18001
transform 1 0 20424 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1467_
timestamp 18001
transform -1 0 21160 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 18001
transform 1 0 20240 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1469_
timestamp 18001
transform 1 0 23920 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1470_
timestamp 18001
transform 1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1471_
timestamp 18001
transform -1 0 22908 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1472_
timestamp 18001
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1473_
timestamp 18001
transform 1 0 21804 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1474_
timestamp 18001
transform -1 0 22448 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1475_
timestamp 18001
transform -1 0 24380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1476_
timestamp 18001
transform -1 0 25300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1477_
timestamp 18001
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1478_
timestamp 18001
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1479_
timestamp 18001
transform 1 0 23460 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1480_
timestamp 18001
transform 1 0 24380 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1481_
timestamp 18001
transform -1 0 25024 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 18001
transform 1 0 26956 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1483_
timestamp 18001
transform 1 0 27416 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1484_
timestamp 18001
transform -1 0 27508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1485_
timestamp 18001
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1486_
timestamp 18001
transform -1 0 25208 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1487_
timestamp 18001
transform 1 0 25208 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1488_
timestamp 18001
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1489_
timestamp 18001
transform 1 0 24840 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1490_
timestamp 18001
transform -1 0 28520 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1491_
timestamp 18001
transform -1 0 27968 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1492_
timestamp 18001
transform -1 0 30084 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1493_
timestamp 18001
transform 1 0 23920 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1494_
timestamp 18001
transform 1 0 28704 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1495_
timestamp 18001
transform 1 0 28060 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1496_
timestamp 18001
transform -1 0 29348 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1497_
timestamp 18001
transform 1 0 30452 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1498_
timestamp 18001
transform 1 0 30176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1499_
timestamp 18001
transform -1 0 29440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1500_
timestamp 18001
transform -1 0 29532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1501_
timestamp 18001
transform 1 0 28244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1502_
timestamp 18001
transform 1 0 28704 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1503_
timestamp 18001
transform 1 0 28152 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1504_
timestamp 18001
transform 1 0 33212 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1505_
timestamp 18001
transform 1 0 31740 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1506_
timestamp 18001
transform -1 0 31924 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1507_
timestamp 18001
transform -1 0 28704 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 18001
transform 1 0 30452 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1509_
timestamp 18001
transform 1 0 30728 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1510_
timestamp 18001
transform -1 0 31740 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 18001
transform -1 0 33212 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1512_
timestamp 18001
transform -1 0 33488 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1513_
timestamp 18001
transform 1 0 31648 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1514_
timestamp 18001
transform 1 0 32476 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1515_
timestamp 18001
transform 1 0 32108 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1516_
timestamp 18001
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1517_
timestamp 18001
transform -1 0 37536 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1518_
timestamp 18001
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1519_
timestamp 18001
transform -1 0 38456 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1520_
timestamp 18001
transform 1 0 30912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _1521_
timestamp 18001
transform 1 0 33212 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1522_
timestamp 18001
transform 1 0 36064 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1523_
timestamp 18001
transform -1 0 37904 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp 18001
transform 1 0 41676 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1525_
timestamp 18001
transform 1 0 41952 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1526_
timestamp 18001
transform -1 0 41492 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1527_
timestamp 18001
transform -1 0 37444 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1528_
timestamp 18001
transform 1 0 39652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1529_
timestamp 18001
transform -1 0 40480 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1530_
timestamp 18001
transform -1 0 41400 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 18001
transform 1 0 41952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1532_
timestamp 18001
transform 1 0 40020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1533_
timestamp 18001
transform -1 0 40388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1534_
timestamp 18001
transform 1 0 40388 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1535_
timestamp 18001
transform -1 0 39744 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1536_
timestamp 18001
transform 1 0 41768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1537_
timestamp 18001
transform -1 0 40664 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1538_
timestamp 18001
transform 1 0 39836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1539_
timestamp 18001
transform 1 0 41492 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1540_
timestamp 18001
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1541_
timestamp 18001
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1542_
timestamp 18001
transform 1 0 35144 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1543_
timestamp 18001
transform 1 0 40296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1544_
timestamp 18001
transform 1 0 35788 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 18001
transform -1 0 37904 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1546_
timestamp 18001
transform 1 0 14076 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1547_
timestamp 18001
transform -1 0 17112 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1548_
timestamp 18001
transform -1 0 17388 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1549_
timestamp 18001
transform 1 0 16376 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1550_
timestamp 18001
transform 1 0 14904 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1551_
timestamp 18001
transform 1 0 14904 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1552_
timestamp 18001
transform 1 0 15824 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 18001
transform 1 0 15548 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 18001
transform -1 0 35880 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1555_
timestamp 18001
transform 1 0 35880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1556_
timestamp 18001
transform -1 0 34592 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1557_
timestamp 18001
transform -1 0 36432 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1558_
timestamp 18001
transform -1 0 36984 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1559_
timestamp 18001
transform 1 0 36432 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1560_
timestamp 18001
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1561_
timestamp 18001
transform -1 0 38824 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1562_
timestamp 18001
transform 1 0 39192 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1563_
timestamp 18001
transform 1 0 38824 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1564_
timestamp 18001
transform -1 0 38364 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1565_
timestamp 18001
transform 1 0 39928 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1566_
timestamp 18001
transform 1 0 39836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1567_
timestamp 18001
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1568_
timestamp 18001
transform 1 0 40388 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1569_
timestamp 18001
transform -1 0 40388 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 18001
transform -1 0 40388 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1571_
timestamp 18001
transform 1 0 39744 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1572_
timestamp 18001
transform -1 0 39744 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1573_
timestamp 18001
transform -1 0 33212 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1574_
timestamp 18001
transform 1 0 33120 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1575_
timestamp 18001
transform -1 0 32752 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1576_
timestamp 18001
transform 1 0 31372 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1577_
timestamp 18001
transform 1 0 30268 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1578_
timestamp 18001
transform 1 0 30360 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1579_
timestamp 18001
transform -1 0 31096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1580_
timestamp 18001
transform -1 0 33120 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1581_
timestamp 18001
transform -1 0 29072 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1582_
timestamp 18001
transform -1 0 29348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1583_
timestamp 18001
transform -1 0 29256 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1584_
timestamp 18001
transform -1 0 28888 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1585_
timestamp 18001
transform 1 0 27048 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1586_
timestamp 18001
transform 1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1587_
timestamp 18001
transform 1 0 27508 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1588_
timestamp 18001
transform 1 0 27876 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1589_
timestamp 18001
transform -1 0 25668 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1590_
timestamp 18001
transform 1 0 26036 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1591_
timestamp 18001
transform -1 0 26036 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1592_
timestamp 18001
transform -1 0 25484 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1593_
timestamp 18001
transform -1 0 24012 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1594_
timestamp 18001
transform -1 0 24288 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1595_
timestamp 18001
transform 1 0 23552 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1596_
timestamp 18001
transform 1 0 23920 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1597_
timestamp 18001
transform -1 0 21988 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1598_
timestamp 18001
transform -1 0 22632 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1599_
timestamp 18001
transform 1 0 21988 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1600_
timestamp 18001
transform -1 0 21528 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1601_
timestamp 18001
transform 1 0 19136 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1602_
timestamp 18001
transform -1 0 19136 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1603_
timestamp 18001
transform -1 0 19596 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1604_
timestamp 18001
transform 1 0 19596 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1605_
timestamp 18001
transform 1 0 16652 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1606_
timestamp 18001
transform -1 0 17756 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 18001
transform -1 0 15456 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1608_
timestamp 18001
transform -1 0 18308 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1609_
timestamp 18001
transform -1 0 18676 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1610_
timestamp 18001
transform -1 0 19688 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1611_
timestamp 18001
transform 1 0 19228 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1612_
timestamp 18001
transform -1 0 23184 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1613_
timestamp 18001
transform -1 0 24288 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1614_
timestamp 18001
transform -1 0 25116 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1615_
timestamp 18001
transform -1 0 26588 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1616_
timestamp 18001
transform -1 0 27692 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1617_
timestamp 18001
transform 1 0 27140 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1618_
timestamp 18001
transform -1 0 30912 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1619_
timestamp 18001
transform -1 0 32200 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1620_
timestamp 18001
transform 1 0 30820 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1621_
timestamp 18001
transform -1 0 37168 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1622_
timestamp 18001
transform 1 0 38640 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1623_
timestamp 18001
transform 1 0 38272 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1624_
timestamp 18001
transform 1 0 38548 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1625_
timestamp 18001
transform 1 0 37352 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1626_
timestamp 18001
transform 1 0 37168 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1627_
timestamp 18001
transform 1 0 35328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1628_
timestamp 18001
transform 1 0 33764 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1629_
timestamp 18001
transform -1 0 34224 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1630_
timestamp 18001
transform -1 0 35328 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1631_
timestamp 18001
transform -1 0 17940 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1632_
timestamp 18001
transform 1 0 16928 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1633_
timestamp 18001
transform -1 0 19412 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1634_
timestamp 18001
transform 1 0 17388 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1635_
timestamp 18001
transform -1 0 17296 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1636_
timestamp 18001
transform 1 0 17296 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1637_
timestamp 18001
transform 1 0 19412 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1638_
timestamp 18001
transform 1 0 19872 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1639_
timestamp 18001
transform -1 0 19136 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1640_
timestamp 18001
transform 1 0 18860 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1641_
timestamp 18001
transform 1 0 19780 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1642_
timestamp 18001
transform 1 0 20424 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1643_
timestamp 18001
transform 1 0 20056 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1644_
timestamp 18001
transform -1 0 21252 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1645_
timestamp 18001
transform 1 0 19964 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1646_
timestamp 18001
transform -1 0 21160 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1647_
timestamp 18001
transform 1 0 21712 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1648_
timestamp 18001
transform 1 0 20976 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1649_
timestamp 18001
transform 1 0 20516 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1650_
timestamp 18001
transform 1 0 22632 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1651_
timestamp 18001
transform -1 0 23644 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1652_
timestamp 18001
transform 1 0 22908 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1653_
timestamp 18001
transform 1 0 22908 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1654_
timestamp 18001
transform 1 0 23276 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1655_
timestamp 18001
transform 1 0 23552 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1656_
timestamp 18001
transform -1 0 25668 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1657_
timestamp 18001
transform 1 0 24840 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1658_
timestamp 18001
transform 1 0 26036 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1659_
timestamp 18001
transform 1 0 25668 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1660_
timestamp 18001
transform 1 0 25300 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1661_
timestamp 18001
transform 1 0 26956 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1662_
timestamp 18001
transform -1 0 27048 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1663_
timestamp 18001
transform 1 0 26956 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1664_
timestamp 18001
transform 1 0 28428 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1665_
timestamp 18001
transform -1 0 27416 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1666_
timestamp 18001
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1667_
timestamp 18001
transform -1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1668_
timestamp 18001
transform 1 0 27692 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1669_
timestamp 18001
transform 1 0 28796 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1670_
timestamp 18001
transform 1 0 27968 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1671_
timestamp 18001
transform -1 0 28888 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1672_
timestamp 18001
transform 1 0 27416 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1673_
timestamp 18001
transform -1 0 30820 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1674_
timestamp 18001
transform 1 0 30544 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1675_
timestamp 18001
transform -1 0 30820 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1676_
timestamp 18001
transform 1 0 31556 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1677_
timestamp 18001
transform 1 0 30820 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1678_
timestamp 18001
transform 1 0 31556 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1679_
timestamp 18001
transform -1 0 32752 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1680_
timestamp 18001
transform 1 0 32108 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1681_
timestamp 18001
transform -1 0 32476 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1682_
timestamp 18001
transform 1 0 32476 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1683_
timestamp 18001
transform 1 0 32476 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1684_
timestamp 18001
transform 1 0 33120 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1685_
timestamp 18001
transform -1 0 39744 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1686_
timestamp 18001
transform -1 0 38088 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1687_
timestamp 18001
transform -1 0 35328 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1688_
timestamp 18001
transform 1 0 35328 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1689_
timestamp 18001
transform 1 0 35328 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1690_
timestamp 18001
transform -1 0 36984 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1691_
timestamp 18001
transform -1 0 39192 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1692_
timestamp 18001
transform -1 0 38640 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1693_
timestamp 18001
transform 1 0 35972 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1694_
timestamp 18001
transform -1 0 37168 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1695_
timestamp 18001
transform -1 0 36156 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1696_
timestamp 18001
transform -1 0 38456 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1697_
timestamp 18001
transform -1 0 38548 0 1 38080
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1698_
timestamp 18001
transform 1 0 34960 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1699_
timestamp 18001
transform 1 0 35604 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1700_
timestamp 18001
transform 1 0 34684 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1701_
timestamp 18001
transform -1 0 36248 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1702_
timestamp 18001
transform 1 0 35972 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1703_
timestamp 18001
transform -1 0 36616 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1704_
timestamp 18001
transform 1 0 35604 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1705_
timestamp 18001
transform 1 0 37260 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1706_
timestamp 18001
transform -1 0 35880 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1707_
timestamp 18001
transform 1 0 34224 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1708_
timestamp 18001
transform 1 0 34224 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1709_
timestamp 18001
transform -1 0 36064 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1710_
timestamp 18001
transform 1 0 33396 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1711_
timestamp 18001
transform 1 0 18584 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1712_
timestamp 18001
transform 1 0 17388 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1713_
timestamp 18001
transform -1 0 14352 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1714_
timestamp 18001
transform 1 0 14628 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1715_
timestamp 18001
transform 1 0 13156 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1716_
timestamp 18001
transform 1 0 16560 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 18001
transform 1 0 15732 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1718_
timestamp 18001
transform 1 0 19320 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1719_
timestamp 18001
transform 1 0 19228 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1720_
timestamp 18001
transform 1 0 22448 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1721_
timestamp 18001
transform 1 0 21804 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1722_
timestamp 18001
transform 1 0 23460 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 18001
transform 1 0 22908 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1724_
timestamp 18001
transform 1 0 25208 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1725_
timestamp 18001
transform 1 0 24748 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1726_
timestamp 18001
transform 1 0 26956 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 18001
transform 1 0 26956 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1728_
timestamp 18001
transform 1 0 29532 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1729_
timestamp 18001
transform 1 0 28152 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1730_
timestamp 18001
transform 1 0 30820 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1731_
timestamp 18001
transform -1 0 30176 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 18001
transform 1 0 31464 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 18001
transform 1 0 31372 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1734_
timestamp 18001
transform 1 0 41032 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1735_
timestamp 18001
transform 1 0 40664 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 18001
transform 1 0 41216 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1737_
timestamp 18001
transform -1 0 40848 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1738_
timestamp 18001
transform 1 0 38180 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1739_
timestamp 18001
transform 1 0 37904 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 18001
transform 1 0 35788 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1741_
timestamp 18001
transform 1 0 34960 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 18001
transform 1 0 33396 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1743_
timestamp 18001
transform 1 0 32936 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1744_
timestamp 18001
transform 1 0 14628 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1745_
timestamp 18001
transform 1 0 14076 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1746_
timestamp 18001
transform -1 0 17480 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1747_
timestamp 18001
transform 1 0 16652 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 18001
transform 1 0 19780 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1749_
timestamp 18001
transform 1 0 19228 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 18001
transform -1 0 22448 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1751_
timestamp 18001
transform 1 0 21804 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 18001
transform 1 0 23460 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1753_
timestamp 18001
transform 1 0 22448 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 18001
transform 1 0 26036 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1755_
timestamp 18001
transform 1 0 24840 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 18001
transform 1 0 27784 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1757_
timestamp 18001
transform 1 0 26956 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1758_
timestamp 18001
transform 1 0 28612 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 18001
transform 1 0 28244 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1760_
timestamp 18001
transform 1 0 29992 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 18001
transform 1 0 29532 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1762_
timestamp 18001
transform 1 0 31372 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 18001
transform 1 0 31188 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1764_
timestamp 18001
transform 1 0 40940 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 18001
transform 1 0 40480 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1766_
timestamp 18001
transform 1 0 40388 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 18001
transform 1 0 40204 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1768_
timestamp 18001
transform 1 0 39100 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 18001
transform 1 0 37904 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1770_
timestamp 18001
transform 1 0 36616 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1771_
timestamp 18001
transform 1 0 35512 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1772_
timestamp 18001
transform -1 0 34224 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1773_
timestamp 18001
transform 1 0 33764 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1774_
timestamp 18001
transform -1 0 12696 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1775_
timestamp 18001
transform 1 0 11684 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1776_
timestamp 18001
transform 1 0 12696 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1777_
timestamp 18001
transform -1 0 12052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1778_
timestamp 18001
transform -1 0 13432 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1779_
timestamp 18001
transform -1 0 11224 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1780_
timestamp 18001
transform 1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1781_
timestamp 18001
transform 1 0 13432 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1782_
timestamp 18001
transform -1 0 14904 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1783_
timestamp 18001
transform -1 0 14628 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1784_
timestamp 18001
transform 1 0 16192 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 18001
transform 1 0 16652 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1786_
timestamp 18001
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 18001
transform -1 0 18676 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1788_
timestamp 18001
transform 1 0 18216 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 18001
transform -1 0 21528 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1790_
timestamp 18001
transform 1 0 21252 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1791_
timestamp 18001
transform -1 0 23368 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1792_
timestamp 18001
transform 1 0 22356 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 18001
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1794_
timestamp 18001
transform 1 0 23828 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 18001
transform 1 0 23460 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1796_
timestamp 18001
transform -1 0 26588 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1797_
timestamp 18001
transform 1 0 25576 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1798_
timestamp 18001
transform 1 0 27508 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1799_
timestamp 18001
transform 1 0 27324 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 18001
transform 1 0 29716 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 18001
transform -1 0 30084 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 18001
transform 1 0 31280 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1803_
timestamp 18001
transform 1 0 30912 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 18001
transform -1 0 33212 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1805_
timestamp 18001
transform 1 0 32568 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 18001
transform 1 0 38180 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1807_
timestamp 18001
transform 1 0 37720 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 18001
transform 1 0 39836 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1809_
timestamp 18001
transform 1 0 39468 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1810_
timestamp 18001
transform -1 0 38640 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 18001
transform 1 0 39836 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1812_
timestamp 18001
transform -1 0 36616 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 18001
transform 1 0 37996 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1814_
timestamp 18001
transform 1 0 33764 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 18001
transform -1 0 34592 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1816_
timestamp 18001
transform -1 0 15916 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 18001
transform 1 0 15180 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _1818_
timestamp 18001
transform 1 0 11500 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 18001
transform 1 0 12512 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1820_
timestamp 18001
transform 1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1821_
timestamp 18001
transform 1 0 9108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1822_
timestamp 18001
transform 1 0 8004 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1823_
timestamp 18001
transform 1 0 8004 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1824_
timestamp 18001
transform -1 0 9936 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1825_
timestamp 18001
transform 1 0 8924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1826_
timestamp 18001
transform 1 0 9568 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1827_
timestamp 18001
transform 1 0 14904 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1828_
timestamp 18001
transform -1 0 16560 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1829_
timestamp 18001
transform 1 0 20148 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1830_
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1831_
timestamp 18001
transform 1 0 23368 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1832_
timestamp 18001
transform 1 0 25024 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1833_
timestamp 18001
transform -1 0 27324 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1834_
timestamp 18001
transform 1 0 28520 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1835_
timestamp 18001
transform 1 0 29900 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1836_
timestamp 18001
transform 1 0 32108 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1837_
timestamp 18001
transform 1 0 40756 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1838_
timestamp 18001
transform 1 0 39928 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1839_
timestamp 18001
transform 1 0 38272 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1840_
timestamp 18001
transform 1 0 35420 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1841_
timestamp 18001
transform 1 0 33120 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1842_
timestamp 18001
transform 1 0 12788 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1843_
timestamp 18001
transform 1 0 15640 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 18001
transform 1 0 17112 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1845_
timestamp 18001
transform 1 0 19964 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 18001
transform 1 0 21712 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1847_
timestamp 18001
transform 1 0 23368 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1848_
timestamp 18001
transform 1 0 25208 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1849_
timestamp 18001
transform 1 0 26956 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1850_
timestamp 18001
transform 1 0 29716 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1851_
timestamp 18001
transform 1 0 30544 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1852_
timestamp 18001
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1853_
timestamp 18001
transform 1 0 40388 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1854_
timestamp 18001
transform -1 0 39744 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1855_
timestamp 18001
transform 1 0 37812 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1856_
timestamp 18001
transform 1 0 35420 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1857_
timestamp 18001
transform 1 0 33304 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1858_
timestamp 18001
transform 1 0 14076 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1859_
timestamp 18001
transform 1 0 10396 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1860_
timestamp 18001
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1861_
timestamp 18001
transform -1 0 10856 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1862_
timestamp 18001
transform 1 0 10120 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1863_
timestamp 18001
transform 1 0 12328 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1864_
timestamp 18001
transform 1 0 11868 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1865_
timestamp 18001
transform 1 0 11776 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1866_
timestamp 18001
transform 1 0 11592 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1867_
timestamp 18001
transform 1 0 13156 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1868_
timestamp 18001
transform -1 0 14076 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1869_
timestamp 18001
transform -1 0 10672 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1870_
timestamp 18001
transform 1 0 11316 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1871_
timestamp 18001
transform -1 0 11868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1872_
timestamp 18001
transform -1 0 16468 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1873_
timestamp 18001
transform 1 0 15364 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1874_
timestamp 18001
transform -1 0 18308 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1875_
timestamp 18001
transform 1 0 14996 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1876_
timestamp 18001
transform -1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1877_
timestamp 18001
transform 1 0 19412 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1878_
timestamp 18001
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1879_
timestamp 18001
transform -1 0 24380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1880_
timestamp 18001
transform 1 0 17756 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1881_
timestamp 18001
transform -1 0 17480 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1882_
timestamp 18001
transform -1 0 16560 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1883_
timestamp 18001
transform 1 0 16100 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1884_
timestamp 18001
transform -1 0 19872 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1885_
timestamp 18001
transform 1 0 17480 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1886_
timestamp 18001
transform 1 0 18308 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1887_
timestamp 18001
transform -1 0 22448 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1888_
timestamp 18001
transform 1 0 20700 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1889_
timestamp 18001
transform 1 0 21344 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1890_
timestamp 18001
transform 1 0 21896 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1891_
timestamp 18001
transform 1 0 22724 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1892_
timestamp 18001
transform 1 0 24380 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1893_
timestamp 18001
transform -1 0 25024 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1894_
timestamp 18001
transform -1 0 24196 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1895_
timestamp 18001
transform 1 0 23828 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1896_
timestamp 18001
transform -1 0 28060 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1897_
timestamp 18001
transform -1 0 27600 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1898_
timestamp 18001
transform 1 0 26680 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1899_
timestamp 18001
transform -1 0 29072 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1900_
timestamp 18001
transform 1 0 27416 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1901_
timestamp 18001
transform 1 0 28152 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1902_
timestamp 18001
transform 1 0 40112 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1903_
timestamp 18001
transform 1 0 29532 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1904_
timestamp 18001
transform 1 0 40756 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1905_
timestamp 18001
transform 1 0 39744 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 18001
transform 1 0 32108 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1907_
timestamp 18001
transform 1 0 40296 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1908_
timestamp 18001
transform -1 0 40848 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1909_
timestamp 18001
transform 1 0 33212 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1910_
timestamp 18001
transform 1 0 40848 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1911_
timestamp 18001
transform -1 0 39284 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1912_
timestamp 18001
transform 1 0 37904 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1913_
timestamp 18001
transform 1 0 39008 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1914_
timestamp 18001
transform -1 0 40388 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1915_
timestamp 18001
transform 1 0 39008 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1916_
timestamp 18001
transform 1 0 40664 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1917_
timestamp 18001
transform -1 0 35420 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1918_
timestamp 18001
transform 1 0 35788 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1919_
timestamp 18001
transform 1 0 40940 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1920_
timestamp 18001
transform 1 0 39008 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1921_
timestamp 18001
transform 1 0 38180 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1922_
timestamp 18001
transform 1 0 39836 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1923_
timestamp 18001
transform 1 0 32752 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1924_
timestamp 18001
transform 1 0 34684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1925_
timestamp 18001
transform 1 0 40848 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1926_
timestamp 18001
transform -1 0 18860 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1927_
timestamp 18001
transform -1 0 19320 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1928_
timestamp 18001
transform 1 0 17664 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1929_
timestamp 18001
transform 1 0 17756 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1930_
timestamp 18001
transform -1 0 20424 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1931_
timestamp 18001
transform -1 0 19136 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1932_
timestamp 18001
transform -1 0 25024 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1933_
timestamp 18001
transform 1 0 24932 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1934_
timestamp 18001
transform -1 0 26404 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1935_
timestamp 18001
transform -1 0 28980 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1936_
timestamp 18001
transform 1 0 31004 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1937_
timestamp 18001
transform 1 0 32108 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1938_
timestamp 18001
transform -1 0 35328 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1939_
timestamp 18001
transform 1 0 33856 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1940_
timestamp 18001
transform -1 0 35880 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1941_
timestamp 18001
transform 1 0 34684 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1942_
timestamp 18001
transform 1 0 33948 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1943_
timestamp 18001
transform 1 0 13340 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1944_
timestamp 18001
transform 1 0 15364 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1945_
timestamp 18001
transform -1 0 10764 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 18001
transform -1 0 6624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1947_
timestamp 18001
transform -1 0 5612 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1948_
timestamp 18001
transform 1 0 4140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1949_
timestamp 18001
transform 1 0 26404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1950_
timestamp 18001
transform -1 0 16284 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1951_
timestamp 18001
transform 1 0 18584 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1952_
timestamp 18001
transform -1 0 15180 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1953_
timestamp 18001
transform -1 0 20700 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1954_
timestamp 18001
transform 1 0 34684 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1955_
timestamp 18001
transform -1 0 7820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1956_
timestamp 18001
transform 1 0 6992 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1957_
timestamp 18001
transform -1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1958_
timestamp 18001
transform -1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1959_
timestamp 18001
transform 1 0 18400 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1960_
timestamp 18001
transform 1 0 25944 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1961_
timestamp 18001
transform 1 0 2852 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1962_
timestamp 18001
transform -1 0 4416 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1963_
timestamp 18001
transform -1 0 7360 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1964_
timestamp 18001
transform 1 0 5520 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1965_
timestamp 18001
transform 1 0 4324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1966_
timestamp 18001
transform 1 0 2484 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _1967_
timestamp 18001
transform 1 0 2484 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1968_
timestamp 18001
transform -1 0 4140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _1969_
timestamp 18001
transform -1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1970_
timestamp 18001
transform 1 0 5244 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1971_
timestamp 18001
transform -1 0 3496 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1972_
timestamp 18001
transform 1 0 3864 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _1973_
timestamp 18001
transform -1 0 3036 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1974_
timestamp 18001
transform 1 0 5612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1975_
timestamp 18001
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1976_
timestamp 18001
transform 1 0 2392 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1977_
timestamp 18001
transform -1 0 5428 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1978_
timestamp 18001
transform 1 0 2024 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1979_
timestamp 18001
transform 1 0 3312 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1980_
timestamp 18001
transform 1 0 3220 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1981_
timestamp 18001
transform 1 0 3772 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 18001
transform 1 0 2944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1983_
timestamp 18001
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1984_
timestamp 18001
transform 1 0 1840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1985_
timestamp 18001
transform -1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1986_
timestamp 18001
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1987_
timestamp 18001
transform 1 0 25576 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1988_
timestamp 18001
transform 1 0 20516 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1989_
timestamp 18001
transform 1 0 34684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1990_
timestamp 18001
transform -1 0 35236 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1991_
timestamp 18001
transform -1 0 26404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1992_
timestamp 18001
transform -1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1993_
timestamp 18001
transform 1 0 20516 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1994_
timestamp 18001
transform 1 0 22724 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1995_
timestamp 18001
transform -1 0 24656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1996_
timestamp 18001
transform 1 0 26956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1997_
timestamp 18001
transform 1 0 30452 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1998_
timestamp 18001
transform 1 0 33304 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1999_
timestamp 18001
transform 1 0 34224 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2000_
timestamp 18001
transform 1 0 36064 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2001_
timestamp 18001
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2002_
timestamp 18001
transform -1 0 38456 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2003_
timestamp 18001
transform 1 0 35328 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2004_
timestamp 18001
transform -1 0 35788 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2005_
timestamp 18001
transform -1 0 26772 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _2006_
timestamp 18001
transform -1 0 26956 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2007_
timestamp 18001
transform 1 0 23644 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2008_
timestamp 18001
transform 1 0 25576 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2009_
timestamp 18001
transform 1 0 22540 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2010_
timestamp 18001
transform -1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2011_
timestamp 18001
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2012_
timestamp 18001
transform -1 0 23000 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2013_
timestamp 18001
transform 1 0 21712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2014_
timestamp 18001
transform -1 0 19044 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2015_
timestamp 18001
transform 1 0 19964 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2016_
timestamp 18001
transform -1 0 20332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2017_
timestamp 18001
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2018_
timestamp 18001
transform -1 0 24104 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _2019_
timestamp 18001
transform 1 0 23092 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _2020_
timestamp 18001
transform 1 0 24840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2021_
timestamp 18001
transform 1 0 26220 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2022_
timestamp 18001
transform -1 0 28704 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2023_
timestamp 18001
transform -1 0 28336 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2024_
timestamp 18001
transform -1 0 31280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2025_
timestamp 18001
transform 1 0 31464 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2026_
timestamp 18001
transform -1 0 29164 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2027_
timestamp 18001
transform -1 0 28428 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2028_
timestamp 18001
transform 1 0 31556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2029_
timestamp 18001
transform 1 0 32108 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2030_
timestamp 18001
transform -1 0 31924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2031_
timestamp 18001
transform -1 0 34224 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2032_
timestamp 18001
transform -1 0 32752 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2033_
timestamp 18001
transform -1 0 32476 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2034_
timestamp 18001
transform -1 0 34408 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2035_
timestamp 18001
transform 1 0 34684 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _2036_
timestamp 18001
transform -1 0 34500 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2037_
timestamp 18001
transform 1 0 36616 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2038_
timestamp 18001
transform 1 0 35788 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2039_
timestamp 18001
transform -1 0 34500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2040_
timestamp 18001
transform 1 0 37168 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _2041_
timestamp 18001
transform 1 0 37260 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _2042_
timestamp 18001
transform 1 0 36248 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _2043_
timestamp 18001
transform 1 0 26128 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2044_
timestamp 18001
transform 1 0 28612 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2045_
timestamp 18001
transform 1 0 10120 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2046_
timestamp 18001
transform -1 0 6256 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2047_
timestamp 18001
transform 1 0 4416 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _2048_
timestamp 18001
transform 1 0 4784 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2049_
timestamp 18001
transform 1 0 4876 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2050_
timestamp 18001
transform 1 0 2668 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2051_
timestamp 18001
transform 1 0 4692 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2052_
timestamp 18001
transform 1 0 3772 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2053_
timestamp 18001
transform -1 0 5704 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2054_
timestamp 18001
transform 1 0 4048 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2055_
timestamp 18001
transform -1 0 8096 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2056_
timestamp 18001
transform 1 0 6532 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2057_
timestamp 18001
transform 1 0 6900 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2058_
timestamp 18001
transform -1 0 8832 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2059_
timestamp 18001
transform 1 0 7728 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2060_
timestamp 18001
transform 1 0 6992 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2061_
timestamp 18001
transform 1 0 7820 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2062_
timestamp 18001
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2063_
timestamp 18001
transform 1 0 6348 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2064_
timestamp 18001
transform 1 0 5888 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2065_
timestamp 18001
transform -1 0 5520 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2066_
timestamp 18001
transform -1 0 5244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2067_
timestamp 18001
transform 1 0 4232 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2068_
timestamp 18001
transform 1 0 4508 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2069_
timestamp 18001
transform -1 0 3680 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2070_
timestamp 18001
transform -1 0 1840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2071_
timestamp 18001
transform 1 0 2300 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2072_
timestamp 18001
transform 1 0 1840 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2073_
timestamp 18001
transform 1 0 4968 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2074_
timestamp 18001
transform -1 0 3680 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2075_
timestamp 18001
transform 1 0 2484 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2076_
timestamp 18001
transform 1 0 5704 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2077_
timestamp 18001
transform -1 0 3680 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2078_
timestamp 18001
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2079_
timestamp 18001
transform -1 0 4324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2080_
timestamp 18001
transform 1 0 4324 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2081_
timestamp 18001
transform -1 0 4508 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _2082_
timestamp 18001
transform 1 0 4968 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2083_
timestamp 18001
transform 1 0 3956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _2084_
timestamp 18001
transform 1 0 5980 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2085_
timestamp 18001
transform -1 0 6808 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2086_
timestamp 18001
transform 1 0 4784 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2087_
timestamp 18001
transform 1 0 5244 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _2088_
timestamp 18001
transform 1 0 8096 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2089_
timestamp 18001
transform -1 0 7820 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2090_
timestamp 18001
transform 1 0 7452 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _2091_
timestamp 18001
transform 1 0 7636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2092_
timestamp 18001
transform -1 0 8832 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2093_
timestamp 18001
transform 1 0 9660 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2094_
timestamp 18001
transform -1 0 7176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2095_
timestamp 18001
transform 1 0 7360 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2096_
timestamp 18001
transform 1 0 7360 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2097_
timestamp 18001
transform -1 0 9200 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2098_
timestamp 18001
transform 1 0 6348 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2099_
timestamp 18001
transform -1 0 8740 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2100_
timestamp 18001
transform 1 0 7544 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2101_
timestamp 18001
transform 1 0 4324 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2102_
timestamp 18001
transform 1 0 5612 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2103_
timestamp 18001
transform 1 0 4968 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2104_
timestamp 18001
transform 1 0 4692 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2105_
timestamp 18001
transform -1 0 5612 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2106_
timestamp 18001
transform 1 0 5612 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2107_
timestamp 18001
transform 1 0 5612 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _2108_
timestamp 18001
transform -1 0 5612 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _2109_
timestamp 18001
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2110_
timestamp 18001
transform -1 0 4508 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2111_
timestamp 18001
transform -1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2112_
timestamp 18001
transform 1 0 5336 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2113_
timestamp 18001
transform -1 0 4232 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2114_
timestamp 18001
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2115_
timestamp 18001
transform 1 0 3404 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2116_
timestamp 18001
transform 1 0 3220 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2117_
timestamp 18001
transform 1 0 3680 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2118_
timestamp 18001
transform -1 0 3404 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2119_
timestamp 18001
transform -1 0 2576 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2120_
timestamp 18001
transform -1 0 3680 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2121_
timestamp 18001
transform 1 0 2116 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2122_
timestamp 18001
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2123_
timestamp 18001
transform -1 0 3864 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _2124_
timestamp 18001
transform -1 0 3680 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2125_
timestamp 18001
transform 1 0 3864 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2126_
timestamp 18001
transform 1 0 3220 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2127_
timestamp 18001
transform 1 0 2576 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_2  _2128_
timestamp 18001
transform -1 0 4968 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2129_
timestamp 18001
transform -1 0 5244 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2130_
timestamp 18001
transform -1 0 4784 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2131_
timestamp 18001
transform 1 0 4508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2132_
timestamp 18001
transform 1 0 4784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2133_
timestamp 18001
transform 1 0 4876 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2134_
timestamp 18001
transform 1 0 4876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2135_
timestamp 18001
transform -1 0 5152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2136_
timestamp 18001
transform -1 0 6072 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2137_
timestamp 18001
transform -1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2138_
timestamp 18001
transform -1 0 5428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2139_
timestamp 18001
transform 1 0 5336 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2140_
timestamp 18001
transform -1 0 5520 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2141_
timestamp 18001
transform 1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2142_
timestamp 18001
transform 1 0 4508 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _2143_
timestamp 18001
transform -1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2144_
timestamp 18001
transform 1 0 4508 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2145_
timestamp 18001
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2146_
timestamp 18001
transform 1 0 5244 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2147_
timestamp 18001
transform 1 0 4784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _2148_
timestamp 18001
transform 1 0 3772 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _2149_
timestamp 18001
transform -1 0 7544 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2150_
timestamp 18001
transform 1 0 6256 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2151_
timestamp 18001
transform 1 0 7360 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2152_
timestamp 18001
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2153_
timestamp 18001
transform -1 0 16376 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2154_
timestamp 18001
transform -1 0 15640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2155_
timestamp 18001
transform 1 0 14444 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_4  _2156_
timestamp 18001
transform 1 0 17664 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__or4b_2  _2157_
timestamp 18001
transform -1 0 17848 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2158_
timestamp 18001
transform -1 0 13892 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2159_
timestamp 18001
transform -1 0 17480 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2160_
timestamp 18001
transform 1 0 17480 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2161_
timestamp 18001
transform -1 0 15180 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2162_
timestamp 18001
transform -1 0 14352 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2163_
timestamp 18001
transform -1 0 14720 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _2164_
timestamp 18001
transform 1 0 18032 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _2165_
timestamp 18001
transform 1 0 18492 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2166_
timestamp 18001
transform -1 0 10304 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2167_
timestamp 18001
transform -1 0 11224 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2168_
timestamp 18001
transform -1 0 10948 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2169_
timestamp 18001
transform 1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2170_
timestamp 18001
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2171_
timestamp 18001
transform -1 0 17296 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2172_
timestamp 18001
transform 1 0 17940 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2173_
timestamp 18001
transform -1 0 16100 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2174_
timestamp 18001
transform -1 0 17112 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2175_
timestamp 18001
transform 1 0 12512 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _2176_
timestamp 18001
transform 1 0 12052 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2177_
timestamp 18001
transform 1 0 13892 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _2178_
timestamp 18001
transform 1 0 12512 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _2179_
timestamp 18001
transform -1 0 13524 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _2180_
timestamp 18001
transform 1 0 13340 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2181_
timestamp 18001
transform -1 0 12512 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2182_
timestamp 18001
transform -1 0 13432 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2183_
timestamp 18001
transform -1 0 13892 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2184_
timestamp 18001
transform 1 0 12604 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2185_
timestamp 18001
transform 1 0 5060 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2186_
timestamp 18001
transform 1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2187_
timestamp 18001
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2188_
timestamp 18001
transform 1 0 9568 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2189_
timestamp 18001
transform -1 0 10488 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2190_
timestamp 18001
transform 1 0 7912 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _2191_
timestamp 18001
transform -1 0 4508 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2192_
timestamp 18001
transform 1 0 5152 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2193_
timestamp 18001
transform 1 0 7084 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2194_
timestamp 18001
transform -1 0 8096 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2195_
timestamp 18001
transform -1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _2196_
timestamp 18001
transform -1 0 5152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2197_
timestamp 18001
transform -1 0 6992 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2198_
timestamp 18001
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2199_
timestamp 18001
transform 1 0 9660 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2200_
timestamp 18001
transform -1 0 10028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2201_
timestamp 18001
transform 1 0 8372 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2202_
timestamp 18001
transform 1 0 8004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2203_
timestamp 18001
transform 1 0 6624 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2204_
timestamp 18001
transform -1 0 7820 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2205_
timestamp 18001
transform -1 0 9936 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2206_
timestamp 18001
transform -1 0 10764 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2207_
timestamp 18001
transform 1 0 9200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2208_
timestamp 18001
transform 1 0 7268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2209_
timestamp 18001
transform 1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2210_
timestamp 18001
transform 1 0 4048 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2211_
timestamp 18001
transform 1 0 5244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2212_
timestamp 18001
transform 1 0 7176 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _2213_
timestamp 18001
transform -1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2214_
timestamp 18001
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2215_
timestamp 18001
transform -1 0 6256 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2216_
timestamp 18001
transform -1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _2217_
timestamp 18001
transform 1 0 9016 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2218_
timestamp 18001
transform -1 0 9660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2219_
timestamp 18001
transform -1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2220_
timestamp 18001
transform -1 0 8372 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2221_
timestamp 18001
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2222_
timestamp 18001
transform -1 0 8096 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2223_
timestamp 18001
transform 1 0 6348 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2224_
timestamp 18001
transform -1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _2225_
timestamp 18001
transform -1 0 2484 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _2226_
timestamp 18001
transform -1 0 2484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _2227_
timestamp 18001
transform -1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2228_
timestamp 18001
transform 1 0 10580 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2229_
timestamp 18001
transform 1 0 9844 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2230_
timestamp 18001
transform 1 0 30544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2231_
timestamp 18001
transform 1 0 16652 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _2232_
timestamp 18001
transform 1 0 15088 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _2233_
timestamp 18001
transform 1 0 5612 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2234_
timestamp 18001
transform -1 0 6348 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _2235_
timestamp 18001
transform -1 0 14536 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _2236_
timestamp 18001
transform 1 0 12328 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _2237_
timestamp 18001
transform -1 0 9936 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _2238_
timestamp 18001
transform 1 0 9200 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2239_
timestamp 18001
transform 1 0 14076 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2240_
timestamp 18001
transform -1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _2241_
timestamp 18001
transform -1 0 10948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2242_
timestamp 18001
transform -1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2243_
timestamp 18001
transform 1 0 12420 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _2244_
timestamp 18001
transform -1 0 14628 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _2245_
timestamp 18001
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2246_
timestamp 18001
transform -1 0 12972 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _2247_
timestamp 18001
transform 1 0 9016 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _2248_
timestamp 18001
transform -1 0 10120 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _2249_
timestamp 18001
transform 1 0 9752 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _2250_
timestamp 18001
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _2251_
timestamp 18001
transform 1 0 6164 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2252_
timestamp 18001
transform 1 0 8464 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2253_
timestamp 18001
transform -1 0 6256 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2254_
timestamp 18001
transform -1 0 6808 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2255_
timestamp 18001
transform 1 0 6716 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2256_
timestamp 18001
transform -1 0 8188 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2257_
timestamp 18001
transform 1 0 7820 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2258_
timestamp 18001
transform 1 0 6808 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2259_
timestamp 18001
transform 1 0 8004 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2260_
timestamp 18001
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2261_
timestamp 18001
transform 1 0 8004 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2262_
timestamp 18001
transform -1 0 10396 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2263_
timestamp 18001
transform 1 0 9752 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2264_
timestamp 18001
transform 1 0 11132 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2265_
timestamp 18001
transform -1 0 12420 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2266_
timestamp 18001
transform 1 0 10028 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2267_
timestamp 18001
transform -1 0 11408 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2268_
timestamp 18001
transform 1 0 11500 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2269_
timestamp 18001
transform -1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2270_
timestamp 18001
transform 1 0 10948 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2271_
timestamp 18001
transform 1 0 11776 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2272_
timestamp 18001
transform 1 0 13524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2273_
timestamp 18001
transform 1 0 13892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2274_
timestamp 18001
transform 1 0 12972 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2275_
timestamp 18001
transform 1 0 14904 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2276_
timestamp 18001
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2277_
timestamp 18001
transform 1 0 15364 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2278_
timestamp 18001
transform 1 0 14812 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2279_
timestamp 18001
transform 1 0 12972 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2280_
timestamp 18001
transform 1 0 14720 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2281_
timestamp 18001
transform 1 0 13248 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2282_
timestamp 18001
transform 1 0 11592 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2283_
timestamp 18001
transform -1 0 11592 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2284_
timestamp 18001
transform 1 0 12972 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2285_
timestamp 18001
transform 1 0 10948 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2286_
timestamp 18001
transform -1 0 11960 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2287_
timestamp 18001
transform -1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2288_
timestamp 18001
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2289_
timestamp 18001
transform -1 0 12144 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2290_
timestamp 18001
transform 1 0 12696 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2291_
timestamp 18001
transform -1 0 12788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2292_
timestamp 18001
transform -1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2293_
timestamp 18001
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2294_
timestamp 18001
transform 1 0 12788 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2295_
timestamp 18001
transform 1 0 14076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2296_
timestamp 18001
transform 1 0 13340 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2297_
timestamp 18001
transform 1 0 7084 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _2298_
timestamp 18001
transform -1 0 6900 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2299_
timestamp 18001
transform 1 0 7084 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2300_
timestamp 18001
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _2301_
timestamp 18001
transform 1 0 7636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2302_
timestamp 18001
transform 1 0 8924 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2303_
timestamp 18001
transform 1 0 7636 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2304_
timestamp 18001
transform -1 0 8280 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2305_
timestamp 18001
transform 1 0 8280 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a311oi_4  _2306_
timestamp 18001
transform 1 0 4876 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _2307_
timestamp 18001
transform 1 0 6808 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _2308_
timestamp 18001
transform -1 0 7452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2309_
timestamp 18001
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _2310_
timestamp 18001
transform 1 0 7544 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2311_
timestamp 18001
transform 1 0 8188 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2312_
timestamp 18001
transform -1 0 8096 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2313_
timestamp 18001
transform 1 0 6900 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2314_
timestamp 18001
transform -1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2315_
timestamp 18001
transform 1 0 8280 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2316_
timestamp 18001
transform 1 0 9108 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2317_
timestamp 18001
transform -1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2318_
timestamp 18001
transform 1 0 8188 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2319_
timestamp 18001
transform 1 0 9200 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2320_
timestamp 18001
transform -1 0 8556 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2321_
timestamp 18001
transform 1 0 9568 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2322_
timestamp 18001
transform -1 0 9660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2323_
timestamp 18001
transform -1 0 19872 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2324_
timestamp 18001
transform -1 0 20608 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2325_
timestamp 18001
transform -1 0 21528 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2326_
timestamp 18001
transform 1 0 21068 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2327_
timestamp 18001
transform 1 0 24380 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2328_
timestamp 18001
transform -1 0 27600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2329_
timestamp 18001
transform 1 0 26220 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2330_
timestamp 18001
transform -1 0 29348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2331_
timestamp 18001
transform 1 0 28796 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2332_
timestamp 18001
transform -1 0 33488 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2333_
timestamp 18001
transform 1 0 32936 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2334_
timestamp 18001
transform 1 0 33948 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2335_
timestamp 18001
transform 1 0 37168 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2336_
timestamp 18001
transform 1 0 37628 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2337_
timestamp 18001
transform 1 0 38272 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2338_
timestamp 18001
transform 1 0 1932 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2339_
timestamp 18001
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2340_
timestamp 18001
transform 1 0 3588 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2341_
timestamp 18001
transform 1 0 3128 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2342_
timestamp 18001
transform -1 0 2944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2343_
timestamp 18001
transform -1 0 7912 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _2344_
timestamp 18001
transform 1 0 5244 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_1  _2345_
timestamp 18001
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2346_
timestamp 18001
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2347_
timestamp 18001
transform -1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2348_
timestamp 18001
transform -1 0 4968 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2349_
timestamp 18001
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2350_
timestamp 18001
transform -1 0 6348 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2351_
timestamp 18001
transform 1 0 7636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2352_
timestamp 18001
transform -1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2353_
timestamp 18001
transform 1 0 5336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2354_
timestamp 18001
transform 1 0 5612 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2355_
timestamp 18001
transform -1 0 6900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2356_
timestamp 18001
transform 1 0 5152 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2357_
timestamp 18001
transform -1 0 9384 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2358_
timestamp 18001
transform -1 0 6900 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2359_
timestamp 18001
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2360_
timestamp 18001
transform 1 0 9660 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2361_
timestamp 18001
transform -1 0 10396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2362_
timestamp 18001
transform 1 0 8188 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2363_
timestamp 18001
transform -1 0 10304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2364_
timestamp 18001
transform -1 0 11408 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2365_
timestamp 18001
transform 1 0 9936 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2366_
timestamp 18001
transform 1 0 10304 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2367_
timestamp 18001
transform 1 0 9568 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2368_
timestamp 18001
transform -1 0 10396 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2369_
timestamp 18001
transform -1 0 9568 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2370_
timestamp 18001
transform -1 0 10304 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2371_
timestamp 18001
transform -1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2372_
timestamp 18001
transform 1 0 10488 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2373_
timestamp 18001
transform -1 0 11500 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2374_
timestamp 18001
transform 1 0 10948 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2375_
timestamp 18001
transform -1 0 5888 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _2376_
timestamp 18001
transform -1 0 6072 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2377_
timestamp 18001
transform 1 0 4692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2378_
timestamp 18001
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2379_
timestamp 18001
transform 1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2380_
timestamp 18001
transform 1 0 4508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2381_
timestamp 18001
transform -1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2382_
timestamp 18001
transform -1 0 5152 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2383_
timestamp 18001
transform 1 0 2760 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2384_
timestamp 18001
transform 1 0 4324 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2385_
timestamp 18001
transform 1 0 3404 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _2386_
timestamp 18001
transform -1 0 4508 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _2387_
timestamp 18001
transform 1 0 2208 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2388_
timestamp 18001
transform 1 0 3220 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2389_
timestamp 18001
transform 1 0 2024 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2390_
timestamp 18001
transform 1 0 1932 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2391_
timestamp 18001
transform -1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2392_
timestamp 18001
transform -1 0 5060 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2393_
timestamp 18001
transform 1 0 4048 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _2394_
timestamp 18001
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2395_
timestamp 18001
transform 1 0 4968 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2396_
timestamp 18001
transform -1 0 5980 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _2397_
timestamp 18001
transform -1 0 6256 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2398_
timestamp 18001
transform -1 0 5612 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _2399_
timestamp 18001
transform 1 0 4324 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2400_
timestamp 18001
transform 1 0 3036 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2401_
timestamp 18001
transform -1 0 6808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _2402_
timestamp 18001
transform -1 0 7360 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2403_
timestamp 18001
transform -1 0 6808 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2404_
timestamp 18001
transform 1 0 6532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2405_
timestamp 18001
transform -1 0 7544 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2406_
timestamp 18001
transform 1 0 6440 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2407_
timestamp 18001
transform 1 0 6532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2408_
timestamp 18001
transform -1 0 8740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2409_
timestamp 18001
transform -1 0 9384 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2410_
timestamp 18001
transform -1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2411_
timestamp 18001
transform -1 0 9108 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2412_
timestamp 18001
transform 1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2413_
timestamp 18001
transform -1 0 10304 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2414_
timestamp 18001
transform -1 0 11500 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2415_
timestamp 18001
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2416_
timestamp 18001
transform -1 0 10028 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2417_
timestamp 18001
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2418_
timestamp 18001
transform 1 0 10212 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2419_
timestamp 18001
transform -1 0 9292 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2420_
timestamp 18001
transform -1 0 9568 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2421_
timestamp 18001
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2422_
timestamp 18001
transform -1 0 10120 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _2423_
timestamp 18001
transform -1 0 13064 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2424_
timestamp 18001
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2425_
timestamp 18001
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _2426_
timestamp 18001
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _2427_
timestamp 18001
transform -1 0 10672 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _2428_
timestamp 18001
transform 1 0 16652 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _2429_
timestamp 18001
transform -1 0 17112 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2430_
timestamp 18001
transform 1 0 18032 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _2431_
timestamp 18001
transform 1 0 18952 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2432_
timestamp 18001
transform -1 0 20516 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2433_
timestamp 18001
transform 1 0 16100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2434_
timestamp 18001
transform 1 0 6348 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2435_
timestamp 18001
transform 1 0 6348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2436_
timestamp 18001
transform 1 0 7360 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2437_
timestamp 18001
transform 1 0 7360 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2438_
timestamp 18001
transform -1 0 9752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2439_
timestamp 18001
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2440_
timestamp 18001
transform -1 0 11408 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2441_
timestamp 18001
transform 1 0 10580 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2442_
timestamp 18001
transform 1 0 11500 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2443_
timestamp 18001
transform -1 0 13892 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2444_
timestamp 18001
transform 1 0 13616 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2445_
timestamp 18001
transform -1 0 14904 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2446_
timestamp 18001
transform -1 0 14720 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2447_
timestamp 18001
transform 1 0 13616 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2448_
timestamp 18001
transform 1 0 11500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2449_
timestamp 18001
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2450_
timestamp 18001
transform 1 0 11040 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2451_
timestamp 18001
transform -1 0 13984 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2452_
timestamp 18001
transform -1 0 14720 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2453_
timestamp 18001
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2454_
timestamp 18001
transform 1 0 3956 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2455_
timestamp 18001
transform 1 0 4324 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _2456_
timestamp 18001
transform 1 0 5520 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2457_
timestamp 18001
transform 1 0 2944 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2458_
timestamp 18001
transform 1 0 5152 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2459_
timestamp 18001
transform 1 0 6808 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2460_
timestamp 18001
transform 1 0 6808 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2461_
timestamp 18001
transform 1 0 5244 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2462_
timestamp 18001
transform 1 0 3772 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2463_
timestamp 18001
transform 1 0 1656 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2464_
timestamp 18001
transform 1 0 1380 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2465_
timestamp 18001
transform 1 0 1380 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2466_
timestamp 18001
transform 1 0 1840 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2467_
timestamp 18001
transform 1 0 4784 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2468_
timestamp 18001
transform 1 0 6992 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2469_
timestamp 18001
transform 1 0 8096 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2470_
timestamp 18001
transform 1 0 6900 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2471_
timestamp 18001
transform 1 0 4232 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2472_
timestamp 18001
transform -1 0 8188 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2473_
timestamp 18001
transform 1 0 1656 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2474_
timestamp 18001
transform 1 0 1380 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2475_
timestamp 18001
transform 1 0 1380 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2476_
timestamp 18001
transform 1 0 1380 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2477_
timestamp 18001
transform 1 0 6164 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2478_
timestamp 18001
transform 1 0 9660 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2479_
timestamp 18001
transform 1 0 8924 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2480_
timestamp 18001
transform 1 0 8924 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2481_
timestamp 18001
transform 1 0 9108 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2482_
timestamp 18001
transform 1 0 9752 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2483_
timestamp 18001
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2484_
timestamp 18001
transform 1 0 9292 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _2485_
timestamp 18001
transform -1 0 20700 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2486_
timestamp 18001
transform -1 0 20516 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2487_
timestamp 18001
transform 1 0 19596 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2488_
timestamp 18001
transform -1 0 22724 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2489_
timestamp 18001
transform -1 0 25760 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2490_
timestamp 18001
transform -1 0 26680 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2491_
timestamp 18001
transform -1 0 29348 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2492_
timestamp 18001
transform 1 0 28612 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2493_
timestamp 18001
transform 1 0 29532 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2494_
timestamp 18001
transform 1 0 30728 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2495_
timestamp 18001
transform -1 0 35788 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2496_
timestamp 18001
transform -1 0 35052 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2497_
timestamp 18001
transform -1 0 37168 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2498_
timestamp 18001
transform 1 0 39100 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2499_
timestamp 18001
transform -1 0 40204 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2500_
timestamp 18001
transform 1 0 1380 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2501_
timestamp 18001
transform 1 0 1380 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2502_
timestamp 18001
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2503_
timestamp 18001
transform 1 0 1380 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2504_
timestamp 18001
transform 1 0 2392 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2505_
timestamp 18001
transform -1 0 3312 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2506_
timestamp 18001
transform 1 0 1380 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2507_
timestamp 18001
transform 1 0 3772 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2508_
timestamp 18001
transform 1 0 5704 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2509_
timestamp 18001
transform 1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2510_
timestamp 18001
transform -1 0 6808 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2511_
timestamp 18001
transform 1 0 6348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2512_
timestamp 18001
transform -1 0 10028 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2513_
timestamp 18001
transform 1 0 8924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2514_
timestamp 18001
transform 1 0 8096 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2515_
timestamp 18001
transform -1 0 12328 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2516_
timestamp 18001
transform -1 0 10304 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2517_
timestamp 18001
transform 1 0 9384 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2518_
timestamp 18001
transform 1 0 11500 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2519_
timestamp 18001
transform 1 0 11592 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2520_
timestamp 18001
transform 1 0 2852 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2521_
timestamp 18001
transform 1 0 1380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2522_
timestamp 18001
transform -1 0 5980 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2523_
timestamp 18001
transform 1 0 1380 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2524_
timestamp 18001
transform -1 0 3220 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2525_
timestamp 18001
transform -1 0 4324 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2526_
timestamp 18001
transform 1 0 3864 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2527_
timestamp 18001
transform 1 0 3128 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2528_
timestamp 18001
transform 1 0 6348 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2529_
timestamp 18001
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2530_
timestamp 18001
transform 1 0 7636 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2531_
timestamp 18001
transform 1 0 9476 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2532_
timestamp 18001
transform -1 0 12144 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2533_
timestamp 18001
transform 1 0 7636 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2534_
timestamp 18001
transform 1 0 10580 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2535_
timestamp 18001
transform 1 0 10672 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2536_
timestamp 18001
transform -1 0 3220 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2537_
timestamp 18001
transform -1 0 3220 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2538_
timestamp 18001
transform -1 0 3220 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2539_
timestamp 18001
transform 1 0 5428 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2540_
timestamp 18001
transform 1 0 2576 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2541_
timestamp 18001
transform 1 0 2576 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2542_
timestamp 18001
transform 1 0 2208 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2543_
timestamp 18001
transform 1 0 2392 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2544_
timestamp 18001
transform 1 0 14904 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2545_
timestamp 18001
transform 1 0 17020 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2546_
timestamp 18001
transform 1 0 19872 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2547_
timestamp 18001
transform 1 0 21804 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2548_
timestamp 18001
transform 1 0 22908 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2549_
timestamp 18001
transform 1 0 24932 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2550_
timestamp 18001
transform 1 0 26956 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2551_
timestamp 18001
transform 1 0 27600 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2552_
timestamp 18001
transform 1 0 30176 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2553_
timestamp 18001
transform 1 0 31188 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2554_
timestamp 18001
transform 1 0 37352 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2555_
timestamp 18001
transform 1 0 37352 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2556_
timestamp 18001
transform 1 0 35236 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2557_
timestamp 18001
transform 1 0 34684 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2558_
timestamp 18001
transform 1 0 32752 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2559_
timestamp 18001
transform 1 0 17112 0 -1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2560_
timestamp 18001
transform 1 0 16652 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2561_
timestamp 18001
transform -1 0 21344 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2562_
timestamp 18001
transform 1 0 21068 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2563_
timestamp 18001
transform -1 0 25024 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2564_
timestamp 18001
transform 1 0 24012 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2565_
timestamp 18001
transform 1 0 26128 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2566_
timestamp 18001
transform 1 0 27508 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2567_
timestamp 18001
transform 1 0 29440 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2568_
timestamp 18001
transform 1 0 30820 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2569_
timestamp 18001
transform 1 0 38364 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2570_
timestamp 18001
transform 1 0 37720 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2571_
timestamp 18001
transform 1 0 35420 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2572_
timestamp 18001
transform 1 0 34316 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2573_
timestamp 18001
transform 1 0 32384 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _2574_
timestamp 18001
transform 1 0 9200 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2575_
timestamp 18001
transform 1 0 11776 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2576_
timestamp 18001
transform 1 0 10580 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2577_
timestamp 18001
transform 1 0 9568 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2578_
timestamp 18001
transform -1 0 9292 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2579_
timestamp 18001
transform 1 0 16928 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2580_
timestamp 18001
transform 1 0 16836 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2581_
timestamp 18001
transform -1 0 23276 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2582_
timestamp 18001
transform -1 0 22448 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2583_
timestamp 18001
transform 1 0 22448 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2584_
timestamp 18001
transform 1 0 23368 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2585_
timestamp 18001
transform 1 0 25668 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2586_
timestamp 18001
transform 1 0 27140 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2587_
timestamp 18001
transform 1 0 27968 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2588_
timestamp 18001
transform 1 0 30176 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2589_
timestamp 18001
transform 1 0 32108 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2590_
timestamp 18001
transform 1 0 32660 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2591_
timestamp 18001
transform 1 0 35144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2592_
timestamp 18001
transform 1 0 37260 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2593_
timestamp 18001
transform 1 0 37260 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2594_
timestamp 18001
transform 1 0 12880 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2595_
timestamp 18001
transform 1 0 14076 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2596_
timestamp 18001
transform 1 0 15456 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2597_
timestamp 18001
transform 1 0 16652 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2598_
timestamp 18001
transform 1 0 19504 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2599_
timestamp 18001
transform 1 0 21252 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2600_
timestamp 18001
transform 1 0 22356 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 18001
transform 1 0 25300 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2602_
timestamp 18001
transform 1 0 25760 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2603_
timestamp 18001
transform 1 0 27784 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2604_
timestamp 18001
transform -1 0 31464 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2605_
timestamp 18001
transform 1 0 30176 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2606_
timestamp 18001
transform 1 0 36064 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2607_
timestamp 18001
transform -1 0 39928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2608_
timestamp 18001
transform -1 0 38732 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2609_
timestamp 18001
transform 1 0 37536 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2610_
timestamp 18001
transform 1 0 32752 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2611_
timestamp 18001
transform 1 0 14720 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2612_
timestamp 18001
transform -1 0 19872 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 18001
transform -1 0 19136 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2614_
timestamp 18001
transform 1 0 20424 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 18001
transform 1 0 22356 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 18001
transform -1 0 24932 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2617_
timestamp 18001
transform -1 0 27416 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2618_
timestamp 18001
transform -1 0 29164 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2619_
timestamp 18001
transform -1 0 30452 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2620_
timestamp 18001
transform 1 0 30912 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2621_
timestamp 18001
transform 1 0 32752 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2622_
timestamp 18001
transform -1 0 39284 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2623_
timestamp 18001
transform 1 0 40388 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2624_
timestamp 18001
transform 1 0 40388 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2625_
timestamp 18001
transform 1 0 40388 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2626_
timestamp 18001
transform 1 0 34592 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2627_
timestamp 18001
transform -1 0 16744 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2628_
timestamp 18001
transform 1 0 15272 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2629_
timestamp 18001
transform 1 0 17112 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2630_
timestamp 18001
transform 1 0 19872 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2631_
timestamp 18001
transform -1 0 23644 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2632_
timestamp 18001
transform 1 0 23000 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2633_
timestamp 18001
transform 1 0 25024 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2634_
timestamp 18001
transform 1 0 27140 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2635_
timestamp 18001
transform 1 0 28428 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2636_
timestamp 18001
transform 1 0 30084 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2637_
timestamp 18001
transform 1 0 32292 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2638_
timestamp 18001
transform 1 0 37260 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2639_
timestamp 18001
transform 1 0 40296 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2640_
timestamp 18001
transform 1 0 40204 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2641_
timestamp 18001
transform -1 0 39560 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2642_
timestamp 18001
transform 1 0 34684 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 18001
transform 1 0 18216 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2644_
timestamp 18001
transform 1 0 17204 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2645_
timestamp 18001
transform 1 0 19412 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2646_
timestamp 18001
transform 1 0 21252 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2647_
timestamp 18001
transform 1 0 23000 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 18001
transform 1 0 24380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2649_
timestamp 18001
transform 1 0 25760 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2650_
timestamp 18001
transform 1 0 27140 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2651_
timestamp 18001
transform -1 0 31648 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2652_
timestamp 18001
transform 1 0 30728 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2653_
timestamp 18001
transform 1 0 32568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2654_
timestamp 18001
transform 1 0 33028 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2655_
timestamp 18001
transform 1 0 34500 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2656_
timestamp 18001
transform 1 0 35236 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2657_
timestamp 18001
transform 1 0 35328 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2658_
timestamp 18001
transform -1 0 19136 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 18001
transform 1 0 15456 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 18001
transform 1 0 20608 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2661_
timestamp 18001
transform 1 0 21804 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2662_
timestamp 18001
transform -1 0 26772 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2663_
timestamp 18001
transform 1 0 24288 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 18001
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2665_
timestamp 18001
transform 1 0 27416 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2666_
timestamp 18001
transform 1 0 30912 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2667_
timestamp 18001
transform 1 0 30636 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2668_
timestamp 18001
transform 1 0 35328 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2669_
timestamp 18001
transform 1 0 39192 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2670_
timestamp 18001
transform 1 0 38272 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2671_
timestamp 18001
transform 1 0 39652 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2672_
timestamp 18001
transform -1 0 37536 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2673_
timestamp 18001
transform 1 0 13064 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2674_
timestamp 18001
transform 1 0 15272 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2675_
timestamp 18001
transform 1 0 28796 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2676_
timestamp 18001
transform 1 0 26956 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2677_
timestamp 18001
transform 1 0 16652 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2678_
timestamp 18001
transform 1 0 29532 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2679_
timestamp 18001
transform 1 0 14260 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2680_
timestamp 18001
transform 1 0 14812 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2681_
timestamp 18001
transform 1 0 17112 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 18001
transform 1 0 19872 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 18001
transform 1 0 20792 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 18001
transform 1 0 22632 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 18001
transform 1 0 24748 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 18001
transform 1 0 26312 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2687_
timestamp 18001
transform 1 0 28888 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 18001
transform 1 0 30176 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 18001
transform 1 0 32476 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 18001
transform 1 0 35144 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2691_
timestamp 18001
transform 1 0 37260 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 18001
transform 1 0 33764 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 18001
transform -1 0 38088 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 18001
transform 1 0 32384 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 18001
transform 1 0 16008 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 18001
transform 1 0 13248 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2697_
timestamp 18001
transform 1 0 14720 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2698_
timestamp 18001
transform 1 0 17940 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2699_
timestamp 18001
transform 1 0 20332 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2700_
timestamp 18001
transform 1 0 22172 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 18001
transform 1 0 24104 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 18001
transform 1 0 25852 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2703_
timestamp 18001
transform 1 0 27416 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2704_
timestamp 18001
transform -1 0 31372 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2705_
timestamp 18001
transform 1 0 30176 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2706_
timestamp 18001
transform 1 0 40388 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2707_
timestamp 18001
transform -1 0 41952 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2708_
timestamp 18001
transform 1 0 37352 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2709_
timestamp 18001
transform 1 0 34776 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2710_
timestamp 18001
transform 1 0 32384 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2711_
timestamp 18001
transform 1 0 13156 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2712_
timestamp 18001
transform 1 0 15456 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2713_
timestamp 18001
transform 1 0 18124 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2714_
timestamp 18001
transform -1 0 22448 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2715_
timestamp 18001
transform 1 0 22448 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2716_
timestamp 18001
transform 1 0 24380 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2717_
timestamp 18001
transform 1 0 26220 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2718_
timestamp 18001
transform 1 0 27600 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2719_
timestamp 18001
transform 1 0 29532 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2720_
timestamp 18001
transform 1 0 30176 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2721_
timestamp 18001
transform 1 0 40020 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2722_
timestamp 18001
transform 1 0 40112 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2723_
timestamp 18001
transform 1 0 37352 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2724_
timestamp 18001
transform 1 0 34960 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2725_
timestamp 18001
transform 1 0 32476 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2726_
timestamp 18001
transform 1 0 11500 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2727_
timestamp 18001
transform 1 0 14904 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2728_
timestamp 18001
transform 1 0 16744 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2729_
timestamp 18001
transform 1 0 19780 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2730_
timestamp 18001
transform 1 0 20424 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2731_
timestamp 18001
transform 1 0 22908 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2732_
timestamp 18001
transform 1 0 25024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2733_
timestamp 18001
transform 1 0 26956 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2734_
timestamp 18001
transform 1 0 29532 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2735_
timestamp 18001
transform 1 0 30268 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2736_
timestamp 18001
transform 1 0 32108 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2737_
timestamp 18001
transform 1 0 37260 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2738_
timestamp 18001
transform 1 0 39284 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2739_
timestamp 18001
transform 1 0 39376 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2740_
timestamp 18001
transform 1 0 37628 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2741_
timestamp 18001
transform 1 0 34132 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2742_
timestamp 18001
transform -1 0 15548 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2743_
timestamp 18001
transform 1 0 11040 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2744_
timestamp 18001
transform 1 0 8372 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2745_
timestamp 18001
transform 1 0 7360 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2746_
timestamp 18001
transform 1 0 6900 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2747_
timestamp 18001
transform 1 0 9936 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2748_
timestamp 18001
transform 1 0 14076 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2749_
timestamp 18001
transform -1 0 17388 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2750_
timestamp 18001
transform 1 0 18676 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2751_
timestamp 18001
transform 1 0 20884 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2752_
timestamp 18001
transform 1 0 22816 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2753_
timestamp 18001
transform 1 0 24564 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2754_
timestamp 18001
transform 1 0 26956 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2755_
timestamp 18001
transform 1 0 28428 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2756_
timestamp 18001
transform 1 0 29440 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2757_
timestamp 18001
transform 1 0 30820 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2758_
timestamp 18001
transform 1 0 40572 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2759_
timestamp 18001
transform 1 0 39376 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2760_
timestamp 18001
transform 1 0 37352 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2761_
timestamp 18001
transform 1 0 35052 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2762_
timestamp 18001
transform 1 0 32568 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2763_
timestamp 18001
transform 1 0 11960 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2764_
timestamp 18001
transform -1 0 15640 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2765_
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2766_
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2767_
timestamp 18001
transform 1 0 21804 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2768_
timestamp 18001
transform -1 0 24196 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2769_
timestamp 18001
transform 1 0 24748 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2770_
timestamp 18001
transform 1 0 26404 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2771_
timestamp 18001
transform -1 0 29716 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2772_
timestamp 18001
transform 1 0 29532 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2773_
timestamp 18001
transform -1 0 32476 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2774_
timestamp 18001
transform 1 0 40296 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2775_
timestamp 18001
transform 1 0 39836 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2776_
timestamp 18001
transform 1 0 37352 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2777_
timestamp 18001
transform 1 0 35052 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2778_
timestamp 18001
transform 1 0 32568 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2779_
timestamp 18001
transform -1 0 14076 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2780_
timestamp 18001
transform 1 0 9936 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2781_
timestamp 18001
transform 1 0 10856 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2782_
timestamp 18001
transform 1 0 9292 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2783_
timestamp 18001
transform -1 0 11132 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2784_
timestamp 18001
transform 1 0 11868 0 1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2785_
timestamp 18001
transform 1 0 11500 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2786_
timestamp 18001
transform 1 0 11500 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2787_
timestamp 18001
transform 1 0 11500 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2788_
timestamp 18001
transform 1 0 10948 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2789_
timestamp 18001
transform -1 0 15088 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2790_
timestamp 18001
transform 1 0 19228 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2791_
timestamp 18001
transform 1 0 15640 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2792_
timestamp 18001
transform 1 0 17848 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2793_
timestamp 18001
transform 1 0 20976 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2794_
timestamp 18001
transform -1 0 24196 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2795_
timestamp 18001
transform 1 0 24380 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2796_
timestamp 18001
transform 1 0 27140 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2797_
timestamp 18001
transform 1 0 27784 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2798_
timestamp 18001
transform 1 0 40388 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2799_
timestamp 18001
transform 1 0 40388 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2800_
timestamp 18001
transform 1 0 40388 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2801_
timestamp 18001
transform 1 0 38824 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2802_
timestamp 18001
transform 1 0 40388 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2803_
timestamp 18001
transform 1 0 40388 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2804_
timestamp 18001
transform 1 0 39652 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2805_
timestamp 18001
transform 1 0 40388 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2806_
timestamp 18001
transform 1 0 18124 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2807_
timestamp 18001
transform 1 0 14444 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2808_
timestamp 18001
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2809_
timestamp 18001
transform 1 0 13156 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2810_
timestamp 18001
transform 1 0 12696 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _2811_
timestamp 18001
transform 1 0 18308 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2812_
timestamp 18001
transform 1 0 17664 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2813_
timestamp 18001
transform 1 0 19780 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2814_
timestamp 18001
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2815_
timestamp 18001
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2816_
timestamp 18001
transform -1 0 26312 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2817_
timestamp 18001
transform -1 0 27324 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2818_
timestamp 18001
transform -1 0 28428 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2819_
timestamp 18001
transform 1 0 31648 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2820_
timestamp 18001
transform 1 0 33120 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2821_
timestamp 18001
transform -1 0 34868 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2822_
timestamp 18001
transform -1 0 36340 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2823_
timestamp 18001
transform 1 0 34960 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2824_
timestamp 18001
transform -1 0 37076 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2825_
timestamp 18001
transform 1 0 34592 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2826_
timestamp 18001
transform 1 0 13708 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _2827_
timestamp 18001
transform -1 0 3312 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2828_
timestamp 18001
transform 1 0 1380 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2829_
timestamp 18001
transform 1 0 3772 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2830_
timestamp 18001
transform 1 0 15088 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 18001
transform -1 0 28612 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 18001
transform -1 0 29716 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform 1 0 21896 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 18001
transform -1 0 13064 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 18001
transform 1 0 11316 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 18001
transform 1 0 32108 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 18001
transform 1 0 32200 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_clk
timestamp 18001
transform -1 0 4784 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_clk
timestamp 18001
transform 1 0 10120 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_clk
timestamp 18001
transform -1 0 16192 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_clk
timestamp 18001
transform 1 0 17480 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_clk
timestamp 18001
transform 1 0 11408 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_clk
timestamp 18001
transform 1 0 3864 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_clk
timestamp 18001
transform 1 0 6164 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_clk
timestamp 18001
transform 1 0 6624 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_clk
timestamp 18001
transform -1 0 4232 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_clk
timestamp 18001
transform 1 0 12328 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_clk
timestamp 18001
transform 1 0 17940 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_clk
timestamp 18001
transform 1 0 17204 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_clk
timestamp 18001
transform 1 0 18124 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_clk
timestamp 18001
transform -1 0 23644 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_clk
timestamp 18001
transform 1 0 27324 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_clk
timestamp 18001
transform 1 0 23276 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_clk
timestamp 18001
transform -1 0 28428 0 1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_clk
timestamp 18001
transform 1 0 32108 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_clk
timestamp 18001
transform 1 0 38088 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_clk
timestamp 18001
transform 1 0 40848 0 1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_clk
timestamp 18001
transform 1 0 37260 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_21_clk
timestamp 18001
transform 1 0 38732 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_22_clk
timestamp 18001
transform -1 0 35696 0 1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_23_clk
timestamp 18001
transform 1 0 31280 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_24_clk
timestamp 18001
transform -1 0 28336 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_25_clk
timestamp 18001
transform 1 0 32016 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_26_clk
timestamp 18001
transform 1 0 37996 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_27_clk
timestamp 18001
transform 1 0 38272 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_28_clk
timestamp 18001
transform 1 0 35788 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_29_clk
timestamp 18001
transform -1 0 36248 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_30_clk
timestamp 18001
transform -1 0 31464 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_31_clk
timestamp 18001
transform -1 0 25668 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_32_clk
timestamp 18001
transform 1 0 28244 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_33_clk
timestamp 18001
transform 1 0 21252 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_34_clk
timestamp 18001
transform 1 0 17204 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_35_clk
timestamp 18001
transform 1 0 20700 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_36_clk
timestamp 18001
transform -1 0 12328 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_37_clk
timestamp 18001
transform -1 0 6072 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_38_clk
timestamp 18001
transform -1 0 4784 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_39_clk
timestamp 18001
transform 1 0 6808 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 18001
transform 1 0 11500 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload1
timestamp 18001
transform 1 0 11500 0 -1 34816
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinvlp_4  clkload2
timestamp 18001
transform 1 0 32200 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload3
timestamp 18001
transform 1 0 3772 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_4  clkload4
timestamp 18001
transform 1 0 10396 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  clkload5
timestamp 18001
transform 1 0 16376 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 18001
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_12  clkload7
timestamp 18001
transform -1 0 23000 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload8
timestamp 18001
transform 1 0 10672 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload9
timestamp 18001
transform 1 0 5060 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload10
timestamp 18001
transform 1 0 3220 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 18001
transform 1 0 6440 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload12
timestamp 18001
transform 1 0 17480 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload13
timestamp 18001
transform 1 0 3864 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload14
timestamp 18001
transform 1 0 6348 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload15
timestamp 18001
transform 1 0 6624 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload16
timestamp 18001
transform 1 0 3772 0 1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_4  clkload17
timestamp 18001
transform 1 0 12328 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload18
timestamp 18001
transform 1 0 17940 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  clkload19
timestamp 18001
transform 1 0 17388 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__inv_12  clkload20
timestamp 18001
transform 1 0 18124 0 -1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  clkload21
timestamp 18001
transform 1 0 32844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload22
timestamp 18001
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_8  clkload23
timestamp 18001
transform 1 0 38272 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload24
timestamp 18001
transform 1 0 35788 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload25
timestamp 18001
transform 1 0 35236 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_12  clkload26
timestamp 18001
transform 1 0 29532 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload27
timestamp 18001
transform 1 0 24656 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload28
timestamp 18001
transform 1 0 27048 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload29
timestamp 18001
transform 1 0 24380 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload30
timestamp 18001
transform 1 0 22908 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload31
timestamp 18001
transform 1 0 27416 0 -1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload32
timestamp 18001
transform 1 0 31372 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_8  clkload33
timestamp 18001
transform 1 0 38088 0 -1 41344
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload34
timestamp 18001
transform 1 0 40848 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  clkload35
timestamp 18001
transform 1 0 36800 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload36
timestamp 18001
transform 1 0 39836 0 1 26112
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_8  clkload37
timestamp 18001
transform 1 0 34684 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  clkload38
timestamp 18001
transform 1 0 30452 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 18001
transform 1 0 35328 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 18001
transform -1 0 36064 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 18001
transform -1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 18001
transform -1 0 16284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 18001
transform 1 0 28612 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 18001
transform 1 0 5060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 18001
transform -1 0 3404 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout38
timestamp 18001
transform 1 0 3312 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 18001
transform -1 0 13984 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 18001
transform -1 0 28796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 18001
transform 1 0 33304 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 18001
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 18001
transform -1 0 16100 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout44
timestamp 18001
transform 1 0 32200 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 18001
transform -1 0 24196 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 18001
transform 1 0 38824 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 18001
transform -1 0 21068 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 18001
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 18001
transform -1 0 24472 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout50
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 18001
transform 1 0 21068 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 18001
transform 1 0 32292 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 18001
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout54
timestamp 18001
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 18001
transform 1 0 18676 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout56
timestamp 18001
transform 1 0 32660 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 18001
transform -1 0 19872 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout58
timestamp 18001
transform 1 0 34316 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout59
timestamp 18001
transform -1 0 13984 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 18001
transform 1 0 20792 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp 18001
transform -1 0 28888 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 18001
transform 1 0 34040 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 18001
transform -1 0 16560 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp 18001
transform 1 0 25392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 18001
transform -1 0 13800 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout66
timestamp 18001
transform -1 0 29348 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 18001
transform -1 0 15732 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout68
timestamp 18001
transform 1 0 29256 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout69
timestamp 18001
transform 1 0 39836 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 18001
transform 1 0 15456 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 18001
transform 1 0 20332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 18001
transform 1 0 20700 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 18001
transform -1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 18001
transform 1 0 29624 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 18001
transform -1 0 17296 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 18001
transform -1 0 17296 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 18001
transform 1 0 29532 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout78
timestamp 18001
transform -1 0 18676 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 18001
transform 1 0 19872 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout80
timestamp 18001
transform 1 0 28244 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 18001
transform -1 0 18860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 18001
transform 1 0 3312 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 18001
transform -1 0 32476 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout85
timestamp 18001
transform -1 0 36340 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout86
timestamp 18001
transform -1 0 19044 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout87
timestamp 18001
transform 1 0 29624 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 18001
transform -1 0 29716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp 18001
transform -1 0 29900 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 18001
transform 1 0 38456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 18001
transform -1 0 39468 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout92
timestamp 18001
transform -1 0 4968 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 18001
transform -1 0 29348 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout94
timestamp 18001
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout95
timestamp 18001
transform 1 0 33212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout96
timestamp 18001
transform 1 0 32844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 18001
transform -1 0 18216 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 18001
transform -1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout99
timestamp 18001
transform -1 0 32016 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout100
timestamp 18001
transform 1 0 34960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 18001
transform -1 0 29624 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 18001
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout103
timestamp 18001
transform -1 0 28336 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout104
timestamp 18001
transform 1 0 31464 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout105
timestamp 18001
transform 1 0 15364 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout106
timestamp 18001
transform 1 0 28796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout107
timestamp 18001
transform 1 0 34592 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout108
timestamp 18001
transform 1 0 14996 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout109
timestamp 18001
transform -1 0 12328 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout110
timestamp 18001
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 18001
transform 1 0 26312 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout112
timestamp 18001
transform 1 0 36340 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout113
timestamp 18001
transform -1 0 13984 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout114
timestamp 18001
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout115
timestamp 18001
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout116
timestamp 18001
transform 1 0 13984 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout117
timestamp 18001
transform -1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout118
timestamp 18001
transform -1 0 7636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 18001
transform -1 0 12696 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout120
timestamp 18001
transform -1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout121
timestamp 18001
transform -1 0 6164 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout122
timestamp 18001
transform -1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout123
timestamp 18001
transform -1 0 10672 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout124
timestamp 18001
transform 1 0 22540 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout125
timestamp 18001
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout126
timestamp 18001
transform 1 0 22724 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout127
timestamp 18001
transform -1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout128
timestamp 18001
transform 1 0 6808 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout129
timestamp 18001
transform -1 0 6900 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout130
timestamp 18001
transform -1 0 9200 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout131
timestamp 18001
transform -1 0 13708 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout132
timestamp 18001
transform -1 0 16560 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout133
timestamp 18001
transform -1 0 21712 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout134
timestamp 18001
transform -1 0 19872 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout135
timestamp 18001
transform -1 0 16008 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout136
timestamp 18001
transform 1 0 21068 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout137
timestamp 18001
transform -1 0 23552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout138
timestamp 18001
transform -1 0 27600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout139
timestamp 18001
transform -1 0 32660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout140
timestamp 18001
transform 1 0 25852 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout141
timestamp 18001
transform -1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout142
timestamp 18001
transform 1 0 30636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout143
timestamp 18001
transform 1 0 39192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout144
timestamp 18001
transform -1 0 38456 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout145
timestamp 18001
transform 1 0 41676 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout146
timestamp 18001
transform 1 0 41768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout147
timestamp 18001
transform 1 0 40572 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout148
timestamp 18001
transform -1 0 32660 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout149
timestamp 18001
transform -1 0 32752 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout150
timestamp 18001
transform 1 0 32752 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout151
timestamp 18001
transform -1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout152
timestamp 18001
transform -1 0 42228 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout153
timestamp 18001
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout154
timestamp 18001
transform 1 0 37260 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout155
timestamp 18001
transform -1 0 42044 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout156
timestamp 18001
transform 1 0 41124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout157
timestamp 18001
transform -1 0 39744 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636986456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 18001
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 18001
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_119
timestamp 1636986456
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 18001
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 18001
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636986456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636986456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636986456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636986456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636986456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636986456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 18001
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636986456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636986456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 18001
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636986456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636986456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 18001
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636986456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636986456
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 18001
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636986456
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1636986456
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 18001
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1636986456
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1636986456
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 18001
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1636986456
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_405
timestamp 1636986456
transform 1 0 38364 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 18001
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1636986456
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1636986456
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_445
timestamp 18001
transform 1 0 42044 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_15
timestamp 18001
transform 1 0 2484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_21
timestamp 18001
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 18001
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_69
timestamp 18001
transform 1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 18001
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 18001
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_56
timestamp 1636986456
transform 1 0 6256 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_68
timestamp 18001
transform 1 0 7360 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 18001
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 18001
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_98
timestamp 18001
transform 1 0 10120 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_113
timestamp 1636986456
transform 1 0 11500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_125
timestamp 1636986456
transform 1 0 12604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 18001
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 18001
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 18001
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 18001
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 18001
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 18001
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_100
timestamp 18001
transform 1 0 10304 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_109
timestamp 18001
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 18001
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_50
timestamp 18001
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_71
timestamp 18001
transform 1 0 7636 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 18001
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_126
timestamp 1636986456
transform 1 0 12696 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 18001
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636986456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636986456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636986456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 18001
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636986456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636986456
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 18001
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 18001
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1636986456
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1636986456
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 18001
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 18001
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1636986456
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1636986456
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 18001
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 18001
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636986456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_445
timestamp 18001
transform 1 0 42044 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 18001
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 18001
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 18001
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_77
timestamp 18001
transform 1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 18001
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 18001
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 18001
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_119
timestamp 1636986456
transform 1 0 12052 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_131
timestamp 1636986456
transform 1 0 13156 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_143
timestamp 1636986456
transform 1 0 14260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_155
timestamp 1636986456
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636986456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636986456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636986456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636986456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 18001
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 18001
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636986456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636986456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636986456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 18001
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 18001
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636986456
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636986456
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636986456
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 18001
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1636986456
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1636986456
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1636986456
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 18001
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 18001
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1636986456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1636986456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 18001
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 18001
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 18001
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 18001
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_49
timestamp 18001
transform 1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 18001
transform 1 0 6348 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_70
timestamp 1636986456
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 18001
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_89
timestamp 18001
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_98
timestamp 18001
transform 1 0 10120 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_102
timestamp 18001
transform 1 0 10488 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_123
timestamp 1636986456
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 18001
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 18001
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636986456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636986456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636986456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636986456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 18001
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 18001
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636986456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636986456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636986456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636986456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 18001
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 18001
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636986456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636986456
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636986456
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 18001
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 18001
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636986456
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1636986456
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1636986456
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1636986456
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 18001
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 18001
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1636986456
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1636986456
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1636986456
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1636986456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 18001
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 18001
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1636986456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636986456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_445
timestamp 18001
transform 1 0 42044 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636986456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 18001
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636986456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_69
timestamp 18001
transform 1 0 7452 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_104
timestamp 18001
transform 1 0 10672 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_120
timestamp 1636986456
transform 1 0 12144 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_132
timestamp 1636986456
transform 1 0 13248 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_144
timestamp 1636986456
transform 1 0 14352 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_156
timestamp 1636986456
transform 1 0 15456 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636986456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636986456
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636986456
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636986456
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 18001
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 18001
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636986456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636986456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636986456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636986456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 18001
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 18001
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636986456
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636986456
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636986456
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636986456
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 18001
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 18001
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1636986456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1636986456
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1636986456
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1636986456
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 18001
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 18001
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1636986456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636986456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636986456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636986456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 18001
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp 18001
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 18001
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_67
timestamp 1636986456
transform 1 0 7268 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp 18001
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_101
timestamp 18001
transform 1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 18001
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 18001
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636986456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636986456
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636986456
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636986456
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 18001
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 18001
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636986456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636986456
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636986456
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636986456
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 18001
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 18001
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636986456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636986456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636986456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636986456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 18001
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636986456
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1636986456
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1636986456
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1636986456
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 18001
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 18001
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1636986456
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1636986456
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1636986456
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1636986456
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 18001
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 18001
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1636986456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636986456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_445
timestamp 18001
transform 1 0 42044 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 18001
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 18001
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 18001
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 18001
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_80
timestamp 18001
transform 1 0 8464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp 18001
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_92
timestamp 1636986456
transform 1 0 9568 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_104
timestamp 18001
transform 1 0 10672 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_122
timestamp 1636986456
transform 1 0 12328 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_134
timestamp 1636986456
transform 1 0 13432 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_146
timestamp 1636986456
transform 1 0 14536 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 18001
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 18001
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636986456
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636986456
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 18001
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636986456
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_241
timestamp 18001
transform 1 0 23276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_247
timestamp 18001
transform 1 0 23828 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_268
timestamp 1636986456
transform 1 0 25760 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_281
timestamp 18001
transform 1 0 26956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_288
timestamp 18001
transform 1 0 27600 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_320
timestamp 1636986456
transform 1 0 30544 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 18001
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1636986456
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_369
timestamp 18001
transform 1 0 35052 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1636986456
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636986456
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1636986456
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1636986456
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 18001
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 18001
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_44
timestamp 18001
transform 1 0 5152 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_53
timestamp 18001
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 18001
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_92
timestamp 1636986456
transform 1 0 9568 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_122
timestamp 1636986456
transform 1 0 12328 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_134
timestamp 18001
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636986456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636986456
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636986456
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636986456
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 18001
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 18001
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 18001
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_206
timestamp 18001
transform 1 0 20056 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 18001
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_263
timestamp 18001
transform 1 0 25300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 18001
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 18001
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 18001
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_369
timestamp 18001
transform 1 0 35052 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_398
timestamp 1636986456
transform 1 0 37720 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_410
timestamp 18001
transform 1 0 38824 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 18001
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1636986456
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1636986456
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_445
timestamp 18001
transform 1 0 42044 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 18001
transform 1 0 3956 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 18001
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 18001
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 18001
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 18001
transform 1 0 6808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_68
timestamp 18001
transform 1 0 7360 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 18001
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_87
timestamp 1636986456
transform 1 0 9108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_99
timestamp 1636986456
transform 1 0 10212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 18001
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636986456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636986456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636986456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636986456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 18001
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 18001
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_238
timestamp 18001
transform 1 0 23000 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_242
timestamp 18001
transform 1 0 23368 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_251
timestamp 18001
transform 1 0 24196 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_260
timestamp 1636986456
transform 1 0 25024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_272
timestamp 18001
transform 1 0 26128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_297
timestamp 18001
transform 1 0 28428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_307
timestamp 18001
transform 1 0 29348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_368
timestamp 18001
transform 1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 18001
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_401
timestamp 1636986456
transform 1 0 37996 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_413
timestamp 1636986456
transform 1 0 39100 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_425
timestamp 1636986456
transform 1 0 40204 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_437
timestamp 18001
transform 1 0 41308 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_445
timestamp 18001
transform 1 0 42044 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_42
timestamp 18001
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_46
timestamp 18001
transform 1 0 5336 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_52
timestamp 18001
transform 1 0 5888 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_56
timestamp 1636986456
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_68
timestamp 1636986456
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 18001
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 18001
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 18001
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_113
timestamp 1636986456
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_125
timestamp 1636986456
transform 1 0 12604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 18001
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636986456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636986456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636986456
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 18001
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 18001
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_204
timestamp 18001
transform 1 0 19872 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_212
timestamp 18001
transform 1 0 20608 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_241
timestamp 18001
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 18001
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_256
timestamp 1636986456
transform 1 0 24656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_268
timestamp 18001
transform 1 0 25760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_281
timestamp 18001
transform 1 0 26956 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_355
timestamp 18001
transform 1 0 33764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_365
timestamp 18001
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_399
timestamp 1636986456
transform 1 0 37812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_411
timestamp 18001
transform 1 0 38916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 18001
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1636986456
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636986456
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_445
timestamp 18001
transform 1 0 42044 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 18001
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 18001
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_66
timestamp 18001
transform 1 0 7176 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_73
timestamp 1636986456
transform 1 0 7820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_85
timestamp 18001
transform 1 0 8924 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_133
timestamp 1636986456
transform 1 0 13340 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_145
timestamp 1636986456
transform 1 0 14444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_157
timestamp 18001
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 18001
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636986456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1636986456
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636986456
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1636986456
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 18001
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 18001
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 18001
transform 1 0 23184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_262
timestamp 18001
transform 1 0 25208 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_270
timestamp 18001
transform 1 0 25944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 18001
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_288
timestamp 18001
transform 1 0 27600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 18001
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_342
timestamp 18001
transform 1 0 32568 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_370
timestamp 18001
transform 1 0 35144 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_379
timestamp 18001
transform 1 0 35972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 18001
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 18001
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_433
timestamp 1636986456
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_445
timestamp 18001
transform 1 0 42044 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 18001
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 18001
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_40
timestamp 18001
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_50
timestamp 18001
transform 1 0 5704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 18001
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 18001
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 18001
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636986456
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636986456
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636986456
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_177
timestamp 18001
transform 1 0 17388 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 18001
transform 1 0 18124 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 18001
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_212
timestamp 1636986456
transform 1 0 20608 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 18001
transform 1 0 21712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 18001
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_234
timestamp 18001
transform 1 0 22632 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 18001
transform 1 0 23552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 18001
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_257
timestamp 18001
transform 1 0 24748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_278
timestamp 18001
transform 1 0 26680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_282
timestamp 18001
transform 1 0 27048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 18001
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_317
timestamp 18001
transform 1 0 30268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_328
timestamp 18001
transform 1 0 31280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_334
timestamp 18001
transform 1 0 31832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_345
timestamp 18001
transform 1 0 32844 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_349
timestamp 18001
transform 1 0 33212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_362
timestamp 18001
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1636986456
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 18001
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_385
timestamp 18001
transform 1 0 36524 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_401
timestamp 18001
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_405
timestamp 18001
transform 1 0 38364 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1636986456
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_445
timestamp 18001
transform 1 0 42044 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_36
timestamp 18001
transform 1 0 4416 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_44
timestamp 18001
transform 1 0 5152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 18001
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 18001
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_64
timestamp 18001
transform 1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 18001
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp 18001
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 18001
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 18001
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 18001
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636986456
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636986456
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 18001
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 18001
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 18001
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 18001
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_241
timestamp 18001
transform 1 0 23276 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 18001
transform 1 0 23828 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 18001
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 18001
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_288
timestamp 18001
transform 1 0 27600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_292
timestamp 18001
transform 1 0 27968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_311
timestamp 18001
transform 1 0 29716 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_320
timestamp 1636986456
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 18001
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_384
timestamp 18001
transform 1 0 36432 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_396
timestamp 18001
transform 1 0 37536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_411
timestamp 18001
transform 1 0 38916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_415
timestamp 18001
transform 1 0 39284 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_420
timestamp 1636986456
transform 1 0 39744 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_432
timestamp 1636986456
transform 1 0 40848 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_444
timestamp 18001
transform 1 0 41952 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_19
timestamp 18001
transform 1 0 2852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_33
timestamp 18001
transform 1 0 4140 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 18001
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 18001
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_64
timestamp 18001
transform 1 0 6992 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 18001
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 18001
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 18001
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 18001
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_126
timestamp 18001
transform 1 0 12696 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_132
timestamp 18001
transform 1 0 13248 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636986456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636986456
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636986456
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_177
timestamp 18001
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_185
timestamp 18001
transform 1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 18001
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 18001
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 18001
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 18001
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_253
timestamp 18001
transform 1 0 24380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_265
timestamp 18001
transform 1 0 25484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_288
timestamp 18001
transform 1 0 27600 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_296
timestamp 1636986456
transform 1 0 28336 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1636986456
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_321
timestamp 18001
transform 1 0 30636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_327
timestamp 18001
transform 1 0 31188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_341
timestamp 18001
transform 1 0 32476 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_353
timestamp 18001
transform 1 0 33580 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 18001
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_365
timestamp 18001
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 18001
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_381
timestamp 18001
transform 1 0 36156 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_406
timestamp 18001
transform 1 0 38456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_410
timestamp 18001
transform 1 0 38824 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 18001
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636986456
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636986456
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_445
timestamp 18001
transform 1 0 42044 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_16
timestamp 18001
transform 1 0 2576 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 18001
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_57
timestamp 18001
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636986456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 18001
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_89
timestamp 18001
transform 1 0 9292 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_98
timestamp 18001
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 18001
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_124
timestamp 18001
transform 1 0 12512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 18001
transform 1 0 13156 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_148
timestamp 1636986456
transform 1 0 14720 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 18001
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636986456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636986456
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 18001
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_233
timestamp 18001
transform 1 0 22540 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_237
timestamp 18001
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_271
timestamp 18001
transform 1 0 26036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 18001
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_297
timestamp 18001
transform 1 0 28428 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_305
timestamp 18001
transform 1 0 29164 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_311
timestamp 18001
transform 1 0 29716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 18001
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_344
timestamp 1636986456
transform 1 0 32752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_356
timestamp 18001
transform 1 0 33856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 18001
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_393
timestamp 18001
transform 1 0 37260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_404
timestamp 18001
transform 1 0 38272 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_433
timestamp 1636986456
transform 1 0 40940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_445
timestamp 18001
transform 1 0 42044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 18001
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_29
timestamp 18001
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_42
timestamp 18001
transform 1 0 4968 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_70
timestamp 1636986456
transform 1 0 7544 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 18001
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 18001
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_107
timestamp 18001
transform 1 0 10948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 18001
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_157
timestamp 1636986456
transform 1 0 15548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_169
timestamp 18001
transform 1 0 16652 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 18001
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 18001
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_230
timestamp 18001
transform 1 0 22264 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_238
timestamp 18001
transform 1 0 23000 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 18001
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_282
timestamp 18001
transform 1 0 27048 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_288
timestamp 18001
transform 1 0 27600 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 18001
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_338
timestamp 1636986456
transform 1 0 32200 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_350
timestamp 1636986456
transform 1 0 33304 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 18001
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 18001
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_375
timestamp 18001
transform 1 0 35604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_390
timestamp 18001
transform 1 0 36984 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1636986456
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1636986456
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_445
timestamp 18001
transform 1 0 42044 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_7
timestamp 18001
transform 1 0 1748 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_20
timestamp 18001
transform 1 0 2944 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_26
timestamp 18001
transform 1 0 3496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_31
timestamp 18001
transform 1 0 3956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 18001
transform 1 0 4324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_70
timestamp 18001
transform 1 0 7544 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_120
timestamp 18001
transform 1 0 12144 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_154
timestamp 1636986456
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 18001
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_174
timestamp 18001
transform 1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_209
timestamp 18001
transform 1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 18001
transform 1 0 21436 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_239
timestamp 18001
transform 1 0 23092 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_254
timestamp 18001
transform 1 0 24472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_264
timestamp 18001
transform 1 0 25392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 18001
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 18001
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_303
timestamp 18001
transform 1 0 28980 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 18001
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 18001
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_346
timestamp 18001
transform 1 0 32936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_367
timestamp 18001
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 18001
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_410
timestamp 1636986456
transform 1 0 38824 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_422
timestamp 1636986456
transform 1 0 39928 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_434
timestamp 1636986456
transform 1 0 41032 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_446
timestamp 18001
transform 1 0 42136 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_24
timestamp 18001
transform 1 0 3312 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_57
timestamp 18001
transform 1 0 6348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 18001
transform 1 0 8096 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_105
timestamp 18001
transform 1 0 10764 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_146
timestamp 18001
transform 1 0 14536 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 18001
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 18001
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_239
timestamp 1636986456
transform 1 0 23092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 18001
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_253
timestamp 18001
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_262
timestamp 18001
transform 1 0 25208 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_270
timestamp 18001
transform 1 0 25944 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_278
timestamp 18001
transform 1 0 26680 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_286
timestamp 18001
transform 1 0 27416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 18001
transform 1 0 28336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 18001
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_321
timestamp 18001
transform 1 0 30636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 18001
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_371
timestamp 18001
transform 1 0 35236 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_400
timestamp 18001
transform 1 0 37904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 18001
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 18001
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_429
timestamp 1636986456
transform 1 0 40572 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_3
timestamp 18001
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_11
timestamp 18001
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_37
timestamp 18001
transform 1 0 4508 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_45
timestamp 18001
transform 1 0 5244 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 18001
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 18001
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_75
timestamp 1636986456
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_87
timestamp 18001
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_91
timestamp 18001
transform 1 0 9476 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 18001
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 18001
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 18001
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_138
timestamp 1636986456
transform 1 0 13800 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 18001
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_193
timestamp 18001
transform 1 0 18860 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_217
timestamp 18001
transform 1 0 21068 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_242
timestamp 18001
transform 1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_250
timestamp 18001
transform 1 0 24104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_260
timestamp 18001
transform 1 0 25024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 18001
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_327
timestamp 18001
transform 1 0 31188 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 18001
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 18001
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_393
timestamp 18001
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_417
timestamp 18001
transform 1 0 39468 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 18001
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_16
timestamp 1636986456
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636986456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 18001
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_101
timestamp 1636986456
transform 1 0 10396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_118
timestamp 18001
transform 1 0 11960 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_126
timestamp 18001
transform 1 0 12696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 18001
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 18001
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_179
timestamp 18001
transform 1 0 17572 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 18001
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636986456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 18001
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_230
timestamp 18001
transform 1 0 22264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 18001
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_279
timestamp 18001
transform 1 0 26772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 18001
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_313
timestamp 18001
transform 1 0 29900 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_321
timestamp 18001
transform 1 0 30636 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_353
timestamp 18001
transform 1 0 33580 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_373
timestamp 18001
transform 1 0 35420 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_394
timestamp 18001
transform 1 0 37352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_417
timestamp 18001
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_425
timestamp 18001
transform 1 0 40204 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_24
timestamp 1636986456
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_36
timestamp 18001
transform 1 0 4416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_44
timestamp 18001
transform 1 0 5152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 18001
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1636986456
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_129
timestamp 18001
transform 1 0 12972 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_135
timestamp 18001
transform 1 0 13524 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_152
timestamp 1636986456
transform 1 0 15088 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 18001
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636986456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_181
timestamp 18001
transform 1 0 17756 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 18001
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 18001
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_233
timestamp 18001
transform 1 0 22540 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 18001
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 18001
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_309
timestamp 18001
transform 1 0 29532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_357
timestamp 18001
transform 1 0 33948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_375
timestamp 18001
transform 1 0 35604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 18001
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_397
timestamp 18001
transform 1 0 37628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_445
timestamp 18001
transform 1 0 42044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 18001
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_37
timestamp 1636986456
transform 1 0 4508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 18001
transform 1 0 6256 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_63
timestamp 1636986456
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 18001
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 18001
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_93
timestamp 1636986456
transform 1 0 9660 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 18001
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 18001
transform 1 0 15272 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_202
timestamp 18001
transform 1 0 19688 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_211
timestamp 18001
transform 1 0 20516 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_232
timestamp 18001
transform 1 0 22448 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 18001
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 18001
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_253
timestamp 18001
transform 1 0 24380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_257
timestamp 18001
transform 1 0 24748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_266
timestamp 18001
transform 1 0 25576 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_296
timestamp 18001
transform 1 0 28336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 18001
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_352
timestamp 18001
transform 1 0 33488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 18001
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_365
timestamp 18001
transform 1 0 34684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_374
timestamp 18001
transform 1 0 35512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_396
timestamp 18001
transform 1 0 37536 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_415
timestamp 18001
transform 1 0 39284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 18001
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_421
timestamp 18001
transform 1 0 39836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_430
timestamp 18001
transform 1 0 40664 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_438
timestamp 18001
transform 1 0 41400 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_9
timestamp 18001
transform 1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 18001
transform 1 0 2484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_42
timestamp 1636986456
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 18001
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636986456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 18001
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_73
timestamp 18001
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_82
timestamp 1636986456
transform 1 0 8648 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_94
timestamp 1636986456
transform 1 0 9752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_106
timestamp 18001
transform 1 0 10856 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1636986456
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 18001
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 18001
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_194
timestamp 18001
transform 1 0 18952 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 18001
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636986456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636986456
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_249
timestamp 18001
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_260
timestamp 1636986456
transform 1 0 25024 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 18001
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_316
timestamp 18001
transform 1 0 30176 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_324
timestamp 18001
transform 1 0 30912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 18001
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_337
timestamp 18001
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_400
timestamp 18001
transform 1 0 37904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_444
timestamp 18001
transform 1 0 41952 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_37
timestamp 18001
transform 1 0 4508 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_47
timestamp 1636986456
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 18001
transform 1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_85
timestamp 18001
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_98
timestamp 1636986456
transform 1 0 10120 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_110
timestamp 1636986456
transform 1 0 11224 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 18001
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 18001
transform 1 0 14628 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 18001
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 18001
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636986456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 18001
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_218
timestamp 1636986456
transform 1 0 21160 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_230
timestamp 1636986456
transform 1 0 22264 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_242
timestamp 18001
transform 1 0 23368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_263
timestamp 18001
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_267
timestamp 18001
transform 1 0 25668 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_275
timestamp 1636986456
transform 1 0 26404 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_287
timestamp 18001
transform 1 0 27508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 18001
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_315
timestamp 18001
transform 1 0 30084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_323
timestamp 18001
transform 1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_336
timestamp 18001
transform 1 0 32016 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_352
timestamp 1636986456
transform 1 0 33488 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 18001
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_369
timestamp 18001
transform 1 0 35052 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1636986456
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_417
timestamp 18001
transform 1 0 39468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_6
timestamp 18001
transform 1 0 1656 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 18001
transform 1 0 2392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_50
timestamp 18001
transform 1 0 5704 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_83
timestamp 18001
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_87
timestamp 18001
transform 1 0 9108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 18001
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 18001
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 18001
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 18001
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 18001
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp 18001
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 18001
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 18001
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 18001
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 18001
transform 1 0 17848 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_228
timestamp 1636986456
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_240
timestamp 18001
transform 1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_267
timestamp 18001
transform 1 0 25668 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 18001
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_286
timestamp 18001
transform 1 0 27416 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_309
timestamp 1636986456
transform 1 0 29532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_321
timestamp 18001
transform 1 0 30636 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 18001
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_343
timestamp 18001
transform 1 0 32660 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1636986456
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_361
timestamp 18001
transform 1 0 34316 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_374
timestamp 1636986456
transform 1 0 35512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_386
timestamp 18001
transform 1 0 36616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_393
timestamp 18001
transform 1 0 37260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_408
timestamp 18001
transform 1 0 38640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_420
timestamp 18001
transform 1 0 39744 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_433
timestamp 18001
transform 1 0 40940 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 18001
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_37
timestamp 18001
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_54
timestamp 18001
transform 1 0 6072 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 18001
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_107
timestamp 1636986456
transform 1 0 10948 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_119
timestamp 18001
transform 1 0 12052 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_131
timestamp 18001
transform 1 0 13156 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_202
timestamp 18001
transform 1 0 19688 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_210
timestamp 18001
transform 1 0 20424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 18001
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_241
timestamp 18001
transform 1 0 23276 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 18001
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 18001
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 18001
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_289
timestamp 18001
transform 1 0 27692 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_298
timestamp 18001
transform 1 0 28520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 18001
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_347
timestamp 18001
transform 1 0 33028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_355
timestamp 18001
transform 1 0 33764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 18001
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_406
timestamp 1636986456
transform 1 0 38456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 18001
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1636986456
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_438
timestamp 18001
transform 1 0 41400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_446
timestamp 18001
transform 1 0 42136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_6
timestamp 18001
transform 1 0 1656 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 18001
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636986456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_69
timestamp 18001
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_77
timestamp 18001
transform 1 0 8188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp 18001
transform 1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_121
timestamp 18001
transform 1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_156
timestamp 1636986456
transform 1 0 15456 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 18001
transform 1 0 17388 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1636986456
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 18001
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 18001
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_232
timestamp 18001
transform 1 0 22448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_251
timestamp 18001
transform 1 0 24196 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_287
timestamp 18001
transform 1 0 27508 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_324
timestamp 18001
transform 1 0 30912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 18001
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_364
timestamp 18001
transform 1 0 34592 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_393
timestamp 18001
transform 1 0 37260 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_402
timestamp 18001
transform 1 0 38088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_414
timestamp 18001
transform 1 0 39192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_418
timestamp 18001
transform 1 0 39560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_426
timestamp 18001
transform 1 0 40296 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 18001
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_54
timestamp 18001
transform 1 0 6072 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_62
timestamp 1636986456
transform 1 0 6808 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 18001
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 18001
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_112
timestamp 18001
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_128
timestamp 1636986456
transform 1 0 12880 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_149
timestamp 18001
transform 1 0 14812 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_161
timestamp 1636986456
transform 1 0 15916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_173
timestamp 18001
transform 1 0 17020 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_184
timestamp 1636986456
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 18001
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_205
timestamp 18001
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 18001
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_230
timestamp 18001
transform 1 0 22264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 18001
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_261
timestamp 1636986456
transform 1 0 25116 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_273
timestamp 1636986456
transform 1 0 26220 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_285
timestamp 18001
transform 1 0 27324 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_293
timestamp 18001
transform 1 0 28060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_302
timestamp 18001
transform 1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_317
timestamp 18001
transform 1 0 30268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_349
timestamp 18001
transform 1 0 33212 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 18001
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 18001
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_365
timestamp 18001
transform 1 0 34684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_374
timestamp 18001
transform 1 0 35512 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_387
timestamp 18001
transform 1 0 36708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_415
timestamp 18001
transform 1 0 39284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 18001
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_421
timestamp 18001
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 18001
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 18001
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_43
timestamp 18001
transform 1 0 5060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_73
timestamp 18001
transform 1 0 7820 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_94
timestamp 18001
transform 1 0 9752 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 18001
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 18001
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_142
timestamp 18001
transform 1 0 14168 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_150
timestamp 18001
transform 1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_189
timestamp 18001
transform 1 0 18492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_197
timestamp 18001
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 18001
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_253
timestamp 1636986456
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 18001
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 18001
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 18001
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 18001
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_285
timestamp 18001
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_314
timestamp 18001
transform 1 0 29992 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_324
timestamp 1636986456
transform 1 0 30912 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 18001
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_352
timestamp 18001
transform 1 0 33488 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_356
timestamp 18001
transform 1 0 33856 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_388
timestamp 18001
transform 1 0 36800 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_404
timestamp 18001
transform 1 0 38272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_446
timestamp 18001
transform 1 0 42136 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636986456
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636986456
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_40
timestamp 18001
transform 1 0 4784 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp 18001
transform 1 0 5520 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_61
timestamp 1636986456
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 18001
transform 1 0 7820 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 18001
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 18001
transform 1 0 10396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_122
timestamp 18001
transform 1 0 12328 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 18001
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_141
timestamp 18001
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_149
timestamp 18001
transform 1 0 14812 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_177
timestamp 18001
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_213
timestamp 1636986456
transform 1 0 20700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_225
timestamp 1636986456
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_237
timestamp 1636986456
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 18001
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 18001
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_261
timestamp 18001
transform 1 0 25116 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_291
timestamp 18001
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 18001
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636986456
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_321
timestamp 18001
transform 1 0 30636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_336
timestamp 18001
transform 1 0 32016 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_353
timestamp 18001
transform 1 0 33580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 18001
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_375
timestamp 18001
transform 1 0 35604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_379
timestamp 18001
transform 1 0 35972 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_407
timestamp 18001
transform 1 0 38548 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_417
timestamp 18001
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_428
timestamp 18001
transform 1 0 40480 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_437
timestamp 18001
transform 1 0 41308 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 18001
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_19
timestamp 18001
transform 1 0 2852 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 18001
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636986456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636986456
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 18001
transform 1 0 8556 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_129
timestamp 1636986456
transform 1 0 12972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 18001
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_178
timestamp 18001
transform 1 0 17480 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 18001
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_235
timestamp 18001
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 18001
transform 1 0 24840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_310
timestamp 18001
transform 1 0 29624 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 18001
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 18001
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_422
timestamp 18001
transform 1 0 39928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 18001
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_36
timestamp 18001
transform 1 0 4416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_40
timestamp 18001
transform 1 0 4784 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_69
timestamp 1636986456
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 18001
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636986456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_97
timestamp 18001
transform 1 0 10028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_105
timestamp 18001
transform 1 0 10764 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_112
timestamp 1636986456
transform 1 0 11408 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_124
timestamp 1636986456
transform 1 0 12512 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 18001
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_169
timestamp 18001
transform 1 0 16652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_178
timestamp 18001
transform 1 0 17480 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_197
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 18001
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 18001
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 18001
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_303
timestamp 18001
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 18001
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_309
timestamp 18001
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_343
timestamp 18001
transform 1 0 32660 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_349
timestamp 18001
transform 1 0 33212 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 18001
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_380
timestamp 1636986456
transform 1 0 36064 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_427
timestamp 18001
transform 1 0 40388 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_445
timestamp 18001
transform 1 0 42044 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_11
timestamp 1636986456
transform 1 0 2116 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_23
timestamp 1636986456
transform 1 0 3220 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1636986456
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 18001
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1636986456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_73
timestamp 1636986456
transform 1 0 7820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_85
timestamp 18001
transform 1 0 8924 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_91
timestamp 18001
transform 1 0 9476 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1636986456
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 18001
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_121
timestamp 18001
transform 1 0 12236 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_131
timestamp 18001
transform 1 0 13156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_139
timestamp 18001
transform 1 0 13892 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 18001
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 18001
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_210
timestamp 18001
transform 1 0 20424 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_233
timestamp 18001
transform 1 0 22540 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 18001
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_306
timestamp 18001
transform 1 0 29256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_314
timestamp 18001
transform 1 0 29992 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 18001
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_353
timestamp 18001
transform 1 0 33580 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_378
timestamp 1636986456
transform 1 0 35880 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 18001
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_413
timestamp 18001
transform 1 0 39100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_446
timestamp 18001
transform 1 0 42136 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 18001
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 18001
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_51
timestamp 18001
transform 1 0 5796 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_59
timestamp 18001
transform 1 0 6532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_69
timestamp 18001
transform 1 0 7452 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 18001
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_103
timestamp 1636986456
transform 1 0 10580 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_115
timestamp 18001
transform 1 0 11684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 18001
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_167
timestamp 18001
transform 1 0 16468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 18001
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 18001
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_228
timestamp 18001
transform 1 0 22080 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 18001
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 18001
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_283
timestamp 18001
transform 1 0 27140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_302
timestamp 18001
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_318
timestamp 18001
transform 1 0 30360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_341
timestamp 18001
transform 1 0 32476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_359
timestamp 18001
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 18001
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_365
timestamp 18001
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_392
timestamp 18001
transform 1 0 37168 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_415
timestamp 18001
transform 1 0 39284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 18001
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 18001
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_445
timestamp 18001
transform 1 0 42044 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_23
timestamp 1636986456
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_35
timestamp 18001
transform 1 0 4324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 18001
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 18001
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_76
timestamp 18001
transform 1 0 8096 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_85
timestamp 18001
transform 1 0 8924 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 18001
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_134
timestamp 1636986456
transform 1 0 13432 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_153
timestamp 1636986456
transform 1 0 15180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 18001
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_177
timestamp 18001
transform 1 0 17388 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 18001
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 18001
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_253
timestamp 18001
transform 1 0 24380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_257
timestamp 18001
transform 1 0 24748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_274
timestamp 18001
transform 1 0 26312 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_37_333
timestamp 18001
transform 1 0 31740 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_345
timestamp 18001
transform 1 0 32844 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 18001
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_409
timestamp 18001
transform 1 0 38732 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_440
timestamp 18001
transform 1 0 41584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_7
timestamp 18001
transform 1 0 1748 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_13
timestamp 18001
transform 1 0 2300 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_32
timestamp 18001
transform 1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_63
timestamp 18001
transform 1 0 6900 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_70
timestamp 18001
transform 1 0 7544 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 18001
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_95
timestamp 18001
transform 1 0 9844 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_126
timestamp 1636986456
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 18001
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636986456
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_177
timestamp 18001
transform 1 0 17388 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 18001
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 18001
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 18001
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_209
timestamp 18001
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 18001
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 18001
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 18001
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_394
timestamp 18001
transform 1 0 37352 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 18001
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 18001
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_430
timestamp 18001
transform 1 0 40664 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636986456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1636986456
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_44
timestamp 1636986456
transform 1 0 5152 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_73
timestamp 1636986456
transform 1 0 7820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_93
timestamp 18001
transform 1 0 9660 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 18001
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 18001
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1636986456
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_195
timestamp 18001
transform 1 0 19044 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_210
timestamp 18001
transform 1 0 20424 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 18001
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_236
timestamp 18001
transform 1 0 22816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_268
timestamp 18001
transform 1 0 25760 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 18001
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_305
timestamp 18001
transform 1 0 29164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_315
timestamp 18001
transform 1 0 30084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_325
timestamp 18001
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 18001
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_344
timestamp 18001
transform 1 0 32752 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_350
timestamp 18001
transform 1 0 33304 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_359
timestamp 18001
transform 1 0 34132 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_372
timestamp 1636986456
transform 1 0 35328 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 18001
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 18001
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_39_410
timestamp 18001
transform 1 0 38824 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_432
timestamp 18001
transform 1 0 40848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_442
timestamp 18001
transform 1 0 41768 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_446
timestamp 18001
transform 1 0 42136 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 18001
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp 18001
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 18001
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636986456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_73
timestamp 18001
transform 1 0 7820 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_81
timestamp 18001
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 18001
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 18001
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 18001
transform 1 0 14444 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_168
timestamp 18001
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 18001
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_204
timestamp 18001
transform 1 0 19872 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_211
timestamp 18001
transform 1 0 20516 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_217
timestamp 18001
transform 1 0 21068 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_226
timestamp 1636986456
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_238
timestamp 1636986456
transform 1 0 23000 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 18001
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 18001
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_266
timestamp 18001
transform 1 0 25576 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_275
timestamp 1636986456
transform 1 0 26404 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_287
timestamp 18001
transform 1 0 27508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_295
timestamp 18001
transform 1 0 28244 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 18001
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 18001
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_314
timestamp 1636986456
transform 1 0 29992 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_326
timestamp 18001
transform 1 0 31096 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_335
timestamp 1636986456
transform 1 0 31924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_347
timestamp 1636986456
transform 1 0 33028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 18001
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 18001
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_365
timestamp 18001
transform 1 0 34684 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_369
timestamp 18001
transform 1 0 35052 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_388
timestamp 18001
transform 1 0 36800 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_398
timestamp 1636986456
transform 1 0 37720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_410
timestamp 18001
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 18001
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_421
timestamp 18001
transform 1 0 39836 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_28
timestamp 18001
transform 1 0 3680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_42
timestamp 1636986456
transform 1 0 4968 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 18001
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_78
timestamp 18001
transform 1 0 8280 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_84
timestamp 18001
transform 1 0 8832 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_97
timestamp 1636986456
transform 1 0 10028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_109
timestamp 18001
transform 1 0 11132 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_140
timestamp 18001
transform 1 0 13984 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_174
timestamp 18001
transform 1 0 17112 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_182
timestamp 18001
transform 1 0 17848 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_193
timestamp 18001
transform 1 0 18860 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_199
timestamp 18001
transform 1 0 19412 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_233
timestamp 1636986456
transform 1 0 22540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_257
timestamp 18001
transform 1 0 24748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_263
timestamp 18001
transform 1 0 25300 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_268
timestamp 1636986456
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_348
timestamp 18001
transform 1 0 33120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_360
timestamp 18001
transform 1 0 34224 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_375
timestamp 18001
transform 1 0 35604 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_384
timestamp 18001
transform 1 0 36432 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636986456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_15
timestamp 18001
transform 1 0 2484 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_49
timestamp 18001
transform 1 0 5612 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_71
timestamp 1636986456
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 18001
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_101
timestamp 1636986456
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_113
timestamp 18001
transform 1 0 11500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_123
timestamp 1636986456
transform 1 0 12420 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_135
timestamp 18001
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 18001
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 18001
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_149
timestamp 18001
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_157
timestamp 18001
transform 1 0 15548 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 18001
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 18001
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_197
timestamp 18001
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_205
timestamp 18001
transform 1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_211
timestamp 18001
transform 1 0 20516 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_219
timestamp 18001
transform 1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_233
timestamp 18001
transform 1 0 22540 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 18001
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_264
timestamp 18001
transform 1 0 25392 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_271
timestamp 18001
transform 1 0 26036 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 18001
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 18001
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 18001
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_384
timestamp 18001
transform 1 0 36432 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_388
timestamp 18001
transform 1 0 36800 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 18001
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_421
timestamp 18001
transform 1 0 39836 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_3
timestamp 18001
transform 1 0 1380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_9
timestamp 18001
transform 1 0 1932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_29
timestamp 18001
transform 1 0 3772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 18001
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 18001
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_63
timestamp 18001
transform 1 0 6900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_67
timestamp 18001
transform 1 0 7268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 18001
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1636986456
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_125
timestamp 18001
transform 1 0 12604 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_152
timestamp 1636986456
transform 1 0 15088 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 18001
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_169
timestamp 18001
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_173
timestamp 18001
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_197
timestamp 18001
transform 1 0 19228 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_205
timestamp 18001
transform 1 0 19964 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_214
timestamp 18001
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 18001
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_234
timestamp 18001
transform 1 0 22632 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_242
timestamp 18001
transform 1 0 23368 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_249
timestamp 18001
transform 1 0 24012 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_254
timestamp 18001
transform 1 0 24472 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 18001
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_285
timestamp 1636986456
transform 1 0 27324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_297
timestamp 18001
transform 1 0 28428 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_319
timestamp 18001
transform 1 0 30452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_381
timestamp 18001
transform 1 0 36156 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_401
timestamp 18001
transform 1 0 37996 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_407
timestamp 18001
transform 1 0 38548 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_415
timestamp 18001
transform 1 0 39284 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 18001
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_29
timestamp 18001
transform 1 0 3772 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 18001
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_101
timestamp 18001
transform 1 0 10396 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 18001
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 18001
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_158
timestamp 1636986456
transform 1 0 15640 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_170
timestamp 18001
transform 1 0 16744 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_176
timestamp 18001
transform 1 0 17296 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_188
timestamp 18001
transform 1 0 18400 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 18001
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_202
timestamp 18001
transform 1 0 19688 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_215
timestamp 18001
transform 1 0 20884 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_238
timestamp 18001
transform 1 0 23000 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 18001
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 18001
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 18001
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_263
timestamp 18001
transform 1 0 25300 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_270
timestamp 1636986456
transform 1 0 25944 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_282
timestamp 1636986456
transform 1 0 27048 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_294
timestamp 1636986456
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 18001
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_312
timestamp 1636986456
transform 1 0 29808 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_324
timestamp 1636986456
transform 1 0 30912 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_336
timestamp 18001
transform 1 0 32016 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_344
timestamp 18001
transform 1 0 32752 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_355
timestamp 18001
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 18001
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_378
timestamp 18001
transform 1 0 35880 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_386
timestamp 1636986456
transform 1 0 36616 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_398
timestamp 18001
transform 1 0 37720 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_407
timestamp 18001
transform 1 0 38548 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_445
timestamp 18001
transform 1 0 42044 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_7
timestamp 18001
transform 1 0 1748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_22
timestamp 18001
transform 1 0 3128 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_28
timestamp 18001
transform 1 0 3680 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 18001
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 18001
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 18001
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 18001
transform 1 0 7084 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 18001
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 18001
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_117
timestamp 18001
transform 1 0 11868 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_123
timestamp 18001
transform 1 0 12420 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_134
timestamp 18001
transform 1 0 13432 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636986456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 18001
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_188
timestamp 18001
transform 1 0 18400 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_195
timestamp 18001
transform 1 0 19044 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_199
timestamp 18001
transform 1 0 19412 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636986456
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636986456
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 18001
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_288
timestamp 1636986456
transform 1 0 27600 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_300
timestamp 18001
transform 1 0 28704 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_308
timestamp 18001
transform 1 0 29440 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_316
timestamp 1636986456
transform 1 0 30176 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_328
timestamp 18001
transform 1 0 31280 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1636986456
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1636986456
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1636986456
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1636986456
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 18001
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 18001
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 18001
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_408
timestamp 18001
transform 1 0 38640 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_430
timestamp 18001
transform 1 0 40664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_434
timestamp 18001
transform 1 0 41032 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp 18001
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_33
timestamp 18001
transform 1 0 4140 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_39
timestamp 18001
transform 1 0 4692 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_47
timestamp 1636986456
transform 1 0 5428 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_59
timestamp 1636986456
transform 1 0 6532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_71
timestamp 1636986456
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 18001
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 18001
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 18001
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_134
timestamp 18001
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636986456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_153
timestamp 18001
transform 1 0 15180 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_167
timestamp 18001
transform 1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 18001
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 18001
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636986456
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_209
timestamp 18001
transform 1 0 20332 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 18001
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 18001
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 18001
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_256
timestamp 1636986456
transform 1 0 24656 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_277
timestamp 18001
transform 1 0 26588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 18001
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 18001
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 18001
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_320
timestamp 18001
transform 1 0 30544 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_344
timestamp 18001
transform 1 0 32752 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_352
timestamp 18001
transform 1 0 33488 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_385
timestamp 1636986456
transform 1 0 36524 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_397
timestamp 18001
transform 1 0 37628 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 18001
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_421
timestamp 18001
transform 1 0 39836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_436
timestamp 18001
transform 1 0 41216 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_445
timestamp 18001
transform 1 0 42044 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636986456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636986456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_27
timestamp 18001
transform 1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_35
timestamp 18001
transform 1 0 4324 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_60
timestamp 1636986456
transform 1 0 6624 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_72
timestamp 18001
transform 1 0 7728 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_81
timestamp 18001
transform 1 0 8556 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_96
timestamp 1636986456
transform 1 0 9936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 18001
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_113
timestamp 18001
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_144
timestamp 18001
transform 1 0 14352 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 18001
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_174
timestamp 18001
transform 1 0 17112 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_193
timestamp 18001
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_206
timestamp 18001
transform 1 0 20056 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 18001
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 18001
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_246
timestamp 18001
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_258
timestamp 18001
transform 1 0 24840 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 18001
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 18001
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_285
timestamp 18001
transform 1 0 27324 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_293
timestamp 18001
transform 1 0 28060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_301
timestamp 18001
transform 1 0 28796 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_314
timestamp 18001
transform 1 0 29992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_343
timestamp 18001
transform 1 0 32660 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_359
timestamp 18001
transform 1 0 34132 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_401
timestamp 18001
transform 1 0 37996 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_409
timestamp 18001
transform 1 0 38732 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_414
timestamp 18001
transform 1 0 39192 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_15
timestamp 18001
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 18001
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_48_29
timestamp 18001
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_42
timestamp 18001
transform 1 0 4968 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_65
timestamp 18001
transform 1 0 7084 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 18001
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_99
timestamp 18001
transform 1 0 10212 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_110
timestamp 18001
transform 1 0 11224 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 18001
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_182
timestamp 18001
transform 1 0 17848 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 18001
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 18001
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_260
timestamp 18001
transform 1 0 25024 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_276
timestamp 1636986456
transform 1 0 26496 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_316
timestamp 18001
transform 1 0 30176 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_343
timestamp 18001
transform 1 0 32660 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_365
timestamp 18001
transform 1 0 34684 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_388
timestamp 18001
transform 1 0 36800 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_415
timestamp 18001
transform 1 0 39284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 18001
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_421
timestamp 18001
transform 1 0 39836 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_425
timestamp 18001
transform 1 0 40204 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_431
timestamp 18001
transform 1 0 40756 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_36
timestamp 18001
transform 1 0 4416 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_44
timestamp 18001
transform 1 0 5152 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 18001
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_57
timestamp 18001
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 18001
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636986456
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_139
timestamp 18001
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_165
timestamp 18001
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1636986456
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_205
timestamp 18001
transform 1 0 19964 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_211
timestamp 1636986456
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 18001
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_225
timestamp 18001
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_233
timestamp 18001
transform 1 0 22540 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_251
timestamp 1636986456
transform 1 0 24196 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_263
timestamp 18001
transform 1 0 25300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_267
timestamp 18001
transform 1 0 25668 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_271
timestamp 18001
transform 1 0 26036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 18001
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 18001
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 18001
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1636986456
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_305
timestamp 18001
transform 1 0 29164 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_311
timestamp 18001
transform 1 0 29716 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 18001
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_337
timestamp 18001
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_363
timestamp 18001
transform 1 0 34500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_371
timestamp 18001
transform 1 0 35236 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_375
timestamp 1636986456
transform 1 0 35604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_387
timestamp 18001
transform 1 0 36708 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 18001
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_404
timestamp 18001
transform 1 0 38272 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_439
timestamp 18001
transform 1 0 41492 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1636986456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_15
timestamp 18001
transform 1 0 2484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_36
timestamp 18001
transform 1 0 4416 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_44
timestamp 18001
transform 1 0 5152 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_51
timestamp 1636986456
transform 1 0 5796 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_63
timestamp 1636986456
transform 1 0 6900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_105
timestamp 1636986456
transform 1 0 10764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_117
timestamp 18001
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_125
timestamp 18001
transform 1 0 12604 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 18001
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 18001
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1636986456
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1636986456
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1636986456
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1636986456
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 18001
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 18001
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1636986456
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_217
timestamp 18001
transform 1 0 21068 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_230
timestamp 18001
transform 1 0 22264 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_234
timestamp 18001
transform 1 0 22632 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 18001
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 18001
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_253
timestamp 18001
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_262
timestamp 18001
transform 1 0 25208 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_273
timestamp 18001
transform 1 0 26220 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_279
timestamp 18001
transform 1 0 26772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_296
timestamp 18001
transform 1 0 28336 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_309
timestamp 18001
transform 1 0 29532 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_315
timestamp 18001
transform 1 0 30084 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_326
timestamp 18001
transform 1 0 31096 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_355
timestamp 18001
transform 1 0 33764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 18001
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_365
timestamp 18001
transform 1 0 34684 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_370
timestamp 18001
transform 1 0 35144 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_376
timestamp 18001
transform 1 0 35696 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_386
timestamp 18001
transform 1 0 36616 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_401
timestamp 18001
transform 1 0 37996 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_410
timestamp 18001
transform 1 0 38824 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 18001
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_426
timestamp 18001
transform 1 0 40296 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_15
timestamp 18001
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_30
timestamp 18001
transform 1 0 3864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 18001
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_77
timestamp 18001
transform 1 0 8188 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_83
timestamp 18001
transform 1 0 8740 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_92
timestamp 18001
transform 1 0 9568 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 18001
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_122
timestamp 18001
transform 1 0 12328 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 18001
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_169
timestamp 18001
transform 1 0 16652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_175
timestamp 18001
transform 1 0 17204 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_181
timestamp 18001
transform 1 0 17756 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 18001
transform 1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_207
timestamp 18001
transform 1 0 20148 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_218
timestamp 18001
transform 1 0 21160 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_245
timestamp 18001
transform 1 0 23644 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_256
timestamp 18001
transform 1 0 24656 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_313
timestamp 18001
transform 1 0 29900 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_327
timestamp 18001
transform 1 0 31188 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_337
timestamp 18001
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_380
timestamp 18001
transform 1 0 36064 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_390
timestamp 18001
transform 1 0 36984 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_406
timestamp 18001
transform 1 0 38456 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_419
timestamp 18001
transform 1 0 39652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_437
timestamp 18001
transform 1 0 41308 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_33
timestamp 18001
transform 1 0 4140 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_41
timestamp 18001
transform 1 0 4876 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_66
timestamp 1636986456
transform 1 0 7176 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 18001
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1636986456
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_97
timestamp 18001
transform 1 0 10028 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_137
timestamp 18001
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 18001
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_152
timestamp 18001
transform 1 0 15088 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_161
timestamp 18001
transform 1 0 15916 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_176
timestamp 18001
transform 1 0 17296 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_230
timestamp 1636986456
transform 1 0 22264 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_242
timestamp 18001
transform 1 0 23368 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 18001
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_264
timestamp 1636986456
transform 1 0 25392 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_276
timestamp 18001
transform 1 0 26496 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_282
timestamp 18001
transform 1 0 27048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_291
timestamp 18001
transform 1 0 27876 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 18001
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_311
timestamp 18001
transform 1 0 29716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_315
timestamp 18001
transform 1 0 30084 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_333
timestamp 18001
transform 1 0 31740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_337
timestamp 18001
transform 1 0 32108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_346
timestamp 1636986456
transform 1 0 32936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 18001
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_385
timestamp 18001
transform 1 0 36524 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_414
timestamp 18001
transform 1 0 39192 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_435
timestamp 1636986456
transform 1 0 41124 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 18001
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_33
timestamp 18001
transform 1 0 4140 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_41
timestamp 18001
transform 1 0 4876 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 18001
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_78
timestamp 18001
transform 1 0 8280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_86
timestamp 18001
transform 1 0 9016 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_109
timestamp 18001
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_124
timestamp 18001
transform 1 0 12512 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_204
timestamp 18001
transform 1 0 19872 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_212
timestamp 18001
transform 1 0 20608 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_221
timestamp 18001
transform 1 0 21436 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1636986456
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_264
timestamp 18001
transform 1 0 25392 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_290
timestamp 18001
transform 1 0 27784 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_294
timestamp 18001
transform 1 0 28152 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 18001
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 18001
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_346
timestamp 18001
transform 1 0 32936 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_359
timestamp 18001
transform 1 0 34132 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_374
timestamp 1636986456
transform 1 0 35512 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_386
timestamp 18001
transform 1 0 36616 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_400
timestamp 1636986456
transform 1 0 37904 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_412
timestamp 18001
transform 1 0 39008 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_15
timestamp 18001
transform 1 0 2484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 18001
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_29
timestamp 18001
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_37
timestamp 18001
transform 1 0 4508 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_52
timestamp 18001
transform 1 0 5888 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_56
timestamp 18001
transform 1 0 6256 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 18001
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 18001
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_125
timestamp 18001
transform 1 0 12604 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_133
timestamp 18001
transform 1 0 13340 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1636986456
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 18001
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_157
timestamp 18001
transform 1 0 15548 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_179
timestamp 18001
transform 1 0 17572 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_183
timestamp 18001
transform 1 0 17940 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 18001
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1636986456
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 18001
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_227
timestamp 1636986456
transform 1 0 21988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_239
timestamp 18001
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_243
timestamp 18001
transform 1 0 23460 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 18001
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_253
timestamp 18001
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_261
timestamp 18001
transform 1 0 25116 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 18001
transform 1 0 26036 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_291
timestamp 18001
transform 1 0 27876 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_297
timestamp 18001
transform 1 0 28428 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 18001
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_341
timestamp 18001
transform 1 0 32476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_362
timestamp 18001
transform 1 0 34408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_390
timestamp 18001
transform 1 0 36984 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_398
timestamp 18001
transform 1 0 37720 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_408
timestamp 18001
transform 1 0 38640 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_445
timestamp 18001
transform 1 0 42044 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 18001
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_16
timestamp 18001
transform 1 0 2576 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_31
timestamp 18001
transform 1 0 3956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_54
timestamp 18001
transform 1 0 6072 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 18001
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_65
timestamp 18001
transform 1 0 7084 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_88
timestamp 18001
transform 1 0 9200 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_104
timestamp 18001
transform 1 0 10672 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1636986456
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_150
timestamp 1636986456
transform 1 0 14904 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_162
timestamp 18001
transform 1 0 16008 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1636986456
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1636986456
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 18001
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_241
timestamp 18001
transform 1 0 23276 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_251
timestamp 18001
transform 1 0 24196 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 18001
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 18001
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 18001
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 18001
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_345
timestamp 18001
transform 1 0 32844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_365
timestamp 18001
transform 1 0 34684 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 18001
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 18001
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_393
timestamp 18001
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_418
timestamp 18001
transform 1 0 39560 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_442
timestamp 18001
transform 1 0 41768 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 18001
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_26
timestamp 18001
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_41
timestamp 18001
transform 1 0 4876 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_54
timestamp 18001
transform 1 0 6072 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_66
timestamp 18001
transform 1 0 7176 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_75
timestamp 18001
transform 1 0 8004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 18001
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 18001
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 18001
transform 1 0 9476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_124
timestamp 18001
transform 1 0 12512 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 18001
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_149
timestamp 18001
transform 1 0 14812 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_170
timestamp 18001
transform 1 0 16744 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_193
timestamp 18001
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 18001
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_208
timestamp 18001
transform 1 0 20240 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_218
timestamp 18001
transform 1 0 21160 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_233
timestamp 18001
transform 1 0 22540 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 18001
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_261
timestamp 18001
transform 1 0 25116 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_267
timestamp 18001
transform 1 0 25668 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 18001
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_309
timestamp 18001
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_322
timestamp 18001
transform 1 0 30728 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_339
timestamp 18001
transform 1 0 32292 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_358
timestamp 18001
transform 1 0 34040 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp 18001
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_385
timestamp 18001
transform 1 0 36524 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_418
timestamp 18001
transform 1 0 39560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_421
timestamp 18001
transform 1 0 39836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_436
timestamp 18001
transform 1 0 41216 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_445
timestamp 18001
transform 1 0 42044 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_34
timestamp 18001
transform 1 0 4232 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_42
timestamp 18001
transform 1 0 4968 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 18001
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 18001
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_113
timestamp 18001
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_117
timestamp 18001
transform 1 0 11868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 18001
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 18001
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 18001
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_183
timestamp 18001
transform 1 0 17940 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 18001
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_241
timestamp 18001
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_259
timestamp 18001
transform 1 0 24932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 18001
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 18001
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1636986456
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_293
timestamp 18001
transform 1 0 28060 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_302
timestamp 18001
transform 1 0 28888 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 18001
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_346
timestamp 18001
transform 1 0 32936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_350
timestamp 18001
transform 1 0 33304 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_360
timestamp 1636986456
transform 1 0 34224 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_372
timestamp 18001
transform 1 0 35328 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 18001
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_440
timestamp 18001
transform 1 0 41584 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_446
timestamp 18001
transform 1 0 42136 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1636986456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_41
timestamp 18001
transform 1 0 4876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_59
timestamp 18001
transform 1 0 6532 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 18001
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 18001
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 18001
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_148
timestamp 18001
transform 1 0 14720 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_186
timestamp 18001
transform 1 0 18216 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_213
timestamp 18001
transform 1 0 20700 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_231
timestamp 18001
transform 1 0 22356 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_235
timestamp 18001
transform 1 0 22724 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 18001
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_279
timestamp 18001
transform 1 0 26772 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_318
timestamp 1636986456
transform 1 0 30360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_339
timestamp 18001
transform 1 0 32292 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_348
timestamp 18001
transform 1 0 33120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 18001
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_365
timestamp 18001
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_395
timestamp 18001
transform 1 0 37444 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_445
timestamp 18001
transform 1 0 42044 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_15
timestamp 18001
transform 1 0 2484 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_23
timestamp 18001
transform 1 0 3220 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_28
timestamp 18001
transform 1 0 3680 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_59_37
timestamp 18001
transform 1 0 4508 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_57
timestamp 18001
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_84
timestamp 1636986456
transform 1 0 8832 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_96
timestamp 18001
transform 1 0 9936 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_102
timestamp 18001
transform 1 0 10488 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 18001
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_157
timestamp 18001
transform 1 0 15548 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_185
timestamp 18001
transform 1 0 18124 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_216
timestamp 18001
transform 1 0 20976 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_242
timestamp 18001
transform 1 0 23368 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_260
timestamp 18001
transform 1 0 25024 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 18001
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_285
timestamp 18001
transform 1 0 27324 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_312
timestamp 18001
transform 1 0 29808 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 18001
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_337
timestamp 18001
transform 1 0 32108 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_360
timestamp 18001
transform 1 0 34224 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_386
timestamp 18001
transform 1 0 36616 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 18001
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_414
timestamp 18001
transform 1 0 39192 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_432
timestamp 18001
transform 1 0 40848 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_442
timestamp 18001
transform 1 0 41768 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_446
timestamp 18001
transform 1 0 42136 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 18001
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_7
timestamp 18001
transform 1 0 1748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_60
timestamp 18001
transform 1 0 6624 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 18001
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 18001
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_124
timestamp 18001
transform 1 0 12512 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_132
timestamp 18001
transform 1 0 13248 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_144
timestamp 18001
transform 1 0 14352 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_156
timestamp 18001
transform 1 0 15456 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_160
timestamp 18001
transform 1 0 15824 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 18001
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_197
timestamp 18001
transform 1 0 19228 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_207
timestamp 18001
transform 1 0 20148 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_217
timestamp 18001
transform 1 0 21068 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_241
timestamp 18001
transform 1 0 23276 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_266
timestamp 18001
transform 1 0 25576 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_289
timestamp 18001
transform 1 0 27692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_293
timestamp 18001
transform 1 0 28060 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 18001
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 18001
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_317
timestamp 1636986456
transform 1 0 30268 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 18001
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_365
timestamp 18001
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_396
timestamp 18001
transform 1 0 37536 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_417
timestamp 18001
transform 1 0 39468 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_425
timestamp 18001
transform 1 0 40204 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_445
timestamp 18001
transform 1 0 42044 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_23
timestamp 18001
transform 1 0 3220 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 18001
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1636986456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_69
timestamp 18001
transform 1 0 7452 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_73
timestamp 1636986456
transform 1 0 7820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_85
timestamp 18001
transform 1 0 8924 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_109
timestamp 18001
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_133
timestamp 18001
transform 1 0 13340 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_140
timestamp 18001
transform 1 0 13984 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_146
timestamp 18001
transform 1 0 14536 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_178
timestamp 18001
transform 1 0 17480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 18001
transform 1 0 17848 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_212
timestamp 1636986456
transform 1 0 20608 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_234
timestamp 18001
transform 1 0 22632 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_246
timestamp 18001
transform 1 0 23736 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 18001
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 18001
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_294
timestamp 18001
transform 1 0 28152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_304
timestamp 18001
transform 1 0 29072 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 18001
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_369
timestamp 18001
transform 1 0 35052 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_373
timestamp 18001
transform 1 0 35420 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 18001
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_399
timestamp 18001
transform 1 0 37812 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_417
timestamp 18001
transform 1 0 39468 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_443
timestamp 18001
transform 1 0 41860 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_15
timestamp 18001
transform 1 0 2484 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_26
timestamp 18001
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_36
timestamp 1636986456
transform 1 0 4416 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_48
timestamp 1636986456
transform 1 0 5520 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_60
timestamp 18001
transform 1 0 6624 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_76
timestamp 18001
transform 1 0 8096 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_85
timestamp 18001
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 18001
transform 1 0 9476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_112
timestamp 18001
transform 1 0 11408 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_124
timestamp 18001
transform 1 0 12512 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_150
timestamp 18001
transform 1 0 14904 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1636986456
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 18001
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 18001
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_206
timestamp 18001
transform 1 0 20056 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 18001
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_269
timestamp 18001
transform 1 0 25852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_273
timestamp 18001
transform 1 0 26220 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_381
timestamp 18001
transform 1 0 36156 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_390
timestamp 18001
transform 1 0 36984 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_417
timestamp 18001
transform 1 0 39468 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_421
timestamp 18001
transform 1 0 39836 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_443
timestamp 18001
transform 1 0 41860 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 18001
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 18001
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 18001
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_88
timestamp 18001
transform 1 0 9200 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_96
timestamp 18001
transform 1 0 9936 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_126
timestamp 18001
transform 1 0 12696 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_184
timestamp 18001
transform 1 0 18032 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_213
timestamp 18001
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 18001
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_229
timestamp 18001
transform 1 0 22172 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_252
timestamp 18001
transform 1 0 24288 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_267
timestamp 18001
transform 1 0 25668 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 18001
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_293
timestamp 18001
transform 1 0 28060 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_301
timestamp 18001
transform 1 0 28796 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_312
timestamp 18001
transform 1 0 29808 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_337
timestamp 18001
transform 1 0 32108 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_350
timestamp 18001
transform 1 0 33304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_354
timestamp 18001
transform 1 0 33672 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_368
timestamp 18001
transform 1 0 34960 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_376
timestamp 18001
transform 1 0 35696 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 18001
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_414
timestamp 18001
transform 1 0 39192 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_444
timestamp 18001
transform 1 0 41952 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_88
timestamp 1636986456
transform 1 0 9200 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_100
timestamp 1636986456
transform 1 0 10304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_112
timestamp 18001
transform 1 0 11408 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 18001
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_155
timestamp 18001
transform 1 0 15364 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_206
timestamp 18001
transform 1 0 20056 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 18001
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_309
timestamp 18001
transform 1 0 29532 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_318
timestamp 18001
transform 1 0 30360 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_326
timestamp 18001
transform 1 0 31096 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_349
timestamp 18001
transform 1 0 33212 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 18001
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_375
timestamp 18001
transform 1 0 35604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_385
timestamp 18001
transform 1 0 36524 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_391
timestamp 18001
transform 1 0 37076 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_400
timestamp 1636986456
transform 1 0 37904 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_412
timestamp 18001
transform 1 0 39008 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_444
timestamp 18001
transform 1 0 41952 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 18001
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 18001
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 18001
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_78
timestamp 1636986456
transform 1 0 8280 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_90
timestamp 1636986456
transform 1 0 9384 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_102
timestamp 18001
transform 1 0 10488 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_110
timestamp 18001
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_113
timestamp 18001
transform 1 0 11500 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_121
timestamp 18001
transform 1 0 12236 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_129
timestamp 18001
transform 1 0 12972 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_150
timestamp 18001
transform 1 0 14904 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_159
timestamp 18001
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 18001
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_176
timestamp 1636986456
transform 1 0 17296 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_191
timestamp 18001
transform 1 0 18676 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_201
timestamp 18001
transform 1 0 19596 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_211
timestamp 18001
transform 1 0 20516 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_215
timestamp 18001
transform 1 0 20884 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_234
timestamp 18001
transform 1 0 22632 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_252
timestamp 1636986456
transform 1 0 24288 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_264
timestamp 1636986456
transform 1 0 25392 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 18001
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_281
timestamp 18001
transform 1 0 26956 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_295
timestamp 18001
transform 1 0 28244 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_307
timestamp 18001
transform 1 0 29348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_321
timestamp 18001
transform 1 0 30636 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_367
timestamp 1636986456
transform 1 0 34868 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_386
timestamp 18001
transform 1 0 36616 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_393
timestamp 18001
transform 1 0 37260 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_406
timestamp 1636986456
transform 1 0 38456 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_418
timestamp 18001
transform 1 0 39560 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_431
timestamp 18001
transform 1 0 40756 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_445
timestamp 18001
transform 1 0 42044 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp 18001
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 18001
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_48
timestamp 18001
transform 1 0 5520 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_60
timestamp 18001
transform 1 0 6624 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 18001
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_93
timestamp 1636986456
transform 1 0 9660 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_105
timestamp 18001
transform 1 0 10764 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_113
timestamp 18001
transform 1 0 11500 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_137
timestamp 18001
transform 1 0 13708 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_150
timestamp 1636986456
transform 1 0 14904 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_162
timestamp 1636986456
transform 1 0 16008 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_174
timestamp 1636986456
transform 1 0 17112 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_186
timestamp 18001
transform 1 0 18216 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_194
timestamp 18001
transform 1 0 18952 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_205
timestamp 1636986456
transform 1 0 19964 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_217
timestamp 18001
transform 1 0 21068 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_234
timestamp 18001
transform 1 0 22632 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_242
timestamp 18001
transform 1 0 23368 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 18001
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_261
timestamp 18001
transform 1 0 25116 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_274
timestamp 1636986456
transform 1 0 26312 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_286
timestamp 1636986456
transform 1 0 27416 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 18001
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_337
timestamp 18001
transform 1 0 32108 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 18001
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_380
timestamp 1636986456
transform 1 0 36064 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_392
timestamp 18001
transform 1 0 37168 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_410
timestamp 18001
transform 1 0 38824 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_418
timestamp 18001
transform 1 0 39560 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_421
timestamp 18001
transform 1 0 39836 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_427
timestamp 18001
transform 1 0 40388 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_445
timestamp 18001
transform 1 0 42044 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1636986456
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_15
timestamp 18001
transform 1 0 2484 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_23
timestamp 18001
transform 1 0 3220 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_28
timestamp 1636986456
transform 1 0 3680 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_40
timestamp 1636986456
transform 1 0 4784 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 18001
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1636986456
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1636986456
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1636986456
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1636986456
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 18001
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 18001
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1636986456
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_125
timestamp 18001
transform 1 0 12604 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_159
timestamp 18001
transform 1 0 15732 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 18001
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1636986456
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_193
timestamp 18001
transform 1 0 18860 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_202
timestamp 1636986456
transform 1 0 19688 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_219
timestamp 18001
transform 1 0 21252 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 18001
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1636986456
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_237
timestamp 18001
transform 1 0 22908 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_243
timestamp 18001
transform 1 0 23460 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_252
timestamp 18001
transform 1 0 24288 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_260
timestamp 18001
transform 1 0 25024 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_265
timestamp 1636986456
transform 1 0 25484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_277
timestamp 18001
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 18001
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_291
timestamp 1636986456
transform 1 0 27876 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_303
timestamp 1636986456
transform 1 0 28980 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_315
timestamp 18001
transform 1 0 30084 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_326
timestamp 18001
transform 1 0 31096 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_333
timestamp 18001
transform 1 0 31740 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_348
timestamp 1636986456
transform 1 0 33120 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_360
timestamp 18001
transform 1 0 34224 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_368
timestamp 18001
transform 1 0 34960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_382
timestamp 18001
transform 1 0 36248 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 18001
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_402
timestamp 18001
transform 1 0 38088 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_414
timestamp 18001
transform 1 0 39192 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_67_427
timestamp 18001
transform 1 0 40388 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1636986456
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1636986456
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 18001
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1636986456
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1636986456
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1636986456
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1636986456
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 18001
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 18001
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1636986456
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1636986456
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1636986456
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_121
timestamp 18001
transform 1 0 12236 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_129
timestamp 18001
transform 1 0 12972 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_141
timestamp 18001
transform 1 0 14076 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_187
timestamp 18001
transform 1 0 18308 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_212
timestamp 18001
transform 1 0 20608 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_234
timestamp 18001
transform 1 0 22632 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_267
timestamp 18001
transform 1 0 25668 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_273
timestamp 18001
transform 1 0 26220 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_302
timestamp 18001
transform 1 0 28888 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_309
timestamp 18001
transform 1 0 29532 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_317
timestamp 18001
transform 1 0 30268 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_344
timestamp 1636986456
transform 1 0 32752 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_356
timestamp 18001
transform 1 0 33856 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_373
timestamp 18001
transform 1 0 35420 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_402
timestamp 18001
transform 1 0 38088 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_412
timestamp 18001
transform 1 0 39008 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_421
timestamp 18001
transform 1 0 39836 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1636986456
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1636986456
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1636986456
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1636986456
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 18001
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 18001
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1636986456
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1636986456
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1636986456
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1636986456
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 18001
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 18001
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1636986456
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_125
timestamp 18001
transform 1 0 12604 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_131
timestamp 18001
transform 1 0 13156 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 18001
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_169
timestamp 18001
transform 1 0 16652 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_179
timestamp 1636986456
transform 1 0 17572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_191
timestamp 18001
transform 1 0 18676 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_200
timestamp 1636986456
transform 1 0 19504 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_212
timestamp 18001
transform 1 0 20608 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_218
timestamp 18001
transform 1 0 21160 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1636986456
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_244
timestamp 1636986456
transform 1 0 23552 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_256
timestamp 18001
transform 1 0 24656 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_265
timestamp 1636986456
transform 1 0 25484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_277
timestamp 18001
transform 1 0 26588 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_288
timestamp 1636986456
transform 1 0 27600 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_300
timestamp 1636986456
transform 1 0 28704 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_312
timestamp 18001
transform 1 0 29808 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_320
timestamp 18001
transform 1 0 30544 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_324
timestamp 1636986456
transform 1 0 30912 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_344
timestamp 18001
transform 1 0 32752 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_352
timestamp 18001
transform 1 0 33488 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_382
timestamp 18001
transform 1 0 36248 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_388
timestamp 18001
transform 1 0 36800 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_420
timestamp 18001
transform 1 0 39744 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_443
timestamp 18001
transform 1 0 41860 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1636986456
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1636986456
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1636986456
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1636986456
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1636986456
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1636986456
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 18001
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 18001
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1636986456
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1636986456
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1636986456
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1636986456
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 18001
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 18001
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1636986456
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1636986456
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_165
timestamp 18001
transform 1 0 16284 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_171
timestamp 18001
transform 1 0 16836 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 18001
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_197
timestamp 18001
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_205
timestamp 18001
transform 1 0 19964 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_231
timestamp 1636986456
transform 1 0 22356 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_243
timestamp 18001
transform 1 0 23460 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 18001
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 18001
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_261
timestamp 18001
transform 1 0 25116 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_275
timestamp 18001
transform 1 0 26404 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_283
timestamp 18001
transform 1 0 27140 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 18001
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 18001
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_309
timestamp 18001
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_317
timestamp 18001
transform 1 0 30268 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_327
timestamp 1636986456
transform 1 0 31188 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_339
timestamp 18001
transform 1 0 32292 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_349
timestamp 1636986456
transform 1 0 33212 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_361
timestamp 18001
transform 1 0 34316 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_365
timestamp 18001
transform 1 0 34684 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_380
timestamp 1636986456
transform 1 0 36064 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_392
timestamp 18001
transform 1 0 37168 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 18001
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 18001
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1636986456
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_433
timestamp 18001
transform 1 0 40940 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636986456
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636986456
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1636986456
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1636986456
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 18001
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 18001
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1636986456
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1636986456
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1636986456
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1636986456
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 18001
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 18001
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1636986456
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1636986456
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1636986456
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_149
timestamp 18001
transform 1 0 14812 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_166
timestamp 18001
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_182
timestamp 18001
transform 1 0 17848 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_207
timestamp 1636986456
transform 1 0 20148 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_219
timestamp 18001
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 18001
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_225
timestamp 18001
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_233
timestamp 18001
transform 1 0 22540 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 18001
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_277
timestamp 18001
transform 1 0 26588 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_323
timestamp 18001
transform 1 0 30820 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1636986456
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_373
timestamp 18001
transform 1 0 35420 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_381
timestamp 18001
transform 1 0 36156 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_389
timestamp 18001
transform 1 0 36892 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_393
timestamp 18001
transform 1 0 37260 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_401
timestamp 18001
transform 1 0 37996 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_415
timestamp 1636986456
transform 1 0 39284 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_427
timestamp 1636986456
transform 1 0 40388 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_439
timestamp 18001
transform 1 0 41492 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1636986456
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1636986456
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 18001
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1636986456
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1636986456
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1636986456
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1636986456
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 18001
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 18001
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1636986456
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1636986456
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1636986456
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1636986456
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 18001
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 18001
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_141
timestamp 18001
transform 1 0 14076 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_169
timestamp 18001
transform 1 0 16652 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_173
timestamp 18001
transform 1 0 17020 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 18001
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_197
timestamp 18001
transform 1 0 19228 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_219
timestamp 18001
transform 1 0 21252 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_232
timestamp 18001
transform 1 0 22448 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_240
timestamp 18001
transform 1 0 23184 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 18001
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1636986456
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_265
timestamp 18001
transform 1 0 25484 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_274
timestamp 18001
transform 1 0 26312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_278
timestamp 18001
transform 1 0 26680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_305
timestamp 18001
transform 1 0 29164 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_309
timestamp 18001
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_317
timestamp 18001
transform 1 0 30268 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_72_338
timestamp 18001
transform 1 0 32200 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_353
timestamp 18001
transform 1 0 33580 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 18001
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_390
timestamp 1636986456
transform 1 0 36984 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_402
timestamp 1636986456
transform 1 0 38088 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_414
timestamp 18001
transform 1 0 39192 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1636986456
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1636986456
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_445
timestamp 18001
transform 1 0 42044 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1636986456
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1636986456
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1636986456
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1636986456
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 18001
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 18001
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1636986456
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1636986456
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1636986456
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1636986456
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 18001
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 18001
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1636986456
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1636986456
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1636986456
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1636986456
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_161
timestamp 18001
transform 1 0 15916 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_169
timestamp 18001
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_178
timestamp 18001
transform 1 0 17480 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_202
timestamp 18001
transform 1 0 19688 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_233
timestamp 18001
transform 1 0 22540 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_254
timestamp 1636986456
transform 1 0 24472 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_266
timestamp 1636986456
transform 1 0 25576 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 18001
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_289
timestamp 18001
transform 1 0 27692 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_310
timestamp 18001
transform 1 0 29624 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_341
timestamp 1636986456
transform 1 0 32476 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_353
timestamp 1636986456
transform 1 0 33580 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_365
timestamp 18001
transform 1 0 34684 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_371
timestamp 18001
transform 1 0 35236 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_413
timestamp 1636986456
transform 1 0 39100 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_425
timestamp 1636986456
transform 1 0 40204 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_437
timestamp 18001
transform 1 0 41308 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_445
timestamp 18001
transform 1 0 42044 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636986456
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636986456
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 18001
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1636986456
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1636986456
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1636986456
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1636986456
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 18001
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 18001
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1636986456
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1636986456
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1636986456
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1636986456
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 18001
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 18001
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1636986456
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_153
timestamp 18001
transform 1 0 15180 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_157
timestamp 18001
transform 1 0 15548 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_178
timestamp 18001
transform 1 0 17480 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_186
timestamp 18001
transform 1 0 18216 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 18001
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_204
timestamp 1636986456
transform 1 0 19872 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_236
timestamp 18001
transform 1 0 22816 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_244
timestamp 18001
transform 1 0 23552 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_273
timestamp 18001
transform 1 0 26220 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_294
timestamp 18001
transform 1 0 28152 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_304
timestamp 18001
transform 1 0 29072 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1636986456
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1636986456
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1636986456
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1636986456
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 18001
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 18001
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_365
timestamp 18001
transform 1 0 34684 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_369
timestamp 18001
transform 1 0 35052 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_390
timestamp 1636986456
transform 1 0 36984 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_402
timestamp 1636986456
transform 1 0 38088 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_414
timestamp 18001
transform 1 0 39192 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1636986456
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1636986456
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_445
timestamp 18001
transform 1 0 42044 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1636986456
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1636986456
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_27
timestamp 18001
transform 1 0 3588 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_29
timestamp 1636986456
transform 1 0 3772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_41
timestamp 1636986456
transform 1 0 4876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 18001
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1636986456
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1636986456
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_81
timestamp 18001
transform 1 0 8556 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_85
timestamp 1636986456
transform 1 0 8924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_97
timestamp 1636986456
transform 1 0 10028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_109
timestamp 18001
transform 1 0 11132 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1636986456
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1636986456
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_137
timestamp 18001
transform 1 0 13708 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_141
timestamp 1636986456
transform 1 0 14076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_153
timestamp 1636986456
transform 1 0 15180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_165
timestamp 18001
transform 1 0 16284 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_169
timestamp 18001
transform 1 0 16652 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_177
timestamp 18001
transform 1 0 17388 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_182
timestamp 1636986456
transform 1 0 17848 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_194
timestamp 18001
transform 1 0 18952 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_197
timestamp 18001
transform 1 0 19228 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_203
timestamp 18001
transform 1 0 19780 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_75_210
timestamp 18001
transform 1 0 20424 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 18001
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 18001
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_225
timestamp 18001
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_233
timestamp 18001
transform 1 0 22540 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_238
timestamp 18001
transform 1 0 23000 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_245
timestamp 18001
transform 1 0 23644 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_251
timestamp 18001
transform 1 0 24196 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_260
timestamp 18001
transform 1 0 25024 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_266
timestamp 1636986456
transform 1 0 25576 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 18001
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1636986456
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_293
timestamp 18001
transform 1 0 28060 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_299
timestamp 18001
transform 1 0 28612 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_303
timestamp 18001
transform 1 0 28980 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_309
timestamp 1636986456
transform 1 0 29532 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_321
timestamp 1636986456
transform 1 0 30636 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_333
timestamp 18001
transform 1 0 31740 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1636986456
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1636986456
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_361
timestamp 18001
transform 1 0 34316 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_365
timestamp 1636986456
transform 1 0 34684 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_377
timestamp 1636986456
transform 1 0 35788 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_389
timestamp 18001
transform 1 0 36892 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1636986456
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1636986456
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_417
timestamp 18001
transform 1 0 39468 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_421
timestamp 1636986456
transform 1 0 39836 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_433
timestamp 1636986456
transform 1 0 40940 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_445
timestamp 18001
transform 1 0 42044 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform -1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform -1 0 5060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform -1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform 1 0 40756 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 18001
transform -1 0 13984 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 18001
transform 1 0 14536 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 18001
transform 1 0 2208 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 18001
transform -1 0 26404 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 18001
transform -1 0 3772 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 18001
transform -1 0 10488 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 18001
transform -1 0 19688 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 18001
transform -1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 18001
transform -1 0 28888 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 18001
transform -1 0 32476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 18001
transform -1 0 21712 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 18001
transform -1 0 23736 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 18001
transform -1 0 24380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 18001
transform -1 0 39284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 18001
transform -1 0 20424 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 18001
transform 1 0 8832 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 18001
transform -1 0 41032 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 18001
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 18001
transform -1 0 34132 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 18001
transform -1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 18001
transform 1 0 10764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 18001
transform -1 0 9384 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 18001
transform -1 0 27140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 18001
transform -1 0 32660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 18001
transform -1 0 29256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 18001
transform -1 0 13524 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 18001
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 18001
transform -1 0 42228 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 18001
transform 1 0 16744 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 18001
transform -1 0 39744 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 18001
transform -1 0 34408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 18001
transform -1 0 35604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 18001
transform -1 0 25024 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 18001
transform -1 0 15272 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 18001
transform -1 0 19136 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 18001
transform 1 0 27140 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 18001
transform -1 0 30820 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 18001
transform 1 0 39008 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 18001
transform -1 0 17848 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 18001
transform -1 0 26772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 18001
transform -1 0 35420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 18001
transform -1 0 40572 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 18001
transform -1 0 39560 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 18001
transform -1 0 34684 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 18001
transform -1 0 19872 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 18001
transform 1 0 19320 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 18001
transform -1 0 23368 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 18001
transform -1 0 17204 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 18001
transform 1 0 20332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 18001
transform -1 0 31648 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 18001
transform -1 0 37260 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 18001
transform -1 0 12972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 18001
transform -1 0 16560 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 18001
transform -1 0 36984 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 18001
transform -1 0 25116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 18001
transform 1 0 32384 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 18001
transform -1 0 21528 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 18001
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 18001
transform -1 0 29072 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 18001
transform -1 0 39560 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 18001
transform -1 0 29532 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 18001
transform -1 0 26864 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 18001
transform 1 0 15916 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 18001
transform -1 0 24932 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 18001
transform -1 0 31372 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 18001
transform -1 0 26496 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 18001
transform 1 0 15732 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 18001
transform -1 0 36984 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 18001
transform -1 0 42044 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 18001
transform -1 0 42228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 18001
transform -1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 18001
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 18001
transform 1 0 14720 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 18001
transform -1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 18001
transform 1 0 32108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 18001
transform -1 0 32936 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 18001
transform -1 0 18584 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 18001
transform -1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 18001
transform -1 0 42228 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 18001
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 18001
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 18001
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 18001
transform -1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 18001
transform 1 0 29900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 18001
transform -1 0 39192 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 18001
transform -1 0 40296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 18001
transform -1 0 14168 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 18001
transform -1 0 30544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 18001
transform 1 0 29440 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 18001
transform -1 0 34960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 18001
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 18001
transform -1 0 33304 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 18001
transform -1 0 21712 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 18001
transform 1 0 24564 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 18001
transform -1 0 36984 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 18001
transform 1 0 36984 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 18001
transform 1 0 36432 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 18001
transform -1 0 39652 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 18001
transform -1 0 40940 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 18001
transform -1 0 12972 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 18001
transform -1 0 34040 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 18001
transform -1 0 11040 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 18001
transform -1 0 42044 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 18001
transform -1 0 39192 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 18001
transform -1 0 30268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 18001
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 18001
transform -1 0 20516 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 18001
transform -1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 18001
transform 1 0 27508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 18001
transform 1 0 25668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 18001
transform -1 0 40572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 18001
transform -1 0 30544 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 18001
transform -1 0 13892 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 18001
transform 1 0 10580 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 18001
transform 1 0 36064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 18001
transform 1 0 34776 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 18001
transform -1 0 7820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 18001
transform -1 0 10304 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 18001
transform -1 0 11408 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 18001
transform 1 0 10396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 18001
transform -1 0 26864 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 18001
transform -1 0 42228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 18001
transform -1 0 41768 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 18001
transform 1 0 35328 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 18001
transform -1 0 30912 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 18001
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 18001
transform -1 0 42228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 18001
transform -1 0 41952 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 18001
transform -1 0 41492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 18001
transform -1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 18001
transform 1 0 9936 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 18001
transform -1 0 29992 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 18001
transform -1 0 35420 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 18001
transform -1 0 39468 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 18001
transform -1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 18001
transform -1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 18001
transform -1 0 23276 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 18001
transform 1 0 34684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 18001
transform 1 0 17480 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 18001
transform 1 0 19320 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 18001
transform -1 0 33212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 18001
transform -1 0 26496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 18001
transform -1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 18001
transform -1 0 42228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 18001
transform -1 0 41768 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 18001
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 18001
transform -1 0 12236 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 18001
transform -1 0 25668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 18001
transform -1 0 27140 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 18001
transform -1 0 42228 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 18001
transform 1 0 39376 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 18001
transform -1 0 37168 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 18001
transform 1 0 34776 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 18001
transform -1 0 35236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 18001
transform -1 0 37076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 18001
transform -1 0 39192 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 18001
transform 1 0 37536 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 18001
transform -1 0 15364 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 18001
transform -1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 18001
transform -1 0 25852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 18001
transform -1 0 39468 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 18001
transform -1 0 32936 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 18001
transform -1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 18001
transform -1 0 26312 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 18001
transform -1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 18001
transform -1 0 18584 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 18001
transform -1 0 35052 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 18001
transform -1 0 21528 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 18001
transform -1 0 28796 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 18001
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 18001
transform -1 0 37076 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 18001
transform -1 0 35604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 18001
transform -1 0 30360 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 18001
transform -1 0 19596 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 18001
transform -1 0 37536 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 18001
transform -1 0 37168 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 18001
transform 1 0 26864 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 18001
transform 1 0 17940 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 18001
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 18001
transform -1 0 32108 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 18001
transform -1 0 30268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 18001
transform -1 0 17388 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 18001
transform -1 0 25116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 18001
transform -1 0 26680 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 18001
transform -1 0 22540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 18001
transform -1 0 21436 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 18001
transform -1 0 11408 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 18001
transform 1 0 20976 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 18001
transform 1 0 27600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 18001
transform -1 0 30268 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 18001
transform -1 0 25852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 18001
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 18001
transform -1 0 37076 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 18001
transform -1 0 39468 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 18001
transform -1 0 33488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 18001
transform 1 0 31096 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 18001
transform -1 0 32844 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 18001
transform -1 0 34132 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 18001
transform -1 0 22540 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 18001
transform -1 0 10028 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 18001
transform -1 0 26496 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 18001
transform -1 0 20516 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 18001
transform -1 0 24288 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 18001
transform 1 0 12696 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 18001
transform -1 0 27876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 18001
transform -1 0 29808 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 18001
transform -1 0 11224 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 18001
transform -1 0 10304 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 18001
transform -1 0 13432 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 18001
transform -1 0 8648 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 18001
transform -1 0 35604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 18001
transform 1 0 12788 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 18001
transform -1 0 41308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 18001
transform -1 0 25760 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 18001
transform -1 0 29256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 18001
transform -1 0 28336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 18001
transform -1 0 42228 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 18001
transform 1 0 30820 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 18001
transform -1 0 29256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 18001
transform -1 0 42044 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 18001
transform 1 0 32292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 18001
transform -1 0 25208 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 18001
transform -1 0 3772 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 18001
transform -1 0 24380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 18001
transform -1 0 23368 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 18001
transform -1 0 37168 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 18001
transform -1 0 38088 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 18001
transform -1 0 8556 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 18001
transform -1 0 13892 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 18001
transform -1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 18001
transform -1 0 25576 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 18001
transform -1 0 21620 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 18001
transform -1 0 20516 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 18001
transform -1 0 35420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 18001
transform 1 0 17940 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 18001
transform -1 0 34132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 18001
transform -1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 18001
transform -1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 18001
transform -1 0 34592 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 18001
transform 1 0 32108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 18001
transform -1 0 5704 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 18001
transform -1 0 16560 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 18001
transform 1 0 4232 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 18001
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 18001
transform -1 0 20240 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 18001
transform -1 0 15732 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 18001
transform -1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 18001
transform -1 0 37904 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 18001
transform -1 0 10028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 18001
transform -1 0 32752 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 18001
transform -1 0 3680 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 18001
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 18001
transform -1 0 16376 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 18001
transform -1 0 11408 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 18001
transform 1 0 14352 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 18001
transform -1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 18001
transform -1 0 18584 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 18001
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 18001
transform -1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 18001
transform -1 0 10948 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 18001
transform 1 0 6900 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 18001
transform -1 0 17388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 18001
transform 1 0 7268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 18001
transform -1 0 4508 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 18001
transform -1 0 13984 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 18001
transform -1 0 21068 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 18001
transform -1 0 15824 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 18001
transform -1 0 7544 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 18001
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 18001
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 18001
transform -1 0 26680 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 18001
transform -1 0 9660 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 18001
transform -1 0 35420 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 18001
transform 1 0 5520 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 18001
transform -1 0 9844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 18001
transform -1 0 17388 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 18001
transform -1 0 22540 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 18001
transform 1 0 37260 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 18001
transform -1 0 33856 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 18001
transform 1 0 13340 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 18001
transform -1 0 16008 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 18001
transform -1 0 14996 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 18001
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 18001
transform -1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 18001
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 18001
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 18001
transform -1 0 42228 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 18001
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 18001
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 18001
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 18001
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 18001
transform -1 0 21068 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 18001
transform 1 0 17480 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 18001
transform 1 0 41676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 18001
transform 1 0 41860 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 18001
transform -1 0 40848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 18001
transform 1 0 41860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 18001
transform -1 0 40388 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 18001
transform 1 0 20056 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 18001
transform -1 0 19780 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 18001
transform 1 0 22632 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 18001
transform -1 0 23644 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 18001
transform -1 0 25576 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 18001
transform 1 0 41860 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 18001
transform -1 0 29440 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 18001
transform 1 0 41308 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 18001
transform 1 0 41492 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 18001
transform 1 0 41860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 18001
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 18001
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 18001
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 18001
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_76
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 42504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_77
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 42504 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_78
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 42504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_79
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 42504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_80
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 42504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_81
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 42504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_82
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 42504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_83
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 42504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_84
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 42504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_85
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 42504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_86
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 42504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_87
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 42504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_88
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 42504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_89
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 42504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_90
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 42504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_91
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 42504 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_92
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 42504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_93
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 42504 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_94
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 42504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_95
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 42504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_96
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 42504 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_97
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 42504 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_98
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 42504 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_99
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 42504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_100
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 42504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_101
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 42504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_102
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 42504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_103
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 42504 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_104
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 42504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_105
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 42504 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_106
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 42504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_107
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 42504 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_108
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 42504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_109
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 42504 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_110
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 42504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_111
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 42504 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_112
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 42504 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_113
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 42504 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_114
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 42504 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_115
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 42504 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_116
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 42504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_117
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 42504 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_118
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 42504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_119
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 42504 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_120
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 42504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_121
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 42504 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_122
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 42504 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_123
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 42504 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_124
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 42504 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_125
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 42504 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_126
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 42504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_127
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 42504 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_128
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 42504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_129
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 42504 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_130
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 42504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_131
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 42504 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_132
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 42504 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_133
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 42504 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_134
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 42504 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_135
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 42504 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_136
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 42504 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_137
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 42504 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_138
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 42504 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_139
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 42504 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_140
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 42504 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_141
timestamp 18001
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 18001
transform -1 0 42504 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_142
timestamp 18001
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 18001
transform -1 0 42504 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_143
timestamp 18001
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 18001
transform -1 0 42504 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_144
timestamp 18001
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 18001
transform -1 0 42504 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_145
timestamp 18001
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 18001
transform -1 0 42504 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_146
timestamp 18001
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 18001
transform -1 0 42504 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_147
timestamp 18001
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 18001
transform -1 0 42504 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_148
timestamp 18001
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 18001
transform -1 0 42504 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_149
timestamp 18001
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 18001
transform -1 0 42504 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_150
timestamp 18001
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 18001
transform -1 0 42504 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_151
timestamp 18001
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 18001
transform -1 0 42504 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_152
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_153
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_154
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_155
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_159
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_160
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_161
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_162
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_163
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_164
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_165
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_166
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_167
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_168
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_169
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_170
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_171
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_172
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_173
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_174
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_175
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_176
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_177
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_178
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_179
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_180
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_181
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_182
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_183
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_184
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_185
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_186
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_187
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_188
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_189
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_190
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_191
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_192
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_193
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_194
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_195
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_196
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_197
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_198
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_199
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_200
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_201
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_202
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_203
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_204
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_205
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_206
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_207
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_208
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_209
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_210
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_211
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_212
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_213
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_214
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_215
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_216
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_217
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_218
timestamp 18001
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_219
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_220
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_221
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_222
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_223
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_224
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_225
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_226
timestamp 18001
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_227
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_228
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_229
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_230
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_231
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_232
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_233
timestamp 18001
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_234
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_235
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_236
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_237
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_238
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_239
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_240
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_241
timestamp 18001
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_242
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_243
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_244
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_245
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_246
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_247
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_248
timestamp 18001
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_249
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_250
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_251
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_252
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_253
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_254
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_255
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_256
timestamp 18001
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_257
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_258
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_259
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_260
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_261
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_262
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_263
timestamp 18001
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_264
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_265
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_266
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_267
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_268
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_269
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_270
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_271
timestamp 18001
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_272
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_273
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_274
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_275
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_276
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_277
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_278
timestamp 18001
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_279
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_280
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_281
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_282
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_283
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_284
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_285
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_286
timestamp 18001
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_287
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_288
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_289
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_290
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_291
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_292
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_293
timestamp 18001
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_294
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_295
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_296
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_297
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_298
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_299
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_300
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_301
timestamp 18001
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_302
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_303
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_304
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_305
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_306
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_307
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_308
timestamp 18001
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_309
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_310
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_311
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_312
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_313
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_314
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_315
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_316
timestamp 18001
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_317
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_318
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_319
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_320
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_321
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_322
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_323
timestamp 18001
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_324
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_325
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_326
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_327
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_328
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_329
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_330
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_331
timestamp 18001
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_332
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_333
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_334
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_335
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_336
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_337
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_338
timestamp 18001
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_339
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_340
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_341
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_342
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_343
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_344
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_345
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_346
timestamp 18001
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_347
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_348
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_349
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_350
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_351
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_352
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_353
timestamp 18001
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_354
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_355
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_356
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_357
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_358
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_359
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_360
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_361
timestamp 18001
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_362
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_363
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_364
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_365
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_366
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_367
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_368
timestamp 18001
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_369
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_370
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_371
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_372
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_373
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_374
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_375
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_376
timestamp 18001
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_377
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_378
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_379
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_380
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_381
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_382
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_383
timestamp 18001
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_384
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_385
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_386
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_387
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_388
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_389
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_390
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_391
timestamp 18001
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_392
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_393
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_394
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_395
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_396
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_397
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_398
timestamp 18001
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_399
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_400
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_401
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_402
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_403
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_404
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_405
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_406
timestamp 18001
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_407
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_408
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_409
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_410
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_411
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_412
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_413
timestamp 18001
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_414
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_415
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_416
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_417
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_418
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_419
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_420
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_421
timestamp 18001
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_422
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_423
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_424
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_425
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_426
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_427
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_428
timestamp 18001
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_429
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_430
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_431
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_432
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_433
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_434
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_435
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_436
timestamp 18001
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_437
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_438
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_439
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_440
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_441
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_442
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_443
timestamp 18001
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_444
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_445
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_446
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_447
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_448
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_449
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_450
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_451
timestamp 18001
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_452
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_453
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_454
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_455
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_456
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_457
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_458
timestamp 18001
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_459
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_460
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_461
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_462
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_463
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_464
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_465
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_466
timestamp 18001
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_467
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_468
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_469
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_470
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_471
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_472
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_473
timestamp 18001
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_474
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_475
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_476
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_477
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_478
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_479
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_480
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_481
timestamp 18001
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_482
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_483
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_484
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_485
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_486
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_487
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_488
timestamp 18001
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_489
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_490
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_491
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_492
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_493
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_494
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_495
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_496
timestamp 18001
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_497
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_498
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_499
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_500
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_501
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_502
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_503
timestamp 18001
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_504
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_505
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_506
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_507
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_508
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_509
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_510
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_511
timestamp 18001
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_512
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_513
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_514
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_515
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_516
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_517
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_518
timestamp 18001
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_519
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_520
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_521
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_522
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_523
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_524
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_525
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_526
timestamp 18001
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_527
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_528
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_529
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_530
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_531
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_532
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_533
timestamp 18001
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_534
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_535
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_536
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_537
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_538
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_539
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_540
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_541
timestamp 18001
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_542
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_543
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_544
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_545
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_546
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_547
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_548
timestamp 18001
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_549
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_550
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_551
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_552
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_553
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_554
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_555
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_556
timestamp 18001
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_557
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_558
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_559
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_560
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_561
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_562
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_563
timestamp 18001
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_564
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_565
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_566
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_567
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_568
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_569
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_570
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_571
timestamp 18001
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_572
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_573
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_574
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_575
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_576
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_577
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_578
timestamp 18001
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_579
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_580
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_581
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_582
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_583
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_584
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_585
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_586
timestamp 18001
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_587
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_588
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_589
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_590
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_591
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_592
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_593
timestamp 18001
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_594
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_595
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_596
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_597
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_598
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_599
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_600
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_601
timestamp 18001
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_602
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_603
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_604
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_605
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_606
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_607
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_608
timestamp 18001
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_609
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_610
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_611
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_612
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_613
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_614
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_615
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_616
timestamp 18001
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_617
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_618
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_619
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_620
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_621
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_622
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_623
timestamp 18001
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_624
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_625
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_626
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_627
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_628
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_629
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_630
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_631
timestamp 18001
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_632
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_633
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_634
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_635
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_636
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_637
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_638
timestamp 18001
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_639
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_640
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_641
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_642
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_643
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_644
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_645
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_646
timestamp 18001
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_647
timestamp 18001
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_648
timestamp 18001
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_649
timestamp 18001
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_650
timestamp 18001
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_651
timestamp 18001
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_652
timestamp 18001
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_653
timestamp 18001
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_654
timestamp 18001
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_655
timestamp 18001
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_656
timestamp 18001
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_657
timestamp 18001
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_658
timestamp 18001
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_659
timestamp 18001
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_660
timestamp 18001
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_661
timestamp 18001
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_662
timestamp 18001
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_663
timestamp 18001
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_664
timestamp 18001
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_665
timestamp 18001
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_666
timestamp 18001
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_667
timestamp 18001
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_668
timestamp 18001
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_669
timestamp 18001
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_670
timestamp 18001
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_671
timestamp 18001
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_672
timestamp 18001
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_673
timestamp 18001
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_674
timestamp 18001
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_675
timestamp 18001
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_676
timestamp 18001
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_677
timestamp 18001
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_678
timestamp 18001
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_679
timestamp 18001
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_680
timestamp 18001
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_681
timestamp 18001
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_682
timestamp 18001
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_683
timestamp 18001
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_684
timestamp 18001
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_685
timestamp 18001
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_686
timestamp 18001
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_687
timestamp 18001
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_688
timestamp 18001
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_689
timestamp 18001
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_690
timestamp 18001
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_691
timestamp 18001
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_692
timestamp 18001
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_693
timestamp 18001
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_694
timestamp 18001
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_695
timestamp 18001
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_696
timestamp 18001
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_697
timestamp 18001
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_698
timestamp 18001
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_699
timestamp 18001
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_700
timestamp 18001
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_701
timestamp 18001
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_702
timestamp 18001
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_703
timestamp 18001
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_704
timestamp 18001
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_705
timestamp 18001
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_706
timestamp 18001
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_707
timestamp 18001
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_708
timestamp 18001
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_709
timestamp 18001
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_710
timestamp 18001
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_711
timestamp 18001
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_712
timestamp 18001
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_713
timestamp 18001
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_714
timestamp 18001
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_715
timestamp 18001
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_716
timestamp 18001
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_717
timestamp 18001
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_718
timestamp 18001
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_719
timestamp 18001
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_720
timestamp 18001
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_721
timestamp 18001
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_722
timestamp 18001
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_723
timestamp 18001
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_724
timestamp 18001
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_725
timestamp 18001
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_726
timestamp 18001
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_727
timestamp 18001
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_728
timestamp 18001
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_729
timestamp 18001
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_730
timestamp 18001
transform 1 0 24288 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_731
timestamp 18001
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_732
timestamp 18001
transform 1 0 29440 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_733
timestamp 18001
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_734
timestamp 18001
transform 1 0 34592 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_735
timestamp 18001
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_736
timestamp 18001
transform 1 0 39744 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire83
timestamp 18001
transform 1 0 3772 0 1 22848
box -38 -48 314 592
<< labels >>
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 ColOut[0]
port 0 nsew signal output
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 ColOut[1]
port 1 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 ColOut[2]
port 2 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 ColOut[3]
port 3 nsew signal output
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 RowIn[0]
port 4 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 RowIn[1]
port 5 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 RowIn[2]
port 6 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 RowIn[3]
port 7 nsew signal input
flabel metal4 s 4868 2128 5188 43568 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 43568 0 FreeSans 1920 90 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 6006 42552 6326 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal5 s 1056 36642 42552 36962 0 FreeSans 2560 0 0 0 VGND
port 8 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 43568 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal4 s 34928 2128 35248 43568 0 FreeSans 1920 90 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 5346 42552 5666 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal5 s 1056 35982 42552 36302 0 FreeSans 2560 0 0 0 VPWR
port 9 nsew power bidirectional
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 clk
port 10 nsew signal input
flabel metal2 s 20626 44987 20682 45787 0 FreeSans 224 90 0 0 complete
port 11 nsew signal output
flabel metal2 s 17406 44987 17462 45787 0 FreeSans 224 90 0 0 display_output[0]
port 12 nsew signal output
flabel metal3 s 42843 26528 43643 26648 0 FreeSans 480 0 0 0 display_output[10]
port 13 nsew signal output
flabel metal3 s 42843 31288 43643 31408 0 FreeSans 480 0 0 0 display_output[11]
port 14 nsew signal output
flabel metal3 s 42843 24488 43643 24608 0 FreeSans 480 0 0 0 display_output[12]
port 15 nsew signal output
flabel metal3 s 42843 28568 43643 28688 0 FreeSans 480 0 0 0 display_output[13]
port 16 nsew signal output
flabel metal3 s 42843 25168 43643 25288 0 FreeSans 480 0 0 0 display_output[14]
port 17 nsew signal output
flabel metal2 s 19982 44987 20038 45787 0 FreeSans 224 90 0 0 display_output[15]
port 18 nsew signal output
flabel metal2 s 19338 44987 19394 45787 0 FreeSans 224 90 0 0 display_output[1]
port 19 nsew signal output
flabel metal2 s 22558 44987 22614 45787 0 FreeSans 224 90 0 0 display_output[2]
port 20 nsew signal output
flabel metal2 s 23202 44987 23258 45787 0 FreeSans 224 90 0 0 display_output[3]
port 21 nsew signal output
flabel metal2 s 25134 44987 25190 45787 0 FreeSans 224 90 0 0 display_output[4]
port 22 nsew signal output
flabel metal3 s 42843 25848 43643 25968 0 FreeSans 480 0 0 0 display_output[5]
port 23 nsew signal output
flabel metal2 s 28998 44987 29054 45787 0 FreeSans 224 90 0 0 display_output[6]
port 24 nsew signal output
flabel metal3 s 42843 27208 43643 27328 0 FreeSans 480 0 0 0 display_output[7]
port 25 nsew signal output
flabel metal3 s 42843 27888 43643 28008 0 FreeSans 480 0 0 0 display_output[8]
port 26 nsew signal output
flabel metal3 s 42843 29248 43643 29368 0 FreeSans 480 0 0 0 display_output[9]
port 27 nsew signal output
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 input_state_FPGA[0]
port 28 nsew signal output
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 input_state_FPGA[1]
port 29 nsew signal output
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 input_state_FPGA[2]
port 30 nsew signal output
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 key_pressed
port 31 nsew signal output
flabel metal3 s 42843 3408 43643 3528 0 FreeSans 480 0 0 0 nRST
port 32 nsew signal input
rlabel metal1 21804 43520 21804 43520 0 VGND
rlabel metal1 21804 42976 21804 42976 0 VPWR
rlabel metal2 11638 1520 11638 1520 0 ColOut[0]
rlabel metal3 1096 12308 1096 12308 0 ColOut[1]
rlabel metal3 1096 10948 1096 10948 0 ColOut[2]
rlabel metal3 751 11628 751 11628 0 ColOut[3]
rlabel metal3 751 15708 751 15708 0 RowIn[0]
rlabel metal3 1188 15028 1188 15028 0 RowIn[1]
rlabel metal3 751 17068 751 17068 0 RowIn[2]
rlabel metal3 1096 17748 1096 17748 0 RowIn[3]
rlabel metal2 9890 35428 9890 35428 0 _0000_
rlabel metal2 10994 34816 10994 34816 0 _0001_
rlabel metal1 15548 13294 15548 13294 0 _0002_
rlabel metal1 17020 12954 17020 12954 0 _0003_
rlabel metal1 30222 12274 30222 12274 0 _0004_
rlabel metal2 9890 36380 9890 36380 0 _0005_
rlabel metal1 28796 13498 28796 13498 0 _0006_
rlabel metal1 27002 14518 27002 14518 0 _0007_
rlabel metal2 5566 28322 5566 28322 0 _0008_
rlabel metal1 7682 34476 7682 34476 0 _0009_
rlabel metal1 8234 33558 8234 33558 0 _0010_
rlabel metal1 7406 31450 7406 31450 0 _0011_
rlabel metal2 4738 32147 4738 32147 0 _0012_
rlabel metal1 6808 29818 6808 29818 0 _0013_
rlabel metal1 1978 32776 1978 32776 0 _0014_
rlabel metal2 2162 32980 2162 32980 0 _0015_
rlabel metal2 1702 30872 1702 30872 0 _0016_
rlabel metal1 2162 28730 2162 28730 0 _0017_
rlabel metal1 7084 36346 7084 36346 0 _0018_
rlabel metal2 7038 38114 7038 38114 0 _0019_
rlabel metal1 5743 37434 5743 37434 0 _0020_
rlabel metal1 4462 36890 4462 36890 0 _0021_
rlabel metal1 2162 37978 2162 37978 0 _0022_
rlabel metal1 2116 36890 2116 36890 0 _0023_
rlabel metal2 2898 35802 2898 35802 0 _0024_
rlabel metal2 2162 35292 2162 35292 0 _0025_
rlabel metal2 5290 34544 5290 34544 0 _0026_
rlabel metal1 4554 21386 4554 21386 0 _0027_
rlabel metal1 4876 23154 4876 23154 0 _0028_
rlabel metal1 5704 20910 5704 20910 0 _0029_
rlabel metal2 3358 20604 3358 20604 0 _0030_
rlabel metal1 6072 26010 6072 26010 0 _0031_
rlabel metal1 6716 18938 6716 18938 0 _0032_
rlabel metal1 6568 17170 6568 17170 0 _0033_
rlabel metal1 7482 16490 7482 16490 0 _0034_
rlabel metal1 7482 17578 7482 17578 0 _0035_
rlabel metal2 9706 19108 9706 19108 0 _0036_
rlabel metal1 8908 19754 8908 19754 0 _0037_
rlabel metal1 11561 18326 11561 18326 0 _0038_
rlabel metal1 10800 19822 10800 19822 0 _0039_
rlabel metal1 11576 20502 11576 20502 0 _0040_
rlabel metal2 13938 19482 13938 19482 0 _0041_
rlabel metal1 13662 18190 13662 18190 0 _0042_
rlabel metal1 14735 17238 14735 17238 0 _0043_
rlabel metal1 14643 16150 14643 16150 0 _0044_
rlabel via1 13933 14994 13933 14994 0 _0045_
rlabel metal1 11576 16150 11576 16150 0 _0046_
rlabel metal1 11530 15062 11530 15062 0 _0047_
rlabel metal2 11546 12988 11546 12988 0 _0048_
rlabel via1 13666 13294 13666 13294 0 _0049_
rlabel metal1 14444 13158 14444 13158 0 _0050_
rlabel metal1 14260 11254 14260 11254 0 _0051_
rlabel metal1 6440 24922 6440 24922 0 _0052_
rlabel metal1 9660 24582 9660 24582 0 _0053_
rlabel metal1 8372 26010 8372 26010 0 _0054_
rlabel metal1 9046 25194 9046 25194 0 _0055_
rlabel metal1 8786 21896 8786 21896 0 _0056_
rlabel metal1 9874 22678 9874 22678 0 _0057_
rlabel metal1 9844 23290 9844 23290 0 _0058_
rlabel metal2 9614 23970 9614 23970 0 _0059_
rlabel metal2 20378 8670 20378 8670 0 _0060_
rlabel metal1 20102 10234 20102 10234 0 _0061_
rlabel metal2 20930 10863 20930 10863 0 _0062_
rlabel metal1 21758 7514 21758 7514 0 _0063_
rlabel metal2 25438 7854 25438 7854 0 _0064_
rlabel metal1 26689 10234 26689 10234 0 _0065_
rlabel metal1 28980 7922 28980 7922 0 _0066_
rlabel metal2 28934 10030 28934 10030 0 _0067_
rlabel metal2 29486 8636 29486 8636 0 _0068_
rlabel metal2 32890 8772 32890 8772 0 _0069_
rlabel metal1 33994 9418 33994 9418 0 _0070_
rlabel metal2 34730 8126 34730 8126 0 _0071_
rlabel metal1 37306 7310 37306 7310 0 _0072_
rlabel metal2 39422 10064 39422 10064 0 _0073_
rlabel metal1 39836 10778 39836 10778 0 _0074_
rlabel metal2 2714 14110 2714 14110 0 _0075_
rlabel metal1 2898 12954 2898 12954 0 _0076_
rlabel metal2 2530 11016 2530 11016 0 _0077_
rlabel metal1 3634 13362 3634 13362 0 _0078_
rlabel metal1 5888 13498 5888 13498 0 _0079_
rlabel metal2 4738 13294 4738 13294 0 _0080_
rlabel metal2 6486 14926 6486 14926 0 _0081_
rlabel metal2 6670 15130 6670 15130 0 _0082_
rlabel metal2 10350 14722 10350 14722 0 _0083_
rlabel metal1 9006 13498 9006 13498 0 _0084_
rlabel metal1 9246 12750 9246 12750 0 _0085_
rlabel metal1 11960 11050 11960 11050 0 _0086_
rlabel metal2 9982 11016 9982 11016 0 _0087_
rlabel metal2 9706 9112 9706 9112 0 _0088_
rlabel metal1 11638 9146 11638 9146 0 _0089_
rlabel metal1 11730 10098 11730 10098 0 _0090_
rlabel metal1 3956 9486 3956 9486 0 _0091_
rlabel metal1 2231 7922 2231 7922 0 _0092_
rlabel metal1 5296 6970 5296 6970 0 _0093_
rlabel metal1 1702 8568 1702 8568 0 _0094_
rlabel metal1 2944 4522 2944 4522 0 _0095_
rlabel metal1 4830 4250 4830 4250 0 _0096_
rlabel metal1 4600 3162 4600 3162 0 _0097_
rlabel metal2 3450 3230 3450 3230 0 _0098_
rlabel metal2 7222 7038 7222 7038 0 _0099_
rlabel metal1 6624 5270 6624 5270 0 _0100_
rlabel metal2 7958 3536 7958 3536 0 _0101_
rlabel metal2 9798 3230 9798 3230 0 _0102_
rlabel metal1 10902 3706 10902 3706 0 _0103_
rlabel metal2 9522 6052 9522 6052 0 _0104_
rlabel metal2 10902 5848 10902 5848 0 _0105_
rlabel metal2 10626 6494 10626 6494 0 _0106_
rlabel metal1 15456 31994 15456 31994 0 _0107_
rlabel metal1 17572 32538 17572 32538 0 _0108_
rlabel metal1 21298 31790 21298 31790 0 _0109_
rlabel metal1 22218 27642 22218 27642 0 _0110_
rlabel metal1 23552 31654 23552 31654 0 _0111_
rlabel metal2 25254 28254 25254 28254 0 _0112_
rlabel metal2 26910 30056 26910 30056 0 _0113_
rlabel metal1 28750 28594 28750 28594 0 _0114_
rlabel metal2 30498 28492 30498 28492 0 _0115_
rlabel metal2 31510 29852 31510 29852 0 _0116_
rlabel metal2 37674 28764 37674 28764 0 _0117_
rlabel metal2 37674 30940 37674 30940 0 _0118_
rlabel metal1 35558 28152 35558 28152 0 _0119_
rlabel metal1 34914 30770 34914 30770 0 _0120_
rlabel metal1 33212 28458 33212 28458 0 _0121_
rlabel metal2 17434 26078 17434 26078 0 _0122_
rlabel metal2 16974 23902 16974 23902 0 _0123_
rlabel metal1 20930 26554 20930 26554 0 _0124_
rlabel metal1 21620 26010 21620 26010 0 _0125_
rlabel metal1 24656 23766 24656 23766 0 _0126_
rlabel metal1 24472 26554 24472 26554 0 _0127_
rlabel metal1 26726 24922 26726 24922 0 _0128_
rlabel metal1 27968 24854 27968 24854 0 _0129_
rlabel metal2 29762 25262 29762 25262 0 _0130_
rlabel metal1 31188 25194 31188 25194 0 _0131_
rlabel metal1 38502 24718 38502 24718 0 _0132_
rlabel metal1 37950 25330 37950 25330 0 _0133_
rlabel metal1 35604 23018 35604 23018 0 _0134_
rlabel metal1 34730 24922 34730 24922 0 _0135_
rlabel metal1 32844 25942 32844 25942 0 _0136_
rlabel metal2 8602 26724 8602 26724 0 _0137_
rlabel metal1 19228 7514 19228 7514 0 _0138_
rlabel metal2 18354 10404 18354 10404 0 _0139_
rlabel metal2 21666 11628 21666 11628 0 _0140_
rlabel metal1 22356 7514 22356 7514 0 _0141_
rlabel metal1 22770 7752 22770 7752 0 _0142_
rlabel metal1 23828 9622 23828 9622 0 _0143_
rlabel metal1 26174 7922 26174 7922 0 _0144_
rlabel metal1 27830 9690 27830 9690 0 _0145_
rlabel metal2 28290 7786 28290 7786 0 _0146_
rlabel metal1 30958 8058 30958 8058 0 _0147_
rlabel metal1 32292 10234 32292 10234 0 _0148_
rlabel metal1 33120 7786 33120 7786 0 _0149_
rlabel metal1 35689 8058 35689 8058 0 _0150_
rlabel metal2 37582 9758 37582 9758 0 _0151_
rlabel metal2 37582 11866 37582 11866 0 _0152_
rlabel metal1 13662 36346 13662 36346 0 _0153_
rlabel metal2 14858 21420 14858 21420 0 _0154_
rlabel metal2 15778 15640 15778 15640 0 _0155_
rlabel metal1 17112 18938 17112 18938 0 _0156_
rlabel metal2 20286 19108 20286 19108 0 _0157_
rlabel metal1 21758 20298 21758 20298 0 _0158_
rlabel metal2 22678 14824 22678 14824 0 _0159_
rlabel metal2 25622 19618 25622 19618 0 _0160_
rlabel metal2 26082 15640 26082 15640 0 _0161_
rlabel metal2 28474 20196 28474 20196 0 _0162_
rlabel metal2 32798 14756 32798 14756 0 _0163_
rlabel metal2 31234 20196 31234 20196 0 _0164_
rlabel metal2 36386 19992 36386 19992 0 _0165_
rlabel metal1 39146 20026 39146 20026 0 _0166_
rlabel metal2 38410 16796 38410 16796 0 _0167_
rlabel metal1 38088 13498 38088 13498 0 _0168_
rlabel metal2 33626 15844 33626 15844 0 _0169_
rlabel metal1 15502 21862 15502 21862 0 _0170_
rlabel metal2 19550 15470 19550 15470 0 _0171_
rlabel metal2 18814 17884 18814 17884 0 _0172_
rlabel metal1 21022 14926 21022 14926 0 _0173_
rlabel metal1 23230 18156 23230 18156 0 _0174_
rlabel metal2 24426 14212 24426 14212 0 _0175_
rlabel metal1 26726 16762 26726 16762 0 _0176_
rlabel metal1 30222 15436 30222 15436 0 _0177_
rlabel metal2 29578 18292 29578 18292 0 _0178_
rlabel metal1 31142 15980 31142 15980 0 _0179_
rlabel metal1 33074 18360 33074 18360 0 _0180_
rlabel metal1 37812 19346 37812 19346 0 _0181_
rlabel metal2 41630 18836 41630 18836 0 _0182_
rlabel metal1 41354 15980 41354 15980 0 _0183_
rlabel metal1 41538 14994 41538 14994 0 _0184_
rlabel metal1 34776 14858 34776 14858 0 _0185_
rlabel metal1 16422 14280 16422 14280 0 _0186_
rlabel metal2 15594 16796 15594 16796 0 _0187_
rlabel metal1 17572 21114 17572 21114 0 _0188_
rlabel metal1 20332 20502 20332 20502 0 _0189_
rlabel metal1 23598 21862 23598 21862 0 _0190_
rlabel metal1 23690 20366 23690 20366 0 _0191_
rlabel metal1 26174 20366 26174 20366 0 _0192_
rlabel metal1 27600 20842 27600 20842 0 _0193_
rlabel metal1 29532 22202 29532 22202 0 _0194_
rlabel metal2 30406 21148 30406 21148 0 _0195_
rlabel metal1 32706 20026 32706 20026 0 _0196_
rlabel metal1 37398 21114 37398 21114 0 _0197_
rlabel metal1 40572 21114 40572 21114 0 _0198_
rlabel metal1 41722 20978 41722 20978 0 _0199_
rlabel metal1 39192 14586 39192 14586 0 _0200_
rlabel metal1 34868 17306 34868 17306 0 _0201_
rlabel metal1 19412 14042 19412 14042 0 _0202_
rlabel metal1 17894 12070 17894 12070 0 _0203_
rlabel metal1 20332 12954 20332 12954 0 _0204_
rlabel metal2 21574 13532 21574 13532 0 _0205_
rlabel metal1 23644 12614 23644 12614 0 _0206_
rlabel via1 24695 12410 24695 12410 0 _0207_
rlabel metal1 26128 11186 26128 11186 0 _0208_
rlabel metal1 27968 12410 27968 12410 0 _0209_
rlabel metal1 31372 11798 31372 11798 0 _0210_
rlabel metal2 31050 13090 31050 13090 0 _0211_
rlabel metal2 32890 13566 32890 13566 0 _0212_
rlabel metal1 33396 12886 33396 12886 0 _0213_
rlabel metal1 34868 11322 34868 11322 0 _0214_
rlabel metal1 35512 13974 35512 13974 0 _0215_
rlabel metal1 35972 13362 35972 13362 0 _0216_
rlabel metal2 18814 15640 18814 15640 0 _0217_
rlabel metal2 18722 17510 18722 17510 0 _0218_
rlabel metal1 20884 15402 20884 15402 0 _0219_
rlabel metal2 21850 18802 21850 18802 0 _0220_
rlabel metal2 26450 15436 26450 15436 0 _0221_
rlabel metal2 24886 18088 24886 18088 0 _0222_
rlabel metal1 28697 15878 28697 15878 0 _0223_
rlabel metal2 28198 19108 28198 19108 0 _0224_
rlabel metal1 31188 14314 31188 14314 0 _0225_
rlabel metal2 31234 18530 31234 18530 0 _0226_
rlabel metal2 37306 18020 37306 18020 0 _0227_
rlabel metal2 39514 19550 39514 19550 0 _0228_
rlabel metal1 38640 16150 38640 16150 0 _0229_
rlabel metal1 39928 13498 39928 13498 0 _0230_
rlabel metal2 37214 15708 37214 15708 0 _0231_
rlabel metal2 14122 37604 14122 37604 0 _0232_
rlabel metal2 14582 24990 14582 24990 0 _0233_
rlabel metal1 15272 41514 15272 41514 0 _0234_
rlabel metal1 17388 40698 17388 40698 0 _0235_
rlabel metal1 20332 41786 20332 41786 0 _0236_
rlabel metal2 21114 40086 21114 40086 0 _0237_
rlabel metal2 23322 41956 23322 41956 0 _0238_
rlabel metal1 25208 40698 25208 40698 0 _0239_
rlabel metal1 26818 42330 26818 42330 0 _0240_
rlabel metal1 29210 41208 29210 41208 0 _0241_
rlabel metal2 30866 41956 30866 41956 0 _0242_
rlabel metal1 32706 40698 32706 40698 0 _0243_
rlabel metal1 35420 42330 35420 42330 0 _0244_
rlabel metal1 37352 42126 37352 42126 0 _0245_
rlabel metal2 34730 39780 34730 39780 0 _0246_
rlabel metal1 37398 39066 37398 39066 0 _0247_
rlabel metal1 33074 37978 33074 37978 0 _0248_
rlabel metal1 17388 36890 17388 36890 0 _0249_
rlabel metal1 13386 39610 13386 39610 0 _0250_
rlabel metal2 15778 36516 15778 36516 0 _0251_
rlabel metal2 18262 35870 18262 35870 0 _0252_
rlabel metal1 21390 35802 21390 35802 0 _0253_
rlabel metal1 22724 35802 22724 35802 0 _0254_
rlabel metal2 24794 35428 24794 35428 0 _0255_
rlabel metal2 26174 35224 26174 35224 0 _0256_
rlabel metal2 27738 34782 27738 34782 0 _0257_
rlabel metal1 30590 35462 30590 35462 0 _0258_
rlabel metal1 30636 35734 30636 35734 0 _0259_
rlabel metal2 40710 39202 40710 39202 0 _0260_
rlabel metal1 41216 36346 41216 36346 0 _0261_
rlabel metal1 37812 34646 37812 34646 0 _0262_
rlabel metal1 34914 34170 34914 34170 0 _0263_
rlabel metal1 32844 36006 32844 36006 0 _0264_
rlabel metal2 14122 38692 14122 38692 0 _0265_
rlabel metal1 16238 39066 16238 39066 0 _0266_
rlabel metal1 18446 36856 18446 36856 0 _0267_
rlabel metal2 22126 37468 22126 37468 0 _0268_
rlabel metal1 22632 36890 22632 36890 0 _0269_
rlabel metal1 24978 36890 24978 36890 0 _0270_
rlabel metal1 26772 36890 26772 36890 0 _0271_
rlabel metal1 28106 35802 28106 35802 0 _0272_
rlabel metal2 29578 38114 29578 38114 0 _0273_
rlabel metal2 30498 36958 30498 36958 0 _0274_
rlabel metal1 40434 38522 40434 38522 0 _0275_
rlabel metal1 40342 35802 40342 35802 0 _0276_
rlabel metal1 37812 35802 37812 35802 0 _0277_
rlabel metal1 35420 34986 35420 34986 0 _0278_
rlabel metal1 33304 35598 33304 35598 0 _0279_
rlabel metal1 11776 35734 11776 35734 0 _0280_
rlabel metal1 15865 19754 15865 19754 0 _0281_
rlabel metal1 18262 21896 18262 21896 0 _0282_
rlabel metal1 21298 21896 21298 21896 0 _0283_
rlabel metal1 21385 23018 21385 23018 0 _0284_
rlabel metal2 23506 21318 23506 21318 0 _0285_
rlabel metal2 25622 21148 25622 21148 0 _0286_
rlabel metal1 27324 22202 27324 22202 0 _0287_
rlabel metal1 29941 23018 29941 23018 0 _0288_
rlabel metal2 30958 22406 30958 22406 0 _0289_
rlabel metal2 32614 21726 32614 21726 0 _0290_
rlabel metal1 37674 22202 37674 22202 0 _0291_
rlabel metal1 39560 21658 39560 21658 0 _0292_
rlabel metal1 39790 23290 39790 23290 0 _0293_
rlabel via1 37945 23086 37945 23086 0 _0294_
rlabel metal1 34500 20026 34500 20026 0 _0295_
rlabel via1 15230 23086 15230 23086 0 _0296_
rlabel metal1 11178 34034 11178 34034 0 _0297_
rlabel metal2 9154 28934 9154 28934 0 _0298_
rlabel metal1 7861 28458 7861 28458 0 _0299_
rlabel metal1 7631 29206 7631 29206 0 _0300_
rlabel metal2 10258 33286 10258 33286 0 _0301_
rlabel metal2 14950 34374 14950 34374 0 _0302_
rlabel metal2 16514 34850 16514 34850 0 _0303_
rlabel metal1 19591 34646 19591 34646 0 _0304_
rlabel via1 21201 33966 21201 33966 0 _0305_
rlabel metal1 23276 33626 23276 33626 0 _0306_
rlabel metal2 25070 33762 25070 33762 0 _0307_
rlabel via1 27273 32402 27273 32402 0 _0308_
rlabel metal2 28566 32198 28566 32198 0 _0309_
rlabel metal1 29854 33082 29854 33082 0 _0310_
rlabel metal2 32154 33082 32154 33082 0 _0311_
rlabel metal1 40848 33626 40848 33626 0 _0312_
rlabel metal2 39974 34102 39974 34102 0 _0313_
rlabel via1 37669 32878 37669 32878 0 _0314_
rlabel metal1 35415 32470 35415 32470 0 _0315_
rlabel metal2 33166 32674 33166 32674 0 _0316_
rlabel metal2 12834 33286 12834 33286 0 _0317_
rlabel metal1 15517 33558 15517 33558 0 _0318_
rlabel metal1 17066 33626 17066 33626 0 _0319_
rlabel metal1 19274 33626 19274 33626 0 _0320_
rlabel metal2 22126 33286 22126 33286 0 _0321_
rlabel metal2 23414 32674 23414 32674 0 _0322_
rlabel metal1 25162 31994 25162 31994 0 _0323_
rlabel metal1 26818 31212 26818 31212 0 _0324_
rlabel metal1 29593 31382 29593 31382 0 _0325_
rlabel metal1 30125 31790 30125 31790 0 _0326_
rlabel metal2 32798 30940 32798 30940 0 _0327_
rlabel via1 40613 32470 40613 32470 0 _0328_
rlabel metal1 39698 31688 39698 31688 0 _0329_
rlabel metal1 37766 31994 37766 31994 0 _0330_
rlabel metal1 35420 31994 35420 31994 0 _0331_
rlabel metal1 33115 31790 33115 31790 0 _0332_
rlabel metal1 13953 32470 13953 32470 0 _0333_
rlabel metal2 10442 27234 10442 27234 0 _0334_
rlabel metal1 11362 30362 11362 30362 0 _0335_
rlabel metal2 10166 30770 10166 30770 0 _0336_
rlabel metal2 10810 31314 10810 31314 0 _0337_
rlabel metal1 12282 21658 12282 21658 0 _0338_
rlabel metal1 11868 22678 11868 22678 0 _0339_
rlabel metal2 11822 23970 11822 23970 0 _0340_
rlabel metal2 11822 24990 11822 24990 0 _0341_
rlabel metal2 11270 26588 11270 26588 0 _0342_
rlabel metal2 15502 30668 15502 30668 0 _0343_
rlabel metal2 19458 28322 19458 28322 0 _0344_
rlabel metal1 16376 42194 16376 42194 0 _0345_
rlabel metal2 18170 42398 18170 42398 0 _0346_
rlabel metal1 21666 41786 21666 41786 0 _0347_
rlabel metal2 24794 28322 24794 28322 0 _0348_
rlabel metal1 24472 42602 24472 42602 0 _0349_
rlabel metal2 27462 27234 27462 27234 0 _0350_
rlabel metal2 28106 42670 28106 42670 0 _0351_
rlabel metal1 40940 25806 40940 25806 0 _0352_
rlabel metal2 40710 28254 40710 28254 0 _0353_
rlabel metal2 40710 29852 40710 29852 0 _0354_
rlabel metal1 39284 27030 39284 27030 0 _0355_
rlabel metal2 41078 31076 41078 31076 0 _0356_
rlabel metal2 40986 23970 40986 23970 0 _0357_
rlabel metal1 40112 29206 40112 29206 0 _0358_
rlabel metal1 40802 24922 40802 24922 0 _0359_
rlabel metal1 18538 32538 18538 32538 0 _0360_
rlabel metal1 18528 22610 18528 22610 0 _0361_
rlabel metal2 17802 20230 17802 20230 0 _0362_
rlabel via1 20097 22610 20097 22610 0 _0363_
rlabel metal1 19228 20910 19228 20910 0 _0364_
rlabel metal1 24472 21658 24472 21658 0 _0365_
rlabel metal2 26956 22746 26956 22746 0 _0366_
rlabel via1 27006 23086 27006 23086 0 _0367_
rlabel metal1 28336 23290 28336 23290 0 _0368_
rlabel metal1 31839 23018 31839 23018 0 _0369_
rlabel viali 33437 23086 33437 23086 0 _0370_
rlabel metal1 34653 22678 34653 22678 0 _0371_
rlabel metal1 35696 21386 35696 21386 0 _0372_
rlabel metal2 35282 21794 35282 21794 0 _0373_
rlabel via1 36758 20502 36758 20502 0 _0374_
rlabel metal1 34684 18802 34684 18802 0 _0375_
rlabel via1 14025 23698 14025 23698 0 _0376_
rlabel metal2 15410 19142 15410 19142 0 _0377_
rlabel metal2 14674 27438 14674 27438 0 _0378_
rlabel metal1 19182 28084 19182 28084 0 _0379_
rlabel metal2 18814 28866 18814 28866 0 _0380_
rlabel via2 15686 29053 15686 29053 0 _0381_
rlabel metal1 11040 30226 11040 30226 0 _0382_
rlabel metal1 10810 30226 10810 30226 0 _0383_
rlabel metal1 12098 30192 12098 30192 0 _0384_
rlabel metal1 17204 27438 17204 27438 0 _0385_
rlabel metal2 18722 26163 18722 26163 0 _0386_
rlabel metal1 18400 26282 18400 26282 0 _0387_
rlabel metal1 14030 29138 14030 29138 0 _0388_
rlabel metal2 13662 28832 13662 28832 0 _0389_
rlabel metal1 12328 27982 12328 27982 0 _0390_
rlabel metal2 13938 27353 13938 27353 0 _0391_
rlabel metal1 13064 27098 13064 27098 0 _0392_
rlabel metal2 12834 28458 12834 28458 0 _0393_
rlabel metal2 13754 27744 13754 27744 0 _0394_
rlabel metal1 13846 26316 13846 26316 0 _0395_
rlabel metal1 5658 5882 5658 5882 0 _0396_
rlabel metal1 5934 8432 5934 8432 0 _0397_
rlabel metal2 6670 9044 6670 9044 0 _0398_
rlabel metal2 10442 10778 10442 10778 0 _0399_
rlabel metal1 7958 10098 7958 10098 0 _0400_
rlabel metal1 7820 9622 7820 9622 0 _0401_
rlabel via2 6762 11645 6762 11645 0 _0402_
rlabel metal1 6164 11186 6164 11186 0 _0403_
rlabel metal1 7498 11730 7498 11730 0 _0404_
rlabel metal1 7866 9554 7866 9554 0 _0405_
rlabel metal2 8326 8908 8326 8908 0 _0406_
rlabel metal1 6670 11832 6670 11832 0 _0407_
rlabel metal1 6256 10030 6256 10030 0 _0408_
rlabel metal1 8280 7514 8280 7514 0 _0409_
rlabel metal1 10074 5338 10074 5338 0 _0410_
rlabel metal2 8326 7140 8326 7140 0 _0411_
rlabel metal1 8740 8058 8740 8058 0 _0412_
rlabel metal1 7222 11118 7222 11118 0 _0413_
rlabel metal2 7590 10812 7590 10812 0 _0414_
rlabel metal1 9430 10098 9430 10098 0 _0415_
rlabel metal2 9614 10268 9614 10268 0 _0416_
rlabel metal2 9890 10404 9890 10404 0 _0417_
rlabel metal2 7866 10200 7866 10200 0 _0418_
rlabel metal1 5244 4794 5244 4794 0 _0419_
rlabel metal1 4976 8602 4976 8602 0 _0420_
rlabel metal2 5658 9010 5658 9010 0 _0421_
rlabel metal1 7038 11186 7038 11186 0 _0422_
rlabel metal2 6578 9690 6578 9690 0 _0423_
rlabel metal2 7130 9962 7130 9962 0 _0424_
rlabel metal1 6164 9146 6164 9146 0 _0425_
rlabel via2 9062 7939 9062 7939 0 _0426_
rlabel metal1 9292 7174 9292 7174 0 _0427_
rlabel metal1 9292 6970 9292 6970 0 _0428_
rlabel metal1 9292 8058 9292 8058 0 _0429_
rlabel metal1 7820 7718 7820 7718 0 _0430_
rlabel metal1 7912 8602 7912 8602 0 _0431_
rlabel metal2 7544 11084 7544 11084 0 _0432_
rlabel metal1 5888 11322 5888 11322 0 _0433_
rlabel metal2 2070 11866 2070 11866 0 _0434_
rlabel metal2 6210 19006 6210 19006 0 _0435_
rlabel metal1 6440 18938 6440 18938 0 _0436_
rlabel metal1 12880 17102 12880 17102 0 _0437_
rlabel metal1 13110 16456 13110 16456 0 _0438_
rlabel metal1 9200 17238 9200 17238 0 _0439_
rlabel metal1 10212 17306 10212 17306 0 _0440_
rlabel metal1 12834 17748 12834 17748 0 _0441_
rlabel metal1 10902 17544 10902 17544 0 _0442_
rlabel metal1 12466 18632 12466 18632 0 _0443_
rlabel metal1 9706 15334 9706 15334 0 _0444_
rlabel metal1 8602 18802 8602 18802 0 _0445_
rlabel metal1 13984 16762 13984 16762 0 _0446_
rlabel metal2 12926 17612 12926 17612 0 _0447_
rlabel metal1 11224 17034 11224 17034 0 _0448_
rlabel metal1 9825 17102 9825 17102 0 _0449_
rlabel metal1 9614 16422 9614 16422 0 _0450_
rlabel metal1 7774 14484 7774 14484 0 _0451_
rlabel metal2 2714 12818 2714 12818 0 _0452_
rlabel metal1 6762 17782 6762 17782 0 _0453_
rlabel metal1 6210 17306 6210 17306 0 _0454_
rlabel metal1 7452 18054 7452 18054 0 _0455_
rlabel metal1 7544 17306 7544 17306 0 _0456_
rlabel metal1 8280 19482 8280 19482 0 _0457_
rlabel metal1 11270 17782 11270 17782 0 _0458_
rlabel metal2 10350 19652 10350 19652 0 _0459_
rlabel metal1 12128 18666 12128 18666 0 _0460_
rlabel metal1 11270 18938 11270 18938 0 _0461_
rlabel metal2 11914 19074 11914 19074 0 _0462_
rlabel metal2 12190 20434 12190 20434 0 _0463_
rlabel metal2 13110 18666 13110 18666 0 _0464_
rlabel metal1 13938 19380 13938 19380 0 _0465_
rlabel metal1 13018 16116 13018 16116 0 _0466_
rlabel metal1 15088 17646 15088 17646 0 _0467_
rlabel metal1 13110 15538 13110 15538 0 _0468_
rlabel metal1 14352 16082 14352 16082 0 _0469_
rlabel metal1 11546 15674 11546 15674 0 _0470_
rlabel metal1 13018 15402 13018 15402 0 _0471_
rlabel metal1 13018 15674 13018 15674 0 _0472_
rlabel metal1 11454 14586 11454 14586 0 _0473_
rlabel metal1 11132 14994 11132 14994 0 _0474_
rlabel metal2 13018 13362 13018 13362 0 _0475_
rlabel metal1 12830 14042 12830 14042 0 _0476_
rlabel metal2 13202 13090 13202 13090 0 _0477_
rlabel metal1 13754 11322 13754 11322 0 _0478_
rlabel metal1 7866 23290 7866 23290 0 _0479_
rlabel metal1 6670 23834 6670 23834 0 _0480_
rlabel metal1 7084 24786 7084 24786 0 _0481_
rlabel metal1 8326 24922 8326 24922 0 _0482_
rlabel metal1 8280 24650 8280 24650 0 _0483_
rlabel metal1 8924 23698 8924 23698 0 _0484_
rlabel metal1 7452 21998 7452 21998 0 _0485_
rlabel metal1 7406 21896 7406 21896 0 _0486_
rlabel metal1 7820 21658 7820 21658 0 _0487_
rlabel metal1 8234 21930 8234 21930 0 _0488_
rlabel metal1 8510 22576 8510 22576 0 _0489_
rlabel metal1 6900 22610 6900 22610 0 _0490_
rlabel metal1 8326 22644 8326 22644 0 _0491_
rlabel metal1 9016 22610 9016 22610 0 _0492_
rlabel metal1 8188 23086 8188 23086 0 _0493_
rlabel metal1 9016 23086 9016 23086 0 _0494_
rlabel metal2 9338 23902 9338 23902 0 _0495_
rlabel metal1 9476 23698 9476 23698 0 _0496_
rlabel metal1 2714 12784 2714 12784 0 _0497_
rlabel metal1 5625 10982 5625 10982 0 _0498_
rlabel metal1 3588 12818 3588 12818 0 _0499_
rlabel metal1 7498 9928 7498 9928 0 _0500_
rlabel metal2 6118 10948 6118 10948 0 _0501_
rlabel metal1 2530 11152 2530 11152 0 _0502_
rlabel metal1 3630 12954 3630 12954 0 _0503_
rlabel metal1 6486 13362 6486 13362 0 _0504_
rlabel metal1 5566 13940 5566 13940 0 _0505_
rlabel metal1 5382 13974 5382 13974 0 _0506_
rlabel via1 6758 14042 6758 14042 0 _0507_
rlabel metal1 9576 14246 9576 14246 0 _0508_
rlabel metal1 7912 15470 7912 15470 0 _0509_
rlabel metal1 10166 14416 10166 14416 0 _0510_
rlabel metal1 8510 13260 8510 13260 0 _0511_
rlabel metal1 10212 12410 10212 12410 0 _0512_
rlabel metal1 9982 12852 9982 12852 0 _0513_
rlabel metal1 9384 11118 9384 11118 0 _0514_
rlabel metal1 9890 9486 9890 9486 0 _0515_
rlabel metal1 11224 8942 11224 8942 0 _0516_
rlabel metal1 11316 10098 11316 10098 0 _0517_
rlabel metal2 5474 9384 5474 9384 0 _0518_
rlabel metal1 5428 9486 5428 9486 0 _0519_
rlabel metal1 3956 7922 3956 7922 0 _0520_
rlabel metal1 4232 7174 4232 7174 0 _0521_
rlabel metal1 4922 7888 4922 7888 0 _0522_
rlabel metal2 13018 6460 13018 6460 0 _0523_
rlabel metal1 3864 7514 3864 7514 0 _0524_
rlabel metal1 2438 7310 2438 7310 0 _0525_
rlabel metal2 2346 7718 2346 7718 0 _0526_
rlabel metal2 2714 7956 2714 7956 0 _0527_
rlabel metal1 2852 5678 2852 5678 0 _0528_
rlabel metal1 2622 5712 2622 5712 0 _0529_
rlabel metal2 3818 4794 3818 4794 0 _0530_
rlabel metal1 4140 4794 4140 4794 0 _0531_
rlabel metal1 4784 4114 4784 4114 0 _0532_
rlabel metal2 5382 3502 5382 3502 0 _0533_
rlabel metal1 5014 3570 5014 3570 0 _0534_
rlabel metal2 3542 3740 3542 3740 0 _0535_
rlabel metal2 6670 8092 6670 8092 0 _0536_
rlabel metal1 6808 7854 6808 7854 0 _0537_
rlabel metal2 6578 7208 6578 7208 0 _0538_
rlabel metal1 6762 5712 6762 5712 0 _0539_
rlabel metal2 7038 5236 7038 5236 0 _0540_
rlabel metal1 8280 4114 8280 4114 0 _0541_
rlabel metal1 8786 4454 8786 4454 0 _0542_
rlabel metal1 9154 4114 9154 4114 0 _0543_
rlabel metal2 11178 4012 11178 4012 0 _0544_
rlabel metal1 10580 3978 10580 3978 0 _0545_
rlabel metal1 8142 3604 8142 3604 0 _0546_
rlabel metal1 10028 4794 10028 4794 0 _0547_
rlabel metal2 10258 4250 10258 4250 0 _0548_
rlabel metal2 8970 6324 8970 6324 0 _0549_
rlabel metal1 12489 6766 12489 6766 0 _0550_
rlabel metal2 10074 5916 10074 5916 0 _0551_
rlabel metal1 12742 6664 12742 6664 0 _0552_
rlabel metal1 11040 6290 11040 6290 0 _0553_
rlabel metal1 10166 6256 10166 6256 0 _0554_
rlabel metal1 17204 31790 17204 31790 0 _0555_
rlabel metal1 17848 30702 17848 30702 0 _0556_
rlabel metal1 19918 27914 19918 27914 0 _0557_
rlabel metal2 20838 28832 20838 28832 0 _0558_
rlabel metal2 21206 28764 21206 28764 0 _0559_
rlabel metal1 16192 29206 16192 29206 0 _0560_
rlabel metal2 15962 30107 15962 30107 0 _0561_
rlabel metal2 17710 31178 17710 31178 0 _0562_
rlabel metal1 17204 30294 17204 30294 0 _0563_
rlabel metal1 16008 30906 16008 30906 0 _0564_
rlabel metal1 16008 31790 16008 31790 0 _0565_
rlabel metal1 20148 31314 20148 31314 0 _0566_
rlabel metal2 18722 30464 18722 30464 0 _0567_
rlabel metal1 19228 31790 19228 31790 0 _0568_
rlabel metal1 18446 30906 18446 30906 0 _0569_
rlabel metal1 18722 31824 18722 31824 0 _0570_
rlabel metal2 18078 32164 18078 32164 0 _0571_
rlabel viali 20194 30700 20194 30700 0 _0572_
rlabel metal2 21758 30430 21758 30430 0 _0573_
rlabel metal1 20148 30906 20148 30906 0 _0574_
rlabel metal1 20608 30362 20608 30362 0 _0575_
rlabel metal1 20470 30226 20470 30226 0 _0576_
rlabel metal3 21390 31756 21390 31756 0 _0577_
rlabel metal1 21528 31450 21528 31450 0 _0578_
rlabel metal1 24978 30260 24978 30260 0 _0579_
rlabel metal1 22034 30192 22034 30192 0 _0580_
rlabel metal2 21850 30396 21850 30396 0 _0581_
rlabel metal1 22816 30158 22816 30158 0 _0582_
rlabel metal1 22494 29818 22494 29818 0 _0583_
rlabel metal1 22172 27438 22172 27438 0 _0584_
rlabel metal1 21988 27438 21988 27438 0 _0585_
rlabel metal2 25990 30396 25990 30396 0 _0586_
rlabel metal1 24794 29818 24794 29818 0 _0587_
rlabel metal1 24104 30906 24104 30906 0 _0588_
rlabel metal1 24334 31450 24334 31450 0 _0589_
rlabel metal2 25806 29308 25806 29308 0 _0590_
rlabel metal2 25346 28730 25346 28730 0 _0591_
rlabel metal1 25438 28492 25438 28492 0 _0592_
rlabel metal1 26174 30090 26174 30090 0 _0593_
rlabel metal1 26496 30226 26496 30226 0 _0594_
rlabel metal2 27094 29818 27094 29818 0 _0595_
rlabel metal2 27186 30090 27186 30090 0 _0596_
rlabel metal1 30038 29682 30038 29682 0 _0597_
rlabel metal2 29486 29308 29486 29308 0 _0598_
rlabel metal2 29762 28730 29762 28730 0 _0599_
rlabel metal1 29716 28186 29716 28186 0 _0600_
rlabel metal1 30544 30362 30544 30362 0 _0601_
rlabel metal1 30590 29648 30590 29648 0 _0602_
rlabel metal2 30544 29138 30544 29138 0 _0603_
rlabel metal1 30636 29138 30636 29138 0 _0604_
rlabel metal1 37293 29478 37293 29478 0 _0605_
rlabel metal1 30774 30668 30774 30668 0 _0606_
rlabel metal2 31602 30396 31602 30396 0 _0607_
rlabel metal2 31694 30022 31694 30022 0 _0608_
rlabel metal2 37950 29342 37950 29342 0 _0609_
rlabel metal1 37812 29138 37812 29138 0 _0610_
rlabel metal1 37766 28186 37766 28186 0 _0611_
rlabel metal1 35834 30192 35834 30192 0 _0612_
rlabel metal1 37812 30022 37812 30022 0 _0613_
rlabel metal2 37858 30838 37858 30838 0 _0614_
rlabel metal1 37398 30906 37398 30906 0 _0615_
rlabel viali 35355 30294 35355 30294 0 _0616_
rlabel metal1 35512 29138 35512 29138 0 _0617_
rlabel metal2 36386 28764 36386 28764 0 _0618_
rlabel metal1 36478 28560 36478 28560 0 _0619_
rlabel metal2 34914 29410 34914 29410 0 _0620_
rlabel metal1 34868 31314 34868 31314 0 _0621_
rlabel metal2 36294 30804 36294 30804 0 _0622_
rlabel metal2 16146 30039 16146 30039 0 _0623_
rlabel metal1 34316 30022 34316 30022 0 _0624_
rlabel metal1 33994 29138 33994 29138 0 _0625_
rlabel metal1 34132 27914 34132 27914 0 _0626_
rlabel metal1 32154 25908 32154 25908 0 _0627_
rlabel metal1 19366 26316 19366 26316 0 _0628_
rlabel metal1 20286 27370 20286 27370 0 _0629_
rlabel metal1 17710 25398 17710 25398 0 _0630_
rlabel metal2 18170 25874 18170 25874 0 _0631_
rlabel metal1 17802 25466 17802 25466 0 _0632_
rlabel metal1 20010 24718 20010 24718 0 _0633_
rlabel metal2 18998 24276 18998 24276 0 _0634_
rlabel viali 18630 24106 18630 24106 0 _0635_
rlabel metal1 19872 24786 19872 24786 0 _0636_
rlabel metal1 17526 24038 17526 24038 0 _0637_
rlabel metal1 21252 24786 21252 24786 0 _0638_
rlabel metal2 20102 24854 20102 24854 0 _0639_
rlabel metal2 21022 25058 21022 25058 0 _0640_
rlabel metal1 20378 24922 20378 24922 0 _0641_
rlabel metal2 20286 25670 20286 25670 0 _0642_
rlabel metal2 20746 26146 20746 26146 0 _0643_
rlabel metal2 23874 25568 23874 25568 0 _0644_
rlabel metal1 22034 24752 22034 24752 0 _0645_
rlabel metal2 21482 24582 21482 24582 0 _0646_
rlabel metal2 22494 25092 22494 25092 0 _0647_
rlabel metal1 21850 25160 21850 25160 0 _0648_
rlabel metal1 21712 24922 21712 24922 0 _0649_
rlabel metal2 21574 25636 21574 25636 0 _0650_
rlabel metal1 24564 24718 24564 24718 0 _0651_
rlabel metal1 23736 25194 23736 25194 0 _0652_
rlabel metal2 23690 25466 23690 25466 0 _0653_
rlabel metal1 24012 24786 24012 24786 0 _0654_
rlabel metal1 25208 26486 25208 26486 0 _0655_
rlabel metal1 25208 26010 25208 26010 0 _0656_
rlabel metal1 25024 25738 25024 25738 0 _0657_
rlabel metal1 26082 25466 26082 25466 0 _0658_
rlabel metal2 31786 24412 31786 24412 0 _0659_
rlabel viali 26082 25874 26082 25874 0 _0660_
rlabel metal1 26910 24786 26910 24786 0 _0661_
rlabel metal1 28888 25466 28888 25466 0 _0662_
rlabel metal2 29578 25092 29578 25092 0 _0663_
rlabel metal2 28750 26078 28750 26078 0 _0664_
rlabel metal2 28566 25500 28566 25500 0 _0665_
rlabel metal2 30038 25500 30038 25500 0 _0666_
rlabel metal2 30406 25602 30406 25602 0 _0667_
rlabel metal2 33074 24582 33074 24582 0 _0668_
rlabel metal1 32430 24718 32430 24718 0 _0669_
rlabel metal1 32338 24752 32338 24752 0 _0670_
rlabel metal1 32108 24786 32108 24786 0 _0671_
rlabel metal2 37306 24378 37306 24378 0 _0672_
rlabel metal2 37122 24922 37122 24922 0 _0673_
rlabel metal1 37766 24378 37766 24378 0 _0674_
rlabel metal1 36654 26214 36654 26214 0 _0675_
rlabel metal1 37306 25942 37306 25942 0 _0676_
rlabel metal1 37260 24718 37260 24718 0 _0677_
rlabel metal1 37260 25330 37260 25330 0 _0678_
rlabel metal1 35696 24786 35696 24786 0 _0679_
rlabel metal2 36570 24582 36570 24582 0 _0680_
rlabel metal1 35880 24242 35880 24242 0 _0681_
rlabel metal1 36064 25330 36064 25330 0 _0682_
rlabel metal2 36018 25772 36018 25772 0 _0683_
rlabel metal2 35282 25024 35282 25024 0 _0684_
rlabel metal2 33810 24412 33810 24412 0 _0685_
rlabel metal2 33902 25092 33902 25092 0 _0686_
rlabel metal1 33534 25466 33534 25466 0 _0687_
rlabel metal1 39468 12138 39468 12138 0 _0688_
rlabel metal1 14168 34034 14168 34034 0 _0689_
rlabel metal2 14306 35360 14306 35360 0 _0690_
rlabel metal1 14674 36176 14674 36176 0 _0691_
rlabel metal1 15226 22134 15226 22134 0 _0692_
rlabel metal2 17434 13702 17434 13702 0 _0693_
rlabel metal2 18814 16218 18814 16218 0 _0694_
rlabel metal1 18860 15674 18860 15674 0 _0695_
rlabel metal1 19918 17510 19918 17510 0 _0696_
rlabel metal1 19688 18190 19688 18190 0 _0697_
rlabel metal1 18998 17102 18998 17102 0 _0698_
rlabel metal1 18906 17204 18906 17204 0 _0699_
rlabel metal2 21482 17714 21482 17714 0 _0700_
rlabel metal1 21344 17034 21344 17034 0 _0701_
rlabel metal2 20930 16762 20930 16762 0 _0702_
rlabel metal1 20746 17170 20746 17170 0 _0703_
rlabel metal2 20838 17578 20838 17578 0 _0704_
rlabel metal2 20470 16286 20470 16286 0 _0705_
rlabel metal2 24150 17646 24150 17646 0 _0706_
rlabel metal1 21942 17612 21942 17612 0 _0707_
rlabel metal1 22264 17646 22264 17646 0 _0708_
rlabel metal1 21942 17748 21942 17748 0 _0709_
rlabel metal1 22264 17850 22264 17850 0 _0710_
rlabel metal1 24288 17034 24288 17034 0 _0711_
rlabel metal2 24978 16966 24978 16966 0 _0712_
rlabel metal1 24518 16558 24518 16558 0 _0713_
rlabel metal1 21850 17544 21850 17544 0 _0714_
rlabel metal1 24794 17204 24794 17204 0 _0715_
rlabel metal1 24840 16150 24840 16150 0 _0716_
rlabel metal1 27462 17578 27462 17578 0 _0717_
rlabel via2 28474 17187 28474 17187 0 _0718_
rlabel metal1 26496 18258 26496 18258 0 _0719_
rlabel metal1 25576 17238 25576 17238 0 _0720_
rlabel metal1 25116 17238 25116 17238 0 _0721_
rlabel metal1 25392 17306 25392 17306 0 _0722_
rlabel metal1 25070 17612 25070 17612 0 _0723_
rlabel metal2 29486 16898 29486 16898 0 _0724_
rlabel metal2 29210 16898 29210 16898 0 _0725_
rlabel metal1 28520 16558 28520 16558 0 _0726_
rlabel metal1 27600 17034 27600 17034 0 _0727_
rlabel metal2 29118 16898 29118 16898 0 _0728_
rlabel metal2 28842 16745 28842 16745 0 _0729_
rlabel metal1 30268 17646 30268 17646 0 _0730_
rlabel metal1 30682 17714 30682 17714 0 _0731_
rlabel metal2 29210 18122 29210 18122 0 _0732_
rlabel metal2 28934 17850 28934 17850 0 _0733_
rlabel metal2 28474 18530 28474 18530 0 _0734_
rlabel metal1 28566 17850 28566 17850 0 _0735_
rlabel metal1 32568 17102 32568 17102 0 _0736_
rlabel metal1 31694 17034 31694 17034 0 _0737_
rlabel metal1 30958 17136 30958 17136 0 _0738_
rlabel metal1 30498 17646 30498 17646 0 _0739_
rlabel metal2 30866 17442 30866 17442 0 _0740_
rlabel metal2 31510 16762 31510 16762 0 _0741_
rlabel metal1 32752 17306 32752 17306 0 _0742_
rlabel metal1 32706 19448 32706 19448 0 _0743_
rlabel metal1 32016 17782 32016 17782 0 _0744_
rlabel metal2 31510 18734 31510 18734 0 _0745_
rlabel metal1 32062 17306 32062 17306 0 _0746_
rlabel metal1 37720 19142 37720 19142 0 _0747_
rlabel metal2 37214 18258 37214 18258 0 _0748_
rlabel metal1 37766 17850 37766 17850 0 _0749_
rlabel metal1 32108 17850 32108 17850 0 _0750_
rlabel metal2 36202 18326 36202 18326 0 _0751_
rlabel metal2 37674 18258 37674 18258 0 _0752_
rlabel metal2 41814 19414 41814 19414 0 _0753_
rlabel metal2 40342 19584 40342 19584 0 _0754_
rlabel metal1 39974 18258 39974 18258 0 _0755_
rlabel metal1 39652 18870 39652 18870 0 _0756_
rlabel metal2 40250 18972 40250 18972 0 _0757_
rlabel metal2 40802 17374 40802 17374 0 _0758_
rlabel metal1 40020 17238 40020 17238 0 _0759_
rlabel metal2 40342 17918 40342 17918 0 _0760_
rlabel metal1 39422 17272 39422 17272 0 _0761_
rlabel metal1 39514 17136 39514 17136 0 _0762_
rlabel metal2 41630 15436 41630 15436 0 _0763_
rlabel metal2 40250 15776 40250 15776 0 _0764_
rlabel metal2 40618 16252 40618 16252 0 _0765_
rlabel metal2 41722 14518 41722 14518 0 _0766_
rlabel metal2 40066 13770 40066 13770 0 _0767_
rlabel metal1 36064 14994 36064 14994 0 _0768_
rlabel metal1 35926 14892 35926 14892 0 _0769_
rlabel metal1 36984 14790 36984 14790 0 _0770_
rlabel metal2 16698 25058 16698 25058 0 _0771_
rlabel metal2 16606 25313 16606 25313 0 _0772_
rlabel metal1 15916 25330 15916 25330 0 _0773_
rlabel metal2 15134 25738 15134 25738 0 _0774_
rlabel metal1 17434 41208 17434 41208 0 _0775_
rlabel via1 34362 36550 34362 36550 0 _0776_
rlabel metal1 34270 36788 34270 36788 0 _0777_
rlabel metal1 34454 37196 34454 37196 0 _0778_
rlabel metal1 36340 36822 36340 36822 0 _0779_
rlabel metal2 36846 36550 36846 36550 0 _0780_
rlabel metal2 36018 36890 36018 36890 0 _0781_
rlabel metal2 36938 37128 36938 37128 0 _0782_
rlabel metal1 38732 36822 38732 36822 0 _0783_
rlabel metal2 39146 36550 39146 36550 0 _0784_
rlabel metal1 38456 37842 38456 37842 0 _0785_
rlabel metal2 37674 37060 37674 37060 0 _0786_
rlabel metal2 40342 37400 40342 37400 0 _0787_
rlabel metal1 39928 37434 39928 37434 0 _0788_
rlabel metal1 39100 38318 39100 38318 0 _0789_
rlabel metal1 38870 38760 38870 38760 0 _0790_
rlabel metal1 39744 39406 39744 39406 0 _0791_
rlabel metal1 40112 39066 40112 39066 0 _0792_
rlabel metal2 39698 39406 39698 39406 0 _0793_
rlabel via1 39605 40018 39605 40018 0 _0794_
rlabel metal2 32522 38012 32522 38012 0 _0795_
rlabel metal1 33120 37910 33120 37910 0 _0796_
rlabel metal1 36938 39950 36938 39950 0 _0797_
rlabel metal2 32338 39304 32338 39304 0 _0798_
rlabel metal1 32890 38964 32890 38964 0 _0799_
rlabel metal1 30636 37910 30636 37910 0 _0800_
rlabel metal2 31050 39508 31050 39508 0 _0801_
rlabel metal2 31694 39338 31694 39338 0 _0802_
rlabel metal2 28658 38114 28658 38114 0 _0803_
rlabel metal2 28934 38148 28934 38148 0 _0804_
rlabel metal1 29026 39338 29026 39338 0 _0805_
rlabel metal2 28566 39032 28566 39032 0 _0806_
rlabel metal1 27600 37910 27600 37910 0 _0807_
rlabel metal2 27922 37366 27922 37366 0 _0808_
rlabel metal1 27462 38930 27462 38930 0 _0809_
rlabel metal1 27646 38896 27646 38896 0 _0810_
rlabel metal2 25254 38726 25254 38726 0 _0811_
rlabel metal2 25714 38624 25714 38624 0 _0812_
rlabel metal1 25806 39338 25806 39338 0 _0813_
rlabel metal2 25254 39304 25254 39304 0 _0814_
rlabel metal2 23782 38726 23782 38726 0 _0815_
rlabel metal2 23966 38726 23966 38726 0 _0816_
rlabel metal2 24058 39338 24058 39338 0 _0817_
rlabel metal1 24426 39066 24426 39066 0 _0818_
rlabel metal1 21758 38522 21758 38522 0 _0819_
rlabel metal2 22310 38369 22310 38369 0 _0820_
rlabel metal1 24150 39474 24150 39474 0 _0821_
rlabel via1 21037 38930 21037 38930 0 _0822_
rlabel metal1 19596 38318 19596 38318 0 _0823_
rlabel metal2 19274 38148 19274 38148 0 _0824_
rlabel metal1 19504 38930 19504 38930 0 _0825_
rlabel metal2 19734 38964 19734 38964 0 _0826_
rlabel metal2 17710 38352 17710 38352 0 _0827_
rlabel metal2 18446 39236 18446 39236 0 _0828_
rlabel metal2 17158 39644 17158 39644 0 _0829_
rlabel metal1 18630 39440 18630 39440 0 _0830_
rlabel metal2 18630 39780 18630 39780 0 _0831_
rlabel metal1 19918 39066 19918 39066 0 _0832_
rlabel metal1 23138 39338 23138 39338 0 _0833_
rlabel metal2 23138 39814 23138 39814 0 _0834_
rlabel metal1 24656 39610 24656 39610 0 _0835_
rlabel metal1 26542 39440 26542 39440 0 _0836_
rlabel metal2 26542 39814 26542 39814 0 _0837_
rlabel metal1 27784 39406 27784 39406 0 _0838_
rlabel via2 31786 39389 31786 39389 0 _0839_
rlabel metal2 30774 40324 30774 40324 0 _0840_
rlabel metal1 32108 39610 32108 39610 0 _0841_
rlabel metal1 37122 39916 37122 39916 0 _0842_
rlabel metal1 37444 40154 37444 40154 0 _0843_
rlabel metal1 38548 40018 38548 40018 0 _0844_
rlabel metal1 38456 38318 38456 38318 0 _0845_
rlabel metal1 38226 38352 38226 38352 0 _0846_
rlabel metal1 36892 37842 36892 37842 0 _0847_
rlabel metal1 36547 37298 36547 37298 0 _0848_
rlabel metal2 35466 37502 35466 37502 0 _0849_
rlabel metal2 34178 36924 34178 36924 0 _0850_
rlabel metal1 34822 37264 34822 37264 0 _0851_
rlabel metal2 35282 37349 35282 37349 0 _0852_
rlabel metal2 17342 39746 17342 39746 0 _0853_
rlabel metal1 19550 41072 19550 41072 0 _0854_
rlabel metal1 17848 40494 17848 40494 0 _0855_
rlabel metal1 17710 40562 17710 40562 0 _0856_
rlabel metal1 17480 40630 17480 40630 0 _0857_
rlabel metal1 20286 40528 20286 40528 0 _0858_
rlabel metal2 20010 41412 20010 41412 0 _0859_
rlabel metal2 18722 39746 18722 39746 0 _0860_
rlabel metal2 20102 40290 20102 40290 0 _0861_
rlabel metal1 20654 41514 20654 41514 0 _0862_
rlabel metal1 21252 40630 21252 40630 0 _0863_
rlabel metal1 20562 39066 20562 39066 0 _0864_
rlabel metal1 20562 40460 20562 40460 0 _0865_
rlabel metal1 21156 40154 21156 40154 0 _0866_
rlabel metal1 21482 40562 21482 40562 0 _0867_
rlabel metal1 21804 41106 21804 41106 0 _0868_
rlabel metal1 23138 41072 23138 41072 0 _0869_
rlabel metal2 23230 39746 23230 39746 0 _0870_
rlabel metal1 23506 41106 23506 41106 0 _0871_
rlabel metal1 23644 41242 23644 41242 0 _0872_
rlabel metal1 26266 40494 26266 40494 0 _0873_
rlabel metal2 25162 39780 25162 39780 0 _0874_
rlabel metal2 26082 40290 26082 40290 0 _0875_
rlabel metal1 25852 40494 25852 40494 0 _0876_
rlabel metal1 25622 40562 25622 40562 0 _0877_
rlabel metal2 27370 41321 27370 41321 0 _0878_
rlabel metal2 26818 39780 26818 39780 0 _0879_
rlabel metal1 27738 40562 27738 40562 0 _0880_
rlabel metal1 27370 42194 27370 42194 0 _0881_
rlabel metal2 27370 41956 27370 41956 0 _0882_
rlabel metal1 28198 39474 28198 39474 0 _0883_
rlabel metal2 28198 40052 28198 40052 0 _0884_
rlabel metal1 28704 40562 28704 40562 0 _0885_
rlabel metal1 28428 40698 28428 40698 0 _0886_
rlabel metal2 30498 41106 30498 41106 0 _0887_
rlabel metal1 30636 39610 30636 39610 0 _0888_
rlabel metal1 31786 41548 31786 41548 0 _0889_
rlabel metal2 31142 41650 31142 41650 0 _0890_
rlabel metal1 31050 41514 31050 41514 0 _0891_
rlabel metal1 32154 41140 32154 41140 0 _0892_
rlabel metal2 32246 39780 32246 39780 0 _0893_
rlabel metal2 32430 40630 32430 40630 0 _0894_
rlabel metal2 32798 40698 32798 40698 0 _0895_
rlabel metal2 32706 41004 32706 41004 0 _0896_
rlabel metal1 36478 41038 36478 41038 0 _0897_
rlabel metal2 39330 40222 39330 40222 0 _0898_
rlabel metal2 36846 41106 36846 41106 0 _0899_
rlabel metal2 35650 41956 35650 41956 0 _0900_
rlabel metal2 35374 41956 35374 41956 0 _0901_
rlabel metal1 36202 41548 36202 41548 0 _0902_
rlabel metal1 38594 39066 38594 39066 0 _0903_
rlabel metal1 36662 41106 36662 41106 0 _0904_
rlabel metal1 36570 41786 36570 41786 0 _0905_
rlabel metal1 36202 38964 36202 38964 0 _0906_
rlabel metal1 37996 37978 37996 37978 0 _0907_
rlabel metal1 36754 38726 36754 38726 0 _0908_
rlabel metal1 35006 39440 35006 39440 0 _0909_
rlabel metal1 34914 39372 34914 39372 0 _0910_
rlabel metal1 35972 39066 35972 39066 0 _0911_
rlabel metal2 36478 37604 36478 37604 0 _0912_
rlabel metal2 36018 38454 36018 38454 0 _0913_
rlabel metal1 37398 38998 37398 38998 0 _0914_
rlabel metal2 35834 38692 35834 38692 0 _0915_
rlabel metal2 34270 37604 34270 37604 0 _0916_
rlabel metal2 34822 38182 34822 38182 0 _0917_
rlabel metal1 34684 37910 34684 37910 0 _0918_
rlabel metal2 17710 37026 17710 37026 0 _0919_
rlabel metal2 15502 35462 15502 35462 0 _0920_
rlabel metal1 14352 35190 14352 35190 0 _0921_
rlabel metal1 16422 36006 16422 36006 0 _0922_
rlabel metal1 19550 35258 19550 35258 0 _0923_
rlabel metal1 22402 35258 22402 35258 0 _0924_
rlabel metal1 23414 35258 23414 35258 0 _0925_
rlabel metal2 25254 34816 25254 34816 0 _0926_
rlabel metal2 27002 34850 27002 34850 0 _0927_
rlabel metal1 29532 34170 29532 34170 0 _0928_
rlabel metal2 30866 34986 30866 34986 0 _0929_
rlabel metal2 31510 35190 31510 35190 0 _0930_
rlabel metal1 41124 35802 41124 35802 0 _0931_
rlabel metal1 40802 36006 40802 36006 0 _0932_
rlabel metal1 38318 34170 38318 34170 0 _0933_
rlabel metal1 35650 33830 35650 33830 0 _0934_
rlabel metal2 33442 34816 33442 34816 0 _0935_
rlabel metal2 14674 36992 14674 36992 0 _0936_
rlabel metal1 17296 35802 17296 35802 0 _0937_
rlabel metal2 19826 36312 19826 36312 0 _0938_
rlabel metal2 22402 36550 22402 36550 0 _0939_
rlabel metal2 23506 35666 23506 35666 0 _0940_
rlabel metal2 26082 35768 26082 35768 0 _0941_
rlabel metal1 27738 34170 27738 34170 0 _0942_
rlabel metal1 28704 34170 28704 34170 0 _0943_
rlabel metal2 30038 36244 30038 36244 0 _0944_
rlabel metal1 31556 35258 31556 35258 0 _0945_
rlabel metal2 40986 36448 40986 36448 0 _0946_
rlabel metal2 40434 35428 40434 35428 0 _0947_
rlabel metal2 39146 34544 39146 34544 0 _0948_
rlabel metal1 36340 34170 36340 34170 0 _0949_
rlabel metal1 34224 34170 34224 34170 0 _0950_
rlabel metal2 12282 36380 12282 36380 0 _0951_
rlabel metal1 13156 29682 13156 29682 0 _0952_
rlabel metal2 11638 28356 11638 28356 0 _0953_
rlabel metal2 13018 20944 13018 20944 0 _0954_
rlabel metal1 11040 28390 11040 28390 0 _0955_
rlabel metal1 13018 31654 13018 31654 0 _0956_
rlabel metal2 16422 24752 16422 24752 0 _0957_
rlabel metal1 18446 20026 18446 20026 0 _0958_
rlabel metal1 14674 20434 14674 20434 0 _0959_
rlabel metal2 16330 19516 16330 19516 0 _0960_
rlabel metal1 16974 20570 16974 20570 0 _0961_
rlabel via2 18630 21981 18630 21981 0 _0962_
rlabel via2 21666 21981 21666 21981 0 _0963_
rlabel metal1 22862 27574 22862 27574 0 _0964_
rlabel metal2 22402 25636 22402 25636 0 _0965_
rlabel metal1 23828 20910 23828 20910 0 _0966_
rlabel metal1 26404 20910 26404 20910 0 _0967_
rlabel metal2 27784 29138 27784 29138 0 _0968_
rlabel metal2 29946 25398 29946 25398 0 _0969_
rlabel metal1 32246 27404 32246 27404 0 _0970_
rlabel metal2 33166 25568 33166 25568 0 _0971_
rlabel metal1 38088 21998 38088 21998 0 _0972_
rlabel metal1 39836 21658 39836 21658 0 _0973_
rlabel metal1 40158 23086 40158 23086 0 _0974_
rlabel metal2 38226 26724 38226 26724 0 _0975_
rlabel metal2 34178 20951 34178 20951 0 _0976_
rlabel metal1 18607 32402 18607 32402 0 _0977_
rlabel metal2 33442 32130 33442 32130 0 _0978_
rlabel metal1 9844 28390 9844 28390 0 _0979_
rlabel metal2 8510 28832 8510 28832 0 _0980_
rlabel metal2 9430 28832 9430 28832 0 _0981_
rlabel metal1 13662 27574 13662 27574 0 _0982_
rlabel metal1 13294 28186 13294 28186 0 _0983_
rlabel metal1 11730 28560 11730 28560 0 _0984_
rlabel metal2 11546 27642 11546 27642 0 _0985_
rlabel metal1 16008 30090 16008 30090 0 _0986_
rlabel metal2 15226 30396 15226 30396 0 _0987_
rlabel metal1 17664 29274 17664 29274 0 _0988_
rlabel metal1 14950 29274 14950 29274 0 _0989_
rlabel via1 35192 27438 35192 27438 0 _0990_
rlabel metal2 38962 27999 38962 27999 0 _0991_
rlabel metal2 17802 27744 17802 27744 0 _0992_
rlabel metal1 16330 42296 16330 42296 0 _0993_
rlabel metal1 16054 42194 16054 42194 0 _0994_
rlabel metal1 18906 42602 18906 42602 0 _0995_
rlabel metal1 18722 42670 18722 42670 0 _0996_
rlabel metal1 21712 41514 21712 41514 0 _0997_
rlabel metal2 21390 41457 21390 41457 0 _0998_
rlabel metal2 24610 28560 24610 28560 0 _0999_
rlabel metal2 24426 28798 24426 28798 0 _1000_
rlabel metal2 24058 42874 24058 42874 0 _1001_
rlabel metal1 23644 30906 23644 30906 0 _1002_
rlabel metal2 26910 27642 26910 27642 0 _1003_
rlabel metal1 26864 27098 26864 27098 0 _1004_
rlabel metal1 28428 42874 28428 42874 0 _1005_
rlabel metal1 28244 29274 28244 29274 0 _1006_
rlabel metal1 40986 27336 40986 27336 0 _1007_
rlabel metal2 40802 27098 40802 27098 0 _1008_
rlabel metal1 40434 28186 40434 28186 0 _1009_
rlabel metal2 39882 28016 39882 28016 0 _1010_
rlabel metal1 41078 30192 41078 30192 0 _1011_
rlabel metal1 33902 28934 33902 28934 0 _1012_
rlabel metal1 38962 26010 38962 26010 0 _1013_
rlabel metal2 38962 26928 38962 26928 0 _1014_
rlabel metal2 40894 30906 40894 30906 0 _1015_
rlabel metal1 39836 30090 39836 30090 0 _1016_
rlabel metal1 35834 27472 35834 27472 0 _1017_
rlabel metal2 41354 25126 41354 25126 0 _1018_
rlabel metal1 39836 29274 39836 29274 0 _1019_
rlabel metal1 39882 29512 39882 29512 0 _1020_
rlabel metal2 34730 27642 34730 27642 0 _1021_
rlabel metal1 41170 24922 41170 24922 0 _1022_
rlabel metal1 19044 29274 19044 29274 0 _1023_
rlabel metal2 10074 29308 10074 29308 0 _1024_
rlabel metal1 5336 28050 5336 28050 0 _1025_
rlabel metal1 5290 31858 5290 31858 0 _1026_
rlabel metal2 4278 18530 4278 18530 0 _1027_
rlabel metal2 26542 13872 26542 13872 0 _1028_
rlabel metal1 16054 28390 16054 28390 0 _1029_
rlabel metal1 19090 28016 19090 28016 0 _1030_
rlabel metal1 14812 20570 14812 20570 0 _1031_
rlabel metal1 19734 14246 19734 14246 0 _1032_
rlabel metal1 36087 42194 36087 42194 0 _1033_
rlabel metal1 7958 24786 7958 24786 0 _1034_
rlabel metal1 7590 26010 7590 26010 0 _1035_
rlabel metal2 3266 3706 3266 3706 0 _1036_
rlabel metal1 10442 6324 10442 6324 0 _1037_
rlabel via2 33994 37213 33994 37213 0 _1038_
rlabel metal1 25530 29648 25530 29648 0 _1039_
rlabel metal2 4278 30158 4278 30158 0 _1040_
rlabel metal1 5704 32946 5704 32946 0 _1041_
rlabel metal1 6394 33082 6394 33082 0 _1042_
rlabel metal1 5152 30838 5152 30838 0 _1043_
rlabel metal2 4922 28730 4922 28730 0 _1044_
rlabel metal1 5612 30090 5612 30090 0 _1045_
rlabel metal2 4094 26690 4094 26690 0 _1046_
rlabel metal1 5428 29138 5428 29138 0 _1047_
rlabel metal2 4692 18700 4692 18700 0 _1048_
rlabel metal1 4876 24174 4876 24174 0 _1049_
rlabel metal1 4646 24786 4646 24786 0 _1050_
rlabel metal1 3404 23562 3404 23562 0 _1051_
rlabel metal2 10626 18479 10626 18479 0 _1052_
rlabel metal1 5336 18870 5336 18870 0 _1053_
rlabel metal1 8326 24174 8326 24174 0 _1054_
rlabel metal1 4278 26928 4278 26928 0 _1055_
rlabel metal2 3542 26452 3542 26452 0 _1056_
rlabel metal1 8464 33966 8464 33966 0 _1057_
rlabel metal1 4968 27506 4968 27506 0 _1058_
rlabel metal1 3312 24378 3312 24378 0 _1059_
rlabel metal1 1886 24208 1886 24208 0 _1060_
rlabel metal1 20010 12614 20010 12614 0 _1061_
rlabel metal2 26082 13532 26082 13532 0 _1062_
rlabel metal1 21551 14042 21551 14042 0 _1063_
rlabel metal1 35374 13226 35374 13226 0 _1064_
rlabel metal1 29026 13464 29026 13464 0 _1065_
rlabel metal2 26358 13702 26358 13702 0 _1066_
rlabel metal2 22310 12036 22310 12036 0 _1067_
rlabel metal1 23460 10098 23460 10098 0 _1068_
rlabel metal1 24334 9146 24334 9146 0 _1069_
rlabel metal1 27600 9350 27600 9350 0 _1070_
rlabel metal1 32430 8840 32430 8840 0 _1071_
rlabel metal2 33902 9588 33902 9588 0 _1072_
rlabel metal1 35650 9520 35650 9520 0 _1073_
rlabel metal2 36938 10370 36938 10370 0 _1074_
rlabel metal1 37812 10778 37812 10778 0 _1075_
rlabel metal1 37812 12614 37812 12614 0 _1076_
rlabel metal1 36938 8466 36938 8466 0 _1077_
rlabel metal1 36294 12954 36294 12954 0 _1078_
rlabel via1 26741 8942 26741 8942 0 _1079_
rlabel metal1 26864 8806 26864 8806 0 _1080_
rlabel metal2 24242 10438 24242 10438 0 _1081_
rlabel metal1 26220 11798 26220 11798 0 _1082_
rlabel metal1 22954 9350 22954 9350 0 _1083_
rlabel metal2 22218 11322 22218 11322 0 _1084_
rlabel metal1 21482 12172 21482 12172 0 _1085_
rlabel metal1 22356 10778 22356 10778 0 _1086_
rlabel metal2 21850 11900 21850 11900 0 _1087_
rlabel metal2 18538 11560 18538 11560 0 _1088_
rlabel metal2 20102 11900 20102 11900 0 _1089_
rlabel viali 21942 11730 21942 11730 0 _1090_
rlabel metal2 22494 12036 22494 12036 0 _1091_
rlabel metal1 23644 9146 23644 9146 0 _1092_
rlabel metal1 24886 11798 24886 11798 0 _1093_
rlabel metal1 26266 11696 26266 11696 0 _1094_
rlabel metal1 27416 11866 27416 11866 0 _1095_
rlabel metal1 28428 11118 28428 11118 0 _1096_
rlabel metal1 28106 11322 28106 11322 0 _1097_
rlabel metal2 31510 9860 31510 9860 0 _1098_
rlabel metal1 28934 11832 28934 11832 0 _1099_
rlabel metal1 28382 11730 28382 11730 0 _1100_
rlabel metal2 28382 11288 28382 11288 0 _1101_
rlabel metal2 31970 9758 31970 9758 0 _1102_
rlabel metal1 32200 9350 32200 9350 0 _1103_
rlabel metal1 31924 11118 31924 11118 0 _1104_
rlabel metal1 32476 10030 32476 10030 0 _1105_
rlabel metal2 32246 11322 32246 11322 0 _1106_
rlabel metal1 32522 11322 32522 11322 0 _1107_
rlabel metal2 34730 9894 34730 9894 0 _1108_
rlabel metal1 34822 9350 34822 9350 0 _1109_
rlabel metal1 34224 11322 34224 11322 0 _1110_
rlabel metal1 37582 12750 37582 12750 0 _1111_
rlabel metal1 35558 10438 35558 10438 0 _1112_
rlabel metal1 35926 11050 35926 11050 0 _1113_
rlabel metal1 36570 11186 36570 11186 0 _1114_
rlabel metal1 37352 12614 37352 12614 0 _1115_
rlabel metal1 29118 13260 29118 13260 0 _1116_
rlabel metal2 28842 13498 28842 13498 0 _1117_
rlabel metal1 5382 27948 5382 27948 0 _1118_
rlabel metal2 5290 27642 5290 27642 0 _1119_
rlabel metal1 4876 27642 4876 27642 0 _1120_
rlabel metal1 3468 29614 3468 29614 0 _1121_
rlabel metal1 4094 28594 4094 28594 0 _1122_
rlabel metal1 3404 31790 3404 31790 0 _1123_
rlabel metal2 5474 29920 5474 29920 0 _1124_
rlabel metal1 4968 28730 4968 28730 0 _1125_
rlabel metal1 7222 36040 7222 36040 0 _1126_
rlabel metal2 7130 36346 7130 36346 0 _1127_
rlabel metal2 7314 37638 7314 37638 0 _1128_
rlabel metal1 7222 37876 7222 37876 0 _1129_
rlabel metal1 8694 37094 8694 37094 0 _1130_
rlabel metal1 8510 37366 8510 37366 0 _1131_
rlabel metal1 6256 37978 6256 37978 0 _1132_
rlabel metal2 4646 36754 4646 36754 0 _1133_
rlabel metal2 4462 36924 4462 36924 0 _1134_
rlabel metal2 2622 38012 2622 38012 0 _1135_
rlabel metal2 1886 37638 1886 37638 0 _1136_
rlabel metal1 2530 37808 2530 37808 0 _1137_
rlabel metal2 2898 37264 2898 37264 0 _1138_
rlabel metal1 5750 35768 5750 35768 0 _1139_
rlabel metal1 2714 36720 2714 36720 0 _1140_
rlabel metal2 6118 36006 6118 36006 0 _1141_
rlabel metal1 3220 34714 3220 34714 0 _1142_
rlabel metal1 4508 35190 4508 35190 0 _1143_
rlabel metal1 5106 34612 5106 34612 0 _1144_
rlabel metal1 4508 34714 4508 34714 0 _1145_
rlabel metal1 8924 34170 8924 34170 0 _1146_
rlabel metal1 6164 33830 6164 33830 0 _1147_
rlabel metal1 8402 34646 8402 34646 0 _1148_
rlabel metal2 5566 34340 5566 34340 0 _1149_
rlabel metal1 7682 33864 7682 33864 0 _1150_
rlabel metal2 7866 35020 7866 35020 0 _1151_
rlabel metal1 8004 34170 8004 34170 0 _1152_
rlabel metal1 8188 32878 8188 32878 0 _1153_
rlabel metal1 7590 32844 7590 32844 0 _1154_
rlabel metal1 7866 32912 7866 32912 0 _1155_
rlabel metal2 7406 33252 7406 33252 0 _1156_
rlabel metal1 8280 32266 8280 32266 0 _1157_
rlabel metal1 7038 31994 7038 31994 0 _1158_
rlabel metal1 8280 31450 8280 31450 0 _1159_
rlabel metal2 4830 32640 4830 32640 0 _1160_
rlabel metal1 5520 31994 5520 31994 0 _1161_
rlabel metal1 5244 31790 5244 31790 0 _1162_
rlabel metal1 3680 33490 3680 33490 0 _1163_
rlabel metal1 5566 30600 5566 30600 0 _1164_
rlabel metal1 5474 30906 5474 30906 0 _1165_
rlabel metal1 5290 29682 5290 29682 0 _1166_
rlabel metal2 5566 29920 5566 29920 0 _1167_
rlabel metal1 4830 30260 4830 30260 0 _1168_
rlabel metal2 5382 29818 5382 29818 0 _1169_
rlabel metal2 3818 32844 3818 32844 0 _1170_
rlabel metal2 3634 32572 3634 32572 0 _1171_
rlabel metal2 3266 32844 3266 32844 0 _1172_
rlabel metal2 4094 30906 4094 30906 0 _1173_
rlabel metal1 2346 32436 2346 32436 0 _1174_
rlabel metal2 3266 31110 3266 31110 0 _1175_
rlabel metal2 3818 30566 3818 30566 0 _1176_
rlabel metal1 3358 29648 3358 29648 0 _1177_
rlabel metal1 2898 28526 2898 28526 0 _1178_
rlabel metal1 3818 29070 3818 29070 0 _1179_
rlabel metal1 3128 28730 3128 28730 0 _1180_
rlabel metal2 6026 25568 6026 25568 0 _1181_
rlabel metal2 6578 26316 6578 26316 0 _1182_
rlabel metal2 4370 21862 4370 21862 0 _1183_
rlabel metal1 4692 22406 4692 22406 0 _1184_
rlabel metal2 5244 22508 5244 22508 0 _1185_
rlabel metal1 5244 22746 5244 22746 0 _1186_
rlabel metal1 5244 17714 5244 17714 0 _1187_
rlabel metal2 5382 17170 5382 17170 0 _1188_
rlabel metal2 5382 19142 5382 19142 0 _1189_
rlabel metal1 5428 20570 5428 20570 0 _1190_
rlabel metal1 5658 17782 5658 17782 0 _1191_
rlabel metal1 5106 15878 5106 15878 0 _1192_
rlabel metal1 5520 17306 5520 17306 0 _1193_
rlabel metal1 5198 17306 5198 17306 0 _1194_
rlabel metal1 5704 17850 5704 17850 0 _1195_
rlabel metal2 5290 18564 5290 18564 0 _1196_
rlabel metal2 4830 19924 4830 19924 0 _1197_
rlabel metal2 6946 24106 6946 24106 0 _1198_
rlabel metal1 7682 23120 7682 23120 0 _1199_
rlabel metal1 6946 25806 6946 25806 0 _1200_
rlabel metal1 15686 27438 15686 27438 0 _1201_
rlabel metal1 14720 26350 14720 26350 0 _1202_
rlabel metal1 14536 26554 14536 26554 0 _1203_
rlabel metal1 18538 29070 18538 29070 0 _1204_
rlabel metal2 17158 30379 17158 30379 0 _1205_
rlabel metal1 13892 26758 13892 26758 0 _1206_
rlabel metal2 18262 28832 18262 28832 0 _1207_
rlabel metal1 17802 28016 17802 28016 0 _1208_
rlabel metal1 14720 28050 14720 28050 0 _1209_
rlabel metal1 14122 27846 14122 27846 0 _1210_
rlabel metal3 1004 41548 1004 41548 0 clk
rlabel metal2 32246 34442 32246 34442 0 clknet_0_clk
rlabel metal1 17710 20502 17710 20502 0 clknet_2_0__leaf_clk
rlabel metal1 17250 33864 17250 33864 0 clknet_2_1__leaf_clk
rlabel metal3 38111 20740 38111 20740 0 clknet_2_2__leaf_clk
rlabel metal1 40204 36142 40204 36142 0 clknet_2_3__leaf_clk
rlabel metal2 2438 19550 2438 19550 0 clknet_leaf_0_clk
rlabel metal2 19918 42432 19918 42432 0 clknet_leaf_10_clk
rlabel metal1 14674 32878 14674 32878 0 clknet_leaf_11_clk
rlabel metal1 18998 32300 18998 32300 0 clknet_leaf_12_clk
rlabel metal1 21344 26894 21344 26894 0 clknet_leaf_13_clk
rlabel metal1 28474 32266 28474 32266 0 clknet_leaf_14_clk
rlabel metal1 21850 33524 21850 33524 0 clknet_leaf_15_clk
rlabel metal2 28934 39746 28934 39746 0 clknet_leaf_16_clk
rlabel metal2 32430 38114 32430 38114 0 clknet_leaf_17_clk
rlabel metal2 37306 42466 37306 42466 0 clknet_leaf_18_clk
rlabel metal1 40894 37842 40894 37842 0 clknet_leaf_19_clk
rlabel metal2 11546 15504 11546 15504 0 clknet_leaf_1_clk
rlabel metal2 37398 32606 37398 32606 0 clknet_leaf_20_clk
rlabel metal1 38364 24786 38364 24786 0 clknet_leaf_21_clk
rlabel metal2 35282 28322 35282 28322 0 clknet_leaf_22_clk
rlabel metal1 32522 31790 32522 31790 0 clknet_leaf_23_clk
rlabel metal1 27646 20434 27646 20434 0 clknet_leaf_24_clk
rlabel metal2 32798 16796 32798 16796 0 clknet_leaf_25_clk
rlabel metal2 39238 17680 39238 17680 0 clknet_leaf_26_clk
rlabel via1 35282 13821 35282 13821 0 clknet_leaf_27_clk
rlabel metal1 40158 11798 40158 11798 0 clknet_leaf_28_clk
rlabel metal1 32660 7922 32660 7922 0 clknet_leaf_29_clk
rlabel metal2 13846 20434 13846 20434 0 clknet_leaf_2_clk
rlabel metal1 31142 9622 31142 9622 0 clknet_leaf_30_clk
rlabel metal1 26496 12818 26496 12818 0 clknet_leaf_31_clk
rlabel metal2 24886 14688 24886 14688 0 clknet_leaf_32_clk
rlabel metal1 21482 18292 21482 18292 0 clknet_leaf_33_clk
rlabel metal2 13938 14076 13938 14076 0 clknet_leaf_34_clk
rlabel metal1 21114 8398 21114 8398 0 clknet_leaf_35_clk
rlabel metal1 9522 3094 9522 3094 0 clknet_leaf_36_clk
rlabel metal1 7268 6222 7268 6222 0 clknet_leaf_37_clk
rlabel metal2 1426 8160 1426 8160 0 clknet_leaf_38_clk
rlabel metal1 2852 13362 2852 13362 0 clknet_leaf_39_clk
rlabel metal1 19826 22474 19826 22474 0 clknet_leaf_3_clk
rlabel metal1 12581 30158 12581 30158 0 clknet_leaf_4_clk
rlabel metal1 1426 24650 1426 24650 0 clknet_leaf_5_clk
rlabel metal1 4462 32198 4462 32198 0 clknet_leaf_6_clk
rlabel metal1 1426 33524 1426 33524 0 clknet_leaf_7_clk
rlabel metal2 1426 37842 1426 37842 0 clknet_leaf_8_clk
rlabel metal1 13064 38862 13064 38862 0 clknet_leaf_9_clk
rlabel metal1 20700 43418 20700 43418 0 complete
rlabel metal2 17710 44251 17710 44251 0 display_output[0]
rlabel metal2 41906 26945 41906 26945 0 display_output[10]
rlabel metal3 42512 31348 42512 31348 0 display_output[11]
rlabel via2 40618 24565 40618 24565 0 display_output[12]
rlabel metal2 42090 28815 42090 28815 0 display_output[13]
rlabel metal2 40158 25449 40158 25449 0 display_output[14]
rlabel metal2 20286 44251 20286 44251 0 display_output[15]
rlabel metal2 19550 44251 19550 44251 0 display_output[1]
rlabel metal2 22862 44251 22862 44251 0 display_output[2]
rlabel metal2 23414 44251 23414 44251 0 display_output[3]
rlabel metal2 25346 44251 25346 44251 0 display_output[4]
rlabel metal2 42090 27149 42090 27149 0 display_output[5]
rlabel metal2 29210 44251 29210 44251 0 display_output[6]
rlabel via2 41538 27285 41538 27285 0 display_output[7]
rlabel metal2 41722 28169 41722 28169 0 display_output[8]
rlabel metal2 42090 29665 42090 29665 0 display_output[9]
rlabel metal2 7590 25976 7590 25976 0 equal_input
rlabel metal1 13064 36142 13064 36142 0 gencon_inst.ALU_finish
rlabel metal1 15456 33966 15456 33966 0 gencon_inst.ALU_in1\[0\]
rlabel metal2 41446 35190 41446 35190 0 gencon_inst.ALU_in1\[10\]
rlabel via1 41262 34918 41262 34918 0 gencon_inst.ALU_in1\[11\]
rlabel metal2 39606 33762 39606 33762 0 gencon_inst.ALU_in1\[12\]
rlabel metal1 36662 32742 36662 32742 0 gencon_inst.ALU_in1\[13\]
rlabel metal1 33994 31892 33994 31892 0 gencon_inst.ALU_in1\[14\]
rlabel metal1 14076 32878 14076 32878 0 gencon_inst.ALU_in1\[15\]
rlabel metal2 16974 35904 16974 35904 0 gencon_inst.ALU_in1\[1\]
rlabel metal2 20654 33694 20654 33694 0 gencon_inst.ALU_in1\[2\]
rlabel metal1 24012 33354 24012 33354 0 gencon_inst.ALU_in1\[3\]
rlabel metal1 24978 33014 24978 33014 0 gencon_inst.ALU_in1\[4\]
rlabel metal1 26082 34646 26082 34646 0 gencon_inst.ALU_in1\[5\]
rlabel metal1 28244 31926 28244 31926 0 gencon_inst.ALU_in1\[6\]
rlabel metal1 29532 33830 29532 33830 0 gencon_inst.ALU_in1\[7\]
rlabel metal1 31418 34578 31418 34578 0 gencon_inst.ALU_in1\[8\]
rlabel metal2 32154 32164 32154 32164 0 gencon_inst.ALU_in1\[9\]
rlabel metal1 15778 34374 15778 34374 0 gencon_inst.ALU_in2\[0\]
rlabel metal1 40894 34578 40894 34578 0 gencon_inst.ALU_in2\[10\]
rlabel metal1 41262 34986 41262 34986 0 gencon_inst.ALU_in2\[11\]
rlabel metal1 38732 33082 38732 33082 0 gencon_inst.ALU_in2\[12\]
rlabel metal1 36662 33422 36662 33422 0 gencon_inst.ALU_in2\[13\]
rlabel metal1 34040 32742 34040 32742 0 gencon_inst.ALU_in2\[14\]
rlabel metal1 13478 33626 13478 33626 0 gencon_inst.ALU_in2\[15\]
rlabel metal1 16560 35598 16560 35598 0 gencon_inst.ALU_in2\[1\]
rlabel metal1 20286 35122 20286 35122 0 gencon_inst.ALU_in2\[2\]
rlabel metal2 23230 34782 23230 34782 0 gencon_inst.ALU_in2\[3\]
rlabel metal1 23920 34714 23920 34714 0 gencon_inst.ALU_in2\[4\]
rlabel metal1 25852 34102 25852 34102 0 gencon_inst.ALU_in2\[5\]
rlabel metal1 27830 33830 27830 33830 0 gencon_inst.ALU_in2\[6\]
rlabel metal1 29854 32300 29854 32300 0 gencon_inst.ALU_in2\[7\]
rlabel metal1 30866 34646 30866 34646 0 gencon_inst.ALU_in2\[8\]
rlabel metal1 31878 34034 31878 34034 0 gencon_inst.ALU_in2\[9\]
rlabel metal1 16882 42262 16882 42262 0 gencon_inst.ALU_out\[0\]
rlabel metal1 36984 42534 36984 42534 0 gencon_inst.ALU_out\[10\]
rlabel metal1 36616 42194 36616 42194 0 gencon_inst.ALU_out\[11\]
rlabel metal1 35374 39304 35374 39304 0 gencon_inst.ALU_out\[12\]
rlabel metal1 36708 39270 36708 39270 0 gencon_inst.ALU_out\[13\]
rlabel metal1 33948 38182 33948 38182 0 gencon_inst.ALU_out\[14\]
rlabel metal2 17802 36193 17802 36193 0 gencon_inst.ALU_out\[15\]
rlabel metal1 18630 41446 18630 41446 0 gencon_inst.ALU_out\[1\]
rlabel metal1 21712 41990 21712 41990 0 gencon_inst.ALU_out\[2\]
rlabel metal2 21850 39423 21850 39423 0 gencon_inst.ALU_out\[3\]
rlabel metal1 25346 31416 25346 31416 0 gencon_inst.ALU_out\[4\]
rlabel via2 25990 40579 25990 40579 0 gencon_inst.ALU_out\[5\]
rlabel metal1 27876 30770 27876 30770 0 gencon_inst.ALU_out\[6\]
rlabel metal2 36478 27234 36478 27234 0 gencon_inst.ALU_out\[7\]
rlabel metal3 37743 28900 37743 28900 0 gencon_inst.ALU_out\[8\]
rlabel metal1 33258 40426 33258 40426 0 gencon_inst.ALU_out\[9\]
rlabel metal2 13846 33490 13846 33490 0 gencon_inst.addOrSub
rlabel metal1 15134 37808 15134 37808 0 gencon_inst.add_calc.diffSign
rlabel metal1 41952 38930 41952 38930 0 gencon_inst.add_calc.main.GENERATE_ADDER\[10\].thingy.in1
rlabel metal2 40710 37468 40710 37468 0 gencon_inst.add_calc.main.GENERATE_ADDER\[11\].thingy.in1
rlabel metal1 39238 36006 39238 36006 0 gencon_inst.add_calc.main.GENERATE_ADDER\[12\].thingy.in1
rlabel metal1 37122 36720 37122 36720 0 gencon_inst.add_calc.main.GENERATE_ADDER\[13\].thingy.in1
rlabel metal1 34500 36754 34500 36754 0 gencon_inst.add_calc.main.GENERATE_ADDER\[14\].thingy.in1
rlabel metal1 17710 39372 17710 39372 0 gencon_inst.add_calc.main.GENERATE_ADDER\[1\].thingy.in1
rlabel metal1 20148 37774 20148 37774 0 gencon_inst.add_calc.main.GENERATE_ADDER\[2\].thingy.in1
rlabel metal2 21022 37604 21022 37604 0 gencon_inst.add_calc.main.GENERATE_ADDER\[3\].thingy.in1
rlabel metal1 24242 38896 24242 38896 0 gencon_inst.add_calc.main.GENERATE_ADDER\[4\].thingy.in1
rlabel metal1 26041 38250 26041 38250 0 gencon_inst.add_calc.main.GENERATE_ADDER\[5\].thingy.in1
rlabel metal1 28198 37808 28198 37808 0 gencon_inst.add_calc.main.GENERATE_ADDER\[6\].thingy.in1
rlabel metal1 28980 38250 28980 38250 0 gencon_inst.add_calc.main.GENERATE_ADDER\[7\].thingy.in1
rlabel metal1 32430 38386 32430 38386 0 gencon_inst.add_calc.main.GENERATE_ADDER\[8\].thingy.in1
rlabel metal2 31970 37910 31970 37910 0 gencon_inst.add_calc.main.GENERATE_ADDER\[9\].thingy.in1
rlabel metal1 15870 38930 15870 38930 0 gencon_inst.add_calc.main.a0.in1
rlabel metal1 14950 39814 14950 39814 0 gencon_inst.add_calc.main.in2\[0\]
rlabel metal2 42182 40052 42182 40052 0 gencon_inst.add_calc.main.in2\[10\]
rlabel metal1 39928 37230 39928 37230 0 gencon_inst.add_calc.main.in2\[11\]
rlabel metal2 39238 36414 39238 36414 0 gencon_inst.add_calc.main.in2\[12\]
rlabel metal2 36938 36414 36938 36414 0 gencon_inst.add_calc.main.in2\[13\]
rlabel metal1 35696 36142 35696 36142 0 gencon_inst.add_calc.main.in2\[14\]
rlabel metal1 16698 36890 16698 36890 0 gencon_inst.add_calc.main.in2\[1\]
rlabel metal1 20332 36686 20332 36686 0 gencon_inst.add_calc.main.in2\[2\]
rlabel metal1 22954 36006 22954 36006 0 gencon_inst.add_calc.main.in2\[3\]
rlabel metal1 24840 36210 24840 36210 0 gencon_inst.add_calc.main.in2\[4\]
rlabel metal1 26220 35598 26220 35598 0 gencon_inst.add_calc.main.in2\[5\]
rlabel metal1 27002 36108 27002 36108 0 gencon_inst.add_calc.main.in2\[6\]
rlabel metal1 29670 35054 29670 35054 0 gencon_inst.add_calc.main.in2\[7\]
rlabel metal1 29900 37230 29900 37230 0 gencon_inst.add_calc.main.in2\[8\]
rlabel metal1 32982 37230 32982 37230 0 gencon_inst.add_calc.main.in2\[9\]
rlabel metal2 11362 36516 11362 36516 0 gencon_inst.add_calc.next_finish
rlabel metal1 15318 37230 15318 37230 0 gencon_inst.add_calc.sameSignVal
rlabel via1 10994 32963 10994 32963 0 gencon_inst.add_calc.start
rlabel metal1 11569 35802 11569 35802 0 gencon_inst.add_calc.state\[0\]
rlabel metal1 33994 37706 33994 37706 0 gencon_inst.add_calc.state\[1\]
rlabel metal1 36386 36244 36386 36244 0 gencon_inst.add_calc.state\[2\]
rlabel metal1 17020 29138 17020 29138 0 gencon_inst.gencon_state\[0\]
rlabel metal2 16238 28594 16238 28594 0 gencon_inst.gencon_state\[1\]
rlabel metal1 17020 27370 17020 27370 0 gencon_inst.gencon_state\[2\]
rlabel metal2 14950 29138 14950 29138 0 gencon_inst.gencon_state\[3\]
rlabel metal2 15456 26214 15456 26214 0 gencon_inst.key_read
rlabel metal1 9154 21522 9154 21522 0 gencon_inst.keypad_input\[0\]
rlabel metal1 9890 22406 9890 22406 0 gencon_inst.keypad_input\[1\]
rlabel metal2 10534 23324 10534 23324 0 gencon_inst.keypad_input\[2\]
rlabel metal2 10718 24582 10718 24582 0 gencon_inst.keypad_input\[3\]
rlabel metal1 17480 31790 17480 31790 0 gencon_inst.latched_keypad_input\[0\]
rlabel metal2 13294 22848 13294 22848 0 gencon_inst.latched_keypad_input\[1\]
rlabel metal2 13294 23936 13294 23936 0 gencon_inst.latched_keypad_input\[2\]
rlabel metal1 21206 24072 21206 24072 0 gencon_inst.latched_keypad_input\[3\]
rlabel metal2 12926 33286 12926 33286 0 gencon_inst.latched_operator_input\[0\]
rlabel metal1 11638 31790 11638 31790 0 gencon_inst.latched_operator_input\[1\]
rlabel metal1 11086 32334 11086 32334 0 gencon_inst.latched_operator_input\[2\]
rlabel metal1 16468 20026 16468 20026 0 gencon_inst.mult_calc.INn1\[0\]
rlabel metal1 38916 22066 38916 22066 0 gencon_inst.mult_calc.INn1\[10\]
rlabel metal1 40802 20434 40802 20434 0 gencon_inst.mult_calc.INn1\[11\]
rlabel metal2 40802 23324 40802 23324 0 gencon_inst.mult_calc.INn1\[12\]
rlabel metal2 39054 20604 39054 20604 0 gencon_inst.mult_calc.INn1\[13\]
rlabel metal2 35558 20060 35558 20060 0 gencon_inst.mult_calc.INn1\[14\]
rlabel metal1 15134 22950 15134 22950 0 gencon_inst.mult_calc.INn1\[15\]
rlabel metal2 18170 21658 18170 21658 0 gencon_inst.mult_calc.INn1\[1\]
rlabel metal2 21206 21692 21206 21692 0 gencon_inst.mult_calc.INn1\[2\]
rlabel metal1 23230 22066 23230 22066 0 gencon_inst.mult_calc.INn1\[3\]
rlabel metal2 24334 21794 24334 21794 0 gencon_inst.mult_calc.INn1\[4\]
rlabel metal1 27002 21420 27002 21420 0 gencon_inst.mult_calc.INn1\[5\]
rlabel metal1 28566 22066 28566 22066 0 gencon_inst.mult_calc.INn1\[6\]
rlabel metal2 30958 23460 30958 23460 0 gencon_inst.mult_calc.INn1\[7\]
rlabel metal1 32200 22066 32200 22066 0 gencon_inst.mult_calc.INn1\[8\]
rlabel metal2 33534 21828 33534 21828 0 gencon_inst.mult_calc.INn1\[9\]
rlabel metal1 19780 22746 19780 22746 0 gencon_inst.mult_calc.INn2\[0\]
rlabel metal2 35512 19380 35512 19380 0 gencon_inst.mult_calc.INn2\[10\]
rlabel metal1 34914 21454 34914 21454 0 gencon_inst.mult_calc.INn2\[11\]
rlabel metal1 36248 21862 36248 21862 0 gencon_inst.mult_calc.INn2\[12\]
rlabel metal1 35512 20298 35512 20298 0 gencon_inst.mult_calc.INn2\[13\]
rlabel metal1 36064 19142 36064 19142 0 gencon_inst.mult_calc.INn2\[14\]
rlabel metal1 14950 23494 14950 23494 0 gencon_inst.mult_calc.INn2\[15\]
rlabel metal1 19136 19822 19136 19822 0 gencon_inst.mult_calc.INn2\[1\]
rlabel metal2 20700 18394 20700 18394 0 gencon_inst.mult_calc.INn2\[2\]
rlabel metal1 20792 19686 20792 19686 0 gencon_inst.mult_calc.INn2\[3\]
rlabel via3 25691 13668 25691 13668 0 gencon_inst.mult_calc.INn2\[4\]
rlabel metal1 25714 21998 25714 21998 0 gencon_inst.mult_calc.INn2\[5\]
rlabel metal1 25898 14008 25898 14008 0 gencon_inst.mult_calc.INn2\[6\]
rlabel metal2 25714 14212 25714 14212 0 gencon_inst.mult_calc.INn2\[7\]
rlabel metal3 33879 13804 33879 13804 0 gencon_inst.mult_calc.INn2\[8\]
rlabel metal2 34592 19244 34592 19244 0 gencon_inst.mult_calc.INn2\[9\]
rlabel metal2 17342 15844 17342 15844 0 gencon_inst.mult_calc.adderSave\[0\]
rlabel metal1 38088 18258 38088 18258 0 gencon_inst.mult_calc.adderSave\[10\]
rlabel metal1 41078 19482 41078 19482 0 gencon_inst.mult_calc.adderSave\[11\]
rlabel metal2 40066 16456 40066 16456 0 gencon_inst.mult_calc.adderSave\[12\]
rlabel metal1 41492 14042 41492 14042 0 gencon_inst.mult_calc.adderSave\[13\]
rlabel metal2 35466 15164 35466 15164 0 gencon_inst.mult_calc.adderSave\[14\]
rlabel metal1 17986 17204 17986 17204 0 gencon_inst.mult_calc.adderSave\[1\]
rlabel metal2 21482 15504 21482 15504 0 gencon_inst.mult_calc.adderSave\[2\]
rlabel metal1 23920 19278 23920 19278 0 gencon_inst.mult_calc.adderSave\[3\]
rlabel metal2 24978 15198 24978 15198 0 gencon_inst.mult_calc.adderSave\[4\]
rlabel metal1 26404 18190 26404 18190 0 gencon_inst.mult_calc.adderSave\[5\]
rlabel via2 30498 15453 30498 15453 0 gencon_inst.mult_calc.adderSave\[6\]
rlabel metal1 29808 19278 29808 19278 0 gencon_inst.mult_calc.adderSave\[7\]
rlabel metal1 32292 16626 32292 16626 0 gencon_inst.mult_calc.adderSave\[8\]
rlabel metal1 33074 18836 33074 18836 0 gencon_inst.mult_calc.adderSave\[9\]
rlabel metal1 20102 12750 20102 12750 0 gencon_inst.mult_calc.compCount.in2\[0\]
rlabel metal2 34362 13906 34362 13906 0 gencon_inst.mult_calc.compCount.in2\[10\]
rlabel metal1 34776 12682 34776 12682 0 gencon_inst.mult_calc.compCount.in2\[11\]
rlabel metal1 36248 11866 36248 11866 0 gencon_inst.mult_calc.compCount.in2\[12\]
rlabel metal1 37168 14042 37168 14042 0 gencon_inst.mult_calc.compCount.in2\[13\]
rlabel metal1 37076 13158 37076 13158 0 gencon_inst.mult_calc.compCount.in2\[14\]
rlabel metal1 20010 12104 20010 12104 0 gencon_inst.mult_calc.compCount.in2\[1\]
rlabel metal1 21942 12240 21942 12240 0 gencon_inst.mult_calc.compCount.in2\[2\]
rlabel metal1 23138 13498 23138 13498 0 gencon_inst.mult_calc.compCount.in2\[3\]
rlabel metal2 24794 12478 24794 12478 0 gencon_inst.mult_calc.compCount.in2\[4\]
rlabel metal1 26220 12410 26220 12410 0 gencon_inst.mult_calc.compCount.in2\[5\]
rlabel metal1 27140 11662 27140 11662 0 gencon_inst.mult_calc.compCount.in2\[6\]
rlabel metal1 28888 12614 28888 12614 0 gencon_inst.mult_calc.compCount.in2\[7\]
rlabel metal1 30590 11526 30590 11526 0 gencon_inst.mult_calc.compCount.in2\[8\]
rlabel metal1 32476 13362 32476 13362 0 gencon_inst.mult_calc.compCount.in2\[9\]
rlabel metal1 33994 9588 33994 9588 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[10\].thingy.in1
rlabel metal1 34270 9588 34270 9588 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[11\].thingy.in1
rlabel metal2 35558 9350 35558 9350 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[12\].thingy.in1
rlabel metal1 40618 10098 40618 10098 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[13\].thingy.in1
rlabel metal1 38318 11118 38318 11118 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[14\].thingy.in1
rlabel metal1 19228 8602 19228 8602 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.cIn
rlabel metal2 18814 10948 18814 10948 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[1\].thingy.in1
rlabel metal2 21390 11560 21390 11560 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[2\].thingy.in1
rlabel metal2 20930 9350 20930 9350 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[3\].thingy.in1
rlabel metal1 26450 9452 26450 9452 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[4\].thingy.in1
rlabel metal1 26266 9622 26266 9622 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[5\].thingy.in1
rlabel metal1 27002 9588 27002 9588 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[6\].thingy.in1
rlabel metal1 30406 10676 30406 10676 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[7\].thingy.in1
rlabel metal2 31234 8976 31234 8976 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[8\].thingy.in1
rlabel metal1 32154 9146 32154 9146 0 gencon_inst.mult_calc.count.GENERATE_ADDER\[9\].thingy.in1
rlabel metal2 19366 8126 19366 8126 0 gencon_inst.mult_calc.countSave\[0\]
rlabel metal2 33902 10268 33902 10268 0 gencon_inst.mult_calc.countSave\[10\]
rlabel metal1 34638 8058 34638 8058 0 gencon_inst.mult_calc.countSave\[11\]
rlabel metal1 36984 7922 36984 7922 0 gencon_inst.mult_calc.countSave\[12\]
rlabel metal2 39054 9860 39054 9860 0 gencon_inst.mult_calc.countSave\[13\]
rlabel metal2 39514 11628 39514 11628 0 gencon_inst.mult_calc.countSave\[14\]
rlabel metal1 19320 10098 19320 10098 0 gencon_inst.mult_calc.countSave\[1\]
rlabel metal2 21482 11492 21482 11492 0 gencon_inst.mult_calc.countSave\[2\]
rlabel metal1 21252 7310 21252 7310 0 gencon_inst.mult_calc.countSave\[3\]
rlabel metal1 24426 7854 24426 7854 0 gencon_inst.mult_calc.countSave\[4\]
rlabel metal1 25438 9690 25438 9690 0 gencon_inst.mult_calc.countSave\[5\]
rlabel metal1 27508 8058 27508 8058 0 gencon_inst.mult_calc.countSave\[6\]
rlabel metal1 29532 10098 29532 10098 0 gencon_inst.mult_calc.countSave\[7\]
rlabel metal1 30084 7310 30084 7310 0 gencon_inst.mult_calc.countSave\[8\]
rlabel metal1 32062 8398 32062 8398 0 gencon_inst.mult_calc.countSave\[9\]
rlabel metal1 15916 20978 15916 20978 0 gencon_inst.mult_calc.diffSign
rlabel metal1 14812 14586 14812 14586 0 gencon_inst.mult_calc.finish
rlabel metal1 37490 19380 37490 19380 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in1
rlabel metal1 37306 19312 37306 19312 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[10\].thingy.in2
rlabel metal2 42090 20876 42090 20876 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in1
rlabel metal2 42182 19380 42182 19380 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[11\].thingy.in2
rlabel metal1 41860 22066 41860 22066 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in1
rlabel metal2 41814 17408 41814 17408 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[12\].thingy.in2
rlabel metal1 41814 15062 41814 15062 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in1
rlabel metal1 42090 15572 42090 15572 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[13\].thingy.in2
rlabel metal2 36478 17102 36478 17102 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in1
rlabel metal2 36386 16388 36386 16388 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[14\].thingy.in2
rlabel metal1 20286 21420 20286 21420 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in1
rlabel metal2 18078 18020 18078 18020 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[1\].thingy.in2
rlabel metal2 21666 20910 21666 20910 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in1
rlabel metal1 22034 17204 22034 17204 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[2\].thingy.in2
rlabel metal1 23966 18224 23966 18224 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in1
rlabel metal1 24564 18802 24564 18802 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[3\].thingy.in2
rlabel metal1 24334 16116 24334 16116 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in1
rlabel metal1 25070 16592 25070 16592 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[4\].thingy.in2
rlabel metal2 27186 20026 27186 20026 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in1
rlabel metal1 27232 17238 27232 17238 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[5\].thingy.in2
rlabel metal2 28934 21284 28934 21284 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in1
rlabel metal2 27738 17408 27738 17408 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[6\].thingy.in2
rlabel metal1 30544 18326 30544 18326 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in1
rlabel metal2 30682 18802 30682 18802 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[7\].thingy.in2
rlabel metal1 31832 16558 31832 16558 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in1
rlabel metal1 33442 16524 33442 16524 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[8\].thingy.in2
rlabel metal2 34086 20740 34086 20740 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in1
rlabel metal2 33718 17442 33718 17442 0 gencon_inst.mult_calc.main.GENERATE_ADDER\[9\].thingy.in2
rlabel metal1 17802 16524 17802 16524 0 gencon_inst.mult_calc.main.a0.in1
rlabel metal2 19458 15266 19458 15266 0 gencon_inst.mult_calc.main.a0.in2
rlabel metal1 31096 14042 31096 14042 0 gencon_inst.mult_calc.next_finish
rlabel metal1 17204 16218 17204 16218 0 gencon_inst.mult_calc.out\[0\]
rlabel metal1 37582 20502 37582 20502 0 gencon_inst.mult_calc.out\[10\]
rlabel metal1 39054 19856 39054 19856 0 gencon_inst.mult_calc.out\[11\]
rlabel metal1 36800 16762 36800 16762 0 gencon_inst.mult_calc.out\[12\]
rlabel metal1 39008 13294 39008 13294 0 gencon_inst.mult_calc.out\[13\]
rlabel metal1 34270 16218 34270 16218 0 gencon_inst.mult_calc.out\[14\]
rlabel metal2 17066 25500 17066 25500 0 gencon_inst.mult_calc.out\[15\]
rlabel metal1 18032 18734 18032 18734 0 gencon_inst.mult_calc.out\[1\]
rlabel metal1 21344 19278 21344 19278 0 gencon_inst.mult_calc.out\[2\]
rlabel metal1 22678 21114 22678 21114 0 gencon_inst.mult_calc.out\[3\]
rlabel metal1 24012 15470 24012 15470 0 gencon_inst.mult_calc.out\[4\]
rlabel metal1 26542 19482 26542 19482 0 gencon_inst.mult_calc.out\[5\]
rlabel metal1 26818 16218 26818 16218 0 gencon_inst.mult_calc.out\[6\]
rlabel metal1 29486 20570 29486 20570 0 gencon_inst.mult_calc.out\[7\]
rlabel metal1 32522 14280 32522 14280 0 gencon_inst.mult_calc.out\[8\]
rlabel metal1 32338 20570 32338 20570 0 gencon_inst.mult_calc.out\[9\]
rlabel metal1 18538 16660 18538 16660 0 gencon_inst.mult_calc.start
rlabel metal1 16859 13498 16859 13498 0 gencon_inst.mult_calc.state\[0\]
rlabel metal1 29578 13294 29578 13294 0 gencon_inst.mult_calc.state\[2\]
rlabel metal2 18078 12716 18078 12716 0 gencon_inst.mult_calc.state\[3\]
rlabel metal1 32430 15334 32430 15334 0 gencon_inst.mult_calc.state\[4\]
rlabel metal1 14766 27064 14766 27064 0 gencon_inst.next_state\[0\]
rlabel metal1 13409 28594 13409 28594 0 gencon_inst.next_state\[1\]
rlabel metal2 13478 26078 13478 26078 0 gencon_inst.next_state\[2\]
rlabel metal1 12834 29274 12834 29274 0 gencon_inst.next_state\[3\]
rlabel metal1 16606 33082 16606 33082 0 gencon_inst.operand1\[0\]
rlabel metal1 39836 32810 39836 32810 0 gencon_inst.operand1\[10\]
rlabel metal2 38134 30022 38134 30022 0 gencon_inst.operand1\[11\]
rlabel metal2 37030 27472 37030 27472 0 gencon_inst.operand1\[12\]
rlabel metal1 35742 31314 35742 31314 0 gencon_inst.operand1\[13\]
rlabel metal1 34454 27438 34454 27438 0 gencon_inst.operand1\[14\]
rlabel metal2 14398 30940 14398 30940 0 gencon_inst.operand1\[15\]
rlabel metal1 18124 32538 18124 32538 0 gencon_inst.operand1\[1\]
rlabel metal1 21114 32334 21114 32334 0 gencon_inst.operand1\[2\]
rlabel metal1 21758 27404 21758 27404 0 gencon_inst.operand1\[3\]
rlabel metal2 24150 32062 24150 32062 0 gencon_inst.operand1\[4\]
rlabel metal1 25484 30362 25484 30362 0 gencon_inst.operand1\[5\]
rlabel metal1 26266 30260 26266 30260 0 gencon_inst.operand1\[6\]
rlabel metal1 30176 28526 30176 28526 0 gencon_inst.operand1\[7\]
rlabel metal1 31878 27846 31878 27846 0 gencon_inst.operand1\[8\]
rlabel metal2 32522 31076 32522 31076 0 gencon_inst.operand1\[9\]
rlabel metal1 16192 33286 16192 33286 0 gencon_inst.operand2\[0\]
rlabel metal1 38548 33422 38548 33422 0 gencon_inst.operand2\[10\]
rlabel metal1 40296 30566 40296 30566 0 gencon_inst.operand2\[11\]
rlabel metal1 39008 33558 39008 33558 0 gencon_inst.operand2\[12\]
rlabel metal1 36202 33558 36202 33558 0 gencon_inst.operand2\[13\]
rlabel metal2 33074 28390 33074 28390 0 gencon_inst.operand2\[14\]
rlabel metal1 14950 29172 14950 29172 0 gencon_inst.operand2\[15\]
rlabel metal1 18030 34646 18030 34646 0 gencon_inst.operand2\[1\]
rlabel metal1 20516 34578 20516 34578 0 gencon_inst.operand2\[2\]
rlabel metal1 19780 21114 19780 21114 0 gencon_inst.operand2\[3\]
rlabel metal1 23874 33558 23874 33558 0 gencon_inst.operand2\[4\]
rlabel metal1 25668 33490 25668 33490 0 gencon_inst.operand2\[5\]
rlabel metal1 27416 32878 27416 32878 0 gencon_inst.operand2\[6\]
rlabel metal1 30084 27438 30084 27438 0 gencon_inst.operand2\[7\]
rlabel metal1 31234 32198 31234 32198 0 gencon_inst.operand2\[8\]
rlabel metal1 32568 33490 32568 33490 0 gencon_inst.operand2\[9\]
rlabel via2 15226 26435 15226 26435 0 gencon_inst.operator_input\[0\]
rlabel metal1 10396 26962 10396 26962 0 gencon_inst.operator_input\[1\]
rlabel metal1 10166 27914 10166 27914 0 gencon_inst.operator_input\[2\]
rlabel metal2 10258 29376 10258 29376 0 gencon_inst.prev_operator_input\[0\]
rlabel metal1 9568 28662 9568 28662 0 gencon_inst.prev_operator_input\[1\]
rlabel metal1 8372 29002 8372 29002 0 gencon_inst.prev_operator_input\[2\]
rlabel metal1 13018 27404 13018 27404 0 gencon_inst.prev_read_input
rlabel metal1 8234 26350 8234 26350 0 gencon_inst.read_input
rlabel metal1 3795 15470 3795 15470 0 input_ctrl_inst.RowMid\[0\]
rlabel via1 3243 15130 3243 15130 0 input_ctrl_inst.RowMid\[1\]
rlabel metal1 3795 17646 3795 17646 0 input_ctrl_inst.RowMid\[2\]
rlabel metal1 3427 18938 3427 18938 0 input_ctrl_inst.RowMid\[3\]
rlabel metal2 4830 17680 4830 17680 0 input_ctrl_inst.RowSync\[0\]
rlabel metal1 5336 18326 5336 18326 0 input_ctrl_inst.RowSync\[1\]
rlabel metal1 5060 17646 5060 17646 0 input_ctrl_inst.RowSync\[2\]
rlabel metal2 5014 18938 5014 18938 0 input_ctrl_inst.RowSync\[3\]
rlabel metal1 4370 21522 4370 21522 0 input_ctrl_inst.col_index\[0\]
rlabel metal1 9798 12614 9798 12614 0 input_ctrl_inst.col_index\[10\]
rlabel metal1 10350 11118 10350 11118 0 input_ctrl_inst.col_index\[11\]
rlabel metal1 10166 11288 10166 11288 0 input_ctrl_inst.col_index\[12\]
rlabel metal1 11132 9486 11132 9486 0 input_ctrl_inst.col_index\[13\]
rlabel metal1 13432 9690 13432 9690 0 input_ctrl_inst.col_index\[14\]
rlabel metal2 12926 10404 12926 10404 0 input_ctrl_inst.col_index\[15\]
rlabel metal1 5106 9350 5106 9350 0 input_ctrl_inst.col_index\[16\]
rlabel metal1 4094 8568 4094 8568 0 input_ctrl_inst.col_index\[17\]
rlabel metal1 4646 8466 4646 8466 0 input_ctrl_inst.col_index\[18\]
rlabel metal1 4646 8364 4646 8364 0 input_ctrl_inst.col_index\[19\]
rlabel metal1 3266 20400 3266 20400 0 input_ctrl_inst.col_index\[1\]
rlabel metal1 1748 5134 1748 5134 0 input_ctrl_inst.col_index\[20\]
rlabel metal2 4370 5236 4370 5236 0 input_ctrl_inst.col_index\[21\]
rlabel metal2 4830 5134 4830 5134 0 input_ctrl_inst.col_index\[22\]
rlabel metal1 5014 4522 5014 4522 0 input_ctrl_inst.col_index\[23\]
rlabel metal1 7268 7786 7268 7786 0 input_ctrl_inst.col_index\[24\]
rlabel metal2 7406 5134 7406 5134 0 input_ctrl_inst.col_index\[25\]
rlabel metal1 9568 4046 9568 4046 0 input_ctrl_inst.col_index\[26\]
rlabel metal1 9200 5202 9200 5202 0 input_ctrl_inst.col_index\[27\]
rlabel metal1 9522 5202 9522 5202 0 input_ctrl_inst.col_index\[28\]
rlabel metal1 9522 6086 9522 6086 0 input_ctrl_inst.col_index\[29\]
rlabel metal2 3910 10948 3910 10948 0 input_ctrl_inst.col_index\[2\]
rlabel metal1 9798 6324 9798 6324 0 input_ctrl_inst.col_index\[30\]
rlabel metal1 9660 6970 9660 6970 0 input_ctrl_inst.col_index\[31\]
rlabel metal1 5704 17646 5704 17646 0 input_ctrl_inst.col_index\[3\]
rlabel metal2 7130 13770 7130 13770 0 input_ctrl_inst.col_index\[4\]
rlabel metal1 6762 12920 6762 12920 0 input_ctrl_inst.col_index\[5\]
rlabel metal1 7482 13226 7482 13226 0 input_ctrl_inst.col_index\[6\]
rlabel metal1 8280 14450 8280 14450 0 input_ctrl_inst.col_index\[7\]
rlabel metal2 9614 12580 9614 12580 0 input_ctrl_inst.col_index\[8\]
rlabel metal2 10718 13668 10718 13668 0 input_ctrl_inst.col_index\[9\]
rlabel metal1 8142 36142 8142 36142 0 input_ctrl_inst.debounce_cnt\[0\]
rlabel metal1 7038 33422 7038 33422 0 input_ctrl_inst.debounce_cnt\[10\]
rlabel metal2 7130 33082 7130 33082 0 input_ctrl_inst.debounce_cnt\[11\]
rlabel metal1 7268 32402 7268 32402 0 input_ctrl_inst.debounce_cnt\[12\]
rlabel metal1 5566 31858 5566 31858 0 input_ctrl_inst.debounce_cnt\[13\]
rlabel metal2 6118 30532 6118 30532 0 input_ctrl_inst.debounce_cnt\[14\]
rlabel metal1 3496 32742 3496 32742 0 input_ctrl_inst.debounce_cnt\[15\]
rlabel metal1 3450 31110 3450 31110 0 input_ctrl_inst.debounce_cnt\[16\]
rlabel metal2 3174 31076 3174 31076 0 input_ctrl_inst.debounce_cnt\[17\]
rlabel metal1 3680 30362 3680 30362 0 input_ctrl_inst.debounce_cnt\[18\]
rlabel metal1 6762 36788 6762 36788 0 input_ctrl_inst.debounce_cnt\[1\]
rlabel metal1 9062 38386 9062 38386 0 input_ctrl_inst.debounce_cnt\[2\]
rlabel metal2 7038 37604 7038 37604 0 input_ctrl_inst.debounce_cnt\[3\]
rlabel metal1 5014 37196 5014 37196 0 input_ctrl_inst.debounce_cnt\[4\]
rlabel metal2 3450 37808 3450 37808 0 input_ctrl_inst.debounce_cnt\[5\]
rlabel metal2 2070 37570 2070 37570 0 input_ctrl_inst.debounce_cnt\[6\]
rlabel via2 4370 35003 4370 35003 0 input_ctrl_inst.debounce_cnt\[7\]
rlabel metal1 4094 35666 4094 35666 0 input_ctrl_inst.debounce_cnt\[8\]
rlabel metal1 5566 34476 5566 34476 0 input_ctrl_inst.debounce_cnt\[9\]
rlabel metal2 7038 21760 7038 21760 0 input_ctrl_inst.decoded_key\[0\]
rlabel metal1 6302 23052 6302 23052 0 input_ctrl_inst.decoded_key\[1\]
rlabel metal1 7406 20808 7406 20808 0 input_ctrl_inst.decoded_key\[2\]
rlabel metal1 5129 20298 5129 20298 0 input_ctrl_inst.decoded_key\[3\]
rlabel metal2 2070 26044 2070 26044 0 input_ctrl_inst.input_control_state\[0\]
rlabel metal2 2622 25398 2622 25398 0 input_ctrl_inst.input_control_state\[1\]
rlabel metal1 5612 25126 5612 25126 0 input_ctrl_inst.input_control_state\[2\]
rlabel metal1 3404 26418 3404 26418 0 input_ctrl_inst.next_state\[0\]
rlabel metal2 1702 24548 1702 24548 0 input_ctrl_inst.next_state\[1\]
rlabel metal2 4094 25432 4094 25432 0 input_ctrl_inst.next_state\[2\]
rlabel metal1 7544 26418 7544 26418 0 input_ctrl_inst.read_input_flag
rlabel metal2 9430 16864 9430 16864 0 input_ctrl_inst.scan_timer\[0\]
rlabel metal1 14858 16966 14858 16966 0 input_ctrl_inst.scan_timer\[10\]
rlabel metal1 12972 17646 12972 17646 0 input_ctrl_inst.scan_timer\[11\]
rlabel metal1 13018 15946 13018 15946 0 input_ctrl_inst.scan_timer\[12\]
rlabel metal2 14766 15300 14766 15300 0 input_ctrl_inst.scan_timer\[13\]
rlabel metal2 11362 16116 11362 16116 0 input_ctrl_inst.scan_timer\[14\]
rlabel metal2 12926 14620 12926 14620 0 input_ctrl_inst.scan_timer\[15\]
rlabel metal1 12742 12750 12742 12750 0 input_ctrl_inst.scan_timer\[16\]
rlabel metal1 12650 13158 12650 13158 0 input_ctrl_inst.scan_timer\[17\]
rlabel metal1 13846 12852 13846 12852 0 input_ctrl_inst.scan_timer\[18\]
rlabel metal1 14214 12750 14214 12750 0 input_ctrl_inst.scan_timer\[19\]
rlabel metal1 7728 17034 7728 17034 0 input_ctrl_inst.scan_timer\[1\]
rlabel metal1 8004 17170 8004 17170 0 input_ctrl_inst.scan_timer\[2\]
rlabel metal2 8786 18020 8786 18020 0 input_ctrl_inst.scan_timer\[3\]
rlabel metal1 8280 19346 8280 19346 0 input_ctrl_inst.scan_timer\[4\]
rlabel metal1 10166 20026 10166 20026 0 input_ctrl_inst.scan_timer\[5\]
rlabel metal1 10902 18394 10902 18394 0 input_ctrl_inst.scan_timer\[6\]
rlabel via1 10994 18581 10994 18581 0 input_ctrl_inst.scan_timer\[7\]
rlabel metal2 12926 19856 12926 19856 0 input_ctrl_inst.scan_timer\[8\]
rlabel metal2 14122 18020 14122 18020 0 input_ctrl_inst.scan_timer\[9\]
rlabel metal3 866 21148 866 21148 0 input_state_FPGA[0]
rlabel metal1 1472 21658 1472 21658 0 input_state_FPGA[1]
rlabel metal3 751 22508 751 22508 0 input_state_FPGA[2]
rlabel metal3 751 26588 751 26588 0 key_pressed
rlabel via2 42182 3485 42182 3485 0 nRST
rlabel metal2 1794 15674 1794 15674 0 net1
rlabel via3 21045 42908 21045 42908 0 net10
rlabel metal1 37858 21012 37858 21012 0 net100
rlabel metal2 19090 16626 19090 16626 0 net101
rlabel metal1 37812 16082 37812 16082 0 net102
rlabel metal1 17112 14246 17112 14246 0 net103
rlabel metal1 37996 20366 37996 20366 0 net104
rlabel metal1 18906 37808 18906 37808 0 net105
rlabel metal1 36248 36754 36248 36754 0 net106
rlabel metal1 38594 36720 38594 36720 0 net107
rlabel metal1 31786 36856 31786 36856 0 net108
rlabel metal1 19780 37298 19780 37298 0 net109
rlabel metal1 17480 42874 17480 42874 0 net11
rlabel metal1 25576 36686 25576 36686 0 net110
rlabel via1 31970 36227 31970 36227 0 net111
rlabel metal1 41262 38828 41262 38828 0 net112
rlabel metal1 21114 41684 21114 41684 0 net113
rlabel metal2 5382 11084 5382 11084 0 net114
rlabel via2 12558 18717 12558 18717 0 net115
rlabel metal2 14122 20026 14122 20026 0 net116
rlabel metal1 14168 21590 14168 21590 0 net117
rlabel metal1 7275 12138 7275 12138 0 net118
rlabel metal2 9936 12852 9936 12852 0 net119
rlabel metal1 40434 26826 40434 26826 0 net12
rlabel metal2 12466 7310 12466 7310 0 net120
rlabel metal2 2714 13532 2714 13532 0 net121
rlabel metal1 3273 18666 3273 18666 0 net122
rlabel metal2 6670 20332 6670 20332 0 net123
rlabel metal2 17710 18530 17710 18530 0 net124
rlabel metal2 21666 13396 21666 13396 0 net125
rlabel metal2 21298 14569 21298 14569 0 net126
rlabel metal1 21581 20502 21581 20502 0 net127
rlabel metal1 6033 32470 6033 32470 0 net128
rlabel metal1 10909 31382 10909 31382 0 net129
rlabel metal1 41952 32402 41952 32402 0 net13
rlabel metal1 8517 36822 8517 36822 0 net130
rlabel metal1 9115 34986 9115 34986 0 net131
rlabel metal1 15495 32810 15495 32810 0 net132
rlabel metal1 20371 32470 20371 32470 0 net133
rlabel metal1 19373 41514 19373 41514 0 net134
rlabel metal1 16337 41582 16337 41582 0 net135
rlabel metal1 16054 37162 16054 37162 0 net136
rlabel metal1 13064 37230 13064 37230 0 net137
rlabel metal1 27508 7786 27508 7786 0 net138
rlabel metal1 31878 7820 31878 7820 0 net139
rlabel metal1 40802 24718 40802 24718 0 net14
rlabel metal1 23499 20502 23499 20502 0 net140
rlabel metal1 30130 20502 30130 20502 0 net141
rlabel metal2 25070 18870 25070 18870 0 net142
rlabel metal1 33389 7786 33389 7786 0 net143
rlabel metal1 36754 13335 36754 13335 0 net144
rlabel metal1 41959 14314 41959 14314 0 net145
rlabel metal2 41446 18938 41446 18938 0 net146
rlabel metal1 41768 19346 41768 19346 0 net147
rlabel metal1 22777 26282 22777 26282 0 net148
rlabel metal1 31602 36713 31602 36713 0 net149
rlabel metal2 39974 29121 39974 29121 0 net15
rlabel metal1 32614 36720 32614 36720 0 net150
rlabel metal1 32614 36822 32614 36822 0 net151
rlabel metal1 38923 28458 38923 28458 0 net152
rlabel metal1 42044 24786 42044 24786 0 net153
rlabel metal1 36761 42602 36761 42602 0 net154
rlabel metal1 40526 36713 40526 36713 0 net155
rlabel metal1 41814 37842 41814 37842 0 net156
rlabel metal2 41032 17102 41032 17102 0 net157
rlabel metal2 3818 15844 3818 15844 0 net158
rlabel metal1 2861 19346 2861 19346 0 net159
rlabel metal1 40342 25772 40342 25772 0 net16
rlabel metal2 3818 18020 3818 18020 0 net160
rlabel metal1 3404 16762 3404 16762 0 net161
rlabel metal1 12098 26962 12098 26962 0 net162
rlabel metal2 41078 22848 41078 22848 0 net163
rlabel metal1 41262 21114 41262 21114 0 net164
rlabel metal2 13570 11594 13570 11594 0 net165
rlabel via1 15230 12138 15230 12138 0 net166
rlabel metal2 2898 22508 2898 22508 0 net167
rlabel metal1 24886 21012 24886 21012 0 net168
rlabel metal1 2162 24140 2162 24140 0 net169
rlabel metal1 19734 43214 19734 43214 0 net17
rlabel metal1 9660 28526 9660 28526 0 net170
rlabel metal1 18584 21318 18584 21318 0 net171
rlabel metal1 21528 21318 21528 21318 0 net172
rlabel metal1 28014 21862 28014 21862 0 net173
rlabel metal2 31326 21760 31326 21760 0 net174
rlabel metal2 20838 21114 20838 21114 0 net175
rlabel metal1 22770 21998 22770 21998 0 net176
rlabel metal1 23506 22678 23506 22678 0 net177
rlabel metal1 37950 21862 37950 21862 0 net178
rlabel metal1 18906 20842 18906 20842 0 net179
rlabel metal2 19826 42398 19826 42398 0 net18
rlabel metal2 9338 29818 9338 29818 0 net180
rlabel metal1 40250 20502 40250 20502 0 net181
rlabel metal1 27508 20570 27508 20570 0 net182
rlabel metal1 33166 21862 33166 21862 0 net183
rlabel via1 30038 22073 30038 22073 0 net184
rlabel metal2 11454 23902 11454 23902 0 net185
rlabel metal2 8694 28866 8694 28866 0 net186
rlabel metal1 25622 20842 25622 20842 0 net187
rlabel metal2 31970 21318 31970 21318 0 net188
rlabel metal1 28336 21522 28336 21522 0 net189
rlabel metal2 22770 42058 22770 42058 0 net19
rlabel metal1 12788 13906 12788 13906 0 net190
rlabel metal2 13754 14076 13754 14076 0 net191
rlabel metal2 41538 20706 41538 20706 0 net192
rlabel metal2 17158 18836 17158 18836 0 net193
rlabel metal1 38318 20910 38318 20910 0 net194
rlabel metal1 33396 19822 33396 19822 0 net195
rlabel metal1 34868 19686 34868 19686 0 net196
rlabel metal1 24104 33626 24104 33626 0 net197
rlabel metal1 13386 24208 13386 24208 0 net198
rlabel metal1 18492 19686 18492 19686 0 net199
rlabel metal1 1840 14994 1840 14994 0 net2
rlabel metal1 23138 29648 23138 29648 0 net20
rlabel metal1 27600 20026 27600 20026 0 net200
rlabel metal1 30038 21658 30038 21658 0 net201
rlabel metal1 40480 33558 40480 33558 0 net202
rlabel metal1 17112 16762 17112 16762 0 net203
rlabel metal1 25806 33626 25806 33626 0 net204
rlabel metal1 34178 31450 34178 31450 0 net205
rlabel metal2 40434 33728 40434 33728 0 net206
rlabel metal2 38870 33184 38870 33184 0 net207
rlabel metal1 33810 32402 33810 32402 0 net208
rlabel metal2 19182 20128 19182 20128 0 net209
rlabel metal1 25852 43282 25852 43282 0 net21
rlabel metal1 19775 19822 19775 19822 0 net210
rlabel metal1 22494 34578 22494 34578 0 net211
rlabel metal1 15686 33830 15686 33830 0 net212
rlabel metal2 20654 34816 20654 34816 0 net213
rlabel metal1 30498 32878 30498 32878 0 net214
rlabel metal1 35834 17306 35834 17306 0 net215
rlabel metal2 11178 10234 11178 10234 0 net216
rlabel metal2 16054 35088 16054 35088 0 net217
rlabel metal1 36110 33490 36110 33490 0 net218
rlabel metal1 24150 32538 24150 32538 0 net219
rlabel metal2 28934 28101 28934 28101 0 net22
rlabel metal2 32614 33728 32614 33728 0 net220
rlabel metal1 20654 33490 20654 33490 0 net221
rlabel metal1 19304 33898 19304 33898 0 net222
rlabel metal1 26818 33014 26818 33014 0 net223
rlabel metal2 38318 32028 38318 32028 0 net224
rlabel metal2 28842 30804 28842 30804 0 net225
rlabel metal1 26220 31450 26220 31450 0 net226
rlabel metal1 16376 21862 16376 21862 0 net227
rlabel metal1 22862 32878 22862 32878 0 net228
rlabel metal1 29026 31926 29026 31926 0 net229
rlabel metal1 29302 42670 29302 42670 0 net23
rlabel metal2 25714 32300 25714 32300 0 net230
rlabel metal2 16146 33728 16146 33728 0 net231
rlabel metal1 36110 31790 36110 31790 0 net232
rlabel metal1 41124 32742 41124 32742 0 net233
rlabel metal1 41492 23290 41492 23290 0 net234
rlabel metal1 16376 21998 16376 21998 0 net235
rlabel metal1 14536 17714 14536 17714 0 net236
rlabel metal2 15410 17340 15410 17340 0 net237
rlabel metal2 31050 31076 31050 31076 0 net238
rlabel metal1 32706 31450 32706 31450 0 net239
rlabel metal1 41124 27438 41124 27438 0 net24
rlabel metal1 32200 30906 32200 30906 0 net240
rlabel metal2 17618 34272 17618 34272 0 net241
rlabel metal1 15640 23290 15640 23290 0 net242
rlabel metal2 41538 25772 41538 25772 0 net243
rlabel metal1 19412 10030 19412 10030 0 net244
rlabel metal1 21781 7378 21781 7378 0 net245
rlabel metal2 22402 9180 22402 9180 0 net246
rlabel metal1 10810 31858 10810 31858 0 net247
rlabel metal1 30406 31314 30406 31314 0 net248
rlabel metal1 38456 18394 38456 18394 0 net249
rlabel metal2 39790 28220 39790 28220 0 net25
rlabel metal1 39422 14926 39422 14926 0 net250
rlabel metal1 13386 32878 13386 32878 0 net251
rlabel metal2 29210 7956 29210 7956 0 net252
rlabel metal2 29854 8092 29854 8092 0 net253
rlabel metal1 34316 8602 34316 8602 0 net254
rlabel metal1 32384 8262 32384 8262 0 net255
rlabel metal1 31832 9010 31832 9010 0 net256
rlabel metal1 21068 11526 21068 11526 0 net257
rlabel metal1 25024 8466 25024 8466 0 net258
rlabel metal1 34040 8942 34040 8942 0 net259
rlabel metal1 40802 30260 40802 30260 0 net26
rlabel metal2 37858 8738 37858 8738 0 net260
rlabel metal1 37168 8942 37168 8942 0 net261
rlabel metal1 38916 11322 38916 11322 0 net262
rlabel metal1 40066 11662 40066 11662 0 net263
rlabel metal1 12098 12818 12098 12818 0 net264
rlabel metal1 33028 10030 33028 10030 0 net265
rlabel metal2 10074 35870 10074 35870 0 net266
rlabel metal1 39238 31926 39238 31926 0 net267
rlabel metal1 38180 10098 38180 10098 0 net268
rlabel metal1 29210 10166 29210 10166 0 net269
rlabel metal1 1610 21114 1610 21114 0 net27
rlabel metal1 11638 22950 11638 22950 0 net270
rlabel metal1 19596 13906 19596 13906 0 net271
rlabel metal1 18906 12750 18906 12750 0 net272
rlabel metal1 27462 8534 27462 8534 0 net273
rlabel metal1 25438 10642 25438 10642 0 net274
rlabel metal1 37720 10642 37720 10642 0 net275
rlabel metal1 29302 10608 29302 10608 0 net276
rlabel metal1 13110 34170 13110 34170 0 net277
rlabel metal1 11260 32878 11260 32878 0 net278
rlabel metal2 36754 16864 36754 16864 0 net279
rlabel metal2 1426 21692 1426 21692 0 net28
rlabel metal1 35558 18938 35558 18938 0 net280
rlabel metal2 7130 37808 7130 37808 0 net281
rlabel metal2 8602 21794 8602 21794 0 net282
rlabel metal1 10626 36550 10626 36550 0 net283
rlabel metal2 11086 23494 11086 23494 0 net284
rlabel metal2 26174 17340 26174 17340 0 net285
rlabel metal1 40986 15504 40986 15504 0 net286
rlabel metal2 40710 14620 40710 14620 0 net287
rlabel metal1 36248 14586 36248 14586 0 net288
rlabel metal2 29946 18496 29946 18496 0 net289
rlabel metal2 1426 22916 1426 22916 0 net29
rlabel metal2 30130 18462 30130 18462 0 net290
rlabel metal2 41078 39712 41078 39712 0 net291
rlabel metal1 40802 16150 40802 16150 0 net292
rlabel metal1 40756 16218 40756 16218 0 net293
rlabel metal1 26266 8432 26266 8432 0 net294
rlabel metal1 10580 32198 10580 32198 0 net295
rlabel metal1 29026 19482 29026 19482 0 net296
rlabel metal1 34454 36074 34454 36074 0 net297
rlabel metal2 38778 16932 38778 16932 0 net298
rlabel metal1 21666 10642 21666 10642 0 net299
rlabel metal1 1702 17306 1702 17306 0 net3
rlabel metal1 1748 26962 1748 26962 0 net30
rlabel metal2 23690 18428 23690 18428 0 net300
rlabel metal2 22586 18530 22586 18530 0 net301
rlabel metal2 33534 16626 33534 16626 0 net302
rlabel metal1 17664 16082 17664 16082 0 net303
rlabel metal1 19734 8058 19734 8058 0 net304
rlabel metal2 32522 18428 32522 18428 0 net305
rlabel metal2 25990 16762 25990 16762 0 net306
rlabel metal2 17710 22780 17710 22780 0 net307
rlabel metal1 41492 18326 41492 18326 0 net308
rlabel metal1 40894 18802 40894 18802 0 net309
rlabel metal1 36110 41616 36110 41616 0 net31
rlabel metal1 5980 15130 5980 15130 0 net310
rlabel metal1 10350 34986 10350 34986 0 net311
rlabel via2 24978 21845 24978 21845 0 net312
rlabel metal1 26404 22066 26404 22066 0 net313
rlabel metal1 39100 13226 39100 13226 0 net314
rlabel metal1 40250 36074 40250 36074 0 net315
rlabel metal1 34914 15062 34914 15062 0 net316
rlabel metal2 35466 15844 35466 15844 0 net317
rlabel metal1 34454 21318 34454 21318 0 net318
rlabel metal1 36120 22610 36120 22610 0 net319
rlabel metal2 35374 40324 35374 40324 0 net32
rlabel metal1 38410 19482 38410 19482 0 net320
rlabel metal1 38594 18802 38594 18802 0 net321
rlabel metal2 14582 36652 14582 36652 0 net322
rlabel metal1 19826 36142 19826 36142 0 net323
rlabel metal1 23966 35802 23966 35802 0 net324
rlabel metal1 38548 34986 38548 34986 0 net325
rlabel metal1 32016 36074 32016 36074 0 net326
rlabel metal2 13202 18428 13202 18428 0 net327
rlabel metal1 25300 12818 25300 12818 0 net328
rlabel metal2 7038 26044 7038 26044 0 net329
rlabel metal2 2714 6528 2714 6528 0 net33
rlabel metal2 17894 36890 17894 36890 0 net330
rlabel metal1 33718 36074 33718 36074 0 net331
rlabel metal1 20976 23494 20976 23494 0 net332
rlabel metal1 27738 36822 27738 36822 0 net333
rlabel metal1 13800 15470 13800 15470 0 net334
rlabel metal1 35604 11118 35604 11118 0 net335
rlabel metal2 34822 11934 34822 11934 0 net336
rlabel metal1 29716 35802 29716 35802 0 net337
rlabel metal1 18768 11866 18768 11866 0 net338
rlabel metal1 36370 34034 36370 34034 0 net339
rlabel metal1 16100 31994 16100 31994 0 net34
rlabel metal1 36156 21522 36156 21522 0 net340
rlabel metal1 27462 35802 27462 35802 0 net341
rlabel metal2 18906 18428 18906 18428 0 net342
rlabel metal1 26634 23494 26634 23494 0 net343
rlabel metal1 30682 37978 30682 37978 0 net344
rlabel metal1 29072 34986 29072 34986 0 net345
rlabel metal1 16422 36142 16422 36142 0 net346
rlabel metal1 22218 35598 22218 35598 0 net347
rlabel metal1 25300 35054 25300 35054 0 net348
rlabel metal1 21068 15062 21068 15062 0 net349
rlabel metal1 34868 31178 34868 31178 0 net35
rlabel metal2 20746 14620 20746 14620 0 net350
rlabel metal1 10074 9588 10074 9588 0 net351
rlabel metal1 21942 37842 21942 37842 0 net352
rlabel metal2 30682 15538 30682 15538 0 net353
rlabel metal1 29210 15062 29210 15062 0 net354
rlabel metal1 24978 13974 24978 13974 0 net355
rlabel metal1 24840 14586 24840 14586 0 net356
rlabel metal1 36156 35666 36156 35666 0 net357
rlabel metal1 38548 35666 38548 35666 0 net358
rlabel metal1 32706 15674 32706 15674 0 net359
rlabel metal1 6302 38420 6302 38420 0 net36
rlabel metal2 31510 15640 31510 15640 0 net360
rlabel metal2 32108 21556 32108 21556 0 net361
rlabel metal1 32568 12818 32568 12818 0 net362
rlabel metal1 21436 12818 21436 12818 0 net363
rlabel metal2 8234 20060 8234 20060 0 net364
rlabel metal1 25530 36754 25530 36754 0 net365
rlabel metal2 19642 37434 19642 37434 0 net366
rlabel metal1 23230 36890 23230 36890 0 net367
rlabel metal1 13248 36006 13248 36006 0 net368
rlabel metal2 27186 11934 27186 11934 0 net369
rlabel via1 7511 37842 7511 37842 0 net37
rlabel metal1 28888 35802 28888 35802 0 net370
rlabel metal2 10534 12036 10534 12036 0 net371
rlabel metal2 8418 13498 8418 13498 0 net372
rlabel metal2 12742 30430 12742 30430 0 net373
rlabel metal2 6946 16388 6946 16388 0 net374
rlabel metal2 34914 15198 34914 15198 0 net375
rlabel metal1 13524 19346 13524 19346 0 net376
rlabel metal1 40158 19856 40158 19856 0 net377
rlabel metal2 24978 21148 24978 21148 0 net378
rlabel metal1 28336 12138 28336 12138 0 net379
rlabel metal1 5635 35666 5635 35666 0 net38
rlabel metal2 27462 13022 27462 13022 0 net380
rlabel metal2 40894 38522 40894 38522 0 net381
rlabel metal2 31786 12410 31786 12410 0 net382
rlabel metal1 28198 16218 28198 16218 0 net383
rlabel metal1 40986 38250 40986 38250 0 net384
rlabel metal1 32752 12954 32752 12954 0 net385
rlabel metal2 24058 13056 24058 13056 0 net386
rlabel metal2 3174 37196 3174 37196 0 net387
rlabel metal1 23046 19482 23046 19482 0 net388
rlabel metal1 22448 13906 22448 13906 0 net389
rlabel metal1 17480 20366 17480 20366 0 net39
rlabel metal1 36294 14382 36294 14382 0 net390
rlabel metal1 37582 18394 37582 18394 0 net391
rlabel metal1 7314 13974 7314 13974 0 net392
rlabel metal2 13202 16252 13202 16252 0 net393
rlabel metal2 28934 23290 28934 23290 0 net394
rlabel metal1 24334 15402 24334 15402 0 net395
rlabel metal2 20562 17408 20562 17408 0 net396
rlabel metal1 19734 15674 19734 15674 0 net397
rlabel metal2 33442 14178 33442 14178 0 net398
rlabel metal1 18860 18326 18860 18326 0 net399
rlabel metal1 1702 18394 1702 18394 0 net4
rlabel metal1 34086 21624 34086 21624 0 net40
rlabel metal1 32476 18326 32476 18326 0 net400
rlabel metal1 8786 25942 8786 25942 0 net401
rlabel metal1 11086 15538 11086 15538 0 net402
rlabel metal2 34270 14144 34270 14144 0 net403
rlabel metal1 33028 16422 33028 16422 0 net404
rlabel metal2 5290 9724 5290 9724 0 net405
rlabel metal1 16146 13838 16146 13838 0 net406
rlabel via2 5658 35581 5658 35581 0 net407
rlabel metal2 3634 8636 3634 8636 0 net408
rlabel via1 19181 32402 19181 32402 0 net409
rlabel metal1 39560 23154 39560 23154 0 net41
rlabel metal1 14766 38318 14766 38318 0 net410
rlabel metal1 8970 3570 8970 3570 0 net411
rlabel metal1 37076 13498 37076 13498 0 net412
rlabel metal1 8188 25942 8188 25942 0 net413
rlabel metal1 31832 37162 31832 37162 0 net414
rlabel metal1 2898 31246 2898 31246 0 net415
rlabel metal2 10534 3706 10534 3706 0 net416
rlabel metal1 15226 25228 15226 25228 0 net417
rlabel metal1 10258 20468 10258 20468 0 net418
rlabel metal1 14766 30906 14766 30906 0 net419
rlabel metal1 33442 20944 33442 20944 0 net42
rlabel metal2 11730 10064 11730 10064 0 net420
rlabel metal2 17894 17612 17894 17612 0 net421
rlabel metal2 5382 4624 5382 4624 0 net422
rlabel metal1 7866 33490 7866 33490 0 net423
rlabel metal2 10258 12410 10258 12410 0 net424
rlabel metal1 7636 13906 7636 13906 0 net425
rlabel metal1 15410 13906 15410 13906 0 net426
rlabel metal1 8096 31314 8096 31314 0 net427
rlabel metal2 14582 32640 14582 32640 0 net428
rlabel metal1 3266 37842 3266 37842 0 net429
rlabel metal1 20746 31280 20746 31280 0 net43
rlabel metal1 13248 12818 13248 12818 0 net430
rlabel metal1 20056 28050 20056 28050 0 net431
rlabel metal1 14352 39406 14352 39406 0 net432
rlabel metal2 6854 13124 6854 13124 0 net433
rlabel metal2 9798 6154 9798 6154 0 net434
rlabel metal1 8878 14382 8878 14382 0 net435
rlabel metal1 25530 26418 25530 26418 0 net436
rlabel metal1 7774 37842 7774 37842 0 net437
rlabel metal1 34270 37978 34270 37978 0 net438
rlabel metal2 5934 34204 5934 34204 0 net439
rlabel metal1 33718 29648 33718 29648 0 net44
rlabel metal1 8786 4080 8786 4080 0 net440
rlabel metal1 16330 41106 16330 41106 0 net441
rlabel metal1 21344 41582 21344 41582 0 net442
rlabel metal1 37812 39066 37812 39066 0 net443
rlabel metal1 32568 30226 32568 30226 0 net444
rlabel metal1 14260 34714 14260 34714 0 net445
rlabel metal1 14490 24106 14490 24106 0 net446
rlabel metal1 13754 32742 13754 32742 0 net447
rlabel metal1 19642 42568 19642 42568 0 net45
rlabel metal2 39054 25296 39054 25296 0 net46
rlabel metal1 16514 26486 16514 26486 0 net47
rlabel metal2 27186 26112 27186 26112 0 net48
rlabel metal1 20976 25874 20976 25874 0 net49
rlabel metal2 41906 7106 41906 7106 0 net5
rlabel via1 32627 24854 32627 24854 0 net50
rlabel metal1 16744 31790 16744 31790 0 net51
rlabel metal1 34086 28118 34086 28118 0 net52
rlabel metal1 4968 3026 4968 3026 0 net53
rlabel metal2 11270 6732 11270 6732 0 net54
rlabel metal1 21988 25262 21988 25262 0 net55
rlabel metal1 36708 25874 36708 25874 0 net56
rlabel metal2 32338 27166 32338 27166 0 net57
rlabel metal2 39238 29716 39238 29716 0 net58
rlabel metal1 23552 33422 23552 33422 0 net59
rlabel metal1 10258 2414 10258 2414 0 net6
rlabel metal1 25760 33422 25760 33422 0 net60
rlabel metal2 36018 32640 36018 32640 0 net61
rlabel metal1 38410 31892 38410 31892 0 net62
rlabel metal1 14950 20434 14950 20434 0 net63
rlabel metal2 25346 23970 25346 23970 0 net64
rlabel metal1 18906 32300 18906 32300 0 net65
rlabel metal1 39330 30158 39330 30158 0 net66
rlabel metal1 20010 35156 20010 35156 0 net67
rlabel metal1 36846 34034 36846 34034 0 net68
rlabel metal1 39928 33422 39928 33422 0 net69
rlabel metal1 1748 12410 1748 12410 0 net7
rlabel metal2 38962 34850 38962 34850 0 net70
rlabel metal1 18147 31790 18147 31790 0 net71
rlabel via2 22034 41565 22034 41565 0 net72
rlabel metal1 39422 29614 39422 29614 0 net73
rlabel metal1 39974 31280 39974 31280 0 net74
rlabel metal1 20654 30056 20654 30056 0 net75
rlabel metal2 14996 27540 14996 27540 0 net76
rlabel metal1 38180 26894 38180 26894 0 net77
rlabel metal1 17802 12818 17802 12818 0 net78
rlabel metal1 19826 16116 19826 16116 0 net79
rlabel metal1 1748 11118 1748 11118 0 net8
rlabel metal1 41630 18224 41630 18224 0 net80
rlabel metal2 19918 15708 19918 15708 0 net81
rlabel metal1 3496 24922 3496 24922 0 net82
rlabel metal2 6118 20196 6118 20196 0 net83
rlabel metal1 32246 42092 32246 42092 0 net84
rlabel metal2 36110 39780 36110 39780 0 net85
rlabel metal1 17434 12852 17434 12852 0 net86
rlabel metal2 37490 10506 37490 10506 0 net87
rlabel metal1 18998 9928 18998 9928 0 net88
rlabel metal1 28014 16048 28014 16048 0 net89
rlabel metal1 1748 11730 1748 11730 0 net9
rlabel metal1 37490 17578 37490 17578 0 net90
rlabel metal2 32154 16643 32154 16643 0 net91
rlabel metal2 2714 23868 2714 23868 0 net92
rlabel metal1 19458 8874 19458 8874 0 net93
rlabel metal2 18998 17187 18998 17187 0 net94
rlabel metal2 41354 19142 41354 19142 0 net95
rlabel metal2 29210 13991 29210 13991 0 net96
rlabel metal1 21022 20910 21022 20910 0 net97
rlabel metal1 27416 20366 27416 20366 0 net98
rlabel metal1 36754 14450 36754 14450 0 net99
<< properties >>
string FIXED_BBOX 0 0 43643 45787
<< end >>
