* NGSPICE file created from pwm_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt pwm_wrapper CLK VGND VPWR addr[0] addr[10] addr[11] addr[12] addr[13] addr[14]
+ addr[15] addr[16] addr[17] addr[18] addr[19] addr[1] addr[20] addr[21] addr[22]
+ addr[23] addr[24] addr[25] addr[26] addr[27] addr[28] addr[29] addr[2] addr[30]
+ addr[31] addr[3] addr[4] addr[5] addr[6] addr[7] addr[8] addr[9] error nRST pwm_out[0]
+ pwm_out[1] rdata[0] rdata[10] rdata[11] rdata[12] rdata[13] rdata[14] rdata[15]
+ rdata[16] rdata[17] rdata[18] rdata[19] rdata[1] rdata[20] rdata[21] rdata[22] rdata[23]
+ rdata[24] rdata[25] rdata[26] rdata[27] rdata[28] rdata[29] rdata[2] rdata[30] rdata[31]
+ rdata[3] rdata[4] rdata[5] rdata[6] rdata[7] rdata[8] rdata[9] ren request_stall
+ strobe[0] strobe[1] strobe[2] strobe[3] wdata[0] wdata[10] wdata[11] wdata[12] wdata[13]
+ wdata[14] wdata[15] wdata[16] wdata[17] wdata[18] wdata[19] wdata[1] wdata[20] wdata[21]
+ wdata[22] wdata[23] wdata[24] wdata[25] wdata[26] wdata[27] wdata[28] wdata[29]
+ wdata[2] wdata[30] wdata[31] wdata[3] wdata[4] wdata[5] wdata[6] wdata[7] wdata[8]
+ wdata[9] wen
XFILLER_67_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3155_ _1716_ _0536_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2106_ net251 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] net106 VGND
+ VGND VPWR VPWR _0023_ sky130_fd_sc_hd__mux2_1
X_3086_ net121 _0667_ _0670_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] VGND VGND
+ VPWR VPWR _0671_ sky130_fd_sc_hd__a22oi_1
X_2037_ _1510_ _1513_ _1529_ _1511_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout162_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3988_ clknet_leaf_3_CLK _0180_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_2939_ _0522_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__nand2_1
XFILLER_89_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2304__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3196__A _1656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_6_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3911_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\] net133
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] sky130_fd_sc_hd__dfrtp_4
X_3842_ clknet_leaf_24_CLK _0068_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2214__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3773_ clknet_leaf_21_CLK _0000_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__1924__A_N net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2724_ _1661_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\]
+ _1699_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a22o_1
X_2655_ _1648_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\] VGND VGND VPWR
+ VPWR _0275_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_74_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2586_ net70 _1800_ _1801_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__or3_1
XANTENNA__3553__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout138 net139 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout116 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] VGND VGND VPWR VPWR net116
+ sky130_fd_sc_hd__buf_2
Xfanout105 _1574_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_2
Xfanout127 net128 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_4
Xfanout149 net150 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
XFILLER_74_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3207_ _0515_ _0516_ _0514_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__a21o_1
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3138_ net108 _0721_ _0722_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] VGND VGND
+ VPWR VPWR _0723_ sky130_fd_sc_hd__o22ai_1
XANTENNA__2456__Y _1682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3069_ net118 _0651_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__a21o_1
XFILLER_63_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout78_X net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3407__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2440_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] VGND VGND VPWR VPWR
+ _1666_ sky130_fd_sc_hd__inv_2
XFILLER_96_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2371_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable net34 _1599_ VGND VGND
+ VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_96_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4041_ clknet_leaf_32_CLK _0233_ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_37_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2209__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3825_ clknet_leaf_9_CLK _0051_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3756_ clknet_leaf_18_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[16\]
+ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] sky130_fd_sc_hd__dfrtp_4
X_2707_ _1667_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\]
+ _1674_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a22o_1
X_3687_ _1160_ _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__nand2_1
XANTENNA__3564__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2638_ net112 _1835_ _1837_ net70 VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__a211o_1
XFILLER_99_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2569_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] _1787_ net74 VGND VGND VPWR
+ VPWR _1790_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3800__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3474__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input55_A wdata[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1940_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] _1428_ _1432_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\]
+ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__a22o_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ _1362_ _1363_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__and2_1
X_3610_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__nand2_1
X_3541_ _1612_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\] VGND VGND VPWR
+ VPWR _1125_ sky130_fd_sc_hd__nor2_1
XANTENNA__3384__A _0889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3472_ _1053_ _1054_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2423_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] VGND VGND VPWR VPWR _1649_
+ sky130_fd_sc_hd__inv_2
X_2354_ net212 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] net94 VGND
+ VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2285_ net287 net44 net82 VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
X_4024_ clknet_leaf_6_CLK _0216_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3808_ clknet_leaf_21_CLK _0034_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout128_X net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3739_ _1317_ _1318_ _1625_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2294__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3915__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2312__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_X net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2070_ _1551_ _1562_ _1552_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_6_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2285__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2972_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ _0555_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__a211o_1
X_1923_ _1412_ _1415_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_26_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1854_ _1101_ _1346_ _1100_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__a21o_1
XANTENNA__2222__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3524_ _1099_ _1106_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__a21o_1
XFILLER_89_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3455_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _1700_ _0979_ VGND VGND VPWR
+ VPWR _1040_ sky130_fd_sc_hd__or3_1
X_2406_ net115 VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__inv_2
X_3386_ _0695_ _0720_ _0970_ myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND VGND
+ VPWR VPWR _0971_ sky130_fd_sc_hd__o31ai_1
XFILLER_97_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2458__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2337_ net213 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\] net93 VGND
+ VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2268_ net204 net56 net81 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
X_4007_ clknet_leaf_32_CLK _0199_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2276__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2199_ net305 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\] net101 VGND
+ VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
XFILLER_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2921__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2132__S net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold41 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[19\] VGND VGND VPWR VPWR net244
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[43\] VGND VGND VPWR VPWR net233
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[54\] VGND VGND VPWR VPWR net277
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[22\] VGND VGND VPWR VPWR net255
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold63 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[43\] VGND VGND VPWR VPWR net266
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[61\] VGND VGND VPWR VPWR net299
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input18_A addr[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2267__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold85 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[0\] VGND VGND VPWR VPWR net288
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2307__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3240_ _1698_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _0825_ sky130_fd_sc_hd__nor2_1
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3171_ _0655_ _0754_ _0755_ _0646_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a31o_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2122_ _1579_ _1581_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__nor2_1
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2258__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2053_ _1649_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] _1544_ _1545_
+ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_65_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2217__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2955_ _0528_ _0529_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nor2_1
X_1906_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1394_ _1395_ _1398_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__a32o_1
X_2886_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3507_ _1088_ _1090_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_9_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3438_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _1712_ VGND VGND VPWR VPWR _1023_
+ sky130_fd_sc_hd__and2_1
X_3369_ _0848_ _0852_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nand2_1
XFILLER_85_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2249__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2724__A2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3482__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ _0351_ _0353_ _0355_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__and4_1
X_2671_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[14\]
+ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3223_ _0480_ _0807_ _0806_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__a21o_1
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3154_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__inv_2
X_2105_ net304 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] net106 VGND
+ VGND VPWR VPWR _0022_ sky130_fd_sc_hd__mux2_1
X_3085_ _0668_ _0669_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nand2_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2036_ _1624_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\]
+ _1623_ _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__o221a_1
XANTENNA__2651__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout155_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3987_ clknet_leaf_3_CLK _0179_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_2938_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or2_1
Xclkbuf_2_2__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_2__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_2869_ _1677_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[18\] _0431_ _0452_
+ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__o2111a_1
XANTENNA__1914__B1 _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3803__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3759__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3477__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2320__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input40_X net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2881__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3910_ clknet_leaf_30_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[6\] net133
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_32_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3841_ clknet_leaf_23_CLK _0067_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3772_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag_c net167
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag sky130_fd_sc_hd__dfrtp_2
X_2723_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\]
+ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__nand2_1
X_2654_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] _1838_ VGND VGND VPWR
+ VPWR _0274_ sky130_fd_sc_hd__or2_1
X_2585_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] _1795_ VGND VGND VPWR VPWR _1801_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_74_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout117 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] VGND VGND VPWR VPWR net117
+ sky130_fd_sc_hd__buf_2
Xfanout128 net134 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_4
Xfanout106 _1574_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
Xfanout139 net169 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_2
X_3206_ _1661_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] _0790_ VGND
+ VGND VPWR VPWR _0791_ sky130_fd_sc_hd__o21a_1
XANTENNA__2466__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3137_ _0514_ _0551_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3068_ net119 _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout158_X net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2019_ net116 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] VGND VGND VPWR
+ VPWR _1512_ sky130_fd_sc_hd__and2b_1
XFILLER_23_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2140__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2863__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2315__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3000__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3040__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2370_ _1583_ _1587_ _1593_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__and3_2
XFILLER_96_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4040_ clknet_leaf_31_CLK _0232_ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_37_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2606__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2225__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3824_ clknet_leaf_10_CLK _0050_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_3755_ clknet_leaf_18_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\]
+ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] sky130_fd_sc_hd__dfrtp_4
X_3686_ _1122_ _1129_ _1157_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__a21o_1
X_2706_ _1664_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ _1693_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__a221o_1
X_2637_ net112 _1835_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2568_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\]
+ _1784_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__and3_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2499_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\] VGND VGND VPWR VPWR
+ _1725_ sky130_fd_sc_hd__inv_2
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2135__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout90_X net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A wdata[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2533__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1870_ _1354_ _1355_ _1356_ _1150_ _1147_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__a2111o_1
XANTENNA__3013__A1 _0564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3540_ _1616_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\] VGND VGND VPWR
+ VPWR _1124_ sky130_fd_sc_hd__nor2_1
X_3471_ _1053_ _1054_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2422_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND VPWR VPWR
+ _1648_ sky130_fd_sc_hd__inv_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2353_ net294 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] net94 VGND
+ VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
XFILLER_57_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4023_ clknet_leaf_5_CLK _0215_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_2284_ net217 net43 net82 VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2744__A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3807_ clknet_leaf_22_CLK _0033_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_1999_ _1057_ _1202_ _1491_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__nand3_1
XFILLER_20_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3738_ _1167_ _1317_ _1138_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__a21bo_1
X_3669_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__inv_2
XFILLER_69_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3491__A1 _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2654__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2564__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2971_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and2_1
XFILLER_91_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1922_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1410_ _1411_ _1414_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\]
+ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__a32o_1
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1853_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] _1290_ _1289_ VGND
+ VGND VPWR VPWR _1346_ sky130_fd_sc_hd__a21o_1
X_3523_ _1609_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\] VGND VGND VPWR
+ VPWR _1107_ sky130_fd_sc_hd__nor2_1
X_3454_ _0974_ _1038_ _0977_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__o21ba_1
X_2405_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND VPWR VPWR
+ _1631_ sky130_fd_sc_hd__inv_2
XFILLER_97_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3385_ net111 _0740_ _0744_ _0731_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__o211ai_1
XFILLER_97_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2336_ net310 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\] net92 VGND
+ VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
X_2267_ net215 net45 net81 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4006_ clknet_leaf_31_CLK _0198_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_9_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2198_ net260 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\] net101 VGND
+ VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2736__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold31 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[57\] VGND VGND VPWR VPWR net234
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold20 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[44\] VGND VGND VPWR VPWR net223
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[24\] VGND VGND VPWR VPWR net245
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold53 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[36\] VGND VGND VPWR VPWR net256
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[35\] VGND VGND VPWR VPWR net267
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold97 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[17\] VGND VGND VPWR VPWR net300
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[42\] VGND VGND VPWR VPWR net278
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold86 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[2\] VGND VGND VPWR VPWR net289
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3510__A_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2323__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3170_ net118 _0651_ _0652_ net119 VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__a211o_1
XFILLER_39_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2121_ _1577_ _1578_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__or3_1
XFILLER_39_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2052_ _1651_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _1545_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2954_ _0530_ _0538_ _0529_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a21boi_1
X_1905_ _1385_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__nand2_1
X_2885_ _0428_ _0465_ _0470_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag_c
+ sky130_fd_sc_hd__and3_1
XANTENNA__3877__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2233__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3806__RESET_B net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2718__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2194__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3506_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout100_A _1591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3437_ _1016_ _1019_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__or3b_1
X_3368_ _0949_ _0952_ _0950_ _0902_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__or4bb_2
XFILLER_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2319_ net244 net44 net77 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
X_3299_ _0483_ _0796_ _0800_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__and3b_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2143__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2185__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_10_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3685__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input30_A addr[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_25_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2318__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2842__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[13\]
+ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__nor2_1
XANTENNA__2176__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3222_ _1675_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\] VGND VGND VPWR
+ VPWR _0807_ sky130_fd_sc_hd__nor2_1
XFILLER_79_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3153_ net110 _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__or2_1
X_2104_ net276 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] net106 VGND
+ VGND VPWR VPWR _0021_ sky130_fd_sc_hd__mux2_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3084_ _0587_ _0665_ _0600_ _0574_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__o211ai_1
XFILLER_67_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2228__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4005__RESET_B net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2035_ _1623_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ _1622_ _1527_ VGND VGND VPWR VPWR _1528_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_99_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3986_ clknet_leaf_35_CLK _0178_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_2937_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__nand2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2868_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2167__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2799_ _0399_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[18\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout103_X net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3667__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2927__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2138__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3110__X _0695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2662__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2158__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2330__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3840_ clknet_leaf_21_CLK _0066_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3771_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2722_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\]
+ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__or2_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2149__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2653_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] _1838_ VGND VGND VPWR
+ VPWR _0273_ sky130_fd_sc_hd__nand2_1
X_2584_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] _1799_ VGND VGND VPWR VPWR
+ _1800_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout107 _1574_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
Xfanout118 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[27\] VGND VGND VPWR VPWR net118
+ sky130_fd_sc_hd__buf_2
Xfanout129 net131 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2321__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3205_ _1661_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] _0789_ VGND
+ VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a21bo_1
XANTENNA__2747__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3136_ _0517_ _0550_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3067_ _0621_ _0649_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] net116 VGND VGND VPWR
+ VPWR _1511_ sky130_fd_sc_hd__nand2b_1
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3969_ clknet_leaf_35_CLK myPWM.g_pwm_channel\[1\].CHANNEL.pwm_next net127 VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.pwm_out sky130_fd_sc_hd__dfrtp_1
XFILLER_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout80_A _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2657__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2312__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3909__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3000__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2331__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2303__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3823_ clknet_leaf_10_CLK _0049_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_3754_ clknet_leaf_19_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[14\]
+ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] sky130_fd_sc_hd__dfrtp_4
X_2705_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\]
+ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__xor2_1
X_3685_ net115 _1263_ _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__o21ba_1
X_2636_ _1836_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__2241__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2542__A1 _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2567_ _1787_ _1788_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[5\]
+ sky130_fd_sc_hd__nor2_1
X_2498_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] VGND VGND VPWR VPWR
+ _1724_ sky130_fd_sc_hd__inv_2
XANTENNA__4020__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3580__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3119_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0699_ _0703_ net123 VGND VGND
+ VPWR VPWR _0704_ sky130_fd_sc_hd__o22a_1
XANTENNA__2058__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2151__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2533__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout83_X net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2326__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3470_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2421_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR VPWR _1647_
+ sky130_fd_sc_hd__inv_2
X_2352_ net287 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\] net94 VGND
+ VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2283_ net246 net42 net82 VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_63_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4022_ clknet_leaf_5_CLK _0214_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2236__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_72_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_A net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3806_ clknet_leaf_16_CLK _0032_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1998_ _1382_ _1490_ _1059_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__a21o_1
X_3737_ _1138_ _1167_ _1317_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__nand3b_1
X_3668_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1246_ _1251_ VGND VGND VPWR
+ VPWR _1252_ sky130_fd_sc_hd__o21ai_1
X_2619_ net71 _1822_ _1823_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__or3_1
X_3599_ _1084_ _1091_ _1174_ _1179_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__or4bb_1
XFILLER_87_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2146__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2670__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input60_A wdata[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2506__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2970_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ _0501_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__and3_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1921_ _1374_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1852_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__or2_1
X_3522_ _1102_ _1103_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__a21o_1
X_3453_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[27\] _1702_ _0978_ _0985_ _1037_
+ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o221a_1
X_2404_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR _1630_
+ sky130_fd_sc_hd__inv_2
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3384_ _0889_ _0924_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__nand3_1
X_2335_ net204 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] net92 VGND
+ VGND VPWR VPWR _0229_ sky130_fd_sc_hd__mux2_1
XFILLER_97_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2266_ net272 net34 net81 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4005_ clknet_leaf_31_CLK _0197_ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2197_ net224 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] net101 VGND
+ VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_1
XFILLER_37_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout133_X net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2736__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold32 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[26\] VGND VGND VPWR VPWR net235
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[36\] VGND VGND VPWR VPWR net213
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[32\] VGND VGND VPWR VPWR net224
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[63\] VGND VGND VPWR VPWR net268
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[49\] VGND VGND VPWR VPWR net246
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold54 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[14\] VGND VGND VPWR VPWR net257
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[60\] VGND VGND VPWR VPWR net301
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[56\] VGND VGND VPWR VPWR net279
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2665__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold87 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[1\] VGND VGND VPWR VPWR net290
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_100_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_29_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_61_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input63_X net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2120_ net22 net21 net25 net24 VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__or4_1
X_2051_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] _1718_ _1543_ VGND VGND VPWR
+ VPWR _1544_ sky130_fd_sc_hd__a21o_1
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2953_ _0533_ _0537_ _0532_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a21o_1
X_1904_ _1055_ _1380_ _1384_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__or3_1
X_2884_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] _0426_ _0467_ _0469_
+ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__o211a_1
XANTENNA__2718__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3505_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__nand2_1
X_3436_ _1013_ _1015_ _1018_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__and4_1
XFILLER_97_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3367_ _0908_ _0913_ _0951_ _0948_ _0924_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__a32o_1
X_2318_ net313 net43 net77 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XFILLER_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3298_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _0880_ _0882_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\]
+ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__a22oi_1
X_2249_ net313 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] net97 VGND
+ VGND VPWR VPWR _0148_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2957__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input23_A addr[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2395__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2334__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3221_ _1677_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\] VGND VGND VPWR
+ VPWR _0806_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_9_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_9_CLK sky130_fd_sc_hd__clkbuf_8
X_3152_ _0533_ _0537_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2103_ net322 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] net106 VGND
+ VGND VPWR VPWR _0020_ sky130_fd_sc_hd__mux2_1
X_3083_ _0576_ _0586_ _0665_ _0584_ _0574_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__a311o_1
X_2034_ _1622_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ _1620_ _1526_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__o221a_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3985_ clknet_leaf_3_CLK _0177_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2936_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__inv_2
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2244__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2867_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] _0399_ _0405_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\]
+ _0432_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__o221a_1
XANTENNA__3583__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2798_ net69 _0397_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or3_1
X_3419_ _1659_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] VGND VGND VPWR
+ VPWR _1004_ sky130_fd_sc_hd__or2_1
XFILLER_58_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2154__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2329__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2853__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3770_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[30\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] sky130_fd_sc_hd__dfrtp_4
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2721_ _0322_ _0324_ _0326_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or4_1
X_2652_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[31\]
+ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__xnor2_1
X_2583_ net70 _1798_ _1799_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[10\]
+ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_74_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout119 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] VGND VGND VPWR VPWR net119
+ sky130_fd_sc_hd__buf_2
Xfanout108 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] VGND VGND VPWR VPWR net108
+ sky130_fd_sc_hd__buf_2
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3204_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] _1712_ VGND VGND VPWR
+ VPWR _0789_ sky130_fd_sc_hd__and2_1
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2239__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3135_ _0706_ _0718_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__or3b_1
X_3066_ _0617_ _0650_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2085__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2763__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2017_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1728_ VGND VGND VPWR VPWR
+ _1510_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout160_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3968_ clknet_leaf_8_CLK _0161_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2919_ _0502_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__and2_1
X_3899_ clknet_leaf_14_CLK _0125_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3594__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2149__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2673__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3009__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2848__A _1656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2839__B1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2583__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3822_ clknet_leaf_29_CLK _0048_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2913__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3753_ clknet_leaf_19_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[13\]
+ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] sky130_fd_sc_hd__dfrtp_4
X_2704_ _0318_ _0319_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__or3b_1
X_3684_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1266_ _1267_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__a22oi_1
X_2635_ net70 _1834_ _1835_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__or3_1
XANTENNA__3915__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2566_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1784_ net74 VGND VGND VPWR
+ VPWR _1788_ sky130_fd_sc_hd__o21ai_1
X_2497_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\] VGND VGND VPWR VPWR
+ _1723_ sky130_fd_sc_hd__inv_2
XFILLER_101_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3118_ _0489_ _0559_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3049_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0471_ _0629_ VGND VGND VPWR
+ VPWR _0634_ sky130_fd_sc_hd__and3_1
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3569__A_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout76_X net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2297__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_100_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3499__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout90 net91 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2342__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2420_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] VGND VGND VPWR VPWR _1646_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2351_ net217 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\] net94 VGND
+ VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
Xpwm_wrapper_190 VGND VGND VPWR VPWR pwm_wrapper_190/HI rdata[19] sky130_fd_sc_hd__conb_1
XFILLER_96_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2282_ net307 net41 net82 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
XANTENNA__2288__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4021_ clknet_leaf_4_CLK _0213_ net136 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1997_ _1375_ _1376_ _1378_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__or3b_1
XFILLER_20_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3805_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.pwm_next net167 VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.pwm_out sky130_fd_sc_hd__dfrtp_1
XANTENNA__2252__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3736_ _1313_ _1315_ _1316_ _1319_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__o211a_1
X_3667_ net114 _1247_ _1250_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__o21a_1
X_3598_ _1084_ _1091_ _1180_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__or3b_1
X_2618_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\]
+ _1818_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__and3_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2549_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__nand2_1
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2279__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input53_A wdata[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2337__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3022__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1920_ _1079_ _1371_ _1373_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__nand3_1
XANTENNA__2861__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1851_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__or2_1
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3521_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\]
+ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__and2b_1
X_3452_ net119 _1703_ _0983_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__or3_1
X_3383_ _0927_ _0943_ _0945_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__and4b_1
X_2403_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] VGND VGND VPWR VPWR
+ _1629_ sky130_fd_sc_hd__inv_2
X_2334_ net215 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\] net93 VGND
+ VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3458__B1 _0990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2265_ _1603_ net336 net83 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_68_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4004_ clknet_leaf_1_CLK _0196_ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2196_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[1\]
+ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__nand2_2
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2247__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2681__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2771__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3719_ _1154_ _1302_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__xor2_1
XFILLER_0_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold11 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[28\] VGND VGND VPWR VPWR net214
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[16\] VGND VGND VPWR VPWR net225
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[30\] VGND VGND VPWR VPWR net236
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[31\] VGND VGND VPWR VPWR net247
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[7\] VGND VGND VPWR VPWR net258
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3449__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold66 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[55\] VGND VGND VPWR VPWR net269
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold88 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[37\] VGND VGND VPWR VPWR net291
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[8\] VGND VGND VPWR VPWR net280
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold99 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[13\] VGND VGND VPWR VPWR net302
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2157__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input56_X net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2050_ _1651_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _1543_ sky130_fd_sc_hd__nor2_1
XANTENNA__3304__X _0889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2952_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] _0535_ _0534_ VGND
+ VGND VPWR VPWR _0537_ sky130_fd_sc_hd__a21bo_1
X_1903_ _1394_ _1395_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] VGND VGND VPWR
+ VPWR _1396_ sky130_fd_sc_hd__a21oi_1
X_2883_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] _0426_ _0468_ VGND
+ VGND VPWR VPWR _0469_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_77_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3504_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__and2_1
X_3435_ _1662_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] _1012_ _1017_
+ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__o211a_1
XANTENNA__3923__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3366_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0912_ _0917_ _0921_ _0911_
+ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__o221ai_1
XFILLER_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2317_ net293 net42 net77 VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
X_3297_ _0480_ _0864_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__xnor2_1
X_2248_ net293 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] net97 VGND
+ VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
XFILLER_57_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2179_ net220 net40 net84 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__mux2_1
XFILLER_13_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput67 net67 VGND VGND VPWR VPWR pwm_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2676__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input16_A addr[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2350__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3220_ _1679_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR
+ VPWR _0805_ sky130_fd_sc_hd__nor2_1
XFILLER_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3151_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__inv_2
XANTENNA__2586__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2102_ net263 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] net106 VGND
+ VGND VPWR VPWR _0019_ sky130_fd_sc_hd__mux2_1
XANTENNA__2884__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3082_ _0587_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__xor2_1
X_2033_ _1620_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\] _1524_ _1525_
+ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__a211o_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3984_ clknet_leaf_35_CLK _0176_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_2935_ _0518_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__and2b_1
X_2866_ _0440_ _0444_ _0451_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and3_1
XANTENNA__2260__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2797_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\]
+ _0393_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__and3_1
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3418_ net108 _1713_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__and2_1
XANTENNA_input8_A addr[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3349_ _0788_ _0789_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__nor2_1
XFILLER_97_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2170__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2345__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2720_ _0328_ _0333_ _0335_ _0337_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__or4_1
X_2651_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _0269_ _0271_ VGND VGND VPWR
+ VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[31\] sky130_fd_sc_hd__o21ba_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2582_ net117 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1795_ VGND VGND VPWR
+ VPWR _1799_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_74_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout109 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] VGND VGND VPWR VPWR net109
+ sky130_fd_sc_hd__buf_2
X_3203_ _0787_ _0517_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__and2b_1
X_3134_ _0712_ _0713_ _0715_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__and3_1
XFILLER_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3065_ _0621_ _0649_ _0618_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__a21bo_1
XFILLER_82_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2016_ _1403_ _1494_ _1507_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__or3b_1
XANTENNA__2255__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3967_ clknet_leaf_7_CLK _0160_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2918_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__or2_1
X_3898_ clknet_leaf_13_CLK _0124_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_4
X_2849_ _0360_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable VGND VGND VPWR VPWR
+ _0436_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_96_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold130 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[26\] VGND VGND VPWR VPWR net333
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2165__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3918__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3009__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2536__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3821_ clknet_leaf_29_CLK _0047_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3752_ clknet_leaf_19_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[12\]
+ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\] sky130_fd_sc_hd__dfrtp_1
X_2703_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] _1660_ _1679_ net122
+ _0320_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o221a_1
X_3683_ _1171_ _1174_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__xor2_1
X_2634_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] _1832_ VGND VGND VPWR VPWR
+ _1835_ sky130_fd_sc_hd__and2_1
X_2565_ _1613_ _1785_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__nor2_1
XANTENNA__2527__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2496_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\] VGND VGND VPWR VPWR
+ _1722_ sky130_fd_sc_hd__inv_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3117_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0696_ _0700_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\]
+ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__o22a_1
X_3048_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0632_ _0630_ VGND VGND VPWR
+ VPWR _0633_ sky130_fd_sc_hd__o21a_1
XFILLER_70_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout69_X net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3499__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout80 _1594_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_4
XANTENNA__2757__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout91 _1588_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_4
XFILLER_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2509__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2350_ net246 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\] net94 VGND
+ VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
Xpwm_wrapper_180 VGND VGND VPWR VPWR pwm_wrapper_180/HI rdata[9] sky130_fd_sc_hd__conb_1
X_2281_ net239 net40 net80 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4020_ clknet_leaf_3_CLK _0212_ net136 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xpwm_wrapper_191 VGND VGND VPWR VPWR pwm_wrapper_191/HI rdata[20] sky130_fd_sc_hd__conb_1
XFILLER_37_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3804_ clknet_leaf_14_CLK _0031_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_1996_ _1416_ _1418_ _1420_ _1488_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__o211a_1
X_3735_ _1625_ _1317_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__nand3_1
X_3666_ net114 _1247_ _1249_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND
+ VPWR VPWR _1250_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_93_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2617_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1818_ net114 VGND VGND VPWR
+ VPWR _1822_ sky130_fd_sc_hd__a21oi_1
X_3597_ _1175_ _1179_ _1180_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a21oi_1
X_2548_ net75 VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__inv_2
X_2479_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\] VGND VGND VPWR VPWR
+ _1705_ sky130_fd_sc_hd__inv_2
XFILLER_56_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload0 clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input46_A wdata[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2353__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1850_ _1138_ _1141_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__nand2_1
X_3520_ _1102_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__and2_1
X_3451_ _0988_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nand2b_1
X_3382_ _0929_ _0930_ _0931_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__and4b_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2402_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] VGND VGND VPWR VPWR _1628_
+ sky130_fd_sc_hd__inv_2
XFILLER_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2333_ net272 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] net93 VGND
+ VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
X_2264_ _1583_ _1589_ _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__and3_2
X_2195_ net247 net58 net87 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_1
XFILLER_84_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4003_ clknet_leaf_29_CLK _0195_ net134 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2130__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1979_ _1433_ _1471_ _1431_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3718_ _1130_ _1156_ _1159_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__a21bo_1
X_3649_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] _1232_ VGND VGND VPWR VPWR
+ _1233_ sky130_fd_sc_hd__xnor2_1
XFILLER_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold23 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[27\] VGND VGND VPWR VPWR net226
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[33\] VGND VGND VPWR VPWR net215
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[30\] VGND VGND VPWR VPWR net248
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[23\] VGND VGND VPWR VPWR net237
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[12\] VGND VGND VPWR VPWR net259
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold67 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[27\] VGND VGND VPWR VPWR net270
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold78 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[12\] VGND VGND VPWR VPWR net281
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[16\] VGND VGND VPWR VPWR net292
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_39_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2173__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2188__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input49_X net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2348__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2112__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3033__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2872__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2951_ _0534_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nand2_1
X_1902_ _1053_ _1385_ _1222_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a21o_1
XANTENNA__2083__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2882_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] _0416_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ _1694_ _0429_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__a221o_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2179__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3503_ _1084_ _1085_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_77_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3434_ _1672_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] VGND VGND VPWR
+ VPWR _1019_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0898_ _0896_ VGND VGND VPWR
+ VPWR _0950_ sky130_fd_sc_hd__or3b_1
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3296_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\] _0868_ _0880_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\]
+ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__o22a_1
X_2316_ net225 net41 net77 VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XANTENNA__2258__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2247_ net225 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] net97 VGND
+ VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2103__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2178_ net323 net39 net86 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_1
XANTENNA__2782__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout96_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput68 net68 VGND VGND VPWR VPWR pwm_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__3405__X _0990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2168__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3150_ net109 _0732_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__nand2_1
XFILLER_94_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3081_ _0576_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nand2_1
X_2101_ net228 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] net106 VGND
+ VGND VPWR VPWR _0018_ sky130_fd_sc_hd__mux2_1
XFILLER_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2032_ net117 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__and4bb_1
XFILLER_35_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3983_ clknet_leaf_34_CLK _0175_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2934_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__nand2b_1
X_2865_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] _0385_ _0446_ _0449_
+ _0450_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_CLK_X clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2796_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _0395_ VGND VGND VPWR VPWR
+ _0397_ sky130_fd_sc_hd__nor2_1
X_3417_ _0998_ _1001_ _0997_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2324__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3348_ _0517_ _0787_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__xor2_1
XFILLER_97_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3279_ _0807_ _0863_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__or2_1
XFILLER_45_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout99_X net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2315__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2361__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2650_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _0269_ net71 VGND VGND VPWR
+ VPWR _0271_ sky130_fd_sc_hd__a21o_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2581_ net117 _1795_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] VGND VGND VPWR
+ VPWR _1798_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_74_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2306__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3202_ _0521_ _0525_ _0783_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__o31a_1
XFILLER_94_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3133_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] _0716_ _0717_ VGND VGND VPWR
+ VPWR _0718_ sky130_fd_sc_hd__a21o_1
XFILLER_55_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3064_ _0606_ _0648_ _0607_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a21oi_1
X_2015_ _1403_ _1489_ _1506_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_85_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3966_ clknet_leaf_7_CLK _0159_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_2917_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__nand2_1
X_3897_ clknet_leaf_13_CLK _0123_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2271__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2848_ _1656_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\] VGND VGND VPWR
+ VPWR _0435_ sky130_fd_sc_hd__xnor2_1
X_2779_ _0385_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[12\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold131 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[39\] VGND VGND VPWR VPWR net334
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout101_X net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold120 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[14\] VGND VGND VPWR VPWR net323
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2970__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2181__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_10_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_92_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2356__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2880__A _1688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3820_ clknet_leaf_28_CLK _0046_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3751_ clknet_leaf_19_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[11\]
+ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2091__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2702_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] _1660_ _1689_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\]
+ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3682_ _1179_ _1265_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__xor2_1
X_2633_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] _1832_ VGND VGND VPWR VPWR
+ _1834_ sky130_fd_sc_hd__nor2_1
X_2564_ net74 _1785_ _1786_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[4\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__1916__B1_N net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2495_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] VGND VGND VPWR VPWR
+ _1721_ sky130_fd_sc_hd__inv_2
XFILLER_101_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3116_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0699_ _0700_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\]
+ _0697_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a221o_1
XFILLER_67_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2266__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3047_ _0629_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nand2_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3949_ clknet_leaf_34_CLK _0142_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_21_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2176__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout81 _1594_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_2
Xfanout92 _1597_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_4
Xfanout70 _1774_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_80_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpwm_wrapper_181 VGND VGND VPWR VPWR pwm_wrapper_181/HI rdata[10] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_170 VGND VGND VPWR VPWR pwm_wrapper_170/HI error sky130_fd_sc_hd__conb_1
X_2280_ net298 net39 net82 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
Xpwm_wrapper_192 VGND VGND VPWR VPWR pwm_wrapper_192/HI rdata[21] sky130_fd_sc_hd__conb_1
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2086__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3803_ clknet_leaf_15_CLK _0030_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ _1481_ _1484_ _1486_ _1487_ _1418_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__a2111o_1
X_3734_ _1141_ _1166_ _1278_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__nand3_1
X_3665_ _1069_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2616_ _1821_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[21\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__3809__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3596_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] _1727_ _1179_ _1176_
+ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a31o_1
XANTENNA__3942__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2547_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable _1772_ VGND VGND VPWR VPWR
+ _1773_ sky130_fd_sc_hd__nand2_1
XFILLER_87_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2478_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\] VGND VGND VPWR VPWR
+ _1704_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_50_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4079_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[5\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_54_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2739__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload1 clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_6
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout81_X net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wdata[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3450_ _1687_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] _0990_ _1033_
+ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__a221o_1
X_3381_ net111 _0536_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__or2_1
X_2401_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] VGND VGND VPWR VPWR
+ _1627_ sky130_fd_sc_hd__inv_2
XFILLER_69_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2332_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[1\]
+ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__nand2_2
XFILLER_84_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4002_ clknet_leaf_8_CLK _0194_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_2263_ _1601_ _1575_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__nor2_1
X_2194_ net248 net57 net87 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__mux2_1
XFILLER_37_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3717_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1281_ _1300_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\]
+ _1299_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__o221a_1
X_1978_ _1436_ _1439_ _1469_ _1470_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__o31a_1
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3648_ _1059_ _1197_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__xor2_1
X_3579_ _1151_ _1160_ _1162_ _1146_ _1161_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__o221a_1
Xhold13 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[45\] VGND VGND VPWR VPWR net216
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold24 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[20\] VGND VGND VPWR VPWR net227
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[58\] VGND VGND VPWR VPWR net249
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[31\] VGND VGND VPWR VPWR net238
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3449__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold68 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[51\] VGND VGND VPWR VPWR net271
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[7\] VGND VGND VPWR VPWR net282
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[33\] VGND VGND VPWR VPWR net260
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2950_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__or2_1
X_1901_ _1053_ _1222_ _1385_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__nand3_1
X_2881_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] _0416_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ _1694_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__o221a_1
X_3502_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\]
+ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_77_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3433_ _1665_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] net124 _1710_
+ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_90_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _0896_ _0901_ _0904_ _0905_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__and4_1
X_3295_ _0866_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__or2_1
X_2315_ net296 net40 net76 VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
X_2246_ net296 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] net96 VGND
+ VGND VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2177_ net302 net38 net84 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_1
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2274__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3895__RESET_B net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_X net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout89_A _1588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2184__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input61_X net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3080_ _0603_ _0664_ _0578_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a21o_1
XFILLER_67_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2100_ net300 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] net106 VGND
+ VGND VPWR VPWR _0017_ sky130_fd_sc_hd__mux2_1
XFILLER_94_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2031_ _1619_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ _1618_ _1523_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__o221a_1
XFILLER_54_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2097__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3982_ clknet_leaf_34_CLK _0174_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2094__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2933_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\]
+ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__and2b_1
XFILLER_50_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2864_ _1666_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[11\] _0388_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\]
+ _0439_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__o221a_1
X_2795_ _0395_ _0396_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3416_ _0999_ _1000_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nand2_1
XFILLER_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2269__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3347_ _0929_ _0930_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__o21a_1
XANTENNA__3950__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3278_ _0796_ _0800_ _0483_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__a21boi_1
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2229_ _1602_ net340 net87 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__a21o_1
XFILLER_26_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2260__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2179__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input21_A addr[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2251__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_5 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2580_ net117 _1795_ _1797_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[9\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_74_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2878__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2089__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3201_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] _1714_ _0519_ _0518_
+ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a31oi_1
XFILLER_79_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3132_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] _0714_ _0716_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\]
+ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__o22ai_1
XFILLER_94_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3063_ _0611_ _0647_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__nor2_1
XFILLER_27_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2014_ _1498_ _1503_ _1505_ _1504_ _1501_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__a311o_1
XFILLER_63_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3965_ clknet_leaf_7_CLK _0158_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_3896_ clknet_leaf_13_CLK _0122_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2242__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2916_ _0498_ _0499_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout139_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2847_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\]
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__xnor2_1
Xhold110 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[18\] VGND VGND VPWR VPWR net313
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ net123 _0382_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_96_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold132 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[38\] VGND VGND VPWR VPWR net335
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[11\] VGND VGND VPWR VPWR net324
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3750_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[10\]
+ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2372__S _1599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2701_ _1666_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\]
+ _1676_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a22o_1
X_3681_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] _1727_ _1175_ VGND
+ VGND VPWR VPWR _1265_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2632_ _1833_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[25\]
+ sky130_fd_sc_hd__inv_2
X_2563_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1779_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__a21o_1
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2494_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\] VGND VGND VPWR VPWR
+ _1720_ sky130_fd_sc_hd__inv_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3115_ _0492_ _0565_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__xnor2_1
X_3046_ _0473_ _0628_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nand2_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2282__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3948_ clknet_leaf_34_CLK _0141_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3879_ clknet_leaf_25_CLK _0105_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_21_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_1__f_CLK_X clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2192__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout71 _1774_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xfanout82 _1594_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
XFILLER_80_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout93 _1597_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_2
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpwm_wrapper_171 VGND VGND VPWR VPWR pwm_wrapper_171/HI rdata[0] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_182 VGND VGND VPWR VPWR pwm_wrapper_182/HI rdata[11] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_193 VGND VGND VPWR VPWR pwm_wrapper_193/HI rdata[22] sky130_fd_sc_hd__conb_1
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2367__S _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3761__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3802_ clknet_leaf_14_CLK _0029_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_1994_ _1407_ _1415_ _1485_ _1412_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__or4b_1
X_3733_ _1166_ _1278_ _1141_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__a21o_1
X_3664_ _1078_ _1185_ _1071_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__o21a_1
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload30 clknet_leaf_15_CLK VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_8
X_2615_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1818_ _1820_ net71 VGND VGND
+ VPWR VPWR _1821_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_93_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3595_ _1177_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__nand2_2
X_2546_ _1737_ _1752_ _1771_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__and3_1
X_2477_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\] VGND VGND VPWR VPWR
+ _1703_ sky130_fd_sc_hd__inv_2
XFILLER_87_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2277__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4078_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[4\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] sky130_fd_sc_hd__dfrtp_4
X_3029_ _0611_ _0612_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_leaf_0_CLK VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2187__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout74_X net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2400_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND VPWR VPWR
+ _1626_ sky130_fd_sc_hd__inv_2
X_3380_ _0889_ _0953_ _0958_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a211o_1
X_2331_ net238 net58 net78 VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
XANTENNA__2886__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2262_ net238 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] net98 VGND
+ VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4001_ clknet_leaf_8_CLK _0193_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2097__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2193_ net230 net55 net87 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__mux2_1
XFILLER_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3716_ _1130_ _1156_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1977_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] _1437_ _1438_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\]
+ _1432_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__o32a_1
X_3647_ net112 _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__nand2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3578_ _1621_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\] VGND VGND VPWR
+ VPWR _1162_ sky130_fd_sc_hd__or2_1
X_2529_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\]
+ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__xor2_1
XANTENNA__2796__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_88_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold14 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[50\] VGND VGND VPWR VPWR net217
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[58\] VGND VGND VPWR VPWR net250
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[18\] VGND VGND VPWR VPWR net228
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[47\] VGND VGND VPWR VPWR net239
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3404__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold58 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[56\] VGND VGND VPWR VPWR net261
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[32\] VGND VGND VPWR VPWR net272
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input51_A wdata[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1900_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] _1389_ VGND VGND VPWR VPWR
+ _1393_ sky130_fd_sc_hd__xnor2_1
X_2880_ _1688_ _0411_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3501_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] _1726_ VGND VGND VPWR
+ VPWR _1085_ sky130_fd_sc_hd__nand2_1
XFILLER_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3432_ _1668_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\] _1709_ net123
+ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_90_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _0937_ _0947_ _0946_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__a21o_1
XANTENNA__3505__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3294_ _0591_ _0806_ _0865_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__nor3_1
X_2314_ net257 net39 net77 VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XFILLER_38_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2245_ net257 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] net97 VGND
+ VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
X_2176_ net259 net37 net84 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3948__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2290__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_298 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2566__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input54_X net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ _1619_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] _1521_ _1522_
+ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__a211o_1
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3981_ clknet_leaf_33_CLK _0173_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ _0515_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nand2_2
XFILLER_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2863_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] _0380_ _0435_ _0447_
+ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__2404__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2794_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0393_ net73 VGND VGND VPWR
+ VPWR _0396_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3219__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3415_ net110 _1715_ _1716_ net111 VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a22o_1
X_3346_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0925_ VGND VGND VPWR VPWR _0931_
+ sky130_fd_sc_hd__nand2_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3277_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0859_ _0861_ VGND VGND VPWR
+ VPWR _0862_ sky130_fd_sc_hd__a21oi_1
X_2228_ net268 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] net103 VGND
+ VGND VPWR VPWR _0128_ sky130_fd_sc_hd__mux2_1
XANTENNA__3285__A1 _1682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2159_ net299 net55 net91 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__mux2_1
XFILLER_81_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2285__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2195__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input14_A addr[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2787__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2539__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3200_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] _1714_ _0784_ VGND
+ VGND VPWR VPWR _0785_ sky130_fd_sc_hd__a21o_1
XANTENNA__2894__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3131_ _0513_ _0553_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3062_ _0598_ _0604_ _0614_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__a21oi_1
X_2013_ _1500_ _1501_ _1503_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__or4bb_1
XANTENNA__3502__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3019__A1 _1688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3964_ clknet_leaf_7_CLK _0157_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_3895_ clknet_leaf_13_CLK net262 net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_2915_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__inv_2
X_2846_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\]
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__xnor2_1
Xhold100 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[21\] VGND VGND VPWR VPWR net303
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ net123 _0382_ net73 VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_96_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold111 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[61\] VGND VGND VPWR VPWR net314
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[39\] VGND VGND VPWR VPWR net325
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold133 myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[1\] VGND VGND VPWR VPWR net336
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3961__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input6_A addr[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3329_ _0513_ _0793_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__and2b_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3603__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2700_ _1666_ net124 _1675_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND
+ VPWR VPWR _0318_ sky130_fd_sc_hd__a2bb2o_1
X_3680_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1260_ _1263_ net115 VGND VGND
+ VPWR VPWR _1264_ sky130_fd_sc_hd__a22oi_1
XFILLER_40_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2889__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2631_ net70 _1831_ _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__or3_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2562_ _1784_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__inv_2
X_2493_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] VGND VGND VPWR VPWR
+ _1719_ sky130_fd_sc_hd__inv_2
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2160__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3513__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3114_ _0495_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__xnor2_1
X_3045_ _0471_ _0629_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] VGND VGND VPWR
+ VPWR _0630_ sky130_fd_sc_hd__a21o_1
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout151_A net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3956__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3947_ clknet_leaf_33_CLK _0140_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3878_ clknet_leaf_25_CLK _0104_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2829_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0418_ VGND VGND VPWR VPWR
+ _0420_ sky130_fd_sc_hd__and2_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2151__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_3__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_3__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_279 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout72 net73 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_2
Xfanout83 _1594_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_4
Xfanout94 _1597_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__buf_4
XFILLER_6_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xpwm_wrapper_172 VGND VGND VPWR VPWR pwm_wrapper_172/HI rdata[1] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_183 VGND VGND VPWR VPWR pwm_wrapper_183/HI rdata[12] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_194 VGND VGND VPWR VPWR pwm_wrapper_194/HI rdata[23] sky130_fd_sc_hd__conb_1
XFILLER_77_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2142__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3801_ clknet_leaf_13_CLK _0028_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1483_ VGND VGND VPWR VPWR
+ _1486_ sky130_fd_sc_hd__nor2_1
XFILLER_60_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3732_ _1276_ _1277_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] VGND VGND VPWR
+ VPWR _1316_ sky130_fd_sc_hd__a21o_1
X_3663_ _1063_ _1243_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__xnor2_1
Xclkload20 clknet_leaf_19_CLK VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinv_8
X_2614_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1818_ VGND VGND VPWR VPWR
+ _1820_ sky130_fd_sc_hd__nor2_1
Xclkload31 clknet_leaf_16_CLK VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_93_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3594_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__or2_1
X_2545_ _1761_ _1770_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__nor2_1
X_2476_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] VGND VGND VPWR VPWR
+ _1702_ sky130_fd_sc_hd__inv_2
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2133__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4077_ clknet_leaf_21_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_43_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3028_ _0611_ _0612_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nor2_1
XFILLER_24_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2293__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload3 clknet_leaf_1_CLK VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__2372__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3624__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3624__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2330_ net236 net57 net78 VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
X_2261_ net236 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] net98 VGND
+ VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
X_4000_ clknet_leaf_7_CLK _0192_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_2192_ net206 net54 net87 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__mux2_1
XFILLER_77_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3911__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2407__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1976_ net117 _1442_ _1446_ _1468_ _1443_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__o221a_1
XANTENNA__2413__Y _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3715_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1281_ _1297_ _1298_ _1283_
+ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3646_ _1202_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__xnor2_1
X_3577_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\]
+ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nand2b_1
X_2528_ _1626_ net116 _1650_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _1753_
+ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__o221ai_1
XANTENNA__2288__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2106__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2459_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] VGND VGND VPWR VPWR _1685_
+ sky130_fd_sc_hd__inv_2
Xhold37 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[49\] VGND VGND VPWR VPWR net240
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[5\] VGND VGND VPWR VPWR net229
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold15 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[45\] VGND VGND VPWR VPWR net218
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 _0121_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[23\] VGND VGND VPWR VPWR net251
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_67_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2987__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input44_A wdata[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2198__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3500_ _1081_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nor2_2
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3431_ _1672_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ _1670_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _0939_ _0942_ _0936_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_29_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2313_ net211 net38 net76 VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
X_3293_ _0862_ _0869_ _0875_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__and4_1
X_2244_ net211 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] net96 VGND
+ VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
X_2175_ net232 net36 net84 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__mux2_1
XFILLER_38_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3964__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1959_ _1098_ _1347_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3629_ _1210_ _1211_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR
+ VPWR _1213_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2327__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2318__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_X net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3980_ clknet_leaf_33_CLK _0172_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2931_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__or2_1
XFILLER_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2862_ _1658_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[4\] VGND VGND VPWR
+ VPWR _0448_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_13_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2793_ _1676_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__nor2_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2309__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3414_ _1655_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\] _1715_ net110
+ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_31_CLK sky130_fd_sc_hd__clkbuf_8
X_3345_ net111 _0536_ _0928_ net110 VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a22oi_1
X_3276_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _0860_ VGND VGND VPWR VPWR
+ _0861_ sky130_fd_sc_hd__xnor2_1
X_2227_ net222 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] net103 VGND
+ VGND VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2158_ net301 net54 net91 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_1
XANTENNA__3959__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2089_ net331 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] net105 VGND
+ VGND VPWR VPWR _0006_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout94_A _1597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_22_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_49_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2539__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_13_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_74_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3130_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0709_ _0714_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\]
+ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__a22oi_1
XFILLER_94_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3061_ _0634_ _0635_ _0645_ _0633_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or4b_2
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2012_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1497_ _1504_ VGND VGND VPWR
+ VPWR _1505_ sky130_fd_sc_hd__o21ba_1
XANTENNA__3779__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3963_ clknet_leaf_6_CLK _0156_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_3894_ clknet_leaf_11_CLK _0120_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_4
X_2914_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\]
+ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__nand2b_1
XFILLER_31_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2845_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\]
+ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold101 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[22\] VGND VGND VPWR VPWR net304
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2776_ _0383_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[11\]
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[42\] VGND VGND VPWR VPWR net315
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[4\] VGND VGND VPWR VPWR net326
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[1\] VGND VGND VPWR VPWR net337
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3328_ net124 _0910_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__nand2_1
XFILLER_100_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2296__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3259_ net118 _0838_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__nor2_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout97_X net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_2_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_80_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2630_ net113 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1826_ VGND VGND VPWR
+ VPWR _1832_ sky130_fd_sc_hd__and3_1
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2561_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\]
+ _1779_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__and3_1
XFILLER_99_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2492_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] VGND VGND VPWR VPWR
+ _1718_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_20_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_35_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3113_ _0489_ _0559_ _0487_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__o21a_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3044_ _0473_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__or2_1
XFILLER_55_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3946_ clknet_leaf_33_CLK _0139_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_98_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3877_ clknet_leaf_24_CLK _0103_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2828_ _0419_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[27\]
+ sky130_fd_sc_hd__inv_2
X_2759_ net108 _0370_ net72 VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout73 _0361_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_2
Xfanout95 _1597_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
Xfanout84 _1590_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3173__X _0758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpwm_wrapper_195 VGND VGND VPWR VPWR pwm_wrapper_195/HI rdata[24] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_173 VGND VGND VPWR VPWR pwm_wrapper_173/HI rdata[2] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_184 VGND VGND VPWR VPWR pwm_wrapper_184/HI rdata[13] sky130_fd_sc_hd__conb_1
XFILLER_92_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ clknet_leaf_13_CLK _0027_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1992_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1414_ VGND VGND VPWR VPWR
+ _1485_ sky130_fd_sc_hd__nor2_1
X_3731_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] _1276_ _1277_ _1314_ VGND VGND
+ VPWR VPWR _1315_ sky130_fd_sc_hd__a31o_1
X_3662_ _1060_ _1245_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload10 clknet_leaf_36_CLK VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__3792__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload32 clknet_leaf_17_CLK VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__inv_8
X_3593_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__nand2_1
Xclkload21 clknet_leaf_20_CLK VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__inv_8
X_2613_ _1818_ _1819_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[20\]
+ sky130_fd_sc_hd__nor2_1
X_2544_ _1763_ _1765_ _1767_ _1769_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_93_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2475_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\] VGND VGND VPWR VPWR
+ _1701_ sky130_fd_sc_hd__inv_2
XANTENNA__1934__A1_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3330__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4076_ clknet_leaf_21_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_55_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3027_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__nor2_1
XFILLER_24_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3967__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3929_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[25\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] sky130_fd_sc_hd__dfrtp_4
Xclkload4 clknet_leaf_29_CLK VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_6
XFILLER_3_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3609__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2513__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2260_ net311 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] net98 VGND
+ VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
X_2191_ net270 net53 net87 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__mux2_1
XFILLER_92_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3787__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1975_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1445_ _1463_ _1466_ _1467_
+ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__o221a_1
X_3714_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] _1282_ _1285_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\]
+ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_31_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3645_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] _1720_ _1198_ VGND
+ VGND VPWR VPWR _1229_ sky130_fd_sc_hd__a21o_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout107_A _1574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3576_ _1152_ _1159_ _1153_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2527_ _1607_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\]
+ _1623_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__o22a_1
X_2458_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND VPWR VPWR
+ _1684_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold27 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[29\] VGND VGND VPWR VPWR net230
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[41\] VGND VGND VPWR VPWR net219
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[44\] VGND VGND VPWR VPWR net241
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold49 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[59\] VGND VGND VPWR VPWR net252
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2389_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__inv_2
XFILLER_83_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4059_ clknet_leaf_6_CLK _0251_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_39_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2290__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2987__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input37_A wdata[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1856__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2067__X _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2281__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3430_ _1011_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3361_ _0927_ _0932_ _0943_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__o211a_1
X_2312_ net281 net37 net76 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3292_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0859_ _0871_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\]
+ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__o221a_1
X_2243_ net281 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] net96 VGND
+ VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_1
XFILLER_38_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1847__A1 _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2174_ net253 net35 net84 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__mux2_1
XFILLER_38_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2272__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1958_ _1095_ _1348_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1889_ _1188_ _1194_ _1193_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__a21bo_1
XANTENNA__1992__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3628_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _1210_ _1211_ VGND VGND VPWR
+ VPWR _1212_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_8_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3559_ _1134_ _1138_ _1141_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__or3_1
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3873__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4051__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3890__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2254__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2930_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nand2_1
X_2861_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\]
+ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_13_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ net73 _0392_ _0394_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[16\]
+ sky130_fd_sc_hd__and3_1
XFILLER_7_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3413_ _1657_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ _1655_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__o22a_1
X_3344_ net110 _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__nor2_1
X_3275_ _0573_ _0857_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__xnor2_1
X_2226_ net299 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\] net103 VGND
+ VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ net275 net53 net91 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
X_2088_ net316 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] net105 VGND
+ VGND VPWR VPWR _0005_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_2_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4072__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2611__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout87_A _1590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2236__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_57_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3617__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3060_ _0642_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__nand2_1
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2011_ _1491_ _1502_ _1643_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__a21oi_1
XFILLER_67_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3962_ clknet_leaf_6_CLK _0155_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__3795__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3893_ clknet_leaf_11_CLK _0119_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_4
X_2913_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_75_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2844_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[16\]
+ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_9_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3527__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2775_ net69 _0381_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_96_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold113 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[5\] VGND VGND VPWR VPWR net316
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[41\] VGND VGND VPWR VPWR net327
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[34\] VGND VGND VPWR VPWR net305
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 myPWM.g_pwm_channel\[0\].CHANNEL.polarity VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_84_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3327_ _0505_ _0890_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3258_ _0831_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__nand2_1
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2209_ net241 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\] net100 VGND
+ VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
X_3189_ _1667_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\] VGND VGND VPWR
+ VPWR _0774_ sky130_fd_sc_hd__nor2_1
XFILLER_39_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_93_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3406__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2560_ _1783_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[3\]
+ sky130_fd_sc_hd__inv_2
X_2491_ myPWM.g_pwm_channel\[0\].CHANNEL.polarity VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__inv_2
XFILLER_99_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2696__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2696__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3112_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0696_ VGND VGND VPWR VPWR
+ _0697_ sky130_fd_sc_hd__and2_1
X_3043_ _1696_ _1700_ _0626_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a22o_1
XFILLER_67_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3945_ clknet_leaf_33_CLK _0138_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3876_ clknet_leaf_24_CLK _0102_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2827_ net69 _0417_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__or3_1
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2758_ _0370_ _0371_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[5\]
+ sky130_fd_sc_hd__nor2_1
X_2689_ _1616_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\] _0305_ _0307_
+ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o211a_1
XFILLER_58_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2100__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout74 _1773_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout85 _1590_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xfanout96 net99 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_4
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpwm_wrapper_196 VGND VGND VPWR VPWR pwm_wrapper_196/HI rdata[25] sky130_fd_sc_hd__conb_1
XANTENNA__2678__A1 _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpwm_wrapper_185 VGND VGND VPWR VPWR pwm_wrapper_185/HI rdata[14] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_174 VGND VGND VPWR VPWR pwm_wrapper_174/HI rdata[3] sky130_fd_sc_hd__conb_1
XFILLER_92_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1991_ net115 _1479_ _1483_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND
+ VPWR VPWR _1484_ sky130_fd_sc_hd__a22oi_1
X_3730_ _1274_ _1311_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] VGND VGND VPWR
+ VPWR _1314_ sky130_fd_sc_hd__o21a_1
X_3661_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] _1724_ _1244_ VGND
+ VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a21oi_1
X_3592_ _1631_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\] VGND VGND VPWR
+ VPWR _1176_ sky130_fd_sc_hd__nor2_1
Xclkload22 clknet_leaf_21_CLK VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__bufinv_16
Xclkload33 clknet_leaf_18_CLK VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_8
X_2612_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1816_ net75 VGND VGND VPWR
+ VPWR _1819_ sky130_fd_sc_hd__o21ai_1
Xclkload11 clknet_leaf_2_CLK VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinv_4
X_2543_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1624_ _1648_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\]
+ _1768_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_93_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2474_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] VGND VGND VPWR VPWR
+ _1700_ sky130_fd_sc_hd__inv_2
XFILLER_68_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4075_ clknet_leaf_21_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[1\] net155
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] sky130_fd_sc_hd__dfrtp_1
X_3026_ _1689_ _1704_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3928_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[24\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload5 clknet_leaf_30_CLK VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_6
X_3859_ clknet_leaf_12_CLK _0085_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3893__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2190_ net333 net52 net86 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
XFILLER_65_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1974_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1465_ VGND VGND VPWR VPWR _1467_
+ sky130_fd_sc_hd__or2_1
X_3713_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1285_ _1286_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\]
+ _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3920__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3644_ _1216_ _1225_ _1226_ _1227_ _1212_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a32o_1
X_3575_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\]
+ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__nand2b_1
X_2526_ _1747_ _1749_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__and3b_1
X_2457_ net121 VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__inv_2
Xhold28 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[6\] VGND VGND VPWR VPWR net231
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold17 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[15\] VGND VGND VPWR VPWR net220
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 _0109_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
X_2388_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] VGND VGND VPWR VPWR
+ _1614_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4058_ clknet_leaf_4_CLK _0250_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_2
X_3009_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__nor2_1
XFILLER_71_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout72_X net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2524__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2569__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3360_ _0936_ _0937_ _0942_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__and4_1
X_2311_ net324 net36 net76 VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ _1681_ _0873_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__xnor2_1
X_2242_ net324 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] net96 VGND
+ VGND VPWR VPWR _0141_ sky130_fd_sc_hd__mux2_1
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2173_ net317 net65 net84 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1957_ _1350_ _1449_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] VGND VGND VPWR
+ VPWR _1450_ sky130_fd_sc_hd__o21a_1
X_1888_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ _1201_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__and3_1
X_3627_ _1650_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] VGND VGND VPWR
+ VPWR _1211_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3558_ _1141_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__inv_2
X_2509_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] _1619_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ _1620_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__a22oi_1
XANTENNA__2732__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3489_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] _1725_ _1072_ VGND
+ VGND VPWR VPWR _1073_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3842__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2519__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2860_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] _0380_ _0434_ _0438_
+ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__o2111a_1
XFILLER_62_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__inv_2
X_3412_ _1659_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ _1657_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a22o_1
XANTENNA__2190__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3343_ _0533_ _0778_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__xnor2_1
X_3274_ _0583_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__xnor2_2
X_2225_ net301 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\] net103 VGND
+ VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
XFILLER_66_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2156_ net250 net52 net90 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_1
XFILLER_66_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2087_ net326 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] net104 VGND
+ VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2989_ _0571_ _0572_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout122_X net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2103__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2181__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4041__RESET_B net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input52_X net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2540__A1_N _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2172__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2010_ _1643_ _1491_ _1502_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__nand3_1
XFILLER_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ clknet_leaf_6_CLK _0154_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_85_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2912_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__inv_2
XFILLER_92_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3892_ clknet_leaf_12_CLK _0118_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2843_ _1684_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\] VGND VGND VPWR
+ VPWR _0430_ sky130_fd_sc_hd__nand2_1
XFILLER_31_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2774_ net124 _0379_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__and2_1
XANTENNA__2712__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold125 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[52\] VGND VGND VPWR VPWR net328
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[9\] VGND VGND VPWR VPWR net317
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[9\] VGND VGND VPWR VPWR net306
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 myPWM.g_pwm_channel\[1\].CHANNEL.polarity VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dlygate4sd3_1
X_3326_ net124 _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__or2_1
XFILLER_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3257_ _0835_ _0839_ _0840_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__and4b_1
X_2208_ net266 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\] net100 VGND
+ VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
X_3188_ _1671_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] _0485_ VGND
+ VGND VPWR VPWR _0773_ sky130_fd_sc_hd__or3_1
XFILLER_39_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2139_ net327 net65 net88 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__mux2_1
XFILLER_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1977__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2154__A1 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input12_A addr[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3628__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_99_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2490_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\] VGND VGND VPWR VPWR
+ _1716_ sky130_fd_sc_hd__inv_2
XFILLER_99_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2145__A1 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3111_ _0486_ _0566_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3042_ _1696_ _1700_ _0474_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__o21a_1
XANTENNA__3645__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3944_ clknet_leaf_32_CLK _0137_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_3875_ clknet_leaf_23_CLK _0101_ net155 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_2
X_2826_ net119 net118 _0413_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__and3_1
XFILLER_31_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2757_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0369_ net72 VGND VGND VPWR
+ VPWR _0371_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2688_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] _1781_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[5\]
+ _1612_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__o221a_1
XANTENNA__2136__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A addr[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1895__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3309_ _0492_ _0494_ _0892_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ _1671_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__o32a_1
XFILLER_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout86 net87 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_4
Xfanout75 _1773_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
Xfanout97 net99 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpwm_wrapper_197 VGND VGND VPWR VPWR pwm_wrapper_197/HI rdata[26] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_186 VGND VGND VPWR VPWR pwm_wrapper_186/HI rdata[15] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_175 VGND VGND VPWR VPWR pwm_wrapper_175/HI rdata[4] sky130_fd_sc_hd__conb_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_8_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1990_ _1084_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__xnor2_1
X_3660_ _1063_ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__nor2_1
X_3591_ _1171_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and2b_1
Xclkload23 clknet_leaf_22_CLK VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__clkinv_8
X_2611_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1816_ VGND VGND VPWR VPWR
+ _1818_ sky130_fd_sc_hd__and2_1
Xclkload12 clknet_leaf_3_CLK VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__bufinv_16
X_2542_ _1639_ net113 _1642_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] VGND VGND
+ VPWR VPWR _1768_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2201__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2473_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR _1699_
+ sky130_fd_sc_hd__inv_2
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4074_ clknet_leaf_21_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\] net155
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] sky130_fd_sc_hd__dfrtp_1
X_3025_ _0606_ _0608_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nand2_1
XFILLER_55_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3927_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[23\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_34_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3858_ clknet_leaf_12_CLK _0084_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload6 clknet_leaf_31_CLK VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_4
XFILLER_50_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3789_ clknet_leaf_10_CLK _0016_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_2809_ net121 _0402_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] VGND VGND VPWR
+ VPWR _0406_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2109__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2942__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1973_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] _1462_ _1465_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\]
+ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__a22o_1
X_3712_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] _1286_ _1287_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\]
+ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_31_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3643_ _1649_ _1214_ _1213_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__o21ai_1
X_3574_ _1122_ _1129_ _1143_ _1151_ _1157_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__a2111o_1
X_2525_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] _1610_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\]
+ _1632_ _1750_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__o221a_1
X_2456_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND VPWR VPWR
+ _1682_ sky130_fd_sc_hd__inv_2
Xhold18 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[63\] VGND VGND VPWR VPWR net221
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[11\] VGND VGND VPWR VPWR net232
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2387_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4057_ clknet_leaf_5_CLK _0249_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3008_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__nand2_1
XFILLER_64_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout152_X net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2106__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ net121 _0871_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__nand2_1
X_2310_ net243 net35 net76 VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
X_2241_ net243 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] net96 VGND
+ VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_1
XFILLER_78_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2172_ net280 net64 net84 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1956_ _1345_ _1349_ _1113_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__a21oi_1
X_1887_ _1375_ _1376_ _1378_ _1379_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__and4bb_1
X_3626_ _1052_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_34_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_34_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3557_ _1139_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__and2_1
X_2508_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] _1638_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\]
+ _1646_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__o221a_1
XANTENNA__2732__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3488_ _1069_ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__nor2_1
XFILLER_69_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2439_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] VGND VGND VPWR VPWR _1665_
+ sky130_fd_sc_hd__inv_2
XFILLER_84_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_33_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_25_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_4_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input42_A wdata[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\]
+ _0389_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__and3_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_16_CLK sky130_fd_sc_hd__clkbuf_8
X_3411_ _1680_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] _0992_ _0994_
+ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__o221a_1
XFILLER_98_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3342_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0925_ _0926_ net109 VGND VGND
+ VPWR VPWR _0927_ sky130_fd_sc_hd__o22ai_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3273_ _0573_ _0857_ _0767_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o21a_1
X_2224_ net275 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] net103 VGND
+ VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
X_2155_ net332 net51 net90 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_1
XFILLER_93_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ net320 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] net104 VGND
+ VGND VPWR VPWR _0003_ sky130_fd_sc_hd__mux2_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2988_ _0571_ _0572_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and2_1
XFILLER_21_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1939_ _1132_ _1364_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout115_X net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3609_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__or2_1
XFILLER_1_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input45_X net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_5_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_63_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3960_ clknet_leaf_4_CLK _0153_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2911_ _0489_ _0495_ _0492_ _0486_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or4bb_2
X_3891_ clknet_leaf_12_CLK _0117_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_2
X_2842_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[23\]
+ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__xor2_1
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2773_ net124 _0379_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__nor2_1
XANTENNA__2204__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold115 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[62\] VGND VGND VPWR VPWR net318
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[55\] VGND VGND VPWR VPWR net329
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[48\] VGND VGND VPWR VPWR net307
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold137 myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[0\] VGND VGND VPWR VPWR net340
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3325_ _0509_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__xnor2_1
X_3256_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0832_ VGND VGND VPWR VPWR
+ _0841_ sky130_fd_sc_hd__nand2_1
XFILLER_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2207_ net278 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] net100 VGND
+ VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_1
X_3187_ _0771_ _0505_ _0509_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__and3b_1
X_2138_ net308 net64 net88 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_1
X_2069_ _1635_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] _1561_ VGND
+ VGND VPWR VPWR _1562_ sky130_fd_sc_hd__a21bo_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout92_A _1597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2090__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3110_ _0646_ _0654_ _0662_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or4b_2
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3041_ _0623_ _0625_ _0476_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3914__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3943_ clknet_leaf_32_CLK _0136_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_3874_ clknet_leaf_23_CLK _0100_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2723__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2825_ net118 _0414_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__nor2_1
XFILLER_8_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2756_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0365_ VGND VGND VPWR VPWR _0370_
+ sky130_fd_sc_hd__and4_1
X_2687_ _1612_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[1\]
+ _1605_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3308_ _0492_ _0494_ _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__or3_1
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3239_ _0473_ _0638_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__and3_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout76 net79 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_4
Xfanout87 _1590_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_4
Xfanout98 net99 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_20_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpwm_wrapper_187 VGND VGND VPWR VPWR pwm_wrapper_187/HI rdata[16] sky130_fd_sc_hd__conb_1
XFILLER_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xpwm_wrapper_176 VGND VGND VPWR VPWR pwm_wrapper_176/HI rdata[5] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_198 VGND VGND VPWR VPWR pwm_wrapper_198/HI rdata[27] sky130_fd_sc_hd__conb_1
XFILLER_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload13 clknet_leaf_4_CLK VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__bufinv_16
X_3590_ _1172_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2_2
Xclkload24 clknet_leaf_23_CLK VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_6
X_2610_ _1817_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[19\]
+ sky130_fd_sc_hd__inv_2
X_2541_ _1621_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] _1629_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\]
+ _1766_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_93_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2472_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND VPWR VPWR
+ _1698_ sky130_fd_sc_hd__inv_2
XFILLER_68_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4073_ clknet_leaf_1_CLK _0265_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.alignment
+ sky130_fd_sc_hd__dfrtp_1
X_3024_ _0605_ _0607_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__nor2_1
XFILLER_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout142_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3926_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[22\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2453__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3857_ clknet_leaf_9_CLK _0083_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload7 clknet_leaf_33_CLK VGND VGND VPWR VPWR clkload7/X sky130_fd_sc_hd__clkbuf_8
X_3788_ clknet_leaf_19_CLK _0015_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_2808_ _0405_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[21\]
+ sky130_fd_sc_hd__inv_2
X_2739_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] _1685_ _1690_ net119
+ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__o221a_1
XANTENNA__3284__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1868__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2293__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2302__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2284__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2036__A1 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1972_ _1121_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__xnor2_1
X_3711_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1287_ _1288_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\]
+ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3642_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1224_ VGND VGND VPWR VPWR
+ _1226_ sky130_fd_sc_hd__or2_1
X_3573_ _1154_ _1155_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__or2_1
XANTENNA__2212__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2524_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\]
+ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__xnor2_1
XFILLER_88_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2455_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR _1681_
+ sky130_fd_sc_hd__inv_2
Xhold19 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[62\] VGND VGND VPWR VPWR net222
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2386_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND VPWR VPWR
+ _1612_ sky130_fd_sc_hd__inv_2
XANTENNA__3551__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4056_ clknet_leaf_6_CLK _0248_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3007_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and2_1
XANTENNA__2275__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout145_X net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3909_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[5\] net133
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_7_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2266__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3758__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2240_ net306 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] net96 VGND VGND
+ VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2171_ net282 net63 net84 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_65_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2257__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2207__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1955_ _1092_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__xnor2_1
X_1886_ _1059_ _1202_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__nor2_1
X_3625_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] _1718_ _1207_ _1208_
+ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_8_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3556_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout105_A _1574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2507_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] _1624_ _1645_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__o22a_1
X_3487_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\]
+ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__nand2b_1
X_2438_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND VPWR VPWR
+ _1664_ sky130_fd_sc_hd__inv_2
XFILLER_69_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2369_ myPWM.g_pwm_channel\[0\].CHANNEL.alignment net56 _1598_ VGND VGND VPWR VPWR
+ _0262_ sky130_fd_sc_hd__mux2_1
XFILLER_84_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4039_ clknet_leaf_31_CLK _0231_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_71_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input35_A wdata[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3410_ _1681_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND VPWR
+ VPWR _0995_ sky130_fd_sc_hd__or2_1
XFILLER_98_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3341_ _0528_ _0782_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3272_ _0587_ _0856_ _0765_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__a21boi_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2223_ net250 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\] net102 VGND
+ VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
X_2154_ net261 net50 net90 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
XFILLER_93_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2085_ net289 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] net105 VGND
+ VGND VPWR VPWR _0002_ sky130_fd_sc_hd__mux2_1
XANTENNA__2650__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2987_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__nand2_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] _1428_ _1430_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\]
+ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__o22a_1
X_1869_ _1147_ _1150_ _1361_ _1359_ _1144_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__o311a_1
X_3608_ _1642_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] VGND VGND VPWR
+ VPWR _1192_ sky130_fd_sc_hd__nor2_1
XFILLER_89_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3539_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\]
+ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__nand2b_1
XFILLER_88_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4050__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2310__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input38_X net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2910_ _0493_ _0494_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__nor2_2
X_3890_ clknet_leaf_12_CLK _0116_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2841_ _1698_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\] VGND VGND VPWR
+ VPWR _0428_ sky130_fd_sc_hd__nand2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2772_ _0380_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[10\]
+ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_32_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold116 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[53\] VGND VGND VPWR VPWR net319
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold105 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[40\] VGND VGND VPWR VPWR net308
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[25\] VGND VGND VPWR VPWR net330
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 myPWM.g_pwm_channel\[1\].CHANNEL.alignment VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2220__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3324_ _0505_ _0890_ _0776_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a21bo_1
X_3255_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0834_ VGND VGND VPWR VPWR
+ _0840_ sky130_fd_sc_hd__nand2_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2206_ myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[41\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ net100 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_1
X_3186_ _0493_ _0770_ _0494_ _0489_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__or4b_1
XFILLER_93_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2137_ net325 net63 net88 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2456__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2068_ _1532_ _1540_ _1541_ _1537_ _1539_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__a32o_1
XFILLER_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2462__Y _1688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2130__S net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A _1590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_71_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2305__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3040_ _0617_ _0619_ _0624_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND VPWR VPWR _0625_
+ sky130_fd_sc_hd__a32o_1
XFILLER_48_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3942_ clknet_leaf_32_CLK _0135_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__2605__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3873_ clknet_leaf_22_CLK _0099_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2215__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2824_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[26\] VGND VGND VPWR VPWR
+ _0416_ sky130_fd_sc_hd__inv_2
X_2755_ _0362_ _0368_ _0369_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[4\]
+ sky130_fd_sc_hd__nor3_1
X_2686_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] _1778_ _1783_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\]
+ _0287_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__o221a_1
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3307_ _0489_ _0891_ _0775_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__a21boi_1
X_3238_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] _1700_ _0477_ _0821_
+ _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__a221o_1
XFILLER_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3169_ _0654_ _0659_ _0660_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__or3b_1
XFILLER_66_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout88 _1588_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_4
Xfanout99 _1592_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
Xfanout77 net79 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_20_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpwm_wrapper_177 VGND VGND VPWR VPWR pwm_wrapper_177/HI rdata[6] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_188 VGND VGND VPWR VPWR pwm_wrapper_188/HI rdata[17] sky130_fd_sc_hd__conb_1
XANTENNA_fanout88_X net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2532__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xpwm_wrapper_199 VGND VGND VPWR VPWR pwm_wrapper_199/HI rdata[28] sky130_fd_sc_hd__conb_1
XFILLER_18_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2063__A2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload14 clknet_leaf_5_CLK VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload25 clknet_leaf_24_CLK VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__inv_6
X_2540_ _1639_ net113 _1650_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND
+ VPWR VPWR _1766_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_93_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2471_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] VGND VGND VPWR VPWR _1697_
+ sky130_fd_sc_hd__inv_2
XFILLER_5_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2523__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3079__A1 _0564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4072_ clknet_leaf_1_CLK _0264_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.polarity
+ sky130_fd_sc_hd__dfrtp_1
X_3023_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__or2_1
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3925_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[21\] net136
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout135_A net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3856_ clknet_leaf_10_CLK _0082_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload8 clknet_leaf_34_CLK VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__inv_6
XANTENNA__3565__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3787_ clknet_leaf_18_CLK _0014_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_2807_ net121 _0402_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a21o_1
X_2738_ _1652_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] _1656_ net109
+ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__o22a_1
XFILLER_59_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2669_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[13\]
+ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__and2_1
XFILLER_86_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3801__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_516 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3805__RESET_B net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input65_A wdata[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3194__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3233__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1971_ _1118_ _1344_ _1352_ _1115_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__a31o_1
X_3710_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1288_ _1291_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\]
+ _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_31_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3641_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1218_ _1224_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__a22o_1
X_3572_ _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__inv_2
X_2523_ _1629_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\]
+ _1647_ _1748_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__o221a_1
X_2454_ net122 VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__inv_2
X_2385_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__inv_2
Xinput1 addr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4055_ clknet_leaf_5_CLK _0247_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_67_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3006_ _0589_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__nand2_2
XFILLER_91_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2464__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3908_ clknet_leaf_30_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[4\] net132
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3839_ clknet_leaf_21_CLK _0065_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2735__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4075__RESET_B net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2313__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2170_ net331 net62 net84 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
XFILLER_65_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1954_ _1113_ _1345_ _1349_ _1111_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a31o_1
XANTENNA__2223__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1885_ _1189_ _1195_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__nor2_1
X_3624_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] _1718_ _1719_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\]
+ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__a22o_1
XANTENNA__2193__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3555_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__nand2_1
X_3486_ _1066_ _1068_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2506_ _1614_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] _1633_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\]
+ _1731_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__o221a_1
XFILLER_69_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2437_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__inv_2
X_2368_ net338 net45 _1598_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
X_2299_ _1587_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__and2_1
X_4038_ clknet_leaf_31_CLK _0230_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3445__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_71_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2922__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2133__S net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2708__B1 _1682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2184__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout70_X net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3684__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_101_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input28_A addr[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2308__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2175__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3340_ _0531_ _0780_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__xnor2_1
XFILLER_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1922__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3271_ _0803_ _0810_ _0577_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a21oi_1
X_2222_ net332 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\] net102 VGND
+ VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2153_ net269 net49 net91 VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_1
XFILLER_19_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_6_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2084_ net290 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] net105 VGND
+ VGND VPWR VPWR _0001_ sky130_fd_sc_hd__mux2_1
XANTENNA__2218__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2986_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2_1
X_1937_ _1142_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__xnor2_1
X_1868_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__a21oi_1
X_3607_ _1075_ _1185_ _1186_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__a211oi_1
XANTENNA__2166__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3538_ _1109_ _1118_ _1121_ _1114_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__or4b_2
XFILLER_88_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3469_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nand2_1
XFILLER_69_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2157__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3483__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2827__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2840_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0424_ _0427_ VGND VGND VPWR
+ VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\] sky130_fd_sc_hd__o21ba_1
X_2771_ net69 _0378_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or3_2
Xhold117 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[3\] VGND VGND VPWR VPWR net320
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold106 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[1\] VGND VGND VPWR VPWR net309
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_96_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2148__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold128 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[6\] VGND VGND VPWR VPWR net331
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3323_ _0896_ _0902_ _0905_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and4_1
XFILLER_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3254_ net118 _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__nand2_1
X_2205_ net308 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\] net100 VGND
+ VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_1
XANTENNA__2320__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3185_ _0486_ _0492_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__or2_1
XFILLER_81_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2136_ net335 net62 net89 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_1
XFILLER_93_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2067_ _1511_ _1530_ _1531_ _1559_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__a31o_1
XFILLER_54_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2472__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2969_ _0510_ _0513_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__nand2_1
XANTENNA__2139__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3804__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3639__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout78_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2311__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3478__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2321__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input50_X net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2302__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3941_ clknet_leaf_32_CLK _0134_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_90_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3872_ clknet_leaf_21_CLK _0098_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_2
X_2823_ _0414_ _0415_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[26\]
+ sky130_fd_sc_hd__nor2_1
X_2754_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\]
+ _0365_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and3_1
XANTENNA__2369__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2685_ _0279_ _0281_ _0282_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__or4_1
XANTENNA__2231__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3306_ _0505_ _0509_ _0890_ _0777_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__a31o_1
XANTENNA__2541__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3237_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] _1701_ VGND VGND VPWR
+ VPWR _0822_ sky130_fd_sc_hd__and2_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3168_ _0749_ _0750_ _0752_ _0695_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a31o_1
X_2119_ net18 net17 net20 net19 VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout168_X net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3099_ _0591_ _0663_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__xor2_1
XFILLER_54_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2914__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout89 _1588_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
XFILLER_22_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout78 net79 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2930__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2141__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpwm_wrapper_178 VGND VGND VPWR VPWR pwm_wrapper_178/HI rdata[7] sky130_fd_sc_hd__conb_1
Xpwm_wrapper_189 VGND VGND VPWR VPWR pwm_wrapper_189/HI rdata[18] sky130_fd_sc_hd__conb_1
XFILLER_49_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input10_A addr[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3001__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2316__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_7_CLK VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__clkinv_2
Xclkload26 clknet_leaf_26_CLK VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_93_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2470_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND VPWR VPWR
+ _1696_ sky130_fd_sc_hd__inv_2
XFILLER_5_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4071_ clknet_leaf_29_CLK _0263_ net133 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ sky130_fd_sc_hd__dfrtp_1
X_3022_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__nor2_1
XFILLER_76_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2039__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__2226__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3924_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[20\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload9 clknet_leaf_35_CLK VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__bufinv_16
X_3855_ clknet_leaf_10_CLK _0081_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3786_ clknet_leaf_28_CLK _0013_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout128_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2806_ net121 _0402_ net73 VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__o21ai_1
X_2737_ _1688_ net120 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] _1691_
+ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__o221a_1
X_2668_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[6\]
+ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2599_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ _1806_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__and3_1
XFILLER_101_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A addr[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2136__S net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input58_A wdata[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1970_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1448_ _1462_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\]
+ _1461_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_31_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _1222_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__xnor2_1
X_3571_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__xor2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2522_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] _1628_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\]
+ _1641_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__o22a_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2453_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND VPWR VPWR
+ _1679_ sky130_fd_sc_hd__inv_2
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2384_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__inv_2
XFILLER_83_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4054_ clknet_leaf_5_CLK _0246_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 addr[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3005_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3907_ clknet_leaf_30_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[3\] net132
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] sky130_fd_sc_hd__dfrtp_4
X_3838_ clknet_leaf_15_CLK _0064_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2480__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3769_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[29\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2735__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_28_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1953_ net117 _1442_ _1445_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] VGND VGND
+ VPWR VPWR _1446_ sky130_fd_sc_hd__a22o_1
X_1884_ _1375_ _1376_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_19_CLK sky130_fd_sc_hd__clkbuf_8
X_3623_ _1203_ _1205_ _1206_ _1056_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__o31a_1
XANTENNA__2717__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3554_ _1135_ _1137_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__nor2_1
X_3485_ _1066_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__and2_1
X_2505_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] _1625_ _1627_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__o22a_1
X_2436_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__inv_2
X_2367_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable net34 _1598_ VGND VGND
+ VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
X_2298_ net26 _1576_ _1582_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__and3_1
X_4037_ clknet_leaf_26_CLK _0229_ net131 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3133__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2324__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3270_ net120 _0849_ _0854_ _0844_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__a211oi_1
X_2221_ net261 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\] net103 VGND
+ VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
XFILLER_97_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_8_CLK sky130_fd_sc_hd__clkbuf_8
X_2152_ net284 net48 net90 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2083_ net288 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] net105 VGND
+ VGND VPWR VPWR _0000_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2985_ _0564_ _0567_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a21o_1
XANTENNA__2234__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1936_ _1342_ _1364_ _1367_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__o21a_1
X_1867_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ _1154_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__and3_1
X_3606_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__inv_2
Xinput60 wdata[4] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
X_3537_ _1119_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__and2b_2
X_3468_ _1050_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nand2_1
XFILLER_69_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3399_ net119 _1703_ _1704_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND
+ VPWR VPWR _0984_ sky130_fd_sc_hd__a2bb2o_1
X_2419_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND VPWR VPWR
+ _1645_ sky130_fd_sc_hd__inv_2
XFILLER_29_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2144__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A wdata[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2319__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3004__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2617__B1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2093__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2770_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\]
+ _0375_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__and3_1
Xhold107 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[35\] VGND VGND VPWR VPWR net310
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[57\] VGND VGND VPWR VPWR net332
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[40\] VGND VGND VPWR VPWR net321
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3322_ _0904_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nor2_1
XFILLER_98_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3253_ _0617_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3184_ _0577_ _0766_ _0587_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__or3b_1
X_2204_ net325 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\] net100 VGND
+ VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
X_2135_ net273 net61 net88 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_1
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2066_ _1549_ _1556_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout158_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3568__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2968_ _0548_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nand2_1
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1919_ _1410_ _1411_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR
+ VPWR _1412_ sky130_fd_sc_hd__a21o_1
X_2899_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\]
+ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__and2b_1
XANTENNA__3336__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2139__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2663__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input43_X net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3940_ clknet_leaf_26_CLK _0133_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_51_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3871_ clknet_leaf_22_CLK _0097_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2822_ net119 _0413_ net72 VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__o21ai_1
X_2753_ net109 _0365_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] VGND VGND VPWR
+ VPWR _0368_ sky130_fd_sc_hd__a21oi_1
X_2684_ _0283_ _0300_ _0301_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__or4_1
XFILLER_98_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3305_ _0793_ _0794_ _0795_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a21o_1
XANTENNA__2541__A2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ _0812_ _0814_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__o21bai_2
XFILLER_73_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3167_ net124 _0711_ _0712_ _0751_ _0706_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a221o_1
X_3098_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__inv_2
X_2118_ net9 net8 net11 net10 VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__or4_1
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2049_ net112 _1720_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__nor2_1
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout79 _1596_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout90_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xpwm_wrapper_179 VGND VGND VPWR VPWR pwm_wrapper_179/HI rdata[8] sky130_fd_sc_hd__conb_1
XANTENNA__2658__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2296__A1 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3001__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload16 clknet_leaf_8_CLK VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__inv_6
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2220__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload27 clknet_leaf_28_CLK VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_93_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2523__A2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4070_ clknet_leaf_21_CLK _0262_ net154 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.alignment
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2287__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3021_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nand2_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3923_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[19\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3854_ clknet_leaf_29_CLK _0080_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2805_ _0402_ _0403_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[20\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__2242__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3785_ clknet_leaf_26_CLK _0012_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_2736_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] _1678_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\]
+ _1699_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__o22a_1
X_2667_ _1772_ _1775_ _0286_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_99_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2598_ net74 _1808_ _1809_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[15\]
+ sky130_fd_sc_hd__and3_1
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3219_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\]
+ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2b_1
XANTENNA__2278__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2152__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_68_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout93_X net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2269__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2327__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3570_ _1152_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nand2_1
X_2521_ _1743_ _1744_ _1745_ _1746_ _1742_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__a221o_1
XFILLER_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2452_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR _1678_
+ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2383_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND VPWR VPWR
+ _1609_ sky130_fd_sc_hd__inv_2
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4053_ clknet_leaf_4_CLK _0245_ net136 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3004_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\]
+ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 addr[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2680__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2680__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2237__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3906_ clknet_leaf_29_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[2\] net132
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout140_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3837_ clknet_leaf_15_CLK _0063_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_3768_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_30_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2719_ _1686_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _1688_ net120 _0336_
+ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a221o_1
X_3699_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\] _1282_ VGND VGND VPWR VPWR _1283_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2147__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3007__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2846__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ _1440_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nand2_1
X_1883_ _1341_ _1371_ _1373_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__and3_1
X_3622_ _1059_ _1196_ _1202_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nor2_1
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3484_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__or2_1
X_2504_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] _1615_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ _1620_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__o221a_1
X_2435_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] VGND VGND VPWR VPWR
+ _1661_ sky130_fd_sc_hd__inv_2
XFILLER_69_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2366_ _1589_ _1595_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2297_ net221 net58 net83 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4036_ clknet_leaf_30_CLK _0228_ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_37_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3497__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2340__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2220_ net269 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] net102 VGND
+ VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_1
X_2151_ net319 net47 net90 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
XANTENNA__2883__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2082_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[0\]
+ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__nand2_4
XFILLER_34_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3917__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2984_ _0480_ _0483_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or2_1
XFILLER_61_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1935_ _1133_ _1427_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__xor2_1
X_1866_ _1148_ _1145_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__nand2b_1
Xinput50 wdata[24] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
X_3605_ _1187_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nand2_1
Xinput61 wdata[5] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2250__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_A _1591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3536_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__or2_1
X_3467_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__or2_1
X_2418_ net112 VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__inv_2
X_3398_ _1693_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] VGND VGND VPWR
+ VPWR _0983_ sky130_fd_sc_hd__nor2_1
XFILLER_29_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2349_ net307 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] net94 VGND
+ VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
XANTENNA__2059__A1_N net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4019_ clknet_leaf_3_CLK _0211_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2933__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2160__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input33_A nRST VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2396__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__2865__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3004__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2335__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3020__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold108 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[29\] VGND VGND VPWR VPWR net311
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[20\] VGND VGND VPWR VPWR net322
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_98_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3321_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0900_ _0903_ net123 VGND VGND
+ VPWR VPWR _0906_ sky130_fd_sc_hd__a22o_1
XFILLER_98_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3252_ _0621_ _0836_ _0815_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_13_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3183_ _0765_ _0766_ _0767_ _0581_ _0580_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__o221a_1
X_2203_ net335 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] net101 VGND
+ VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_1
X_2134_ net256 net60 net89 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
XFILLER_66_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2065_ _1532_ _1540_ _1541_ _1557_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__and4b_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2245__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2967_ _0542_ _0544_ _0547_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__a21oi_1
X_1918_ _1076_ _1374_ _1069_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__a21o_1
X_2898_ _0481_ _0482_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nand2_1
X_1849_ _1131_ _1133_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_73_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout106_X net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3519_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__nand2b_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2155__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input36_X net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2854__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3870_ clknet_leaf_14_CLK _0096_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2821_ net119 _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__and2_1
XFILLER_76_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2752_ net109 _0365_ _0367_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[3\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_8_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2683_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[15\]
+ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__xor2_1
XFILLER_98_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3304_ _0843_ _0855_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__and3b_1
X_3235_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] _0816_ _0818_ _0813_
+ _0615_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__a221o_1
XANTENNA__3921__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_100_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3166_ _0715_ _0717_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nand2_1
X_3097_ _0681_ _0677_ _0671_ _0680_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and4b_1
X_2117_ net14 net13 net16 net15 VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__or4_1
X_2048_ _1630_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\] VGND VGND VPWR
+ VPWR _1541_ sky130_fd_sc_hd__nand2_1
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3999_ clknet_leaf_7_CLK _0191_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout69 _0362_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2765__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout83_A _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_9_CLK VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinv_8
Xclkload28 clknet_leaf_13_CLK VGND VGND VPWR VPWR clkload28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2508__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3020_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[58\]
+ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__and2_1
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2584__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3922_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[18\] net136
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[18\] sky130_fd_sc_hd__dfrtp_1
X_3853_ clknet_leaf_1_CLK _0079_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_2804_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] _0400_ net73 VGND VGND VPWR
+ VPWR _0403_ sky130_fd_sc_hd__o21ai_1
X_3784_ clknet_leaf_26_CLK _0011_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_2735_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] _1663_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\]
+ _1693_ _0352_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o221a_1
X_2666_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__or2_1
XFILLER_99_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2597_ net116 _1806_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__nand2_1
XFILLER_99_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3218_ _0796_ _0800_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21o_1
X_3149_ _0531_ _0538_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__xor2_1
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_4_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2941__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2738__B1 _1656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2669__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout86_X net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2343__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2729__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2520_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] net112 VGND VGND VPWR
+ VPWR _1746_ sky130_fd_sc_hd__or2_1
XFILLER_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2451_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND VPWR VPWR
+ _1677_ sky130_fd_sc_hd__inv_2
X_2382_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__inv_2
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4052_ clknet_leaf_3_CLK _0244_ net136 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3003_ _0574_ _0578_ _0582_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_67_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 addr[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3905_ clknet_leaf_1_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[1\] net132
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2253__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3836_ clknet_leaf_14_CLK _0062_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout133_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3767_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[27\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[27\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2718_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] _1663_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\]
+ _1685_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_5_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3698_ _1117_ _1279_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__xnor2_1
X_2649_ _0269_ _0270_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_87_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4053__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2187__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input63_A wdata[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3007__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2111__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3023__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2338__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1951_ _1156_ _1354_ _1355_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__nand3_1
X_1882_ _1070_ _1079_ _1339_ _1341_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__o31a_1
X_3621_ _1075_ _1185_ _1186_ _1204_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a211oi_1
XANTENNA__3776__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3552_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nand2_1
XANTENNA__2178__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1925__A1 _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2503_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\]
+ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__xnor2_1
X_3483_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_1
X_2434_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__inv_2
X_2365_ _1603_ net312 net78 VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__a21o_1
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2296_ net318 net57 net83 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
XANTENNA__2102__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2248__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2638__C1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4035_ clknet_leaf_30_CLK _0227_ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_96_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout136_X net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ clknet_leaf_26_CLK _0045_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2169__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2947__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2158__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3497__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2150_ net328 net46 net90 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
XFILLER_66_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2081_ net339 _1572_ _1573_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.pwm_next
+ sky130_fd_sc_hd__a21oi_1
XFILLER_81_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2592__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2983_ _0564_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__nand2_1
XFILLER_61_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1934_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ _1132_ _1364_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__o2bb2a_1
X_1865_ _1354_ _1355_ _1356_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__a21o_1
Xinput40 wdata[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
Xinput51 wdata[25] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_3604_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__nand2_1
Xinput62 wdata[6] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
X_3535_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__and2_1
XANTENNA__3924__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3466_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nand2_1
X_2417_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] VGND VGND VPWR VPWR _1643_
+ sky130_fd_sc_hd__inv_2
XANTENNA__2323__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3397_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__inv_2
XFILLER_84_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2348_ net239 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] net92 VGND
+ VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
XFILLER_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2279_ net216 net38 net80 VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4018_ clknet_leaf_35_CLK _0210_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2677__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2314__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input26_A addr[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2351__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold109 myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[0\] VGND VGND VPWR VPWR net312
+ sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ _1670_ _0898_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3251_ _0609_ _0613_ _0812_ _0819_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__o31a_1
XANTENNA__2305__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3182_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\]
+ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__nand2b_1
X_2202_ net273 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\] net101 VGND
+ VGND VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2133_ net267 net59 net89 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
XFILLER_66_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2064_ _1533_ _1536_ _1550_ _1551_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__and4b_1
X_2966_ _0517_ _0550_ _0515_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__o21ai_1
X_1917_ _1069_ _1076_ _1374_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nand3_1
X_2897_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__or2_1
XANTENNA__2261__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1848_ _1639_ _1723_ _1338_ _1339_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__o221a_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3518_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__xnor2_2
XFILLER_89_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3449_ _1687_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ _1685_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__o211a_1
XFILLER_94_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2960__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2346__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2820_ net69 _0412_ _0413_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[25\]
+ sky130_fd_sc_hd__nor3_1
X_2751_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[3\] _0365_ net72 VGND VGND VPWR
+ VPWR _0367_ sky130_fd_sc_hd__o21ai_1
X_2682_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] _1796_ VGND VGND VPWR
+ VPWR _0301_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3303_ _0878_ _0881_ _0883_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__and4_1
XFILLER_98_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3234_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__inv_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3165_ _0697_ _0702_ _0704_ _0701_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__o22a_1
XFILLER_81_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3096_ _0678_ _0679_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] VGND VGND VPWR
+ VPWR _0681_ sky130_fd_sc_hd__o21a_1
X_2116_ net27 _1575_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__nor2_1
XFILLER_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2256__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2047_ _1537_ _1538_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout163_A net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3998_ clknet_leaf_7_CLK _0190_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_2949_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__nand2_1
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2765__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout76_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2166__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload29 clknet_leaf_14_CLK VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_6
Xclkload18 clknet_leaf_10_CLK VGND VGND VPWR VPWR clkload18/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__2508__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3921_ clknet_leaf_2_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[17\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] sky130_fd_sc_hd__dfrtp_4
X_3852_ clknet_leaf_30_CLK _0078_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_2803_ net122 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] _0398_ VGND VGND VPWR
+ VPWR _0402_ sky130_fd_sc_hd__and3_1
X_3783_ clknet_leaf_25_CLK _0010_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_2734_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] net110 VGND VGND VPWR
+ VPWR _0352_ sky130_fd_sc_hd__xnor2_1
X_2665_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[4\]
+ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__xnor2_1
X_2596_ net116 _1806_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__or2_1
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3217_ _0801_ _0595_ _0483_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__or3b_1
XANTENNA__2775__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3148_ net109 _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__or2_1
XFILLER_27_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3079_ _0564_ _0567_ _0569_ _0596_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_53_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout79_X net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_74 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2729__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2450_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR _1676_
+ sky130_fd_sc_hd__inv_2
XFILLER_96_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2381_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] VGND VGND VPWR VPWR
+ _1607_ sky130_fd_sc_hd__inv_2
XFILLER_96_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4051_ clknet_leaf_3_CLK _0243_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_4
X_3002_ _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__nand2_2
Xinput5 addr[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3904_ clknet_leaf_1_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[0\] net132
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_51_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3835_ clknet_leaf_13_CLK _0061_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout126_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3766_ clknet_leaf_16_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[26\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] sky130_fd_sc_hd__dfrtp_1
X_2717_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] _1659_ _1689_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\]
+ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__a221o_1
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3697_ _1121_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__xnor2_1
X_2648_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] _0267_ net75 VGND VGND VPWR
+ VPWR _0270_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2579_ net117 _1795_ net74 VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3502__A_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A wdata[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2354__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1950_ _1620_ _1434_ _1435_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__nand3_1
X_1881_ _1371_ _1373_ _1079_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__a21o_1
X_3620_ _1059_ _1189_ _1195_ _1202_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nand4_1
X_3551_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__and2_1
XANTENNA__3182__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2502_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] VGND VGND VPWR VPWR
+ _1728_ sky130_fd_sc_hd__inv_2
X_3482_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__nand2_1
XFILLER_88_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2433_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__inv_2
X_2364_ net221 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\] net95 VGND
+ VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
X_2295_ net314 net55 net83 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
X_4034_ clknet_leaf_8_CLK _0226_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3818_ clknet_leaf_26_CLK _0044_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_3749_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] _1230_ VGND VGND VPWR VPWR
+ _1333_ sky130_fd_sc_hd__or2_1
XFILLER_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2174__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2801__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input59_X net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3034__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2349__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2080_ myPWM.g_pwm_channel\[1\].CHANNEL.polarity _1572_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_49_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2873__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2084__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2982_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ _0497_ _0558_ _0563_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__a221oi_4
X_1933_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] _1423_ _1425_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\]
+ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__a22o_1
X_3603_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__or2_1
Xinput30 addr[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_1864_ _1354_ _1355_ _1356_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__a21oi_1
Xinput52 wdata[26] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_2
Xinput63 wdata[7] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput41 wdata[16] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
X_3534_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__inv_2
XANTENNA__2020__B2 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3465_ _1049_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable _1048_ VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.pwm_next sky130_fd_sc_hd__and3b_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2416_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND VPWR VPWR
+ _1642_ sky130_fd_sc_hd__inv_2
X_3396_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _1700_ _0979_ _0980_ VGND VGND
+ VPWR VPWR _0981_ sky130_fd_sc_hd__a211oi_1
XANTENNA__2259__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3940__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2347_ net298 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] net92 VGND
+ VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2278_ net223 net37 net80 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
XANTENNA__2087__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_4017_ clknet_leaf_3_CLK _0209_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2169__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input19_A addr[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_0__f_CLK_X clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2250__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3250_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0832_ _0834_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__o22ai_1
XFILLER_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3181_ _0574_ _0582_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nand2_1
X_2201_ net256 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] net100 VGND
+ VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_1
XFILLER_78_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2132_ net305 net56 net89 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2063_ _1628_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] _1534_ _1552_
+ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__a2111o_1
XFILLER_47_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2965_ _0521_ _0549_ _0545_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a21oi_1
X_1916_ _1404_ _1408_ net114 VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__a21boi_1
X_2896_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__nand2_1
XANTENNA__2241__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1847_ _1639_ _1723_ _1061_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__a21o_1
XANTENNA__3935__Q myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3760__RESET_B net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3517_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_73_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3448_ _0991_ _0996_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__or3_1
X_3379_ _0843_ _0855_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__and3b_1
XFILLER_85_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_356 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2750_ _0365_ _0366_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[2\]
+ sky130_fd_sc_hd__nor2_1
X_2681_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] _1781_ _1783_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\]
+ _0293_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__a221o_1
XANTENNA__2598__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3302_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] _0885_ _0886_ VGND VGND VPWR
+ VPWR _0887_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3233_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] _1703_ _0817_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\]
+ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a22o_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ _0720_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__or2_1
XFILLER_82_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3095_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0678_ _0679_ VGND VGND VPWR
+ VPWR _0680_ sky130_fd_sc_hd__or3_1
X_2115_ net28 net30 net29 net66 VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__or4b_1
XANTENNA__2764__C myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2046_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1726_ VGND VGND VPWR VPWR
+ _1539_ sky130_fd_sc_hd__or2_1
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout156_A net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3997_ clknet_leaf_6_CLK _0189_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2272__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2948_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_20_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2879_ _1698_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[31\] _0462_ _0463_
+ _0464_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o2111a_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2971__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2182__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload19 clknet_leaf_11_CLK VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__2508__A2 _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input41_X net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2357__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_495 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3920_ clknet_leaf_36_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\]
+ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_17_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3851_ clknet_leaf_26_CLK _0077_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2802_ _0400_ _0401_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__2092__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3782_ clknet_leaf_25_CLK _0009_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2733_ _1654_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _1677_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\]
+ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o221a_1
X_2664_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[9\]
+ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__xnor2_1
X_2595_ _1806_ _1807_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[14\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_59_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3216_ _0480_ _0591_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__nand2_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3147_ _0528_ _0539_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2267__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3078_ _0570_ _0599_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nand2_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2029_ _1618_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ _1617_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1946__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2177__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2380_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__inv_2
XFILLER_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4050_ clknet_leaf_35_CLK _0242_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_3001_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__nand2_1
XANTENNA__2087__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 addr[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3903_ clknet_leaf_16_CLK _0129_ net167 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_mod\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3834_ clknet_leaf_13_CLK _0060_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3765_ clknet_leaf_17_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[25\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3696_ _1117_ _1279_ _1124_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__a21oi_1
X_2716_ _1656_ net109 _1669_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] VGND VGND
+ VPWR VPWR _0334_ sky130_fd_sc_hd__a22o_1
X_2647_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\]
+ _1840_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__and3_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2578_ _1796_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[8\]
+ sky130_fd_sc_hd__inv_2
XFILLER_99_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4062__RESET_B net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout91_X net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input49_A wdata[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1880_ _1083_ _1089_ _1370_ _1372_ _1082_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__o221a_1
X_3550_ _1131_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__or2_1
X_2501_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\] VGND VGND VPWR VPWR
+ _1727_ sky130_fd_sc_hd__inv_2
X_3481_ _1060_ _1063_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or2_1
X_2432_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND VPWR VPWR
+ _1658_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2363_ net318 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] net95 VGND
+ VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
XFILLER_96_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4033_ clknet_leaf_7_CLK _0225_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_2294_ net285 net54 net83 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3230__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3817_ clknet_leaf_25_CLK _0043_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3748_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1218_ VGND VGND VPWR VPWR
+ _1332_ sky130_fd_sc_hd__nor2_1
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2280__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3679_ _1091_ _1181_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2801__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2190__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2981_ _0492_ _0565_ _0490_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__a21bo_1
XANTENNA__3758__Q myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_1932_ _1179_ _1424_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__xor2_1
X_1863_ _1154_ _1155_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__nand2_1
X_3602_ _1075_ _1080_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__and2_1
Xinput20 addr[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 addr[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput53 wdata[27] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput42 wdata[17] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xinput64 wdata[8] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_0_CLK_A CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3533_ _1115_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__or2_1
X_3464_ _1717_ _0973_ _1047_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__and3_1
X_2415_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] VGND VGND VPWR VPWR _1641_
+ sky130_fd_sc_hd__inv_2
X_3395_ _1697_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] _1701_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a22o_1
X_2346_ net216 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\] net92 VGND
+ VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2277_ net233 net36 net80 VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
X_4016_ clknet_leaf_35_CLK _0208_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2128__X _1588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2275__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2185__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_CLK_A clknet_2_1__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2538__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2200_ net267 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\] net101 VGND
+ VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_1
X_3180_ _1684_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] _0764_ _1682_
+ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__o22a_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2131_ net260 net45 net89 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
XFILLER_39_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2710__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2062_ _1635_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] _1542_ _1553_
+ _1554_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__a2111o_1
XANTENNA__2069__A2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2095__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2964_ _0525_ _0542_ _0522_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ _1070_ _1374_ _1338_ _1064_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__o211ai_1
XANTENNA__2777__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2895_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nand2_2
X_1846_ _1060_ _1063_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__nand2_1
XFILLER_89_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3516_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout101_A _1591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ _1027_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__nor2_1
X_3378_ _0878_ _0959_ _0961_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__a211o_1
X_2329_ net311 net55 net78 VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
XFILLER_57_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1991__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1991__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input31_A addr[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2759__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2680_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] _1836_ _0266_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\]
+ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o221a_1
XFILLER_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3301_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0882_ _0885_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__o22ai_1
X_3232_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[57\] _0609_ VGND VGND VPWR
+ VPWR _0817_ sky130_fd_sc_hd__nor2_1
XFILLER_67_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3163_ _0731_ _0747_ _0745_ _0724_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__o2bb2a_1
X_2114_ net247 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] net107 VGND
+ VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_1
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3094_ _0572_ _0668_ _0582_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__a21oi_1
X_2045_ _1632_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\] VGND VGND VPWR
+ VPWR _1538_ sky130_fd_sc_hd__nand2_1
XFILLER_35_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3996_ clknet_leaf_6_CLK _0188_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\]
+ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2878_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[29\]
+ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout104_X net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3910__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2150__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3650__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input34_X net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2141__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2373__S _1599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3850_ clknet_leaf_26_CLK _0076_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3781_ clknet_leaf_25_CLK _0008_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_2801_ net122 _0398_ net73 VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o21ai_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2732_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] _1655_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\]
+ _1697_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o22a_1
X_2663_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[10\]
+ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__xor2_1
X_2594_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1805_ net74 VGND VGND VPWR
+ VPWR _1807_ sky130_fd_sc_hd__o21ai_1
XFILLER_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3215_ _0772_ _0793_ _0794_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a31oi_2
XFILLER_86_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2132__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3146_ _0723_ _0724_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__nor3_1
XFILLER_39_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3077_ _0655_ _0659_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__nand4_1
XFILLER_82_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2028_ _1617_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ _1615_ _1520_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_53_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2283__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3979_ clknet_leaf_32_CLK _0171_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2371__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2039__A2_N myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2193__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2114__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2368__S _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3000_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__or2_1
Xinput7 addr[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3902_ clknet_leaf_15_CLK _0128_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_3833_ clknet_leaf_13_CLK _0059_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3764_ clknet_leaf_17_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[24\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3695_ _1110_ _1114_ _1127_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a21o_1
X_2715_ _0329_ _0330_ _0331_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a22o_1
X_2646_ _0267_ _0268_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2353__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2577_ net70 _1794_ _1795_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__or3_1
XFILLER_99_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2278__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2105__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_66_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3129_ _0501_ _0707_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_38_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3410__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout84_X net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2188__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3480_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__inv_2
X_2500_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR VPWR
+ _1726_ sky130_fd_sc_hd__inv_2
X_2431_ net109 VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__inv_2
XANTENNA__2887__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2362_ net314 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\] net95 VGND
+ VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2293_ net252 net53 net83 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
XANTENNA__2098__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4032_ clknet_leaf_7_CLK _0224_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3816_ clknet_leaf_25_CLK _0042_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout131_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ _1233_ _1236_ _1239_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__and4b_1
XFILLER_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3678_ _1252_ _1255_ _1256_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__or4b_1
XANTENNA__2326__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2629_ _1641_ _1828_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__and2_1
XFILLER_99_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_83_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input61_A wdata[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2317__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_92_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2980_ _0489_ _0495_ _0559_ _0561_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__o31ai_1
X_1931_ _1172_ _1421_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__nand2_1
X_1862_ _1115_ _1120_ _1119_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__a21oi_2
X_3601_ _1087_ _1182_ _1184_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_12_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput10 addr[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 addr[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput54 wdata[28] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
Xinput43 wdata[18] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput32 addr[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput65 wdata[9] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_2
X_3532_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nor2_1
XANTENNA__2308__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3463_ _0973_ _1047_ _1717_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__a21o_1
XANTENNA__3506__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2414_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND VPWR VPWR
+ _1640_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_30_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_30_CLK sky130_fd_sc_hd__clkbuf_8
X_3394_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\]
+ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__and2b_1
XFILLER_96_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2345_ net223 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\] net92 VGND
+ VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
XFILLER_84_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2276_ net315 net35 net80 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
X_4015_ clknet_leaf_34_CLK _0207_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3949__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2291__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_X net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_21_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2990__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input64_X net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_12_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_3_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2130_ net224 net34 net89 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux2_1
XFILLER_39_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2061_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1722_ VGND VGND VPWR VPWR
+ _1554_ sky130_fd_sc_hd__nor2_1
XFILLER_19_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2963_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\]
+ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__nand2_1
X_1914_ _1405_ _1406_ _1638_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2405__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2894_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__or2_1
X_1845_ _1066_ _1076_ _1067_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__a21o_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3515_ _1096_ _1097_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__or2_1
XFILLER_89_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3446_ _0991_ _0993_ _1029_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__or4_1
XFILLER_97_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3377_ _0862_ _0874_ _0875_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__and3_1
X_2328_ net214 net54 net78 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_1
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2286__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2259_ net214 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] net98 VGND
+ VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
XFILLER_72_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A addr[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_1_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_8_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3300_ _0863_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__or2_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3231_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\] _0616_ VGND VGND VPWR
+ VPWR _0816_ sky130_fd_sc_hd__nor2_1
X_3162_ _0739_ _0742_ _0744_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__a211o_1
XFILLER_39_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2113_ net248 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] net107 VGND
+ VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
XFILLER_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3093_ _0572_ _0582_ _0668_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__and3_1
XFILLER_81_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2044_ _1632_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[50\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\]
+ _1726_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3995_ clknet_leaf_6_CLK _0187_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2946_ _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__nand2_1
XFILLER_50_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3411__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2877_ _1692_ _0419_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_20_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3962__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3175__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3429_ net123 _1709_ _1710_ net124 VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_1_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3604__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3780_ clknet_leaf_25_CLK _0007_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2800_ net122 _0398_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and2_1
X_2731_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] _1665_ _1694_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a221o_1
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2662_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] _1817_ VGND VGND VPWR
+ VPWR _0282_ sky130_fd_sc_hd__and2_1
XANTENNA__3782__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2593_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1801_ VGND VGND VPWR VPWR _1806_
+ sky130_fd_sc_hd__and4_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3214_ _0484_ _0773_ _0798_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__nand3b_1
XFILLER_67_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3145_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] _0728_ _0729_ _0726_ VGND VGND
+ VPWR VPWR _0730_ sky130_fd_sc_hd__a211o_1
XANTENNA__1891__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3076_ net120 _0657_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__nand2_1
X_2027_ _1615_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ _1613_ _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__a221o_1
XFILLER_42_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout161_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3957__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3978_ clknet_leaf_32_CLK _0170_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2929_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\]
+ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_33_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 addr[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1873__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3901_ clknet_leaf_15_CLK _0127_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__2822__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3777__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3832_ clknet_leaf_13_CLK _0058_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3763_ clknet_leaf_17_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[23\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2413__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3694_ _1161_ _1273_ _1134_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a21o_1
X_2714_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or2_1
X_2645_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1840_ net75 VGND VGND VPWR
+ VPWR _0268_ sky130_fd_sc_hd__o21ai_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2576_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1791_ VGND VGND VPWR VPWR _1795_
+ sky130_fd_sc_hd__and2_1
XFILLER_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3128_ net124 _0711_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__nand2_1
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2294__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0637_ _0643_ VGND VGND VPWR
+ VPWR _0644_ sky130_fd_sc_hd__a21oi_1
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2813__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout77_X net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2804__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4071__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2280__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2430_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] VGND VGND VPWR VPWR
+ _1656_ sky130_fd_sc_hd__inv_2
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2361_ net285 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] net94 VGND
+ VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
XFILLER_96_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2292_ net249 net52 net83 VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_96_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4031_ clknet_leaf_7_CLK _0223_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2408__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2271__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3815_ clknet_leaf_25_CLK _0041_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3746_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1235_ _1238_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\]
+ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__o22a_1
XFILLER_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3677_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] _1254_ _1260_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\]
+ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_76_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2628_ _1830_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[24\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__2797__B myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2289__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2559_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1779_ _1782_ VGND VGND VPWR
+ VPWR _1783_ sky130_fd_sc_hd__a21o_1
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input54_A wdata[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2199__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3969__D myPWM.g_pwm_channel\[1\].CHANNEL.pwm_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2253__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3450__B1 _0990_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1930_ _1421_ _1422_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__nand2_1
X_1861_ _1118_ _1121_ _1344_ _1352_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__nand4_4
X_3600_ _1158_ _1170_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_12_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 addr[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 addr[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput44 wdata[19] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput55 wdata[29] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput33 nRST VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
X_3531_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__and2_1
Xinput66 wen VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
X_3462_ _1036_ _1040_ _1041_ _1046_ myPWM.g_pwm_channel\[0\].CHANNEL.alignment VGND
+ VGND VPWR VPWR _1047_ sky130_fd_sc_hd__a311o_1
X_3393_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _1704_ _1705_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\]
+ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__o22a_1
X_2413_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND VPWR VPWR
+ _1639_ sky130_fd_sc_hd__inv_2
XFILLER_97_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2344_ net233 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\] net92 VGND
+ VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
XFILLER_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2275_ net219 net65 net80 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
X_4014_ clknet_leaf_33_CLK _0206_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2244__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3965__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3744__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3729_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] _1309_ _1310_ _1307_ _1312_
+ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__o221a_1
XFILLER_79_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2235__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input57_X net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2060_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] _1721_ VGND VGND VPWR VPWR
+ _1553_ sky130_fd_sc_hd__nor2_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2962_ _0545_ _0546_ _0514_ _0516_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o211a_1
X_1913_ _1060_ _1061_ _1404_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__nand3b_1
XFILLER_15_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3785__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2893_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__nand2_1
X_1844_ _1231_ _1334_ _1336_ _1335_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__a31o_1
XANTENNA__3726__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3514_ _1096_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nor2_1
XFILLER_89_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3445_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _1707_ _1708_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\]
+ _0992_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__a221o_1
X_3376_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0859_ _0960_ _1685_ VGND VGND
+ VPWR VPWR _0961_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_97_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2327_ net226 net53 net78 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
XFILLER_69_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2258_ net226 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] net98 VGND
+ VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
XFILLER_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2189_ net330 net51 net86 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_1
XFILLER_25_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2217__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A addr[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3337__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3230_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] _1702_ VGND VGND VPWR
+ VPWR _0815_ sky130_fd_sc_hd__nand2_1
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2695__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3161_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0734_ _0736_ _0733_ VGND VGND
+ VPWR VPWR _0746_ sky130_fd_sc_hd__o31ai_1
XFILLER_39_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2112_ net230 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] net107 VGND
+ VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_1
XFILLER_66_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3092_ _0674_ _0675_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__and3_1
XFILLER_81_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2043_ _1535_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__inv_2
XANTENNA__2416__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3994_ clknet_leaf_4_CLK _0186_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2945_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or2_1
X_2876_ _0430_ _0456_ _0460_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_20_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3428_ _1665_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ _1663_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__o22a_1
XANTENNA__2297__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A addr[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3359_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] _0941_ _0939_ VGND VGND VPWR
+ VPWR _0944_ sky130_fd_sc_hd__a21oi_1
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2686__B2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2332__Y _1597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2730_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\]
+ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__xor2_1
X_2661_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] _1817_ VGND VGND VPWR
+ VPWR _0281_ sky130_fd_sc_hd__nor2_1
X_2592_ net70 _1804_ _1805_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[13\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__2365__B1 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3213_ _0507_ _0776_ _0797_ _0771_ _0506_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__a311o_1
XFILLER_67_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3144_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0725_ _0728_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__o22ai_1
X_3075_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0658_ VGND VGND VPWR VPWR
+ _0660_ sky130_fd_sc_hd__nand2_1
X_2026_ _1613_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ _1611_ _1518_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_53_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout154_A net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3977_ clknet_leaf_32_CLK _0169_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2928_ _0511_ _0512_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__and2_2
XFILLER_31_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2859_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[1\]
+ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_79_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3387__A2 _0758_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3841__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput9 addr[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3900_ clknet_leaf_14_CLK _0126_ net166 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3831_ clknet_leaf_12_CLK _0057_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3762_ clknet_leaf_17_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\]
+ net163 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_0_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3793__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3509__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3693_ _1164_ _1275_ _1133_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a21bo_1
X_2713_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\]
+ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__nand2_1
X_2644_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1840_ VGND VGND VPWR VPWR
+ _0267_ sky130_fd_sc_hd__and2_1
X_2575_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1791_ VGND VGND VPWR VPWR _1794_
+ sky130_fd_sc_hd__nor2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3127_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0709_ _0711_ net124 VGND VGND
+ VPWR VPWR _0712_ sky130_fd_sc_hd__o22a_1
XFILLER_82_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3058_ _0640_ _0641_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] VGND VGND VPWR
+ VPWR _0643_ sky130_fd_sc_hd__o21a_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2009_ _1059_ _1382_ _1490_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__nand3_1
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2163__X _1590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2514__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_CLK_X clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4040__RESET_B net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2360_ net252 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\] net95 VGND
+ VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_69_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2291_ net234 net51 net83 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4030_ clknet_leaf_7_CLK _0222_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3296__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3814_ clknet_leaf_25_CLK _0040_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3745_ _1264_ _1328_ _1262_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3676_ _1084_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_76_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2627_ _1828_ _1829_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__nand2_1
XANTENNA__2430__Y _1656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2558_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1779_ net74 VGND VGND VPWR
+ VPWR _1782_ sky130_fd_sc_hd__o21ai_1
X_2489_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\] VGND VGND VPWR VPWR
+ _1715_ sky130_fd_sc_hd__inv_2
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3039__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A wdata[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ _1344_ _1352_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 addr[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput23 addr[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
X_3530_ _1092_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__nor2_1
Xinput45 wdata[1] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput34 wdata[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput56 wdata[2] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_4
X_3461_ _0988_ _1022_ _1031_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nor4_1
X_2412_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] VGND VGND VPWR VPWR _1638_
+ sky130_fd_sc_hd__inv_2
X_3392_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _1701_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\]
+ _1695_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2343_ net315 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\] net92 VGND
+ VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
XFILLER_69_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4013_ clknet_leaf_33_CLK _0205_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_2274_ net321 net64 net80 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_1
XANTENNA__2419__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__1993__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_1989_ _1090_ _1478_ _1089_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3728_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] _1274_ _1311_ VGND VGND VPWR
+ VPWR _1312_ sky130_fd_sc_hd__or3_1
X_3659_ _1069_ _1078_ _1185_ _1073_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__o31a_1
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2180__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3680__B2 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3680__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2999__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3891__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2171__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3671__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2961_ _0520_ _0522_ _0515_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1912_ _1061_ _1404_ _1060_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a21bo_1
X_2892_ _0474_ _0475_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__nand2_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1843_ _1258_ _1329_ _1331_ _1333_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__o211a_1
XFILLER_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3513_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3444_ _1687_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] _1706_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\]
+ _1028_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__a221o_1
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3375_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0859_ _0860_ VGND VGND VPWR
+ VPWR _0960_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2326_ net235 net52 net78 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XFILLER_85_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2257_ net235 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] net98 VGND
+ VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
XFILLER_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2188_ net264 net50 net86 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_1
XFILLER_53_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout97_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2153__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1898__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_44_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_89_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2144__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3160_ _0727_ _0729_ _0723_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2111_ net206 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] net107 VGND
+ VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
X_3091_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] _0673_ VGND VGND VPWR VPWR
+ _0676_ sky130_fd_sc_hd__nand2_1
Xhold1 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[34\] VGND VGND VPWR VPWR net204
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2042_ net112 _1720_ _1721_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] VGND VGND
+ VPWR VPWR _1535_ sky130_fd_sc_hd__a22o_1
XFILLER_66_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3796__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3993_ clknet_leaf_4_CLK _0185_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_2944_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__nand2_1
X_2875_ _1684_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\] _0458_ _0459_
+ _0457_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__o221a_1
XANTENNA__3528__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2432__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2135__A1 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3427_ _1670_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ _1668_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3358_ net109 _0926_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nand2_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2309_ net306 net65 net76 VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__mux2_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3289_ net121 _0871_ _0873_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] VGND VGND
+ VPWR VPWR _0874_ sky130_fd_sc_hd__o22ai_1
XFILLER_72_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2660_ _1631_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[18\] VGND VGND VPWR
+ VPWR _0280_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2591_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ _1801_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__and3_1
X_3212_ _0505_ _0795_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__nand2_1
XFILLER_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3143_ _0525_ _0542_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__xnor2_1
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3074_ net120 _0657_ _0658_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND
+ VPWR VPWR _0659_ sky130_fd_sc_hd__o22a_1
X_2025_ _1611_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ _1610_ _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_81_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3976_ clknet_leaf_32_CLK _0168_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout147_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2927_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_33_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2858_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] _0383_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[13\]
+ _1667_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__o221a_1
X_2789_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\]
+ _0387_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] VGND VGND VPWR VPWR _0392_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_92_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout102_X net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2101__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2044__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2800__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3810__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3830_ clknet_leaf_11_CLK _0056_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3761_ clknet_leaf_18_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[21\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2712_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] net108 VGND VGND VPWR
+ VPWR _0330_ sky130_fd_sc_hd__or2_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3692_ _1133_ _1164_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__nand3b_1
X_2643_ _0266_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[28\]
+ sky130_fd_sc_hd__inv_2
X_2574_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\] VGND VGND VPWR VPWR
+ _1793_ sky130_fd_sc_hd__inv_2
XFILLER_95_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3126_ _0508_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__xnor2_1
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2510__B2 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0640_ _0641_ _0637_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\]
+ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__o32a_1
XFILLER_82_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2008_ _1492_ _1493_ _1644_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3959_ clknet_leaf_4_CLK _0152_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__2329__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4055__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2265__B1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3894__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2514__B net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2290_ net279 net50 net82 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2264__X _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3813_ clknet_leaf_25_CLK _0039_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_25_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3744_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1266_ _1269_ _1327_ VGND VGND
+ VPWR VPWR _1328_ sky130_fd_sc_hd__o22ai_1
X_3675_ _1091_ _1181_ _1085_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__o21a_1
X_2626_ net113 _1826_ net75 VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_33_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_33_CLK sky130_fd_sc_hd__clkbuf_8
X_2557_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[2\] VGND VGND VPWR VPWR
+ _1781_ sky130_fd_sc_hd__inv_2
XANTENNA__2731__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2488_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[37\] VGND VGND VPWR VPWR
+ _1714_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_34_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3109_ _0682_ _0687_ _0692_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_87_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_24_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout82_X net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_61_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3450__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 addr[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput46 wdata[20] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput24 addr[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 wdata[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xinput57 wdata[30] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_15_CLK sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_70_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3460_ _0997_ _1008_ _1023_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__or4b_1
X_2411_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND VPWR VPWR
+ _1637_ sky130_fd_sc_hd__inv_2
X_3391_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__and2b_1
X_2342_ net219 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\] net92 VGND
+ VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2273_ net334 net63 net81 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
X_4012_ clknet_leaf_33_CLK _0204_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3799__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2229__B1 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3727_ _1131_ _1161_ _1273_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__and3_1
X_1988_ _1426_ _1477_ _1480_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__o21ai_1
X_3658_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] _1230_ _1232_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\]
+ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__a221o_1
XFILLER_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3589_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__or2_1
X_2609_ net71 _1815_ _1816_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__or3_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3913__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2999__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_4_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_4_CLK sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_17_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2960_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__and2_1
X_1911_ _1066_ _1076_ _1374_ _1067_ _1064_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__a311o_1
X_2891_ _0474_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__and2_1
XFILLER_63_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1842_ _1242_ _1333_ _1334_ _1228_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__a31o_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3512_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\]
+ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3443_ _1674_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] _0995_ VGND
+ VGND VPWR VPWR _1028_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3374_ _0883_ _0886_ _0881_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__a21bo_1
X_2325_ net254 net51 net78 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__mux2_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2256_ net254 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] net98 VGND
+ VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2187_ net251 net49 net87 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2104__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3102__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3102__B2 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3405__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2803__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2081__Y myPWM.g_pwm_channel\[1\].CHANNEL.pwm_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input62_X net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2110_ net270 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] net107 VGND
+ VGND VPWR VPWR _0027_ sky130_fd_sc_hd__mux2_1
X_3090_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _0670_ VGND VGND VPWR VPWR
+ _0675_ sky130_fd_sc_hd__or2_1
Xhold2 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[47\] VGND VGND VPWR VPWR net205
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1722_ _1723_ net113 VGND VGND
+ VPWR VPWR _1534_ sky130_fd_sc_hd__a22o_1
XFILLER_66_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3992_ clknet_leaf_5_CLK _0184_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2943_ _0526_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__nor2_2
XANTENNA__3368__X _0953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2874_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[25\]
+ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2713__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3426_ _1663_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[40\]
+ _1662_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a22o_1
XFILLER_97_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3357_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _0938_ _0941_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__o22a_1
X_2308_ net295 net64 net76 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
X_3288_ _0856_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__or2_1
X_2239_ net295 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[8\] net96 VGND VGND
+ VPWR VPWR _0138_ sky130_fd_sc_hd__mux2_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input22_A addr[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2590_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] _1801_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\]
+ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3211_ _0494_ _0770_ _0775_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__or3_1
X_3142_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__inv_2
XFILLER_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3073_ _0610_ _0648_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ _1610_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[35\] _1514_ _1516_
+ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_53_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3975_ clknet_leaf_31_CLK _0167_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2926_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2443__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2857_ _0433_ _0437_ _0441_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__and4_1
X_2788_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0389_ _0391_ VGND VGND VPWR
+ VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[15\] sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_92_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3409_ _1678_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ _1676_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__o221a_1
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2292__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2283__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3760_ clknet_leaf_17_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[20\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] sky130_fd_sc_hd__dfrtp_4
XFILLER_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2711_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] net108 VGND VGND VPWR
+ VPWR _0329_ sky130_fd_sc_hd__nand2_1
X_3691_ _1161_ _1273_ _1131_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__a21o_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2642_ net70 _1839_ _1840_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_78_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2573_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1789_ _1792_ net74 VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[7\] sky130_fd_sc_hd__o211a_1
XANTENNA__2202__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3125_ _0504_ _0708_ _0502_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__a21bo_1
XANTENNA__2438__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3056_ _0474_ _0626_ _0639_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__and3_1
XFILLER_67_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2007_ _1494_ _1498_ _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__or3_1
XFILLER_63_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2274__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3958_ clknet_leaf_6_CLK _0151_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3889_ clknet_leaf_11_CLK _0115_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_4
X_2909_ _1669_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND VPWR
+ VPWR _0494_ sky130_fd_sc_hd__and2_1
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout72_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2811__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2370__X _1599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2256__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3812_ clknet_leaf_24_CLK _0038_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3743_ _1320_ _1324_ _1325_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__o211a_1
X_3674_ _1253_ _1255_ _1256_ _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__a211o_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2625_ net113 _1826_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__nand2_1
X_2556_ _1779_ _1780_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_87_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2487_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[38\] VGND VGND VPWR VPWR
+ _1713_ sky130_fd_sc_hd__inv_2
XFILLER_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3108_ net122 _0686_ _0691_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] _0690_
+ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__a221oi_1
XANTENNA__3772__RESET_B net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_X net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ _0608_ _0611_ _0605_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__a221o_1
XFILLER_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2107__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2631__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3637__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput25 addr[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 addr[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
Xinput36 wdata[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
Xinput58 wdata[31] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
Xinput47 wdata[21] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2410_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR _1636_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3390_ net118 _1702_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__nor2_1
X_2341_ net321 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\] net92 VGND
+ VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
X_2272_ net286 net62 net81 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
X_4011_ clknet_leaf_33_CLK _0203_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3729__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_1987_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1425_ _1479_ net115 VGND VGND
+ VPWR VPWR _1480_ sky130_fd_sc_hd__o22a_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3726_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] _1305_ _1309_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\]
+ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__a22o_1
XANTENNA__3547__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2451__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3657_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1235_ _1240_ VGND VGND VPWR
+ VPWR _1241_ sky130_fd_sc_hd__o21a_1
X_3588_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[49\]
+ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__nand2_1
X_2608_ net115 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1812_ VGND VGND VPWR
+ VPWR _1816_ sky130_fd_sc_hd__and3_1
XFILLER_88_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2539_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] _1610_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\]
+ _1647_ _1764_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__a221o_1
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input52_A wdata[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2300__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2890_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or2_1
X_1910_ _1392_ _1393_ _1396_ _1402_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__or4_1
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1841_ _1332_ _1225_ _1216_ _1226_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_25_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3511_ _1093_ _1094_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_1
X_3442_ _1010_ _1022_ _1023_ _1026_ _1019_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__o32a_1
X_3373_ _0843_ _0955_ _0957_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__o21bai_1
X_2324_ net245 net50 net77 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XANTENNA__2210__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2255_ net245 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] net97 VGND
+ VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2186_ net304 net48 net87 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_1
XFILLER_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2870__A1 _1682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3709_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] _1291_ _1292_ _1104_ VGND VGND
+ VPWR VPWR _1293_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_95_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input55_X net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3875__RESET_B net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2129__B1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[28\] VGND VGND VPWR VPWR net206
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3629__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_94_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2040_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1724_ _1725_ net114 VGND VGND
+ VPWR VPWR _1533_ sky130_fd_sc_hd__a22o_1
XFILLER_62_332 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3991_ clknet_leaf_5_CLK _0183_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2942_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\]
+ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and2b_1
XFILLER_50_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2873_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\]
+ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and2_1
XANTENNA__2205__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3425_ _1002_ _1006_ _1009_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _1007_
+ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__o221a_1
X_3356_ _0784_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nand2b_1
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3287_ _0577_ _0803_ _0810_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__and3_1
X_2307_ net258 net63 net79 VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
X_2238_ net258 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] net99 VGND VGND
+ VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
XANTENNA__3560__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2169_ net316 net61 net84 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2531__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3470__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input15_A addr[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4074__RESET_B net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2062__A2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4003__RESET_B net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] _1711_ _0498_ _0500_
+ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a31o_1
X_3141_ net108 _0721_ _0725_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] VGND VGND
+ VPWR VPWR _0726_ sky130_fd_sc_hd__a22o_1
XANTENNA__2522__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3072_ _0647_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__or2_1
XFILLER_82_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2023_ _1608_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ _1606_ _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__o221a_1
XFILLER_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ clknet_leaf_31_CLK _0166_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2925_ _0501_ _0504_ _0508_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2856_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[8\]
+ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__xnor2_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3555__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2787_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0389_ net73 VGND VGND VPWR
+ VPWR _0391_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_92_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3408_ _1676_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ _1674_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a22o_1
XANTENNA_input7_A addr[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3339_ _0908_ _0921_ _0922_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__and4_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2504__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2710_ _1673_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\]
+ _1687_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3690_ _1161_ _1273_ _1131_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a21oi_1
X_2641_ net112 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] _1835_ VGND VGND VPWR
+ VPWR _1840_ sky130_fd_sc_hd__and3_1
X_2572_ _1791_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__inv_2
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3124_ _0504_ _0708_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__xnor2_1
X_3055_ _0474_ _0626_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_66_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2006_ net113 _1495_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__nor2_1
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2454__A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3957_ clknet_leaf_5_CLK _0150_ net138 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2908_ _1669_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] VGND VGND VPWR
+ VPWR _0493_ sky130_fd_sc_hd__nor2_1
X_3888_ clknet_leaf_10_CLK _0114_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\]
+ sky130_fd_sc_hd__dfrtp_2
X_2839_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\]
+ _0422_ net69 VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a31o_1
XFILLER_78_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2303__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3811_ clknet_leaf_23_CLK _0037_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3742_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[18\] _1263_ _1267_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\]
+ _1268_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__o221a_1
X_3673_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1246_ _1247_ net114 VGND VGND
+ VPWR VPWR _1257_ sky130_fd_sc_hd__o211a_1
XANTENNA__2213__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2624_ _1827_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[23\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__2192__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2555_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1777_ net74 VGND VGND VPWR
+ VPWR _1780_ sky130_fd_sc_hd__o21ai_1
XFILLER_87_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2486_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[39\] VGND VGND VPWR VPWR
+ _1712_ sky130_fd_sc_hd__inv_2
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3552__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3107_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] _0689_ _0691_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\]
+ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__o22a_1
XFILLER_46_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3038_ _0598_ _0604_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__a21oi_1
XFILLER_23_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout155_X net155 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2183__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4082__Q myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 addr[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 addr[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 wdata[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_40_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput48 wdata[22] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
Xinput59 wdata[3] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_75_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2174__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2340_ net334 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\] net93 VGND
+ VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
X_2271_ net291 net61 net80 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4010_ clknet_leaf_32_CLK _0202_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2208__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1986_ _1091_ _1478_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__xor2_1
X_3725_ _1273_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__nand2_1
X_3656_ _1236_ _1239_ _1233_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2165__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2607_ net115 _1812_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR
+ VPWR _1815_ sky130_fd_sc_hd__a21oi_1
X_3587_ _1158_ _1170_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__and2_1
X_2538_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] _1606_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\]
+ _1643_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__a22o_1
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2469_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] VGND VGND VPWR VPWR _1695_
+ sky130_fd_sc_hd__inv_2
XFILLER_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3922__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2642__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_0__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2156__A1 net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wdata[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2552__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3510_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__and2b_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2147__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3441_ _1012_ _1025_ _1016_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a21oi_1
X_3372_ _0831_ _0835_ _0840_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__a31o_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2323_ net237 net49 net77 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2254_ net237 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] net97 VGND
+ VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
X_2185_ net276 net47 net86 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__mux2_1
XFILLER_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1969_ _1118_ _1353_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3708_ _1102_ _1103_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3639_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] _1719_ _1207_ VGND
+ VGND VPWR VPWR _1223_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2138__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2310__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2311__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_X net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[0\] VGND VGND VPWR VPWR net207
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2301__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3990_ clknet_leaf_5_CLK _0182_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2941_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\]
+ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__and2b_1
XFILLER_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2872_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\]
+ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__nor2_1
XANTENNA__2368__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2221__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3424_ _1714_ _1003_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__or2_1
X_3355_ _0525_ _0783_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__nand2_1
X_3286_ _0587_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2540__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_2306_ net231 net62 net79 VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2237_ net231 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] net99 VGND VGND
+ VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_1
XFILLER_72_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2168_ net326 net60 net85 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2099_ net292 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] net106 VGND
+ VGND VPWR VPWR _0016_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2131__S net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout95_A _1597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2531__B2 _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2306__S net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3140_ _0521_ _0549_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3071_ _0598_ _0604_ _0614_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and3_1
X_2022_ _1606_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\]
+ _1604_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__a22o_1
XFILLER_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2216__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3973_ clknet_leaf_31_CLK _0165_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2924_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2855_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\]
+ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__xnor2_1
X_2786_ _0389_ _0390_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[14\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3407_ _1680_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\]
+ _1678_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__a22o_1
X_3338_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0912_ _0913_ _0918_ _0911_
+ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__o2111a_1
XFILLER_100_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3269_ _0853_ _0852_ _0848_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_69_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout98_X net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2640_ net112 _1835_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] VGND VGND VPWR
+ VPWR _1839_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_30_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2571_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[6\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] _1784_ VGND VGND VPWR VPWR _1791_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_78_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3123_ _0501_ _0707_ _0556_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__a21o_1
XFILLER_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3054_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2005_ net113 _1495_ _1497_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] VGND VGND
+ VPWR VPWR _1498_ sky130_fd_sc_hd__a22o_1
XFILLER_48_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout145_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3956_ clknet_leaf_5_CLK _0149_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2907_ _0490_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__and2_1
XFILLER_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2470__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3887_ clknet_leaf_10_CLK _0113_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ sky130_fd_sc_hd__dfrtp_4
X_2838_ _0426_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[30\]
+ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_36_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_36_CLK sky130_fd_sc_hd__clkbuf_8
X_2769_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] _0375_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\]
+ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout100_X net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3880__CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3802__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3476__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2973__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2725__B2 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3810_ clknet_leaf_23_CLK _0036_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3741_ _1321_ _1322_ net116 VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a21o_1
X_3672_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1246_ VGND VGND VPWR VPWR
+ _1256_ sky130_fd_sc_hd__and2_1
XFILLER_9_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_18_CLK sky130_fd_sc_hd__clkbuf_8
X_2623_ net71 _1825_ _1826_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__or3_1
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2554_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__and4_1
XANTENNA__2716__A1 _1656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2485_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\] VGND VGND VPWR VPWR
+ _1711_ sky130_fd_sc_hd__inv_2
XFILLER_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3106_ _0483_ _0568_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__xor2_1
X_3037_ _0610_ _0614_ _0620_ _0617_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__or4b_1
XFILLER_70_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3444__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3939_ clknet_leaf_26_CLK _0132_ net130 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_98_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3380__A1 _0889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3132__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_74_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2078__C _1560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 addr[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput27 addr[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_40_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2314__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput49 wdata[23] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 wdata[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2270_ net213 net60 net80 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_7_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_65_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1985_ _1179_ _1421_ _1372_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__o21a_1
XANTENNA__2224__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3724_ _1146_ _1162_ _1272_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__nand3_1
X_3655_ net113 _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand2_1
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2606_ net115 _1812_ _1814_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[18\]
+ sky130_fd_sc_hd__o21a_1
X_3586_ _1627_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] _1143_ _1163_
+ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__o221a_1
X_2537_ _1605_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\]
+ _1649_ _1762_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__a221o_1
X_2468_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND VPWR VPWR
+ _1694_ sky130_fd_sc_hd__inv_2
X_2399_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] VGND VGND VPWR VPWR _1625_
+ sky130_fd_sc_hd__inv_2
XFILLER_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4069_ clknet_leaf_16_CLK _0261_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.polarity
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2134__S net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout80_X net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3105__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input38_A wdata[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout160 net162 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2309__S net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2092__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3440_ _1014_ _1024_ _1017_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__o21ai_1
X_3371_ _0829_ _0830_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__and2b_1
X_2322_ net255 net48 net77 VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2253_ net255 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] net97 VGND
+ VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2184_ net322 net46 net86 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_1
XFILLER_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2219__S net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2607__B1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_61_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1968_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] _1448_ _1459_ _1460_ _1450_
+ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__a221o_1
X_1899_ _1388_ _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__or2_1
X_3707_ _1604_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_95_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3638_ _1220_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__nor2_1
X_3569_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2196__Y _1591_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2653__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3484__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[2\] VGND VGND VPWR VPWR net208
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_58_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2940_ _0524_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__inv_2
X_2871_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[20\]
+ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3423_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _1714_ VGND VGND VPWR VPWR _1008_
+ sky130_fd_sc_hd__nor2_1
X_3354_ net108 _0933_ _0938_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] VGND VGND
+ VPWR VPWR _0939_ sky130_fd_sc_hd__a22o_1
X_3285_ _1682_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] _0856_ VGND
+ VGND VPWR VPWR _0870_ sky130_fd_sc_hd__o21bai_1
X_2305_ net229 net61 net76 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2236_ net229 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] net99 VGND VGND
+ VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
X_2167_ net320 net59 net85 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
X_2098_ net220 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] net104 VGND
+ VGND VPWR VPWR _0015_ sky130_fd_sc_hd__mux2_1
XFILLER_80_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout88_A _1588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2295__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2383__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2322__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input60_X net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3070_ net118 _0651_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__or2_1
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2021_ _1608_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[34\] VGND VGND VPWR
+ VPWR _1514_ sky130_fd_sc_hd__and2_1
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2286__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3972_ clknet_leaf_29_CLK _0164_ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2923_ _0506_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_33_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2854_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[14\]
+ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__xnor2_1
X_2785_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0387_ net73 VGND VGND VPWR
+ VPWR _0390_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2232__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3406_ _1683_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\]
+ _1681_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__a22o_1
XFILLER_100_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3337_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] _0920_ VGND VGND VPWR VPWR _0922_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__2468__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3268_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0851_ VGND VGND VPWR VPWR
+ _0853_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2219_ net284 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] net102 VGND
+ VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_1
XANTENNA__2277__A1 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3199_ _0525_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_77_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2934__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2931__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2142__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input20_A addr[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_95_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2268__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2317__S net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2570_ _1789_ _1790_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[6\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_78_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3122_ _0513_ _0553_ _0511_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__a21bo_1
XANTENNA__2259__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3053_ _1696_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[62\] VGND VGND VPWR
+ VPWR _0638_ sky130_fd_sc_hd__nand2_1
XFILLER_36_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2004_ _1195_ _1496_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2227__S net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3955_ clknet_leaf_4_CLK _0148_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_2906_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2_1
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3886_ clknet_leaf_28_CLK _0112_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ sky130_fd_sc_hd__dfrtp_2
X_2837_ _0424_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_1
X_2768_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] _0375_ _0377_ VGND VGND VPWR
+ VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[9\] sky130_fd_sc_hd__a21oi_1
X_2699_ _0272_ _0275_ _0295_ _0317_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag_c
+ sky130_fd_sc_hd__and4_1
XANTENNA__3916__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2926__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2137__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2661__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3492__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3740_ net116 _1321_ _1322_ _1323_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_15_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3671_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[21\] _1249_ _1254_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\]
+ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__a22o_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2622_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1823_ VGND VGND VPWR VPWR
+ _1826_ sky130_fd_sc_hd__and2_1
X_2553_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[1\] VGND VGND VPWR VPWR
+ _1778_ sky130_fd_sc_hd__inv_2
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2484_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\] VGND VGND VPWR VPWR
+ _1710_ sky130_fd_sc_hd__inv_2
XFILLER_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3105_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _0684_ _0689_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\]
+ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__a22o_1
XFILLER_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3036_ _0620_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__inv_2
XFILLER_55_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3938_ clknet_leaf_1_CLK _0131_ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3869_ clknet_leaf_15_CLK _0095_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3380__A2 _0953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2656__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 addr[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 addr[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput39 wdata[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2330__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2882__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1984_ _1472_ _1475_ _1476_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__a21oi_1
X_3723_ _1301_ _1304_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__o21a_1
X_3654_ _1191_ _1237_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__or2_1
X_2605_ net115 _1812_ net71 VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2240__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3585_ _1138_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__or2_1
X_2536_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] _1625_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\]
+ _1641_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__a22o_1
X_2467_ net118 VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__inv_2
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2398_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] VGND VGND VPWR VPWR _1624_
+ sky130_fd_sc_hd__inv_2
XFILLER_95_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4068_ clknet_leaf_21_CLK _0260_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable
+ sky130_fd_sc_hd__dfrtp_2
X_3019_ _1688_ _1705_ _0588_ _0603_ _0602_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__o221a_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2150__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_4
Xfanout150 net168 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
XANTENNA_fanout73_X net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2386__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4037__RESET_B net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2325__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3370_ net118 _0838_ _0853_ _0954_ _0846_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__o221a_1
XFILLER_88_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2321_ net303 net47 net77 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
X_2252_ net303 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] net97 VGND
+ VGND VPWR VPWR _0151_ sky130_fd_sc_hd__mux2_1
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2183_ net263 net44 net86 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_38_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2607__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2235__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1967_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\] _1350_ _1449_ _1451_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\]
+ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__o32a_1
X_3706_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__xor2_1
X_1898_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] _1050_ _1387_ VGND VGND VPWR
+ VPWR _1391_ sky130_fd_sc_hd__and3_1
X_3637_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__nor2_1
X_3568_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\]
+ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2519_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] net112 VGND VGND VPWR
+ VPWR _1745_ sky130_fd_sc_hd__nand2_1
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3499_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__nor2_1
XFILLER_76_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2145__S net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input50_A wdata[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold6 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[46\] VGND VGND VPWR VPWR net209
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3005__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2870_ _1682_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[21\] _0453_ _0455_
+ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o211a_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3422_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _1712_ _1713_ net108 VGND VGND
+ VPWR VPWR _1007_ sky130_fd_sc_hd__o22a_1
XANTENNA__2525__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3353_ _0520_ _0785_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__xnor2_1
X_3284_ net122 _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_1
X_2304_ net297 net60 net76 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
X_2235_ net297 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] net96 VGND VGND
+ VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_38_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2166_ net289 net56 net85 VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__mux2_1
XFILLER_26_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout168_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2097_ net323 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] net106 VGND
+ VGND VPWR VPWR _0014_ sky130_fd_sc_hd__mux2_1
XFILLER_80_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2999_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__nor2_1
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3219__A_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input53_X net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4052__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2020_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1728_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ _1624_ _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__a221o_1
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3235__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3971_ clknet_leaf_30_CLK _0163_ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_2922_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] _1709_ VGND VGND VPWR
+ VPWR _0507_ sky130_fd_sc_hd__nand2_1
XFILLER_93_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2853_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[9\]
+ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__xnor2_1
X_2784_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] _0387_ VGND VGND VPWR VPWR
+ _0389_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_92_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3405_ _1687_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ _1683_ _0989_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__o221a_1
XFILLER_58_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3336_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] _0916_ _0920_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\]
+ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__o22a_1
XFILLER_100_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3267_ net120 _0849_ _0851_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND
+ VPWR VPWR _0852_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_69_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ net319 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] net102 VGND
+ VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_1
X_3198_ _0528_ _0782_ _0526_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2149_ net271 net44 net90 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__mux2_1
XANTENNA__3775__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2737__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input13_A addr[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2333__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2728__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3121_ _0701_ _0702_ _0704_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__nand4b_1
X_3052_ _0626_ _0636_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nand2_1
X_2003_ _1189_ _1375_ _1376_ _1188_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_66_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3954_ clknet_leaf_3_CLK _0147_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_2905_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\]
+ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__nand2_1
X_3885_ clknet_leaf_28_CLK _0111_ net150 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_2
X_2836_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0422_ _0361_ VGND VGND VPWR
+ VPWR _0425_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2243__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2719__B1 _1688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2195__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2767_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] _0375_ net73 VGND VGND VPWR
+ VPWR _0377_ sky130_fd_sc_hd__o21ai_1
X_2698_ _1648_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\] _0276_ _0299_
+ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o2111a_1
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input5_A addr[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3319_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0900_ _0903_ net123 VGND VGND
+ VPWR VPWR _0904_ sky130_fd_sc_hd__o22ai_1
XFILLER_100_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2153__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2186__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2328__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2110__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2852__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3670_ _1078_ _1185_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__xnor2_1
X_2621_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] _1823_ VGND VGND VPWR VPWR
+ _1825_ sky130_fd_sc_hd__nor2_1
XANTENNA__2177__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2552_ net70 _1776_ _1777_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[1\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_99_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2483_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\] VGND VGND VPWR VPWR
+ _1709_ sky130_fd_sc_hd__inv_2
XANTENNA__3677__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__3677__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3104_ _0480_ _0688_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__xor2_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3035_ _0618_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__nand2_1
XANTENNA__2238__S net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2101__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout150_A net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3577__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3937_ clknet_leaf_1_CLK _0130_ net132 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3868_ clknet_leaf_14_CLK _0094_ net165 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3799_ clknet_leaf_13_CLK _0026_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_2819_ net120 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] _0408_ VGND VGND VPWR
+ VPWR _0413_ sky130_fd_sc_hd__and3_1
XANTENNA__3593__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2168__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2148__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3487__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput18 addr[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 addr[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2159__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3008__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2847__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2331__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1983_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[16\] _1423_ _1474_ net116 VGND VGND
+ VPWR VPWR _1476_ sky130_fd_sc_hd__o22ai_1
X_3722_ net117 _1303_ _1305_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] VGND VGND
+ VPWR VPWR _1306_ sky130_fd_sc_hd__o22a_1
X_3653_ _1080_ _1185_ _1190_ _1075_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__o211a_1
X_2604_ _1812_ _1813_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[17\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3584_ _1141_ _1166_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__o21a_1
X_2535_ _1754_ _1756_ _1758_ _1760_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__or4_1
X_2466_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND VPWR VPWR
+ _1692_ sky130_fd_sc_hd__inv_2
XANTENNA__2322__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2397_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] VGND VGND VPWR VPWR _1623_
+ sky130_fd_sc_hd__inv_2
XFILLER_95_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4067_ clknet_leaf_10_CLK _0259_ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3018_ _0589_ _0594_ _0596_ _0599_ _0593_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__o221a_1
XFILLER_36_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout140 net145 VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
Xfanout162 net168 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_2
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
XFILLER_19_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2313__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2341__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2320_ net227 net46 net77 VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2251_ net227 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] net97 VGND
+ VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_1
XANTENNA__2577__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2304__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2182_ net228 net43 net86 VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1966_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[3\] _1451_ _1452_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\]
+ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__a221o_1
X_3705_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__and2_1
XANTENNA__2251__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1897_ _1649_ _1388_ _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__or3b_1
X_3636_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__inv_2
X_3567_ _1147_ _1150_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__nand2_1
XFILLER_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2543__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2518_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\]
+ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__nand2_1
X_3498_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nand2_1
XFILLER_75_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2449_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\] VGND VGND VPWR VPWR
+ _1675_ sky130_fd_sc_hd__inv_2
XFILLER_84_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4119_ myPWM.g_pwm_channel\[1\].CHANNEL.pwm_out VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2161__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2534__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__2534__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input43_A wdata[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold7 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[3\] VGND VGND VPWR VPWR net210
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3005__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3021__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2336__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3421_ _1004_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__nand2_1
X_3352_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0935_ VGND VGND VPWR VPWR _0937_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__2525__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2303_ net210 net59 net76 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
X_3283_ _0595_ _0867_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2234_ net210 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] net96 VGND VGND
+ VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
XFILLER_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2165_ net290 net45 net85 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__mux2_1
XFILLER_93_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2096_ net302 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] net104 VGND
+ VGND VPWR VPWR _0013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2246__S net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2998_ _0579_ _0581_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or2_1
X_1949_ _1440_ _1441_ _1357_ _1360_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__a211o_1
X_3619_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] _1720_ _1202_ _1199_
+ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a31o_1
XFILLER_95_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2156__S net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2507__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2398__Y _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input46_X net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3180__B2 _1682_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3970_ clknet_leaf_10_CLK _0162_ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4021__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2921_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] _1709_ VGND VGND VPWR
+ VPWR _0506_ sky130_fd_sc_hd__nor2_1
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2852_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] _0385_ VGND VGND VPWR
+ VPWR _0438_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2783_ _0388_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[13\]
+ sky130_fd_sc_hd__inv_2
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3404_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\]
+ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3335_ _0914_ _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__or2_1
XFILLER_100_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3266_ _0610_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2217_ net328 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] net102 VGND
+ VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3197_ _0531_ _0780_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__a21o_1
XFILLER_26_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2148_ net283 net43 net90 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__mux2_1
XFILLER_54_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2079_ _1337_ _1401_ _1508_ _1509_ _1571_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__a41o_1
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2985__A1 _0564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2737__A1 _1688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout93_A _1597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2675__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2728__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3120_ net123 _0703_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nand2_1
XFILLER_67_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3051_ _0476_ _0623_ _0625_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__or3_1
X_2002_ _1190_ _1377_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3953_ clknet_leaf_3_CLK _0146_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_3884_ clknet_leaf_28_CLK _0110_ net149 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_2
X_2904_ _0487_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__nand2_2
X_2835_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0422_ VGND VGND VPWR VPWR
+ _0424_ sky130_fd_sc_hd__and2_1
X_2766_ _0375_ _0376_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[8\]
+ sky130_fd_sc_hd__nor2_1
X_2697_ _1640_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[25\] _0273_ _0274_
+ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__o2111a_1
X_3318_ _0489_ _0891_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3249_ _0639_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3925__RESET_B net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout96_X net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2344__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2620_ _1824_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[22\]
+ sky130_fd_sc_hd__inv_2
XFILLER_63_5 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2551_ _1606_ _1775_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__nor2_1
XFILLER_99_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2482_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\] VGND VGND VPWR VPWR
+ _1708_ sky130_fd_sc_hd__inv_2
XFILLER_99_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3103_ _0482_ _0568_ _0481_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__a21bo_1
X_4083_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[9\] net150
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\] sky130_fd_sc_hd__dfrtp_4
X_3034_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__or2_1
XANTENNA__3204__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2254__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3936_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag_c net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag sky130_fd_sc_hd__dfrtp_1
X_3867_ clknet_leaf_14_CLK _0093_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_3798_ clknet_leaf_13_CLK _0025_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_2818_ net120 _0408_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[25\] VGND VGND VPWR
+ VPWR _0412_ sky130_fd_sc_hd__a21oi_1
X_2749_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0364_ net72 VGND VGND VPWR
+ VPWR _0366_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2573__C1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2164__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 addr[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3008__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3108__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2339__S net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2095__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1982_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] _1430_ _1474_ net116 VGND VGND
+ VPWR VPWR _1475_ sky130_fd_sc_hd__a22oi_1
X_3721_ _1150_ _1271_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__xnor2_1
X_3652_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[25\] _1235_ VGND VGND VPWR VPWR
+ _1236_ sky130_fd_sc_hd__nand2_1
X_3583_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[47\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\]
+ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__nand2b_1
X_2603_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1810_ net75 VGND VGND VPWR
+ VPWR _1813_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_97_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2534_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] _1613_ _1634_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\]
+ _1759_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__a221o_1
XFILLER_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2465_ net119 VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__inv_2
XFILLER_87_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2396_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR _1622_
+ sky130_fd_sc_hd__inv_2
XANTENNA__2249__S net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4066_ clknet_leaf_11_CLK _0258_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_3017_ _0583_ _0601_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__nand2_1
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3919_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[15\] net133
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1852__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2948__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout130 net131 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2159__S net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout163 net167 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_4
Xfanout141 net145 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__buf_2
Xfanout152 net155 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2683__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__B myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2250_ net244 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] net97 VGND
+ VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_1
XFILLER_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2181_ net300 net42 net86 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_92_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1965_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] _1452_ _1456_ _1457_ VGND VGND
+ VPWR VPWR _1458_ sky130_fd_sc_hd__o22a_1
X_3704_ _1099_ _1106_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__xnor2_1
X_1896_ _1052_ _1386_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3635_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__nand2_1
X_3566_ _1148_ _1149_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout106_A _1574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3497_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__and2_1
XANTENNA__2543__A2 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2517_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\]
+ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__or2_1
X_2448_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[16\] VGND VGND VPWR VPWR _1674_
+ sky130_fd_sc_hd__inv_2
XFILLER_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2379_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] VGND VGND VPWR VPWR
+ _1605_ sky130_fd_sc_hd__inv_2
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4118_ myPWM.g_pwm_channel\[0\].CHANNEL.pwm_out VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4049_ clknet_leaf_35_CLK _0241_ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input36_A wdata[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[13\] VGND VGND VPWR VPWR net211
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2352__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3420_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[5\] _1714_ _1003_ VGND VGND VPWR
+ VPWR _1005_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3351_ net108 _0933_ _0935_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] VGND VGND
+ VPWR VPWR _0936_ sky130_fd_sc_hd__o22a_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2302_ net208 net56 net79 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3282_ _0805_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__nor2_1
XANTENNA__2289__A1 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2233_ net208 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[2\] net96 VGND VGND
+ VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_1
XFILLER_38_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2164_ net288 net34 net85 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__mux2_1
XFILLER_93_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2095_ net259 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] net104 VGND
+ VGND VPWR VPWR _0012_ sky130_fd_sc_hd__mux2_1
XFILLER_34_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2262__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2997_ _0579_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__nor2_1
X_1948_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ _1154_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__a21oi_1
X_1879_ _1172_ _1177_ _1178_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a21bo_1
X_3618_ _1200_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nand2_2
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3549_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__xor2_2
XFILLER_56_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2172__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2507__A2 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3180__A2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_X net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2347__S net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkload1_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2871__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2920_ _0504_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__inv_2
X_2851_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[5\]
+ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2782_ net69 _0386_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or3_1
XFILLER_7_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3403_ _0982_ _0986_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_0_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3334_ _0793_ _0513_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__and2b_1
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3265_ _0613_ _0812_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] _1704_
+ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_37_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2216_ net271 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] net102 VGND
+ VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_1
XFILLER_66_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3196_ _1656_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[35\] VGND VGND VPWR
+ VPWR _0781_ sky130_fd_sc_hd__nor2_1
XFILLER_38_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2257__S net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2147_ net240 net42 net90 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__mux2_1
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2078_ _1569_ _1570_ _1560_ _1567_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__and4b_1
XFILLER_81_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout86_A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2167__S net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_73_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3050_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0632_ VGND VGND VPWR VPWR
+ _0635_ sky130_fd_sc_hd__and2_1
X_2001_ _1644_ _1492_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_82_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3952_ clknet_leaf_35_CLK _0145_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3883_ clknet_leaf_26_CLK net242 net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2903_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or2_1
X_2834_ _0422_ _0423_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[29\]
+ sky130_fd_sc_hd__nor2_1
X_2765_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] _0373_ net72 VGND VGND VPWR
+ VPWR _0376_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_91_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2696_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] _1827_ _1833_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\]
+ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__o221a_1
XFILLER_86_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3317_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0895_ VGND VGND VPWR VPWR
+ _0902_ sky130_fd_sc_hd__or2_1
XFILLER_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3248_ _0477_ _0821_ _0822_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__a21o_1
XFILLER_100_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3179_ _0585_ _0586_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\] VGND
+ VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpwm_wrapper_200 VGND VGND VPWR VPWR pwm_wrapper_200/HI rdata[29] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout89_X net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2550_ _1606_ _1775_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__and2_1
XFILLER_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2481_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\] VGND VGND VPWR VPWR
+ _1707_ sky130_fd_sc_hd__inv_2
XFILLER_99_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3102_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] _0684_ _0686_ net122 VGND VGND
+ VPWR VPWR _0687_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_17_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4082_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[8\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_83_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3033_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__nand2_1
X_3935_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[31\]
+ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] sky130_fd_sc_hd__dfrtp_4
X_3866_ clknet_leaf_13_CLK _0092_ net164 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout136_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3797_ clknet_leaf_12_CLK net265 net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2817_ _0411_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[24\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__2270__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2748_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__and4_1
X_2679_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] _1830_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\]
+ _1642_ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o221a_1
XFILLER_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2180__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input66_A wen VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2867__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2867__B2 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2355__S net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3720_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] _1300_ _1303_ net117 VGND VGND
+ VPWR VPWR _1304_ sky130_fd_sc_hd__a22o_1
X_1981_ _1138_ _1473_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__xnor2_1
X_3651_ _1195_ _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2090__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3582_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] _1728_ _1165_ VGND
+ VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a21oi_1
X_2602_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] _1810_ VGND VGND VPWR VPWR
+ _1812_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_97_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2555__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2533_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] _1623_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\]
+ _1635_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__a22o_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2464_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] VGND VGND VPWR VPWR
+ _1690_ sky130_fd_sc_hd__inv_2
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2395_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] VGND VGND VPWR VPWR
+ _1621_ sky130_fd_sc_hd__inv_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ clknet_leaf_8_CLK _0257_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\]
+ sky130_fd_sc_hd__dfrtp_2
X_3016_ _0574_ _0600_ _0572_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3918_ clknet_leaf_36_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[14\]
+ net128 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[14\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__3586__A2 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3849_ clknet_leaf_25_CLK _0075_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2794__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout120 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] VGND VGND VPWR VPWR net120
+ sky130_fd_sc_hd__buf_2
Xfanout131 net134 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
Xfanout142 net145 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_4
Xfanout164 net166 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2175__S net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2785__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2537__B1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2180_ net292 net41 net86 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__mux2_1
XFILLER_92_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_92_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2085__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1964_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] _1455_ VGND VGND VPWR VPWR _1457_
+ sky130_fd_sc_hd__and2_1
X_3703_ _1095_ _1108_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__xnor2_1
X_1895_ _1050_ _1387_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR
+ VPWR _1388_ sky130_fd_sc_hd__a21oi_1
X_3634_ _1207_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nand2b_1
X_3565_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__or2_1
X_3496_ _1065_ _1069_ _1078_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__or3_1
X_2516_ _1738_ _1739_ _1740_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__a22o_1
XANTENNA__3941__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2447_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] VGND VGND VPWR VPWR
+ _1673_ sky130_fd_sc_hd__inv_2
X_2378_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\] VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__inv_2
X_4048_ clknet_leaf_35_CLK _0240_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2767__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[53\] VGND VGND VPWR VPWR net212
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A addr[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3350_ _0514_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__xnor2_1
X_2301_ net309 net45 net78 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
X_3281_ _0806_ _0865_ _0591_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__o21a_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2232_ net309 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[1\] net98 VGND VGND
+ VPWR VPWR _0131_ sky130_fd_sc_hd__mux2_1
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2163_ _1576_ _1583_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__and3_2
XANTENNA__3238__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2094_ net232 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] net104 VGND
+ VGND VPWR VPWR _0011_ sky130_fd_sc_hd__mux2_1
XFILLER_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2996_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] _1705_ VGND VGND VPWR
+ VPWR _0581_ sky130_fd_sc_hd__nor2_1
XFILLER_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2749__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1947_ _1354_ _1355_ _1156_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__a21o_1
X_1878_ _1365_ _1368_ _1370_ _1179_ _1174_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__a2111o_1
X_3617_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__or2_1
X_3548_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__inv_2
X_3479_ _1061_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__and2_1
XFILLER_88_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3919__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2140__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2850_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable _0436_ net111 VGND VGND
+ VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[0\] sky130_fd_sc_hd__mux2_1
X_2781_ net123 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0382_ VGND VGND VPWR
+ VPWR _0387_ sky130_fd_sc_hd__and3_1
XFILLER_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4030__RESET_B net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3402_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[24\] _1705_ _0976_ _0977_ VGND VGND
+ VPWR VPWR _0987_ sky130_fd_sc_hd__a211o_1
XFILLER_98_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3333_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__inv_2
X_3264_ _0613_ _0812_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2215_ net283 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[50\] net102 VGND
+ VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_1
XFILLER_66_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3195_ _0533_ _0778_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__o21ai_1
XANTENNA__2131__A1 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2146_ net274 net41 net90 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__mux2_1
XFILLER_93_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout166_A net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2077_ _1548_ _1546_ _1547_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__or3b_1
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2273__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_101_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2979_ _0548_ _0552_ _0554_ _0496_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_32_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2183__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2189__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_X net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2113__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2000_ _1057_ _1491_ _1202_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__a21o_1
XANTENNA__2585__C myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3951_ clknet_leaf_3_CLK _0144_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__2093__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2902_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nand2_1
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3882_ clknet_leaf_26_CLK _0108_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_2833_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\] _0420_ _0361_ VGND VGND VPWR
+ VPWR _0423_ sky130_fd_sc_hd__o21ai_1
X_2764_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] _0370_ VGND VGND VPWR VPWR _0375_
+ sky130_fd_sc_hd__and4_1
XANTENNA__1927__A1 _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2695_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] _1827_ _0313_ VGND
+ VGND VPWR VPWR _0314_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3316_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] _0900_ VGND VGND VPWR VPWR
+ _0901_ sky130_fd_sc_hd__nand2_1
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2268__S net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2104__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3247_ _0477_ _0821_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3178_ _0760_ _0762_ _0646_ _0654_ _0662_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_1_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2792__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2129_ _1602_ net337 net91 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__a21o_1
XFILLER_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout169_X net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xpwm_wrapper_201 VGND VGND VPWR VPWR pwm_wrapper_201/HI rdata[30] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2178__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_591 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input11_A addr[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2480_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND VPWR VPWR
+ _1706_ sky130_fd_sc_hd__inv_2
XFILLER_99_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3101_ _0595_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__xnor2_1
XFILLER_68_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2088__S net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4081_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] sky130_fd_sc_hd__dfrtp_4
X_3032_ _0615_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__or2_2
XFILLER_91_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3501__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3220__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3934_ clknet_leaf_10_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[30\]
+ net141 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2117__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3865_ clknet_leaf_13_CLK _0091_ net162 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_2816_ net120 _0408_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__a21o_1
XFILLER_31_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3796_ clknet_leaf_11_CLK _0023_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout129_A net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2747_ net69 _0363_ _0364_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[1\]
+ sky130_fd_sc_hd__nor3_1
X_2678_ _1639_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[24\] _0277_ _0278_
+ _0296_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__o2111a_1
XANTENNA__2325__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input3_A addr[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input59_A wdata[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2316__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input14_X net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1980_ _1142_ _1429_ _1139_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2371__S _1599_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3650_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] _1722_ _1191_ VGND
+ VGND VPWR VPWR _1234_ sky130_fd_sc_hd__a21o_1
X_3581_ _1133_ _1164_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__nor2_1
X_2601_ _1810_ _1811_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2532_ _1607_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[2\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\]
+ _1622_ _1757_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__a221o_1
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2463_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] VGND VGND VPWR VPWR
+ _1689_ sky130_fd_sc_hd__inv_2
XANTENNA__2307__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2394_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] VGND VGND VPWR VPWR _1620_
+ sky130_fd_sc_hd__inv_2
XANTENNA__2400__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_4064_ clknet_leaf_8_CLK _0256_ net144 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[61\]
+ sky130_fd_sc_hd__dfrtp_1
X_3015_ _0576_ _0586_ _0584_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a21o_1
XFILLER_64_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3917_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[13\] net128
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[13\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__2281__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3848_ clknet_leaf_25_CLK _0074_ net148 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3779_ clknet_leaf_24_CLK _0006_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_20_CLK sky130_fd_sc_hd__clkbuf_8
Xfanout110 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[1\] VGND VGND VPWR VPWR net110
+ sky130_fd_sc_hd__buf_2
Xfanout121 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[21\] VGND VGND VPWR VPWR net121
+ sky130_fd_sc_hd__buf_2
Xfanout165 net166 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_4
Xfanout143 net144 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_4
Xfanout154 net155 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2191__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2979__X _0564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_11_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_77_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2890__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ _1453_ _1454_ _1455_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[1\] VGND VGND
+ VPWR VPWR _1456_ sky130_fd_sc_hd__o22a_1
X_1894_ _1053_ _1219_ _1385_ _1221_ _1052_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__a311o_1
X_3702_ _1109_ _1113_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__xnor2_1
X_3633_ _1056_ _1203_ _1205_ _1206_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__or4_1
XANTENNA__2528__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3564_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[11\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__nand2_1
X_3495_ _1076_ _1077_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__nand2_1
X_2515_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] net114 VGND VGND VPWR
+ VPWR _1741_ sky130_fd_sc_hd__nand2_1
X_2446_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] VGND VGND VPWR VPWR _1672_
+ sky130_fd_sc_hd__inv_2
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2377_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag VGND VGND VPWR VPWR _1603_
+ sky130_fd_sc_hd__inv_2
XFILLER_83_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2276__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4047_ clknet_leaf_34_CLK _0239_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2975__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2186__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_0_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_11_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3280_ _0807_ _0863_ _0480_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__o21a_1
X_2300_ net207 net34 net79 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
X_2231_ net207 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\] net99 VGND VGND
+ VPWR VPWR _0130_ sky130_fd_sc_hd__mux2_1
XFILLER_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2162_ net23 _1586_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__nor2_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2093_ net253 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] net104 VGND
+ VGND VPWR VPWR _0010_ sky130_fd_sc_hd__mux2_1
XANTENNA__2096__S net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2995_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__inv_2
XFILLER_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1946_ _1437_ _1438_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] VGND VGND VPWR
+ VPWR _1439_ sky130_fd_sc_hd__o21a_1
X_1877_ _1084_ _1091_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__nand2_1
X_3616_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nand2_1
X_3547_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\]
+ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__xor2_2
XANTENNA__3952__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3478_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__or2_1
X_2429_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__inv_2
XFILLER_84_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input41_A wdata[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2780_ net123 _0382_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] VGND VGND VPWR
+ VPWR _0386_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_2_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_2_1__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2600__B1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3401_ _0974_ _0985_ _0975_ _0978_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__or4b_1
XFILLER_98_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3332_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[10\] _0912_ _0916_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[9\]
+ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__a22o_1
XFILLER_98_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3263_ _0846_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__and2_1
XANTENNA__3504__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2214_ net240 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[49\] net102 VGND
+ VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_1
X_3194_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[34\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\]
+ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__nand2b_1
XFILLER_66_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2145_ net205 net40 net88 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__mux2_1
XFILLER_93_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2076_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] _1568_ _1543_ myPWM.g_pwm_channel\[1\].CHANNEL.alignment
+ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__a211o_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout159_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3947__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2978_ _0490_ _0561_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__a21oi_1
X_1929_ _1174_ _1369_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout114_X net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2830__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3386__A1 _0695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input44_X net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold90 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[17\] VGND VGND VPWR VPWR net293
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3950_ clknet_leaf_35_CLK _0143_ net127 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_2901_ _0484_ _0485_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__or2_2
X_3881_ clknet_leaf_25_CLK _0107_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_84_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2832_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[29\]
+ _0418_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__and3_1
X_2763_ net69 _0373_ _0374_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[7\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_8_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2694_ _0280_ _0292_ _0304_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or4b_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3315_ _0495_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3246_ _1697_ _0828_ _0829_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__o211a_1
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3177_ _0675_ _0680_ _0761_ _0681_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__a31o_1
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _1576_ _1583_ _1587_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_1_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2059_ net114 _1725_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] _1636_
+ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2284__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2040__B2 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xpwm_wrapper_202 VGND VGND VPWR VPWR pwm_wrapper_202/HI rdata[31] sky130_fd_sc_hd__conb_1
XFILLER_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout91_A _1588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3903__RESET_B net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2983__A _0564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2194__S net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2369__S _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3054__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3100_ _0590_ _0663_ _0589_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__a21bo_1
X_4080_ clknet_leaf_20_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\] net154
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] sky130_fd_sc_hd__dfrtp_1
X_3031_ _1694_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\] VGND VGND VPWR
+ VPWR _0616_ sky130_fd_sc_hd__and2_1
XANTENNA__2893__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3933_ clknet_leaf_1_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\] net141
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] sky130_fd_sc_hd__dfrtp_4
X_3864_ clknet_leaf_13_CLK _0090_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2270__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2815_ net120 _0408_ net72 VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__o21ai_1
X_3795_ clknet_leaf_12_CLK _0022_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2746_ net111 net110 myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable VGND VGND
+ VPWR VPWR _0364_ sky130_fd_sc_hd__and3_1
X_2677_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] _1821_ VGND VGND VPWR
+ VPWR _0296_ sky130_fd_sc_hd__xor2_1
XANTENNA__3960__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2279__S net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3229_ _0609_ _0613_ _0617_ _0621_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__or4_1
XANTENNA__2089__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2261__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2189__S net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout94_X net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2252__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3580_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\]
+ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__nand2b_1
X_2600_ _1628_ _1809_ net70 VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2531_ _1612_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\]
+ _1638_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__a22o_1
X_2462_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] VGND VGND VPWR VPWR
+ _1688_ sky130_fd_sc_hd__inv_2
XFILLER_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2099__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3780__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2393_ net117 VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_79_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4063_ clknet_leaf_8_CLK _0255_ net143 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_68_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3014_ _0478_ _0481_ _0479_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a21bo_1
XANTENNA__3512__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout141_A net145 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2243__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3916_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[12\] net128
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_88_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3955__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3847_ clknet_leaf_25_CLK _0073_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3778_ clknet_leaf_24_CLK _0005_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__2798__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2729_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] _1683_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[30\]
+ _1697_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a221o_1
Xfanout122 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR net122
+ sky130_fd_sc_hd__buf_2
Xfanout100 _1591_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__buf_4
Xfanout111 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[0\] VGND VGND VPWR VPWR net111
+ sky130_fd_sc_hd__buf_2
Xfanout144 net145 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
Xfanout133 net134 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_4
Xfanout155 net168 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_2
Xfanout166 net167 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_86_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2234__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[3\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1962_ _1102_ _1346_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1893_ _1053_ _1219_ _1385_ _1221_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__a31o_1
XANTENNA__3775__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3701_ _1092_ _1284_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__xnor2_1
X_3632_ _1212_ _1213_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__and3_1
X_3563_ _1144_ _1145_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nand2_1
X_3494_ _1076_ _1077_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__and2_1
XANTENNA__2411__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2514_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] net114 VGND VGND VPWR
+ VPWR _1740_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2445_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[15\] VGND VGND VPWR VPWR
+ _1671_ sky130_fd_sc_hd__inv_2
X_2376_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.rollover_flag VGND VGND VPWR VPWR _1602_
+ sky130_fd_sc_hd__inv_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4046_ clknet_leaf_34_CLK _0238_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[43\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3666__A1_N net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2292__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2216__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[51\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2991__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2230_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.rollover_flag myPWM.g_pwm_channel\[1\].CHANNEL.data_mod\[0\]
+ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__nand2_1
X_2161_ net268 net58 net91 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__mux2_1
XFILLER_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2092_ net317 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] net104 VGND
+ VGND VPWR VPWR _0009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2994_ _1688_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[56\] VGND VGND VPWR
+ VPWR _0579_ sky130_fd_sc_hd__nor2_1
XANTENNA__2406__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1945_ _1148_ _1434_ _1147_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__a21oi_1
X_1876_ _1365_ _1368_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__and2_1
XANTENNA__3237__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2412__Y _1638_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3615_ _1645_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] VGND VGND VPWR
+ VPWR _1199_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout104_A _1574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3546_ _1122_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__nand2_1
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3477_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\]
+ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__nand2_1
XFILLER_69_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2428_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND VPWR VPWR
+ _1654_ sky130_fd_sc_hd__inv_2
XANTENNA__2287__S net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2359_ net249 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\] net95 VGND
+ VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
XFILLER_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4029_ clknet_leaf_6_CLK _0221_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_15_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2986__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2197__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input34_A wdata[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3610__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3400_ net119 _1703_ _0983_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__a211o_1
XFILLER_98_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3331_ _0501_ _0915_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3262_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] _0845_ VGND VGND VPWR VPWR
+ _0847_ sky130_fd_sc_hd__nand2_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3193_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\]
+ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__and2b_1
XFILLER_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2213_ net274 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\] net102 VGND
+ VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
X_2144_ net209 net39 net88 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__mux2_1
XFILLER_93_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2075_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[62\] _1545_ VGND VGND VPWR
+ VPWR _1568_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_2_2__f_CLK_X clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2977_ _0486_ _0491_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nand2_1
X_1928_ _1174_ _1369_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__or2_1
XANTENNA__3963__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[26\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1859_ _1113_ _1345_ _1349_ _1351_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__a31o_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3529_ _1111_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__nor2_2
XFILLER_69_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2046__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_33_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2594__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_X net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold91 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[52\] VGND VGND VPWR VPWR net294
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[50\] VGND VGND VPWR VPWR net283
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2900_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[16\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[48\]
+ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__and2b_1
X_3880_ clknet_2_2__leaf_CLK _0106_ net146 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2831_ _0420_ _0421_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[28\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_77_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2762_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] _0370_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\]
+ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3783__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2693_ _0309_ _0310_ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__and3_1
XFILLER_98_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3314_ _0489_ _0891_ _0774_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__a21o_1
X_3245_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\] _0826_ VGND VGND VPWR VPWR
+ _0830_ sky130_fd_sc_hd__nand2_1
XFILLER_58_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3176_ _0674_ _0671_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand2b_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ _1600_ _1586_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2058_ _1636_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[52\]
+ _1635_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__o22a_1
XFILLER_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xpwm_wrapper_203 VGND VGND VPWR VPWR pwm_wrapper_203/HI request_stall sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_9_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout84_A _1590_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4049__RESET_B net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3030_ _1694_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\] VGND VGND VPWR
+ VPWR _0615_ sky130_fd_sc_hd__nor2_1
XFILLER_63_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3932_ clknet_leaf_9_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[28\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[28\] sky130_fd_sc_hd__dfrtp_4
X_3863_ clknet_leaf_12_CLK _0089_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2414__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2814_ _0408_ _0409_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[23\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3794_ clknet_leaf_12_CLK _0021_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__2558__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2745_ net111 myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable net110 VGND VGND
+ VPWR VPWR _0363_ sky130_fd_sc_hd__a21oi_1
X_2676_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[29\]
+ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3228_ _0617_ _0621_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__nor2_1
XFILLER_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2295__S net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3159_ net111 _0740_ _0743_ _0739_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__a211oi_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3210__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout87_X net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2994__A _1688_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_416 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ _1626_ net116 _1633_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] _1755_
+ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__a221o_1
XFILLER_5_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2461_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] VGND VGND VPWR VPWR _1687_
+ sky130_fd_sc_hd__inv_2
X_2392_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__inv_2
XANTENNA__3865__RESET_B net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4062_ clknet_leaf_7_CLK _0254_ net145 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_56_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3013_ _0564_ _0567_ _0569_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__a211o_1
XFILLER_76_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2409__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_91_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3915_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[11\] net133
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3846_ clknet_leaf_25_CLK _0072_ net147 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout134_A net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3777_ clknet_leaf_23_CLK _0004_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_2728_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] _1670_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[28\]
+ _1695_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a22o_1
X_2659_ _1629_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[17\] VGND VGND VPWR
+ VPWR _0279_ sky130_fd_sc_hd__xnor2_1
Xfanout101 _1591_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
Xfanout112 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] VGND VGND VPWR VPWR net112
+ sky130_fd_sc_hd__buf_2
XFILLER_101_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout145 net169 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
XFILLER_86_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout156 net158 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout123 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\] VGND VGND VPWR VPWR net123
+ sky130_fd_sc_hd__buf_2
Xfanout134 net169 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_2
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
XFILLER_86_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input64_A wdata[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2170__A1 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3700_ _1109_ _1113_ _1125_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__o21ba_1
X_1961_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] _1290_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[0\]
+ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_99_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1892_ _1380_ _1384_ _1055_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__o21ai_2
X_3631_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[30\] _1214_ VGND VGND VPWR VPWR
+ _1215_ sky130_fd_sc_hd__xnor2_1
X_3562_ _1144_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__and2_1
XANTENNA__3791__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2513_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__nand2_1
X_3493_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__or2_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3489__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2444_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[14\] VGND VGND VPWR VPWR _1670_
+ sky130_fd_sc_hd__inv_2
X_2375_ net27 VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__inv_2
XFILLER_84_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2161__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4045_ clknet_leaf_33_CLK _0237_ net125 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[42\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3661__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3966__Q myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3829_ clknet_leaf_11_CLK _0055_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2602__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2152__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1888__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3168__B1 _0695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2512__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2143__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2160_ net222 net57 net91 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__mux2_1
XFILLER_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2091_ net280 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] net104 VGND
+ VGND VPWR VPWR _0008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2993_ _0575_ _0576_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__nand2_1
XFILLER_34_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1944_ _1147_ _1148_ _1434_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__and3_1
X_3614_ _1197_ _1059_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__and2b_1
X_1875_ _1137_ _1139_ _1343_ _1367_ _1136_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__o221a_1
XANTENNA__2422__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3545_ _1121_ _1128_ _1123_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__o21a_1
X_3476_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\]
+ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__xor2_2
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2427_ net110 VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__inv_2
XANTENNA__2134__A1 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2358_ net234 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\] net95 VGND
+ VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
XFILLER_69_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2289_ net329 net49 net82 VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4028_ clknet_leaf_6_CLK _0220_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2373__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2986__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[55\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A addr[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3625__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3330_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[9\] _1711_ _0914_ VGND
+ VGND VPWR VPWR _0915_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3261_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[26\] _0845_ VGND VGND VPWR VPWR
+ _0846_ sky130_fd_sc_hd__or2_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3192_ _0507_ _0776_ _0506_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a21oi_1
X_2212_ net205 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[47\] net100 VGND
+ VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
X_2143_ net218 net38 net88 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__mux2_1
XFILLER_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2074_ _1542_ _1549_ _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__or3_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2976_ _0487_ _0495_ _0560_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__o21a_1
X_1927_ _1638_ _1405_ _1406_ _1419_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__a31o_1
X_1858_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ _1111_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__a21o_1
XFILLER_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3528_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__nor2_1
XFILLER_39_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3459_ _0998_ _1007_ _1042_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__and4_1
XFILLER_69_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold81 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[54\] VGND VGND VPWR VPWR net284
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[8\] VGND VGND VPWR VPWR net295
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[37\] VGND VGND VPWR VPWR net273
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2830_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[28\] _0418_ net72 VGND VGND VPWR
+ VPWR _0421_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_100_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[6\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\]
+ _0370_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__and3_1
X_2692_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[16\] _1810_ _1811_ _0291_
+ _0294_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_14_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3313_ _0893_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nand2_1
XFILLER_98_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3244_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[30\] _0824_ _0827_ _0826_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[31\]
+ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__o32a_1
XANTENNA_clkbuf_leaf_29_CLK_A clknet_2_0__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3175_ net122 _0686_ _0687_ _0759_ _0683_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__a221o_1
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ net2 net5 _1584_ _1585_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2057_ net113 _1723_ _1724_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[23\] VGND VGND
+ VPWR VPWR _1550_ sky130_fd_sc_hd__o22a_1
XFILLER_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2959_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__inv_2
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2328__A1 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout77_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3912__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2319__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3616__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2520__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3931_ clknet_leaf_1_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[27\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[27\] sky130_fd_sc_hd__dfrtp_1
X_3862_ clknet_leaf_11_CLK _0088_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3794__Q myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2813_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0407_ net72 VGND VGND VPWR
+ VPWR _0409_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3793_ clknet_leaf_12_CLK _0020_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_2744_ net72 VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__inv_2
X_2675_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[12\]
+ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_32_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_32_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_98_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3227_ _0769_ _0803_ _0811_ _0768_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__o211a_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3158_ net110 _0737_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__a21bo_1
X_2109_ net333 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[26\] net107 VGND
+ VGND VPWR VPWR _0026_ sky130_fd_sc_hd__mux2_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout167_X net167 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3089_ net121 _0667_ _0673_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[20\] VGND VGND
+ VPWR VPWR _0674_ sky130_fd_sc_hd__o22a_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_23_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2515__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_14_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_5_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2460_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND VPWR VPWR
+ _1686_ sky130_fd_sc_hd__inv_2
XFILLER_96_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2391_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[7\] VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__inv_2
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4061_ clknet_leaf_6_CLK _0253_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_3012_ _0588_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__or2_1
XANTENNA__3673__C1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2425__A myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3914_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[10\] net128
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3845_ clknet_leaf_24_CLK _0071_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3776_ clknet_leaf_23_CLK _0003_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout127_A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2727_ _0340_ _0341_ _0342_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a211o_1
X_2658_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] _1824_ VGND VGND VPWR
+ VPWR _0278_ sky130_fd_sc_hd__or2_1
XFILLER_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout113 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[24\] VGND VGND VPWR VPWR net113
+ sky130_fd_sc_hd__buf_2
X_2589_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] _1801_ _1803_ VGND VGND VPWR
+ VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[12\] sky130_fd_sc_hd__a21oi_1
XANTENNA__2703__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout102 net103 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout135 net136 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_4
Xfanout146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
Xfanout124 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[11\] VGND VGND VPWR VPWR net124
+ sky130_fd_sc_hd__buf_2
XANTENNA__2703__B2 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout157 net158 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_59_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input1_A addr[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input57_A wdata[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_CLK clknet_2_1__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_3_CLK sky130_fd_sc_hd__clkbuf_8
X_1960_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[32\] _1290_ VGND VGND VPWR
+ VPWR _1453_ sky130_fd_sc_hd__nor2_1
XFILLER_53_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\]
+ _1379_ _1383_ _1381_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__a221o_1
X_3630_ _1052_ _1209_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__xor2_1
X_3561_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\]
+ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__or2_1
X_2512_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[4\]
+ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__or2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3492_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__nand2_1
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2443_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] VGND VGND VPWR VPWR
+ _1669_ sky130_fd_sc_hd__inv_2
X_2374_ net23 VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__inv_2
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4044_ clknet_leaf_33_CLK _0236_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_37_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3828_ clknet_leaf_12_CLK _0054_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3759_ clknet_leaf_17_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[19\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[19\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ net282 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] net104 VGND
+ VGND VPWR VPWR _0007_ sky130_fd_sc_hd__mux2_1
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2992_ _0575_ _0576_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1943_ _1434_ _1435_ _1620_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__a21oi_1
X_3613_ _1191_ _1195_ _1196_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__a21oi_1
X_1874_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__o21ai_1
X_3544_ _1117_ _1127_ _1124_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a21oi_1
X_3475_ _1057_ _1058_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nand2_2
X_2426_ net111 VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__inv_2
X_2357_ net279 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\] net94 VGND
+ VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
X_2288_ net277 net48 net82 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux2_1
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4027_ clknet_leaf_6_CLK _0219_ net139 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3260_ _0621_ _0836_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__xnor2_1
X_3191_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[11\] _1710_ VGND VGND VPWR
+ VPWR _0776_ sky130_fd_sc_hd__nand2_1
X_2211_ net209 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\] net100 VGND
+ VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2142_ net241 net37 net88 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__mux2_1
X_2073_ _1553_ _1554_ _1565_ _1536_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__o31a_1
XFILLER_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2975_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[46\]
+ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__nand2_1
X_1926_ _1407_ _1409_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1857_ _1113_ _1345_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__and3_1
XFILLER_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3527_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[5\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__and2_1
X_3458_ net111 _1716_ _0990_ _1004_ _1005_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__o2111a_1
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3389_ _1695_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[60\] VGND VGND VPWR
+ VPWR _0974_ sky130_fd_sc_hd__nor2_1
X_2409_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR _1635_
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_68_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2608__A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2815__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2291__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold60 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[19\] VGND VGND VPWR VPWR net263
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[60\] VGND VGND VPWR VPWR net285
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[48\] VGND VGND VPWR VPWR net274
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_89_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[15\] VGND VGND VPWR VPWR net296
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2806__B1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2282__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2760_ net108 _0370_ _0372_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[6\]
+ sky130_fd_sc_hd__a21oi_1
X_2691_ _1621_ _1802_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3312_ _0494_ _0892_ _0492_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3243_ _0824_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__nor2_1
XFILLER_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1848__A1 _1639_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3174_ _0690_ _0692_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__or2_1
XFILLER_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ net32 net31 net3 net4 VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_37_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2428__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2056_ _1646_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] _1546_ _1547_
+ _1548_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__a2111o_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2273__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2958_ _0517_ _0520_ _0524_ _0514_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__or4b_1
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1909_ _1646_ _1385_ _1397_ _1399_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__a31o_1
X_2889_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[61\]
+ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2102__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_3__f_CLK_A clknet_0_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input42_X net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2255__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3930_ clknet_leaf_9_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[26\] net140
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[26\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3861_ clknet_leaf_11_CLK _0087_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3792_ clknet_leaf_12_CLK _0019_ net159 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2812_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[23\] _0407_ VGND VGND VPWR VPWR
+ _0408_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_14_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2743_ myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.count_enable _0360_ VGND VGND VPWR VPWR
+ _0361_ sky130_fd_sc_hd__nand2_1
X_2674_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[0\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[0\]
+ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__xor2_1
XANTENNA__2711__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[6\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3226_ _0769_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or2_1
XFILLER_39_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3157_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0734_ _0735_ _0741_ VGND VGND
+ VPWR VPWR _0742_ sky130_fd_sc_hd__o211a_1
X_2108_ net330 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[25\] net107 VGND
+ VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux2_1
X_3088_ _0665_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__nand2_1
X_2039_ _1628_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\]
+ _1727_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2246__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2515__B net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_28_CLK_A clknet_2_2__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2390_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] VGND VGND VPWR VPWR
+ _1616_ sky130_fd_sc_hd__inv_2
X_4060_ clknet_leaf_6_CLK _0252_ net142 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_68_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3011_ _0591_ _0592_ _0594_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__or3_1
XFILLER_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_48_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3913_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[9\] net128
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[9\] sky130_fd_sc_hd__dfrtp_1
X_3844_ clknet_leaf_24_CLK _0070_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3874__RESET_B net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3775_ clknet_leaf_23_CLK _0002_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_2726_ _1658_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[4\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\]
+ _1668_ _0343_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__a221o_1
X_2657_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[22\] _1824_ VGND VGND VPWR
+ VPWR _0277_ sky130_fd_sc_hd__nand2_1
Xfanout103 _1591_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_4
X_2588_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[12\] _1801_ net74 VGND VGND VPWR
+ VPWR _1803_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout136 net169 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_2
Xfanout114 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[22\] VGND VGND VPWR VPWR net114
+ sky130_fd_sc_hd__buf_2
XFILLER_59_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout147 net168 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
Xfanout125 net126 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout169 net33 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_2
Xfanout158 net168 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_2
XFILLER_101_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3209_ _0501_ _0513_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__nor2_1
XFILLER_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2219__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[54\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout92_X net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1890_ _1382_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__inv_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3560_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[44\]
+ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__nand2_1
X_2511_ _1730_ _1732_ _1734_ _1736_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__and4_1
X_3491_ _1639_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[56\] _1065_ _1073_
+ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__o221a_1
XFILLER_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2442_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[13\] VGND VGND VPWR VPWR _1668_
+ sky130_fd_sc_hd__inv_2
XFILLER_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2373_ net341 net56 _1599_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_1
XANTENNA__2200__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4043_ clknet_leaf_33_CLK _0235_ net126 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4073__RESET_B net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2436__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[8\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3827_ clknet_leaf_12_CLK _0053_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3758_ clknet_leaf_18_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[18\]
+ net158 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] sky130_fd_sc_hd__dfrtp_4
X_2709_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[12\]
+ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__xor2_1
X_3689_ _1162_ _1272_ _1146_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_72_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2860__A1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[10\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2612__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[20\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2679__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[24\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2991_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nand2_1
X_1942_ _1150_ _1358_ _1361_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__nand3_1
XANTENNA__2603__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_1873_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[14\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\]
+ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[45\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[13\]
+ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__a22o_1
X_3612_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[25\] _1722_ _1195_ _1192_
+ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__a31o_1
X_3543_ _1614_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\] _1126_ VGND
+ VGND VPWR VPWR _1127_ sky130_fd_sc_hd__a21oi_1
X_3474_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__or2_1
X_2425_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[31\] VGND VGND VPWR VPWR _1651_
+ sky130_fd_sc_hd__inv_2
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2356_ net329 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] net94 VGND
+ VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2287_ net212 net47 net82 VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
X_4026_ clknet_leaf_4_CLK _0218_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2105__S net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2082__Y _1574_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3635__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[30\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2210_ net218 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[45\] net100 VGND
+ VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_59_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3190_ _0493_ _0774_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__nor2_1
X_2141_ net266 net36 net88 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_1
X_2072_ _1534_ _1564_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__nor2_1
XFILLER_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2974_ _0510_ _0513_ _0553_ _0558_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__a31oi_2
XANTENNA__2714__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[29\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_1925_ _1638_ _1405_ _1406_ _1409_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_60_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2588__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1856_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\]
+ _1098_ _1347_ _1096_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__a221o_1
X_3526_ _1095_ _1108_ _1093_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout102_A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3457_ _1653_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[33\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[32\]
+ _1652_ _0999_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__o221a_1
XFILLER_69_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2408_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] VGND VGND VPWR VPWR
+ _1634_ sky130_fd_sc_hd__inv_2
X_3388_ _0965_ _0969_ _0972_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__a21o_1
X_2339_ net286 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\] net93 VGND
+ VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4009_ clknet_leaf_32_CLK _0201_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2608__B myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2579__B1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2751__B1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold50 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[10\] VGND VGND VPWR VPWR net253
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input32_A addr[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[24\] VGND VGND VPWR VPWR net264
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[59\] VGND VGND VPWR VPWR net275
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold83 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[38\] VGND VGND VPWR VPWR net286
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold94 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[4\] VGND VGND VPWR VPWR net297
+ sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_11_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_89_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_8 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2690_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[7\] _1793_ _0284_ _0285_
+ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_20_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3311_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[15\] _0895_ VGND VGND VPWR VPWR
+ _0896_ sky130_fd_sc_hd__nand2_1
XFILLER_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3242_ _0638_ _0823_ _0473_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3298__A1 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3173_ _0633_ _0634_ _0643_ _0757_ _0756_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__o221a_1
XANTENNA__2709__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2124_ net7 net6 net12 net1 VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__or4_1
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2055_ myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\] _1719_ VGND VGND VPWR VPWR
+ _1548_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2957_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[4\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[36\]
+ _0538_ _0541_ _0540_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__a221o_1
X_1908_ _1391_ myPWM.g_pwm_channel\[1\].CHANNEL.alignment _1390_ _1400_ VGND VGND
+ VPWR VPWR _1401_ sky130_fd_sc_hd__and4b_1
X_2888_ _0471_ _0472_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__nand2_1
XFILLER_89_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout105_X net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3509_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[36\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[4\]
+ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__and2b_1
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2724__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_X net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ clknet_leaf_12_CLK _0086_ net161 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3791_ clknet_leaf_11_CLK _0018_ net157 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_2811_ net69 _0406_ _0407_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[22\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ _0339_ _0359_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2203__S net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2673_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[20\] myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[20\]
+ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2191__A1 net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3225_ _0595_ _0809_ _0804_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__o21a_1
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3156_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[2\] _0734_ _0732_ net109 VGND VGND
+ VPWR VPWR _0741_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2107_ net264 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[24\] net106 VGND
+ VGND VPWR VPWR _0024_ sky130_fd_sc_hd__mux2_1
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3087_ _0578_ _0603_ _0664_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__nand3_1
XFILLER_82_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2038_ _1625_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[46\] _1512_ VGND
+ VGND VPWR VPWR _1531_ sky130_fd_sc_hd__or3_1
XFILLER_22_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3989_ clknet_leaf_4_CLK _0181_ net135 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2706__B1 myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2182__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _1594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2173__A1 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3010_ _0592_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__nor2_1
XFILLER_64_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3912_ clknet_leaf_0_CLK myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[8\] net133
+ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[8\] sky130_fd_sc_hd__dfrtp_4
X_3843_ clknet_leaf_24_CLK _0069_ net151 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1987__A1 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[17\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__1987__B2 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2722__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[20\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_3774_ clknet_leaf_21_CLK _0001_ net153 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_2725_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[8\] _1662_ _1679_ net122
+ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a22o_1
X_2656_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[28\] _0266_ VGND VGND VPWR
+ VPWR _0276_ sky130_fd_sc_hd__nand2_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout104 _1574_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_4
X_2587_ _1802_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[11\]
+ sky130_fd_sc_hd__inv_2
XANTENNA__2164__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout137 net139 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_4
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout126 net134 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_4
Xfanout115 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR net115
+ sky130_fd_sc_hd__clkbuf_4
Xfanout159 net162 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net168 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3208_ _0787_ _0792_ _0791_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__o21ai_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3139_ myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[7\] _0722_ VGND VGND VPWR VPWR _0724_
+ sky130_fd_sc_hd__and2_1
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2155__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3182__B myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_X net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2366__X _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3490_ _1637_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[55\] _1060_ VGND
+ VGND VPWR VPWR _1074_ sky130_fd_sc_hd__or3_1
X_2510_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[9\] _1619_ _1631_ net115
+ _1735_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__o221a_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2441_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[13\] VGND VGND VPWR VPWR
+ _1667_ sky130_fd_sc_hd__inv_2
XFILLER_69_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2146__A1 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2372_ net339 net45 _1599_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XFILLER_96_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4042_ clknet_leaf_32_CLK _0234_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[39\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_37_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3826_ clknet_leaf_12_CLK _0052_ net160 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout132_A net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2452__A myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3757_ clknet_leaf_18_CLK myPWM.g_pwm_channel\[0\].CHANNEL.fcnt.next_state\[17\]
+ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[17\] sky130_fd_sc_hd__dfrtp_4
X_2708_ _1652_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[0\] _1682_ net121
+ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_12_CLK_A clknet_2_3__leaf_CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3688_ _1160_ _1270_ _1150_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__a21bo_1
XANTENNA__2137__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2639_ _1838_ VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[27\]
+ sky130_fd_sc_hd__inv_2
XFILLER_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input62_A wdata[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_76_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2301__S net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2300__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2990_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[21\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[53\]
+ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__or2_1
X_1941_ _1358_ _1361_ _1150_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__a21o_1
X_1872_ _1362_ _1363_ _1342_ _1343_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__a211o_1
X_3611_ _1193_ _1194_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__nand2_2
XANTENNA__2367__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3542_ _1614_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\]
+ _1612_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_94_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3473_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[59\]
+ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__nand2_1
XANTENNA__2702__A1_N myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[7\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2424_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[31\] VGND VGND VPWR VPWR
+ _1650_ sky130_fd_sc_hd__inv_2
XANTENNA__2211__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2355_ net277 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[54\] net94 VGND
+ VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2286_ net294 net46 net82 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
XANTENNA__3619__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[27\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_4025_ clknet_leaf_4_CLK _0217_ net137 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3809_ clknet_leaf_22_CLK _0035_ net152 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_69_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2530__B2 myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[19\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_85_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2349__A1 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[48\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2820__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input65_X net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2140_ net278 net35 net88 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
XFILLER_38_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2071_ _1533_ _1563_ _1550_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__o21a_1
XFILLER_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2973_ _0503_ _0508_ _0557_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[44\]
+ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[12\] VGND VGND VPWR VPWR _0558_
+ sky130_fd_sc_hd__a32o_2
XFILLER_34_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1924_ net114 _1404_ _1408_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__and3b_1
XANTENNA__2206__S net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1855_ _1098_ _1347_ _1096_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__a21oi_1
X_3525_ _1095_ _1108_ _1093_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a21oi_1
X_3456_ _0982_ _1039_ _0976_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o21ba_1
XFILLER_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3561__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[12\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_2407_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[19\] VGND VGND VPWR VPWR
+ _1633_ sky130_fd_sc_hd__inv_2
X_3387_ _0753_ _0758_ _0763_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__a31o_1
X_2338_ net291 myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[37\] net93 VGND
+ VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2269_ net310 net59 net80 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_55_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4008_ clknet_leaf_32_CLK _0200_ net129 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold40 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[10\] VGND VGND VPWR VPWR net243
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold51 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[25\] VGND VGND VPWR VPWR net254
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _0024_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 myPWM.g_pwm_channel\[0\].CHANNEL.data_buff\[21\] VGND VGND VPWR VPWR net276
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A addr[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold84 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[51\] VGND VGND VPWR VPWR net287
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 myPWM.g_pwm_channel\[1\].CHANNEL.data_buff\[46\] VGND VGND VPWR VPWR net298
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_71_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3310_ _0486_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3241_ _0473_ _0638_ _0823_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__a31o_1
X_3172_ _0634_ _0635_ _0642_ _0633_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__or4b_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2123_ net26 _1582_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__and2b_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2054_ _1646_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[60\] myPWM.g_pwm_channel\[1\].CHANNEL.f_count\[29\]
+ _1719_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_65_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2956_ _0528_ _0531_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__nor2_1
X_1907_ _1392_ _1393_ _1396_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__or4b_1
X_2887_ myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[31\] myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[63\]
+ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_35_CLK clknet_2_0__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_35_CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__3556__A myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[15\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2460__A myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[23\] VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3508_ myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[6\] myPWM.g_pwm_channel\[1\].CHANNEL.data_double_buff\[38\]
+ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__xor2_2
XANTENNA__2733__B2 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[18\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_3439_ _1011_ _1013_ _1018_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__a21boi_1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__2635__A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_26_CLK clknet_2_2__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_26_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_95_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2810_ net121 myPWM.g_pwm_channel\[0\].CHANNEL.f_count\[22\] _0402_ VGND VGND VPWR
+ VPWR _0407_ sky130_fd_sc_hd__and3_1
X_3790_ clknet_leaf_10_CLK _0017_ net156 VGND VGND VPWR VPWR myPWM.g_pwm_channel\[0\].CHANNEL.data_double_buff\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_70_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _0345_ _0347_ _0349_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_17_CLK clknet_2_3__leaf_CLK VGND VGND VPWR VPWR clknet_leaf_17_CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_68_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_2672_ _1627_ myPWM.g_pwm_channel\[1\].CHANNEL.fcnt.next_state\[16\] _0288_ _0289_
+ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__o221a_1
XFILLER_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3224_ _0591_ _0808_ _0805_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a21oi_1
.ends

