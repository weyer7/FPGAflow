VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpgacell
  CLASS BLOCK ;
  FOREIGN fpgacell ;
  ORIGIN 0.000 0.000 ;
  SIZE 210.000 BY 205.000 ;
  PIN CBeast_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 104.760 210.000 105.360 ;
    END
  END CBeast_in[0]
  PIN CBeast_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 159.160 210.000 159.760 ;
    END
  END CBeast_in[10]
  PIN CBeast_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 164.600 210.000 165.200 ;
    END
  END CBeast_in[11]
  PIN CBeast_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 170.040 210.000 170.640 ;
    END
  END CBeast_in[12]
  PIN CBeast_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 175.480 210.000 176.080 ;
    END
  END CBeast_in[13]
  PIN CBeast_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 180.920 210.000 181.520 ;
    END
  END CBeast_in[14]
  PIN CBeast_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 186.360 210.000 186.960 ;
    END
  END CBeast_in[15]
  PIN CBeast_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 110.200 210.000 110.800 ;
    END
  END CBeast_in[1]
  PIN CBeast_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 115.640 210.000 116.240 ;
    END
  END CBeast_in[2]
  PIN CBeast_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.808400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 206.000 121.080 210.000 121.680 ;
    END
  END CBeast_in[3]
  PIN CBeast_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 126.520 210.000 127.120 ;
    END
  END CBeast_in[4]
  PIN CBeast_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 131.960 210.000 132.560 ;
    END
  END CBeast_in[5]
  PIN CBeast_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 137.400 210.000 138.000 ;
    END
  END CBeast_in[6]
  PIN CBeast_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.808400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 206.000 142.840 210.000 143.440 ;
    END
  END CBeast_in[7]
  PIN CBeast_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 148.280 210.000 148.880 ;
    END
  END CBeast_in[8]
  PIN CBeast_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 206.000 153.720 210.000 154.320 ;
    END
  END CBeast_in[9]
  PIN CBeast_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 17.720 210.000 18.320 ;
    END
  END CBeast_out[0]
  PIN CBeast_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 72.120 210.000 72.720 ;
    END
  END CBeast_out[10]
  PIN CBeast_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 77.560 210.000 78.160 ;
    END
  END CBeast_out[11]
  PIN CBeast_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 83.000 210.000 83.600 ;
    END
  END CBeast_out[12]
  PIN CBeast_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 88.440 210.000 89.040 ;
    END
  END CBeast_out[13]
  PIN CBeast_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 93.880 210.000 94.480 ;
    END
  END CBeast_out[14]
  PIN CBeast_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 99.320 210.000 99.920 ;
    END
  END CBeast_out[15]
  PIN CBeast_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 23.160 210.000 23.760 ;
    END
  END CBeast_out[1]
  PIN CBeast_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 206.000 28.600 210.000 29.200 ;
    END
  END CBeast_out[2]
  PIN CBeast_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 34.040 210.000 34.640 ;
    END
  END CBeast_out[3]
  PIN CBeast_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 39.480 210.000 40.080 ;
    END
  END CBeast_out[4]
  PIN CBeast_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 44.920 210.000 45.520 ;
    END
  END CBeast_out[5]
  PIN CBeast_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 50.360 210.000 50.960 ;
    END
  END CBeast_out[6]
  PIN CBeast_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 55.800 210.000 56.400 ;
    END
  END CBeast_out[7]
  PIN CBeast_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 61.240 210.000 61.840 ;
    END
  END CBeast_out[8]
  PIN CBeast_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 206.000 66.680 210.000 67.280 ;
    END
  END CBeast_out[9]
  PIN CBnorth_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.830 201.000 32.110 205.000 ;
    END
  END CBnorth_in[0]
  PIN CBnorth_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.030 201.000 87.310 205.000 ;
    END
  END CBnorth_in[10]
  PIN CBnorth_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 92.550 201.000 92.830 205.000 ;
    END
  END CBnorth_in[11]
  PIN CBnorth_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 98.070 201.000 98.350 205.000 ;
    END
  END CBnorth_in[12]
  PIN CBnorth_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.590 201.000 103.870 205.000 ;
    END
  END CBnorth_in[13]
  PIN CBnorth_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.110 201.000 109.390 205.000 ;
    END
  END CBnorth_in[14]
  PIN CBnorth_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 114.630 201.000 114.910 205.000 ;
    END
  END CBnorth_in[15]
  PIN CBnorth_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 37.350 201.000 37.630 205.000 ;
    END
  END CBnorth_in[1]
  PIN CBnorth_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 42.870 201.000 43.150 205.000 ;
    END
  END CBnorth_in[2]
  PIN CBnorth_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.390 201.000 48.670 205.000 ;
    END
  END CBnorth_in[3]
  PIN CBnorth_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.910 201.000 54.190 205.000 ;
    END
  END CBnorth_in[4]
  PIN CBnorth_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.430 201.000 59.710 205.000 ;
    END
  END CBnorth_in[5]
  PIN CBnorth_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 64.950 201.000 65.230 205.000 ;
    END
  END CBnorth_in[6]
  PIN CBnorth_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.470 201.000 70.750 205.000 ;
    END
  END CBnorth_in[7]
  PIN CBnorth_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.990 201.000 76.270 205.000 ;
    END
  END CBnorth_in[8]
  PIN CBnorth_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.510 201.000 81.790 205.000 ;
    END
  END CBnorth_in[9]
  PIN CBnorth_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 120.150 201.000 120.430 205.000 ;
    END
  END CBnorth_out[0]
  PIN CBnorth_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 175.350 201.000 175.630 205.000 ;
    END
  END CBnorth_out[10]
  PIN CBnorth_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 180.870 201.000 181.150 205.000 ;
    END
  END CBnorth_out[11]
  PIN CBnorth_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 186.390 201.000 186.670 205.000 ;
    END
  END CBnorth_out[12]
  PIN CBnorth_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 191.910 201.000 192.190 205.000 ;
    END
  END CBnorth_out[13]
  PIN CBnorth_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 197.430 201.000 197.710 205.000 ;
    END
  END CBnorth_out[14]
  PIN CBnorth_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 201.000 203.230 205.000 ;
    END
  END CBnorth_out[15]
  PIN CBnorth_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 201.000 125.950 205.000 ;
    END
  END CBnorth_out[1]
  PIN CBnorth_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 131.190 201.000 131.470 205.000 ;
    END
  END CBnorth_out[2]
  PIN CBnorth_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 136.710 201.000 136.990 205.000 ;
    END
  END CBnorth_out[3]
  PIN CBnorth_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 142.230 201.000 142.510 205.000 ;
    END
  END CBnorth_out[4]
  PIN CBnorth_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 147.750 201.000 148.030 205.000 ;
    END
  END CBnorth_out[5]
  PIN CBnorth_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 153.270 201.000 153.550 205.000 ;
    END
  END CBnorth_out[6]
  PIN CBnorth_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 158.790 201.000 159.070 205.000 ;
    END
  END CBnorth_out[7]
  PIN CBnorth_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 201.000 164.590 205.000 ;
    END
  END CBnorth_out[8]
  PIN CBnorth_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 169.830 201.000 170.110 205.000 ;
    END
  END CBnorth_out[9]
  PIN SBsouth_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END SBsouth_in[0]
  PIN SBsouth_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END SBsouth_in[10]
  PIN SBsouth_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END SBsouth_in[11]
  PIN SBsouth_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END SBsouth_in[12]
  PIN SBsouth_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END SBsouth_in[13]
  PIN SBsouth_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END SBsouth_in[14]
  PIN SBsouth_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END SBsouth_in[15]
  PIN SBsouth_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END SBsouth_in[1]
  PIN SBsouth_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END SBsouth_in[2]
  PIN SBsouth_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END SBsouth_in[3]
  PIN SBsouth_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END SBsouth_in[4]
  PIN SBsouth_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END SBsouth_in[5]
  PIN SBsouth_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END SBsouth_in[6]
  PIN SBsouth_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END SBsouth_in[7]
  PIN SBsouth_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END SBsouth_in[8]
  PIN SBsouth_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END SBsouth_in[9]
  PIN SBsouth_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END SBsouth_out[0]
  PIN SBsouth_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END SBsouth_out[10]
  PIN SBsouth_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END SBsouth_out[11]
  PIN SBsouth_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END SBsouth_out[12]
  PIN SBsouth_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END SBsouth_out[13]
  PIN SBsouth_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END SBsouth_out[14]
  PIN SBsouth_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END SBsouth_out[15]
  PIN SBsouth_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END SBsouth_out[1]
  PIN SBsouth_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END SBsouth_out[2]
  PIN SBsouth_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END SBsouth_out[3]
  PIN SBsouth_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END SBsouth_out[4]
  PIN SBsouth_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END SBsouth_out[5]
  PIN SBsouth_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END SBsouth_out[6]
  PIN SBsouth_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END SBsouth_out[7]
  PIN SBsouth_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END SBsouth_out[8]
  PIN SBsouth_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END SBsouth_out[9]
  PIN SBwest_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END SBwest_in[0]
  PIN SBwest_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END SBwest_in[10]
  PIN SBwest_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END SBwest_in[11]
  PIN SBwest_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END SBwest_in[12]
  PIN SBwest_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END SBwest_in[13]
  PIN SBwest_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END SBwest_in[14]
  PIN SBwest_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END SBwest_in[15]
  PIN SBwest_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END SBwest_in[1]
  PIN SBwest_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END SBwest_in[2]
  PIN SBwest_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END SBwest_in[3]
  PIN SBwest_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END SBwest_in[4]
  PIN SBwest_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END SBwest_in[5]
  PIN SBwest_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END SBwest_in[6]
  PIN SBwest_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.995400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END SBwest_in[7]
  PIN SBwest_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END SBwest_in[8]
  PIN SBwest_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END SBwest_in[9]
  PIN SBwest_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END SBwest_out[0]
  PIN SBwest_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END SBwest_out[10]
  PIN SBwest_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END SBwest_out[11]
  PIN SBwest_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END SBwest_out[12]
  PIN SBwest_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END SBwest_out[13]
  PIN SBwest_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END SBwest_out[14]
  PIN SBwest_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END SBwest_out[15]
  PIN SBwest_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END SBwest_out[1]
  PIN SBwest_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END SBwest_out[2]
  PIN SBwest_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END SBwest_out[3]
  PIN SBwest_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END SBwest_out[4]
  PIN SBwest_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END SBwest_out[5]
  PIN SBwest_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END SBwest_out[6]
  PIN SBwest_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END SBwest_out[7]
  PIN SBwest_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END SBwest_out[8]
  PIN SBwest_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END SBwest_out[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 4.230 201.000 4.510 205.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 26.310 201.000 26.590 205.000 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.790 201.000 21.070 205.000 ;
    END
  END config_en
  PIN en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.750 201.000 10.030 205.000 ;
    END
  END en
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 15.270 201.000 15.550 205.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 193.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 204.480 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 204.480 181.510 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 193.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 193.360 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 204.480 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 204.480 184.810 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 204.430 193.310 ;
      LAYER li1 ;
        RECT 5.520 10.795 204.240 193.205 ;
      LAYER met1 ;
        RECT 4.210 6.500 207.850 195.800 ;
      LAYER met2 ;
        RECT 3.840 200.720 3.950 201.690 ;
        RECT 4.790 200.720 9.470 201.690 ;
        RECT 10.310 200.720 14.990 201.690 ;
        RECT 15.830 200.720 20.510 201.690 ;
        RECT 21.350 200.720 26.030 201.690 ;
        RECT 26.870 200.720 31.550 201.690 ;
        RECT 32.390 200.720 37.070 201.690 ;
        RECT 37.910 200.720 42.590 201.690 ;
        RECT 43.430 200.720 48.110 201.690 ;
        RECT 48.950 200.720 53.630 201.690 ;
        RECT 54.470 200.720 59.150 201.690 ;
        RECT 59.990 200.720 64.670 201.690 ;
        RECT 65.510 200.720 70.190 201.690 ;
        RECT 71.030 200.720 75.710 201.690 ;
        RECT 76.550 200.720 81.230 201.690 ;
        RECT 82.070 200.720 86.750 201.690 ;
        RECT 87.590 200.720 92.270 201.690 ;
        RECT 93.110 200.720 97.790 201.690 ;
        RECT 98.630 200.720 103.310 201.690 ;
        RECT 104.150 200.720 108.830 201.690 ;
        RECT 109.670 200.720 114.350 201.690 ;
        RECT 115.190 200.720 119.870 201.690 ;
        RECT 120.710 200.720 125.390 201.690 ;
        RECT 126.230 200.720 130.910 201.690 ;
        RECT 131.750 200.720 136.430 201.690 ;
        RECT 137.270 200.720 141.950 201.690 ;
        RECT 142.790 200.720 147.470 201.690 ;
        RECT 148.310 200.720 152.990 201.690 ;
        RECT 153.830 200.720 158.510 201.690 ;
        RECT 159.350 200.720 164.030 201.690 ;
        RECT 164.870 200.720 169.550 201.690 ;
        RECT 170.390 200.720 175.070 201.690 ;
        RECT 175.910 200.720 180.590 201.690 ;
        RECT 181.430 200.720 186.110 201.690 ;
        RECT 186.950 200.720 191.630 201.690 ;
        RECT 192.470 200.720 197.150 201.690 ;
        RECT 197.990 200.720 202.670 201.690 ;
        RECT 203.510 200.720 207.830 201.690 ;
        RECT 3.840 4.280 207.830 200.720 ;
        RECT 3.840 3.670 3.950 4.280 ;
        RECT 4.790 3.670 9.470 4.280 ;
        RECT 10.310 3.670 14.990 4.280 ;
        RECT 15.830 3.670 20.510 4.280 ;
        RECT 21.350 3.670 31.550 4.280 ;
        RECT 32.390 3.670 37.070 4.280 ;
        RECT 37.910 3.670 42.590 4.280 ;
        RECT 43.430 3.670 48.110 4.280 ;
        RECT 48.950 3.670 53.630 4.280 ;
        RECT 54.470 3.670 59.150 4.280 ;
        RECT 59.990 3.670 64.670 4.280 ;
        RECT 65.510 3.670 70.190 4.280 ;
        RECT 71.030 3.670 75.710 4.280 ;
        RECT 76.550 3.670 81.230 4.280 ;
        RECT 82.070 3.670 86.750 4.280 ;
        RECT 87.590 3.670 92.270 4.280 ;
        RECT 93.110 3.670 97.790 4.280 ;
        RECT 98.630 3.670 103.310 4.280 ;
        RECT 104.150 3.670 108.830 4.280 ;
        RECT 109.670 3.670 114.350 4.280 ;
        RECT 115.190 3.670 119.870 4.280 ;
        RECT 120.710 3.670 125.390 4.280 ;
        RECT 126.230 3.670 130.910 4.280 ;
        RECT 131.750 3.670 136.430 4.280 ;
        RECT 137.270 3.670 141.950 4.280 ;
        RECT 142.790 3.670 147.470 4.280 ;
        RECT 148.310 3.670 152.990 4.280 ;
        RECT 153.830 3.670 158.510 4.280 ;
        RECT 159.350 3.670 164.030 4.280 ;
        RECT 164.870 3.670 169.550 4.280 ;
        RECT 170.390 3.670 175.070 4.280 ;
        RECT 175.910 3.670 180.590 4.280 ;
        RECT 181.430 3.670 186.110 4.280 ;
        RECT 186.950 3.670 191.630 4.280 ;
        RECT 192.470 3.670 197.150 4.280 ;
        RECT 197.990 3.670 202.670 4.280 ;
        RECT 203.510 3.670 207.830 4.280 ;
      LAYER met3 ;
        RECT 3.990 187.360 207.855 194.985 ;
        RECT 4.400 185.960 205.600 187.360 ;
        RECT 3.990 181.920 207.855 185.960 ;
        RECT 4.400 180.520 205.600 181.920 ;
        RECT 3.990 176.480 207.855 180.520 ;
        RECT 4.400 175.080 205.600 176.480 ;
        RECT 3.990 171.040 207.855 175.080 ;
        RECT 4.400 169.640 205.600 171.040 ;
        RECT 3.990 165.600 207.855 169.640 ;
        RECT 4.400 164.200 205.600 165.600 ;
        RECT 3.990 160.160 207.855 164.200 ;
        RECT 4.400 158.760 205.600 160.160 ;
        RECT 3.990 154.720 207.855 158.760 ;
        RECT 4.400 153.320 205.600 154.720 ;
        RECT 3.990 149.280 207.855 153.320 ;
        RECT 4.400 147.880 205.600 149.280 ;
        RECT 3.990 143.840 207.855 147.880 ;
        RECT 4.400 142.440 205.600 143.840 ;
        RECT 3.990 138.400 207.855 142.440 ;
        RECT 4.400 137.000 205.600 138.400 ;
        RECT 3.990 132.960 207.855 137.000 ;
        RECT 4.400 131.560 205.600 132.960 ;
        RECT 3.990 127.520 207.855 131.560 ;
        RECT 4.400 126.120 205.600 127.520 ;
        RECT 3.990 122.080 207.855 126.120 ;
        RECT 4.400 120.680 205.600 122.080 ;
        RECT 3.990 116.640 207.855 120.680 ;
        RECT 4.400 115.240 205.600 116.640 ;
        RECT 3.990 111.200 207.855 115.240 ;
        RECT 4.400 109.800 205.600 111.200 ;
        RECT 3.990 105.760 207.855 109.800 ;
        RECT 4.400 104.360 205.600 105.760 ;
        RECT 3.990 100.320 207.855 104.360 ;
        RECT 4.400 98.920 205.600 100.320 ;
        RECT 3.990 94.880 207.855 98.920 ;
        RECT 4.400 93.480 205.600 94.880 ;
        RECT 3.990 89.440 207.855 93.480 ;
        RECT 4.400 88.040 205.600 89.440 ;
        RECT 3.990 84.000 207.855 88.040 ;
        RECT 4.400 82.600 205.600 84.000 ;
        RECT 3.990 78.560 207.855 82.600 ;
        RECT 4.400 77.160 205.600 78.560 ;
        RECT 3.990 73.120 207.855 77.160 ;
        RECT 4.400 71.720 205.600 73.120 ;
        RECT 3.990 67.680 207.855 71.720 ;
        RECT 4.400 66.280 205.600 67.680 ;
        RECT 3.990 62.240 207.855 66.280 ;
        RECT 4.400 60.840 205.600 62.240 ;
        RECT 3.990 56.800 207.855 60.840 ;
        RECT 4.400 55.400 205.600 56.800 ;
        RECT 3.990 51.360 207.855 55.400 ;
        RECT 4.400 49.960 205.600 51.360 ;
        RECT 3.990 45.920 207.855 49.960 ;
        RECT 4.400 44.520 205.600 45.920 ;
        RECT 3.990 40.480 207.855 44.520 ;
        RECT 4.400 39.080 205.600 40.480 ;
        RECT 3.990 35.040 207.855 39.080 ;
        RECT 4.400 33.640 205.600 35.040 ;
        RECT 3.990 29.600 207.855 33.640 ;
        RECT 4.400 28.200 205.600 29.600 ;
        RECT 3.990 24.160 207.855 28.200 ;
        RECT 4.400 22.760 205.600 24.160 ;
        RECT 3.990 18.720 207.855 22.760 ;
        RECT 4.400 17.320 205.600 18.720 ;
        RECT 3.990 9.695 207.855 17.320 ;
      LAYER met4 ;
        RECT 6.735 193.760 198.425 194.985 ;
        RECT 6.735 10.375 20.640 193.760 ;
        RECT 23.040 10.375 23.940 193.760 ;
        RECT 26.340 10.375 174.240 193.760 ;
        RECT 176.640 10.375 177.540 193.760 ;
        RECT 179.940 10.375 198.425 193.760 ;
  END
END fpgacell
END LIBRARY

