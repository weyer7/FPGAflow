VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpgacell
  CLASS BLOCK ;
  FOREIGN fpgacell ;
  ORIGIN 0.000 0.000 ;
  SIZE 185.000 BY 185.000 ;
  PIN CBeast_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 93.880 185.000 94.480 ;
    END
  END CBeast_in[0]
  PIN CBeast_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.082400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 181.000 148.280 185.000 148.880 ;
    END
  END CBeast_in[10]
  PIN CBeast_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 153.720 185.000 154.320 ;
    END
  END CBeast_in[11]
  PIN CBeast_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 181.000 159.160 185.000 159.760 ;
    END
  END CBeast_in[12]
  PIN CBeast_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 164.600 185.000 165.200 ;
    END
  END CBeast_in[13]
  PIN CBeast_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 99.320 185.000 99.920 ;
    END
  END CBeast_in[1]
  PIN CBeast_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 104.760 185.000 105.360 ;
    END
  END CBeast_in[2]
  PIN CBeast_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 181.000 110.200 185.000 110.800 ;
    END
  END CBeast_in[3]
  PIN CBeast_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 115.640 185.000 116.240 ;
    END
  END CBeast_in[4]
  PIN CBeast_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 121.080 185.000 121.680 ;
    END
  END CBeast_in[5]
  PIN CBeast_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 126.520 185.000 127.120 ;
    END
  END CBeast_in[6]
  PIN CBeast_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 131.960 185.000 132.560 ;
    END
  END CBeast_in[7]
  PIN CBeast_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 137.400 185.000 138.000 ;
    END
  END CBeast_in[8]
  PIN CBeast_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 142.840 185.000 143.440 ;
    END
  END CBeast_in[9]
  PIN CBeast_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 17.720 185.000 18.320 ;
    END
  END CBeast_out[0]
  PIN CBeast_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 72.120 185.000 72.720 ;
    END
  END CBeast_out[10]
  PIN CBeast_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 77.560 185.000 78.160 ;
    END
  END CBeast_out[11]
  PIN CBeast_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 83.000 185.000 83.600 ;
    END
  END CBeast_out[12]
  PIN CBeast_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 88.440 185.000 89.040 ;
    END
  END CBeast_out[13]
  PIN CBeast_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 23.160 185.000 23.760 ;
    END
  END CBeast_out[1]
  PIN CBeast_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 28.600 185.000 29.200 ;
    END
  END CBeast_out[2]
  PIN CBeast_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 34.040 185.000 34.640 ;
    END
  END CBeast_out[3]
  PIN CBeast_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 39.480 185.000 40.080 ;
    END
  END CBeast_out[4]
  PIN CBeast_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 44.920 185.000 45.520 ;
    END
  END CBeast_out[5]
  PIN CBeast_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 50.360 185.000 50.960 ;
    END
  END CBeast_out[6]
  PIN CBeast_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 55.800 185.000 56.400 ;
    END
  END CBeast_out[7]
  PIN CBeast_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 61.240 185.000 61.840 ;
    END
  END CBeast_out[8]
  PIN CBeast_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 66.680 185.000 67.280 ;
    END
  END CBeast_out[9]
  PIN CBnorth_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 27.690 181.000 27.970 185.000 ;
    END
  END CBnorth_in[0]
  PIN CBnorth_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.890 181.000 83.170 185.000 ;
    END
  END CBnorth_in[10]
  PIN CBnorth_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.410 181.000 88.690 185.000 ;
    END
  END CBnorth_in[11]
  PIN CBnorth_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 93.930 181.000 94.210 185.000 ;
    END
  END CBnorth_in[12]
  PIN CBnorth_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.450 181.000 99.730 185.000 ;
    END
  END CBnorth_in[13]
  PIN CBnorth_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 33.210 181.000 33.490 185.000 ;
    END
  END CBnorth_in[1]
  PIN CBnorth_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 181.000 39.010 185.000 ;
    END
  END CBnorth_in[2]
  PIN CBnorth_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 44.250 181.000 44.530 185.000 ;
    END
  END CBnorth_in[3]
  PIN CBnorth_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 181.000 50.050 185.000 ;
    END
  END CBnorth_in[4]
  PIN CBnorth_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 55.290 181.000 55.570 185.000 ;
    END
  END CBnorth_in[5]
  PIN CBnorth_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 60.810 181.000 61.090 185.000 ;
    END
  END CBnorth_in[6]
  PIN CBnorth_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 66.330 181.000 66.610 185.000 ;
    END
  END CBnorth_in[7]
  PIN CBnorth_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 71.850 181.000 72.130 185.000 ;
    END
  END CBnorth_in[8]
  PIN CBnorth_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 181.000 77.650 185.000 ;
    END
  END CBnorth_in[9]
  PIN CBnorth_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.970 181.000 105.250 185.000 ;
    END
  END CBnorth_out[0]
  PIN CBnorth_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.170 181.000 160.450 185.000 ;
    END
  END CBnorth_out[10]
  PIN CBnorth_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.690 181.000 165.970 185.000 ;
    END
  END CBnorth_out[11]
  PIN CBnorth_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 171.210 181.000 171.490 185.000 ;
    END
  END CBnorth_out[12]
  PIN CBnorth_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 176.730 181.000 177.010 185.000 ;
    END
  END CBnorth_out[13]
  PIN CBnorth_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.490 181.000 110.770 185.000 ;
    END
  END CBnorth_out[1]
  PIN CBnorth_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 181.000 116.290 185.000 ;
    END
  END CBnorth_out[2]
  PIN CBnorth_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.530 181.000 121.810 185.000 ;
    END
  END CBnorth_out[3]
  PIN CBnorth_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.050 181.000 127.330 185.000 ;
    END
  END CBnorth_out[4]
  PIN CBnorth_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.570 181.000 132.850 185.000 ;
    END
  END CBnorth_out[5]
  PIN CBnorth_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.090 181.000 138.370 185.000 ;
    END
  END CBnorth_out[6]
  PIN CBnorth_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.610 181.000 143.890 185.000 ;
    END
  END CBnorth_out[7]
  PIN CBnorth_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.130 181.000 149.410 185.000 ;
    END
  END CBnorth_out[8]
  PIN CBnorth_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 181.000 154.930 185.000 ;
    END
  END CBnorth_out[9]
  PIN SBsouth_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END SBsouth_in[0]
  PIN SBsouth_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END SBsouth_in[10]
  PIN SBsouth_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END SBsouth_in[11]
  PIN SBsouth_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END SBsouth_in[12]
  PIN SBsouth_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END SBsouth_in[13]
  PIN SBsouth_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END SBsouth_in[1]
  PIN SBsouth_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END SBsouth_in[2]
  PIN SBsouth_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END SBsouth_in[3]
  PIN SBsouth_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END SBsouth_in[4]
  PIN SBsouth_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END SBsouth_in[5]
  PIN SBsouth_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END SBsouth_in[6]
  PIN SBsouth_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END SBsouth_in[7]
  PIN SBsouth_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END SBsouth_in[8]
  PIN SBsouth_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END SBsouth_in[9]
  PIN SBsouth_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END SBsouth_out[0]
  PIN SBsouth_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END SBsouth_out[10]
  PIN SBsouth_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END SBsouth_out[11]
  PIN SBsouth_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END SBsouth_out[12]
  PIN SBsouth_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END SBsouth_out[13]
  PIN SBsouth_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END SBsouth_out[1]
  PIN SBsouth_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END SBsouth_out[2]
  PIN SBsouth_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END SBsouth_out[3]
  PIN SBsouth_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END SBsouth_out[4]
  PIN SBsouth_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END SBsouth_out[5]
  PIN SBsouth_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END SBsouth_out[6]
  PIN SBsouth_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END SBsouth_out[7]
  PIN SBsouth_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END SBsouth_out[8]
  PIN SBsouth_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END SBsouth_out[9]
  PIN SBwest_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END SBwest_in[0]
  PIN SBwest_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END SBwest_in[10]
  PIN SBwest_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END SBwest_in[11]
  PIN SBwest_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END SBwest_in[12]
  PIN SBwest_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END SBwest_in[13]
  PIN SBwest_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END SBwest_in[1]
  PIN SBwest_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END SBwest_in[2]
  PIN SBwest_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END SBwest_in[3]
  PIN SBwest_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END SBwest_in[4]
  PIN SBwest_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END SBwest_in[5]
  PIN SBwest_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END SBwest_in[6]
  PIN SBwest_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END SBwest_in[7]
  PIN SBwest_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END SBwest_in[8]
  PIN SBwest_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END SBwest_in[9]
  PIN SBwest_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END SBwest_out[0]
  PIN SBwest_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END SBwest_out[10]
  PIN SBwest_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END SBwest_out[11]
  PIN SBwest_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END SBwest_out[12]
  PIN SBwest_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END SBwest_out[13]
  PIN SBwest_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END SBwest_out[1]
  PIN SBwest_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END SBwest_out[2]
  PIN SBwest_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END SBwest_out[3]
  PIN SBwest_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END SBwest_out[4]
  PIN SBwest_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END SBwest_out[5]
  PIN SBwest_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END SBwest_out[6]
  PIN SBwest_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END SBwest_out[7]
  PIN SBwest_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END SBwest_out[8]
  PIN SBwest_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END SBwest_out[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 5.610 181.000 5.890 185.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.170 181.000 22.450 185.000 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 4.000 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.650 181.000 16.930 185.000 ;
    END
  END config_en
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 11.130 181.000 11.410 185.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2.420 4.640 4.020 179.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 172.420 4.640 174.020 179.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.420 4.640 181.940 6.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.420 174.640 181.940 176.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 5.720 5.200 7.320 179.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.720 5.200 177.320 179.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.980 7.940 181.940 9.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.980 177.940 181.940 179.540 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 3.030 5.355 181.890 179.605 ;
      LAYER li1 ;
        RECT 3.220 5.355 181.700 179.605 ;
      LAYER met1 ;
        RECT 0.070 0.380 183.010 182.880 ;
      LAYER met2 ;
        RECT 0.100 180.720 5.330 182.910 ;
        RECT 6.170 180.720 10.850 182.910 ;
        RECT 11.690 180.720 16.370 182.910 ;
        RECT 17.210 180.720 21.890 182.910 ;
        RECT 22.730 180.720 27.410 182.910 ;
        RECT 28.250 180.720 32.930 182.910 ;
        RECT 33.770 180.720 38.450 182.910 ;
        RECT 39.290 180.720 43.970 182.910 ;
        RECT 44.810 180.720 49.490 182.910 ;
        RECT 50.330 180.720 55.010 182.910 ;
        RECT 55.850 180.720 60.530 182.910 ;
        RECT 61.370 180.720 66.050 182.910 ;
        RECT 66.890 180.720 71.570 182.910 ;
        RECT 72.410 180.720 77.090 182.910 ;
        RECT 77.930 180.720 82.610 182.910 ;
        RECT 83.450 180.720 88.130 182.910 ;
        RECT 88.970 180.720 93.650 182.910 ;
        RECT 94.490 180.720 99.170 182.910 ;
        RECT 100.010 180.720 104.690 182.910 ;
        RECT 105.530 180.720 110.210 182.910 ;
        RECT 111.050 180.720 115.730 182.910 ;
        RECT 116.570 180.720 121.250 182.910 ;
        RECT 122.090 180.720 126.770 182.910 ;
        RECT 127.610 180.720 132.290 182.910 ;
        RECT 133.130 180.720 137.810 182.910 ;
        RECT 138.650 180.720 143.330 182.910 ;
        RECT 144.170 180.720 148.850 182.910 ;
        RECT 149.690 180.720 154.370 182.910 ;
        RECT 155.210 180.720 159.890 182.910 ;
        RECT 160.730 180.720 165.410 182.910 ;
        RECT 166.250 180.720 170.930 182.910 ;
        RECT 171.770 180.720 176.450 182.910 ;
        RECT 177.290 180.720 182.990 182.910 ;
        RECT 0.100 4.280 182.990 180.720 ;
        RECT 0.100 0.350 5.330 4.280 ;
        RECT 6.170 0.350 10.850 4.280 ;
        RECT 11.690 0.350 16.370 4.280 ;
        RECT 17.210 0.350 21.890 4.280 ;
        RECT 22.730 0.350 27.410 4.280 ;
        RECT 28.250 0.350 32.930 4.280 ;
        RECT 33.770 0.350 38.450 4.280 ;
        RECT 39.290 0.350 43.970 4.280 ;
        RECT 44.810 0.350 49.490 4.280 ;
        RECT 50.330 0.350 55.010 4.280 ;
        RECT 55.850 0.350 60.530 4.280 ;
        RECT 61.370 0.350 66.050 4.280 ;
        RECT 66.890 0.350 71.570 4.280 ;
        RECT 72.410 0.350 77.090 4.280 ;
        RECT 77.930 0.350 82.610 4.280 ;
        RECT 83.450 0.350 88.130 4.280 ;
        RECT 88.970 0.350 93.650 4.280 ;
        RECT 94.490 0.350 99.170 4.280 ;
        RECT 100.010 0.350 104.690 4.280 ;
        RECT 105.530 0.350 110.210 4.280 ;
        RECT 111.050 0.350 115.730 4.280 ;
        RECT 116.570 0.350 121.250 4.280 ;
        RECT 122.090 0.350 126.770 4.280 ;
        RECT 127.610 0.350 132.290 4.280 ;
        RECT 133.130 0.350 137.810 4.280 ;
        RECT 138.650 0.350 143.330 4.280 ;
        RECT 144.170 0.350 148.850 4.280 ;
        RECT 149.690 0.350 154.370 4.280 ;
        RECT 155.210 0.350 159.890 4.280 ;
        RECT 160.730 0.350 165.410 4.280 ;
        RECT 166.250 0.350 170.930 4.280 ;
        RECT 171.770 0.350 176.450 4.280 ;
        RECT 177.290 0.350 182.990 4.280 ;
      LAYER met3 ;
        RECT 0.525 165.600 183.015 180.705 ;
        RECT 4.400 164.200 180.600 165.600 ;
        RECT 0.525 160.160 183.015 164.200 ;
        RECT 4.400 158.760 180.600 160.160 ;
        RECT 0.525 154.720 183.015 158.760 ;
        RECT 4.400 153.320 180.600 154.720 ;
        RECT 0.525 149.280 183.015 153.320 ;
        RECT 4.400 147.880 180.600 149.280 ;
        RECT 0.525 143.840 183.015 147.880 ;
        RECT 4.400 142.440 180.600 143.840 ;
        RECT 0.525 138.400 183.015 142.440 ;
        RECT 4.400 137.000 180.600 138.400 ;
        RECT 0.525 132.960 183.015 137.000 ;
        RECT 4.400 131.560 180.600 132.960 ;
        RECT 0.525 127.520 183.015 131.560 ;
        RECT 4.400 126.120 180.600 127.520 ;
        RECT 0.525 122.080 183.015 126.120 ;
        RECT 4.400 120.680 180.600 122.080 ;
        RECT 0.525 116.640 183.015 120.680 ;
        RECT 4.400 115.240 180.600 116.640 ;
        RECT 0.525 111.200 183.015 115.240 ;
        RECT 4.400 109.800 180.600 111.200 ;
        RECT 0.525 105.760 183.015 109.800 ;
        RECT 4.400 104.360 180.600 105.760 ;
        RECT 0.525 100.320 183.015 104.360 ;
        RECT 4.400 98.920 180.600 100.320 ;
        RECT 0.525 94.880 183.015 98.920 ;
        RECT 4.400 93.480 180.600 94.880 ;
        RECT 0.525 89.440 183.015 93.480 ;
        RECT 4.400 88.040 180.600 89.440 ;
        RECT 0.525 84.000 183.015 88.040 ;
        RECT 4.400 82.600 180.600 84.000 ;
        RECT 0.525 78.560 183.015 82.600 ;
        RECT 4.400 77.160 180.600 78.560 ;
        RECT 0.525 73.120 183.015 77.160 ;
        RECT 4.400 71.720 180.600 73.120 ;
        RECT 0.525 67.680 183.015 71.720 ;
        RECT 4.400 66.280 180.600 67.680 ;
        RECT 0.525 62.240 183.015 66.280 ;
        RECT 4.400 60.840 180.600 62.240 ;
        RECT 0.525 56.800 183.015 60.840 ;
        RECT 4.400 55.400 180.600 56.800 ;
        RECT 0.525 51.360 183.015 55.400 ;
        RECT 4.400 49.960 180.600 51.360 ;
        RECT 0.525 45.920 183.015 49.960 ;
        RECT 4.400 44.520 180.600 45.920 ;
        RECT 0.525 40.480 183.015 44.520 ;
        RECT 4.400 39.080 180.600 40.480 ;
        RECT 0.525 35.040 183.015 39.080 ;
        RECT 4.400 33.640 180.600 35.040 ;
        RECT 0.525 29.600 183.015 33.640 ;
        RECT 4.400 28.200 180.600 29.600 ;
        RECT 0.525 24.160 183.015 28.200 ;
        RECT 4.400 22.760 180.600 24.160 ;
        RECT 0.525 18.720 183.015 22.760 ;
        RECT 4.400 17.320 180.600 18.720 ;
        RECT 0.525 4.935 183.015 17.320 ;
      LAYER met4 ;
        RECT 1.215 180.160 171.745 180.705 ;
        RECT 1.215 4.935 2.020 180.160 ;
        RECT 4.420 4.935 5.320 180.160 ;
        RECT 7.720 4.935 171.745 180.160 ;
  END
END fpgacell
END LIBRARY

